// Verilog netlist produced by program LSE :  version Diamond Version 0.0.0
// Netlist written on Wed Jul 29 16:42:05 2020
//
// Verilog Description of module TinyFPGA_B
//

module TinyFPGA_B (CLK, LED, USBPU, ENCODER0_A, ENCODER0_B, ENCODER1_A, 
            ENCODER1_B, HALL1, HALL2, HALL3, FAULT_N, NEOPXL, DE, 
            TX, RX, CS_CLK, CS, CS_MISO, SCL, SDA, INLC, INHC, 
            INLB, INHB, INLA, INHA) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(2[8:18])
    input CLK;   // verilog/TinyFPGA_B.v(3[9:12])
    output LED;   // verilog/TinyFPGA_B.v(4[10:13])
    output USBPU;   // verilog/TinyFPGA_B.v(5[10:15])
    input ENCODER0_A;   // verilog/TinyFPGA_B.v(6[9:19])
    input ENCODER0_B;   // verilog/TinyFPGA_B.v(7[9:19])
    input ENCODER1_A;   // verilog/TinyFPGA_B.v(8[9:19])
    input ENCODER1_B;   // verilog/TinyFPGA_B.v(9[9:19])
    input HALL1 /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(10[9:14])
    input HALL2 /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(11[9:14])
    input HALL3 /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(12[9:14])
    input FAULT_N;   // verilog/TinyFPGA_B.v(13[9:16])
    output NEOPXL;   // verilog/TinyFPGA_B.v(14[10:16])
    output DE;   // verilog/TinyFPGA_B.v(15[10:12])
    output TX /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(16[10:12])
    input RX;   // verilog/TinyFPGA_B.v(17[9:11])
    output CS_CLK;   // verilog/TinyFPGA_B.v(18[10:16])
    output CS;   // verilog/TinyFPGA_B.v(19[10:12])
    input CS_MISO;   // verilog/TinyFPGA_B.v(20[9:16])
    inout SCL /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(21[9:12])
    inout SDA /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(22[9:12])
    output INLC;   // verilog/TinyFPGA_B.v(23[10:14])
    output INHC;   // verilog/TinyFPGA_B.v(24[10:14])
    output INLB;   // verilog/TinyFPGA_B.v(25[10:14])
    output INHB;   // verilog/TinyFPGA_B.v(26[10:14])
    output INLA;   // verilog/TinyFPGA_B.v(27[10:14])
    output INHA;   // verilog/TinyFPGA_B.v(28[10:14])
    
    wire clk16MHz /* synthesis SET_AS_NETWORK=clk16MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[16:24])
    
    wire GND_net, VCC_net, LED_c, ENCODER0_A_N, ENCODER0_B_N, ENCODER1_A_N, 
        ENCODER1_B_N, NEOPXL_c, DE_c, RX_c, CS_CLK_c, CS_c, CS_MISO_c, 
        INLC_c_0, INHC_c_0, INLB_c_0, INHB_c_0, INLA_c_0, INHA_c_0;
    wire [7:0]ID;   // verilog/TinyFPGA_B.v(46[12:14])
    
    wire reset;
    wire [23:0]neopxl_color;   // verilog/TinyFPGA_B.v(49[13:25])
    
    wire hall1, hall2, hall3, pwm_out, dir, GHA, n51002, GHB, 
        GHC;
    wire [23:0]pwm_setpoint;   // verilog/TinyFPGA_B.v(95[20:32])
    wire [23:0]duty;   // verilog/TinyFPGA_B.v(96[21:25])
    
    wire n51926;
    wire [7:0]commutation_state;   // verilog/TinyFPGA_B.v(131[12:29])
    
    wire n51925;
    wire [7:0]commutation_state_prev;   // verilog/TinyFPGA_B.v(132[12:34])
    
    wire dti;
    wire [7:0]dti_counter;   // verilog/TinyFPGA_B.v(141[12:23])
    
    wire tx_o, tx_enable;
    wire [23:0]encoder0_position_scaled;   // verilog/TinyFPGA_B.v(238[21:45])
    wire [23:0]encoder1_position_scaled;   // verilog/TinyFPGA_B.v(240[21:45])
    wire [23:0]displacement;   // verilog/TinyFPGA_B.v(241[21:33])
    wire [23:0]setpoint;   // verilog/TinyFPGA_B.v(242[22:30])
    wire [23:0]Kp;   // verilog/TinyFPGA_B.v(243[22:24])
    wire [23:0]Ki;   // verilog/TinyFPGA_B.v(244[22:24])
    wire [7:0]control_mode;   // verilog/TinyFPGA_B.v(246[14:26])
    wire [23:0]PWMLimit;   // verilog/TinyFPGA_B.v(247[22:30])
    wire [23:0]IntegralLimit;   // verilog/TinyFPGA_B.v(248[22:35])
    wire [23:0]deadband;   // verilog/TinyFPGA_B.v(249[22:30])
    wire [15:0]current;   // verilog/TinyFPGA_B.v(250[22:29])
    wire [15:0]current_limit;   // verilog/TinyFPGA_B.v(251[22:35])
    wire [31:0]baudrate;   // verilog/TinyFPGA_B.v(253[15:23])
    wire [23:0]motor_state;   // verilog/TinyFPGA_B.v(282[22:33])
    
    wire n63351, data_ready, sda_out, sda_enable, scl, scl_enable;
    wire [31:0]delay_counter;   // verilog/TinyFPGA_B.v(351[11:24])
    wire [2:0]\ID_READOUT_FSM.state ;   // verilog/TinyFPGA_B.v(359[15:20])
    
    wire pwm_setpoint_23__N_207, n12171, n12175, n51924, n51364, n51670, 
        n51363, n51923, n6, n260, n51669, n12211, n294, n67828, 
        n51212, n298, n299, n300, n301, n302, n303, n304, n305, 
        n306, n307, n308, n309, n51922, n51921, n15, n4926, 
        n4925, n4924, n4923, n4922, n4921, n4920, n4919, n4918, 
        n4917, n4916, n4915, n4914, n51362, n51001;
    wire [23:0]pwm_setpoint_23__N_3;
    
    wire n51000, n60362, n51211, n69234, n51361;
    wire [7:0]commutation_state_7__N_208;
    
    wire n51920, commutation_state_7__N_216;
    wire [7:0]commutation_state_7__N_27;
    
    wire n29898;
    wire [31:0]encoder0_position;   // verilog/TinyFPGA_B.v(237[11:28])
    
    wire GHA_N_355, GLA_N_372, GHB_N_377, GLB_N_386, GHC_N_391, GLC_N_400, 
        dti_N_404, n29895, n29892, RX_N_2, n4, n67822, n67818, 
        n67816, n67810, n67804, n1744, n1742;
    wire [31:0]motor_state_23__N_91;
    wire [32:0]encoder0_position_scaled_23__N_43;
    wire [23:0]displacement_23__N_67;
    
    wire n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, 
        n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, 
        n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, 
        n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, 
        read_N_409, n7, n36816, n1319, n66810, n29890, n17, n16, 
        n15_adj_5693, n13, n12, n11, n10, n9, n8, n7_adj_5694, 
        n6_adj_5695, n5, n4_adj_5696, n24, n69231, n19, n17_adj_5697, 
        n16_adj_5698, n15_adj_5699, n51919, n1784, n1786, n1788, 
        n1790, n1792, n1794, n1796;
    wire [31:0]encoder1_position;   // verilog/TinyFPGA_B.v(239[11:28])
    
    wire n1822, n1824;
    wire [10:0]timer;   // verilog/neopixel.v(9[12:17])
    wire [1:0]state;   // verilog/neopixel.v(16[11:16])
    wire [4:0]bit_ctr;   // verilog/neopixel.v(17[11:18])
    wire [10:0]\neo_pixel_transmitter.t0 ;   // verilog/neopixel.v(27[14:16])
    wire [5:0]color_bit_N_502;
    
    wire n4913, n4912, n4911, n4910, n4909, n4908, n63339, n50985, 
        n63335, n4938, n4935, n29885, n29881, n43683, n29878, 
        n13_adj_5700, n11_adj_5701, n9_adj_5702, n8_adj_5703, n7_adj_5704, 
        n6_adj_5705, n5_adj_5706, n4_adj_5707, n71090;
    wire [23:0]pwm_counter;   // verilog/pwm.v(11[19:30])
    
    wire n19_adj_5708, n25, n24_adj_5709, n23, n22, n21, n20, 
        n51668, n69232, n51667, n51918, n51917, n51916, n51915, 
        n51666, n51360, n51914, n51913, n51665, n51664, n51663, 
        n51359, n2, n51662, n51912, n625, n51661, n14, n15_adj_5710, 
        n16_adj_5711, n17_adj_5712, n18, n19_adj_5713, n20_adj_5714, 
        n21_adj_5715, n22_adj_5716, n23_adj_5717, n24_adj_5718, n25_adj_5719, 
        n5772, n51911, n51358, rx_data_ready;
    wire [7:0]rx_data;   // verilog/coms.v(94[13:20])
    
    wire n51357;
    wire [7:0]\data_in_frame[23] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[21] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[20] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[18] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[17] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[16] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[12] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[11] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[8] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[7] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[6] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[5] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[4] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[3] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[1] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[0] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_out_frame[27] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[26] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[25] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[24] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[23] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[22] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[21] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[20] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[19] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[18] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[17] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[16] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[15] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[14] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[13] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[12] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[11] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[10] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[9] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[8] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[7] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[6] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[5] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[4] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[3] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[1] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[0] ;   // verilog/coms.v(100[12:26])
    wire [7:0]byte_transmit_counter;   // verilog/coms.v(105[12:33])
    
    wire tx_active, n51660;
    wire [31:0]\FRAME_MATCHER.state ;   // verilog/coms.v(115[11:16])
    wire [31:0]\FRAME_MATCHER.i ;   // verilog/coms.v(118[11:12])
    
    wire \FRAME_MATCHER.rx_data_ready_prev , n51356, n2820, n51910, 
        n51659, n51909, n51355, n51908, n5_adj_5720, n51907, n51658, 
        n51354, n50999, n2873, n51906, n51657, n63329, n51656, 
        n51905, n51655, n63327, n51353, n51654, n51904, n51653, 
        n51903, n4907, n4906, n4905, n3157, n51652, n51902, n51651, 
        n55096, n58627, n58626, n58625, n58624, n58623, n58622, 
        n58621, n58496, n58620, n58619, n58618, n58617, n58616, 
        n58615, n58614, n58613, n58612, n58611, n58610, n58609, 
        n58608, n58607, n58606, n58605, n58604, n58603, n58602, 
        n58601, n58600, n58599, n58598, n58597, n58596, n58595, 
        n58594, n58593, n58592, n58591, n58590, n28975, n58589, 
        n58588, n58587, n58586, n58585, n58584, n58583, n58582, 
        n58581, n58580, n58579, n58578, n58577, n58576, n58575, 
        n28959, n58574, n58573, n58572, n58571, n58570, n58569, 
        n58568, n58567, n58566, n58565, n58497, n28947, n58500, 
        n28945, n58501, n58502, n58504, n58506, n58508, n58509, 
        n58510, n58511, n58512, n58513, n58514, n58515, n58494, 
        n58516, n58517, n28929, n28928, n58518, n58519, n58520, 
        n58521, n58522, n58523, n28921, n58524, n58525, n58526, 
        n58527, n58528, n58529, n58530, n58531, n58532, n58533, 
        n58534, n58535, n58536, n58537, n58493, n58538, n58539, 
        n28903, n58540, n58541, n58495, n58542, n58543, n58544, 
        n58545, n28895, n28894, n58546, n58547, n58548, n58549, 
        n58550, n58551, n58552, n58553, n58505, n58499, n58554, 
        n58555, n58556, n58557, n58558, n58498, n58503, n58559, 
        n58560, n58561, n58562, n58563, n58564, n63321, n54456, 
        n68910, n63319, n42369, n57916, n50984, n51901, n51900, 
        n51899, n51898, n63311, n51897, n51896, n70503, n51895, 
        n51894, n51893, n51892, n51891, n51890, n51335, n51334, 
        n51333, n51332, n51331, n51330, n51889, n51888, n51887, 
        n51886, n51885, n51884, n51883, n51329, n51328, n51882, 
        n51881, n51327, n51326, n51880, n51879, n51878, n50998, 
        n51877, n63301, n68596, n51325, n51324, n51323, n51322, 
        n51876, n50997, n50983, n51875, n51874, n51873, n51872, 
        n51871, n51609, n51608, n51321, n51320, n51607, n51606, 
        n51605, n51319, n51870, n51318, n51869, n51604, n51603, 
        n51868, n51867, n51866, n51602, n51317, n51601, n51865, 
        n51316, n51600, n51864, n50996, n51315, n51314, n51863, 
        n51599, n51598, n51313, n42994, n42941, n68590, n43055, 
        n50982, n42981, n42913, n51862, n51597, n51596, n51595, 
        n51861, n51594, n51312, n51860, n50687, n51593, n51592, 
        n51859, n51311, n51591, n51858, n2076, n51310, n51309, 
        n51857, n51856, n51855, n51854, n42885, n2217, n6_adj_5721, 
        n68576, n63295, n63289, n57918, n71072, n71066, n15_adj_5722, 
        Kp_23__N_748, n63283, n63279, n63277, n29861, n29858, n12209, 
        n25764, n70241, n68906, n63257, n63251, n63245, n63239, 
        n63237, n12173, n29855, n32, n31, n30, n29, n28, n29851, 
        n27, n26, n25_adj_5723, n24_adj_5724, n23_adj_5725, n63229, 
        n22_adj_5726, n21_adj_5727, n20_adj_5728, n19_adj_5729, n18_adj_5730, 
        n17_adj_5731, n16_adj_5732, n63219, \FRAME_MATCHER.i_31__N_2509 , 
        n5_adj_5733, n5_adj_5734, n51308, n50995, n69308, n51307, 
        n63215, n43543, n29786, n63209, n29771, n29765, n29764, 
        n43723, n29756, n29674, n29668, n43719, n15_adj_5735, n43717, 
        n29650, n29649, n29648, n29647, n29643, n29642, n29639, 
        n29638, n29637, n29636, n29635, n29634, n29633, n29632, 
        n29631, n29630, n29629, n29628, n29627, n29626, n29625, 
        n29624, n29623, n29622, n29621, n29618, n29617, n29616, 
        n29615, n29614, n29613, n29612, n43715, n29608, n29607, 
        n29606, n29605, n29604, n29602, n43713, n29595, n43709, 
        n43605, n43601, n29583, n29582, n29581, n29578, n43595, 
        n29575, n29574, n29573, n29570, n29567, n29566, n29565, 
        n29563, n29562, n29560, n29558, n29557, n29556, n43695, 
        n29551, n29550, n29549, n29548, n29547, n29546, n29545, 
        n29542, n29539, n29538, n43747, n29535, n29530, n29529, 
        n29523, n29520, n63207, n43679, n43677, n43691, n43689, 
        n29474, n29468, n57852, n58957, n57874, n57876, n57878, 
        n30_adj_5736, n70477, n14_adj_5737, n13_adj_5738, n12_adj_5739, 
        n11_adj_5740, n69436, n23_adj_5741, n21_adj_5742, n19_adj_5743, 
        n17_adj_5744, n16_adj_5745, n15_adj_5746, n13_adj_5747, n11_adj_5748, 
        n10_adj_5749, n9_adj_5750, n8_adj_5751, n7_adj_5752, n6_adj_5753, 
        n4_adj_5754, n25411, n58492, n51306, n51853, n15_adj_5755, 
        n54620, n4_adj_5756, n4_adj_5757, n63191, n10_adj_5758, n6_adj_5759, 
        n30510, n30494, n522, control_update;
    wire [23:0]\PID_CONTROLLER.integral ;   // verilog/motorControl.v(35[23:31])
    
    wire n6_adj_5760, n30439, n30438, n30437, n63185, n51852, n155, 
        n212, n213, n214, n219, n230;
    wire [23:0]\PID_CONTROLLER.integral_23__N_3715 ;
    
    wire n361, n367, n375, n376, n401, n10_adj_5761, n455, n456, 
        n30424, n30421, n30420, n30416, n6_adj_5762, n30410, n57996, 
        n51305, n30406, n43501, n15_adj_5763, n11_adj_5764, n10_adj_5765, 
        n521;
    wire [1:0]a_new;   // vhdl/quadrature_decoder.vhd(39[9:14])
    wire [1:0]b_new;   // vhdl/quadrature_decoder.vhd(40[9:14])
    
    wire a_prev, b_prev, debounce_cnt_N_3833, n30391, position_31__N_3836, 
        n30387, n520, n519, n518, n63179, n63177, n30386, n9_adj_5766, 
        n30385, n30384, n30383, n30382, n30381, n30380, n30379, 
        n30378, n30377, n30376, n30374, n30372, n30371, n30370, 
        n30369, n30368, n30367, n30366, n61361, n30365, n30364, 
        n30363, n8_adj_5767;
    wire [1:0]a_new_adj_5996;   // vhdl/quadrature_decoder.vhd(39[9:14])
    wire [1:0]b_new_adj_5997;   // vhdl/quadrature_decoder.vhd(40[9:14])
    
    wire a_prev_adj_5770, b_prev_adj_5771, debounce_cnt_N_3833_adj_5772, 
        position_31__N_3836_adj_5773, n405, n404, n403, n402, n7_adj_5774, 
        n63159, n6_adj_5775;
    wire [7:0]data_adj_6007;   // verilog/eeprom.v(23[12:16])
    
    wire ready_prev, rw;
    wire [7:0]state_adj_6008;   // verilog/eeprom.v(27[11:16])
    
    wire n51851;
    wire [7:0]state_7__N_3918;
    
    wire n8_adj_5778, n5_adj_5779, n4_adj_5780, n3, n2_adj_5781, n71060, 
        n71054, n30330, n30329, n30328, n59702, n63153, n30327, 
        n30326, n30325, n30324, n30323, n6615, n30319, n30318, 
        n30317, n63147, n30316, n30315, n30313, n30312, n51850, 
        n30311, n30310, n30309, n30308, n30305, n51849, n63145, 
        n4904, n4903, clk_out;
    wire [15:0]data_adj_6015;   // verilog/tli4970.v(27[14:18])
    wire [7:0]state_adj_6017;   // verilog/tli4970.v(29[13:18])
    
    wire n19_adj_5792, n18_adj_5793, n17_adj_5794, n4_adj_5795, n3_adj_5796, 
        n2_adj_5797, n63135, n30273, n63131, n30255, n12177, n12179, 
        n12181, n12183, n8_adj_5798, state_7__N_4319, n16_adj_5799, 
        n30238, n30237, n30236, n30235, n30234, n30233, n30232, 
        n30231, n30230, n43725, n14_adj_5800, n8_adj_5801, n30224, 
        n59656, n30218, n61472, n59648, n10_adj_5802, r_Rx_Data;
    wire [7:0]r_Clock_Count;   // verilog/uart_rx.v(33[17:30])
    wire [2:0]r_Bit_Index;   // verilog/uart_rx.v(34[17:28])
    wire [2:0]r_SM_Main;   // verilog/uart_rx.v(37[17:26])
    
    wire n59644, n22835, n12185, n12187, n12189, n12191, n12193, 
        n12195, n12197, n12199, n30205, n59638;
    wire [24:0]o_Rx_DV_N_3488;
    
    wire n71048, n12201, n12203, n12205, n12207;
    wire [2:0]r_SM_Main_2__N_3446;
    
    wire n15_adj_5803, n30199, n14_adj_5804, n13_adj_5805, n12_adj_5806, 
        n30198, n63119;
    wire [2:0]r_SM_Main_adj_6027;   // verilog/uart_tx.v(32[16:25])
    wire [8:0]r_Clock_Count_adj_6028;   // verilog/uart_tx.v(33[16:29])
    
    wire n63115, n51848, n51304, n51303, n63113;
    wire [2:0]r_SM_Main_2__N_3536;
    
    wire n58108, n11_adj_5817, n10_adj_5818, n9_adj_5819, n8_adj_5820, 
        n7_adj_5821, n6_adj_5822, n30169, n61577;
    wire [7:0]state_adj_6041;   // verilog/i2c_controller.v(33[12:17])
    
    wire n68341;
    wire [7:0]saved_addr;   // verilog/i2c_controller.v(34[12:22])
    
    wire enable_slow_N_4213, n63109, n5_adj_5824, n30154, n5_adj_5825, 
        n51302;
    wire [7:0]state_7__N_4110;
    
    wire n29432, n6426, n51301, n20181;
    wire [7:0]state_7__N_4126;
    
    wire n30139, n30134, n54490, n29426, n30133, n30132, n30131, 
        n30130, n30129, n30128, n30126, n29423, n29420, n29417, 
        n58978, n30125, n30124, n30123, n30122, n30121, n30120, 
        n63103, n29410, n7447, n7446, n7445, n7444, n7443, n7442, 
        n828, n829, n830, n831, n832, n833, n861, n7_adj_5826, 
        n896, n897, n898, n899, n900, n901, n927, n928, n929, 
        n930, n931, n932, n933, n937, n938, n939, n940, n941, 
        n942, n943, n944, n945, n946, n947, n948, n949, n950, 
        n951, n952, n953, n954, n955, n956, n957, n960, n995, 
        n996, n997, n998, n999, n1000, n1001, n60815, n63085, 
        n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, 
        n1059, n63083, n1093, n1094, n1095, n1096, n1097, n1098, 
        n1099, n1100, n1101, n63079, n1125, n1126, n1127, n1128, 
        n1129, n1130, n1131, n1132, n1133, n12_adj_5827, n1158, 
        n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, 
        n1201, n1224_adj_5828, n1225_adj_5829, n1226_adj_5830, n1227_adj_5831, 
        n1228_adj_5832, n1229_adj_5833, n1230_adj_5834, n1231_adj_5835, 
        n1232_adj_5836, n1233_adj_5837, n18_adj_5838, n17_adj_5839, 
        n1257, n16_adj_5840, n14_adj_5841, n12_adj_5842, n1292, n1293, 
        n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, 
        n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, 
        n1331, n1332, n1333, n41634, n41635, n1356, n1391, n1392, 
        n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, 
        n1401, n1422, n1423, n1424, n1425, n1426, n1427, n1428, 
        n1429, n1430, n1431, n1432, n1433, n1455, n1490, n1491, 
        n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, 
        n1500, n1501, n1521, n1522, n1523, n1524, n1525, n1526, 
        n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1554, 
        n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, 
        n1596, n1597, n1598, n1599, n1600, n1601, n1620, n1621, 
        n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, 
        n1630, n1631, n1632, n1633, n19_adj_5843, n1653, n20_adj_5844, 
        n51847, n1688, n1689, n1690, n1691, n1692, n1693, n1694, 
        n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1719, 
        n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, 
        n1728, n1729, n1730, n1731, n1732, n1733, n1752, n51846, 
        n4_adj_5845, n1787, n1788_adj_5846, n1789, n1790_adj_5847, 
        n1791, n1792_adj_5848, n1793, n1794_adj_5849, n1795, n1796_adj_5850, 
        n1797, n1798, n1799, n1800, n1801, n1818, n1819, n1820, 
        n1821, n1822_adj_5851, n1823, n1824_adj_5852, n1825, n1826, 
        n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1851, 
        n51845, n1885, n1886, n1887, n1888, n1889, n1890, n1891, 
        n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, 
        n1900, n1901, n51571, n71225, n1917, n1918, n1919, n1920, 
        n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, 
        n1929, n1930, n1931, n1932, n1933, n51570, n1950, n1985, 
        n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, 
        n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, 
        n51844, n2016, n2017, n2018, n2019, n2020, n2021, n2022, 
        n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, 
        n2031, n2032, n2033, n51843, n2049, n51569, n51842, n51568, 
        n51567, n67721, n2084, n2085, n2086, n2087, n2088, n2089, 
        n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, 
        n2098, n2099, n2100, n2101, n2115, n2116, n2117, n2118, 
        n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, 
        n2127, n2128, n2129, n2130, n2131, n2132, n2133, n63053, 
        n59516, n2148, n490, n59514, n2182, n2183, n2184, n2185, 
        n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, 
        n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, 
        n36, n2214, n2215, n2216, n2217_adj_5853, n2218, n2219, 
        n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, 
        n2228, n2229, n2230, n2231, n2232, n2233, n2247, n2282, 
        n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, 
        n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, 
        n2299, n2300, n2301, n33, n59512, n2313, n2314, n2315, 
        n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, 
        n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, 
        n2332, n2333, n40820, n40838, n2346, n40853, n87, n63047, 
        n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, 
        n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, 
        n2397, n2398, n2399, n2400, n2401, n2412, n2413, n2414, 
        n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, 
        n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, 
        n2431, n2432, n2433, n2445, n37330, n161, n2480, n2481, 
        n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, 
        n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497, 
        n2498, n2499, n2500, n2501, n2511, n2512, n2513, n2514, 
        n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, 
        n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, 
        n2531, n2532, n2533, n43503, n2544, n164, n63045, n98, 
        n160, n163, n2579, n2580, n2581, n2582, n2583, n2584, 
        n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, 
        n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, 
        n2601, n159, n2610, n2611, n2612, n2613, n2614, n2615, 
        n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, 
        n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, 
        n2632, n2633, n2643, n59510, n2678, n2679, n2680, n2681, 
        n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689, 
        n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, 
        n2698, n2699, n2700, n2701, n2709, n2710, n2711, n2712, 
        n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, 
        n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, 
        n2729, n2730, n2731, n2732, n2733, n4_adj_5854, n70371, 
        n2742, n59507, n28_adj_5855, n63043, n59505, n2777, n2778, 
        n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786, 
        n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, 
        n2795, n2796, n2797, n2798, n2799, n2800, n2801, n51566, 
        n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815, 
        n2816, n2817, n2818, n2819, n2820_adj_5856, n2821, n2822, 
        n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, 
        n2831, n2832, n2833, n2841, n20182, n2876, n2877, n2878, 
        n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886, 
        n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894, 
        n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2907, 
        n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915, 
        n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, 
        n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, 
        n2932, n2933, n75, n2940, n2975, n2976, n2977, n2978, 
        n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, 
        n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994, 
        n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3006, 
        n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014, 
        n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, 
        n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, 
        n3031, n3032, n3033, n3039, n63039, n71222, n3074, n3075, 
        n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, 
        n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, 
        n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099, 
        n3100, n3101, n3105, n3106, n3107, n3108, n3109, n3110, 
        n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, 
        n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, 
        n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3138, 
        n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, 
        n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, 
        n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, 
        n3197, n3198, n3199, n3200, n3201, n3204, n3205, n3206, 
        n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, 
        n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, 
        n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, 
        n3231, n3232, n3233, n70164, n3237, n51841, n51300, n417, 
        n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, 
        n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, 
        n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295, 
        n3296, n71003, n3298, n3301, n51840, n29_adj_5857, n27_adj_5858, 
        n70919, n51565, n51299, n51564, n42812, n61, n24_adj_5859, 
        n23_adj_5860, n60274, n62, n67691, n51563, n22_adj_5861, 
        n51298, n25414, n28_adj_5862, n40, n51297, n51839, n63021, 
        n68200, n69307, n68198, n63553, n68194, n51838, n51837, 
        n4_adj_5863, n51836, n27901, n51562, n51561, n25_adj_5864, 
        n70454, n43, n45, n51560, n51559, n50994, n30110, n51835, 
        n51834, n51558, n43727, n27855, n51557, n51556, n51555, 
        n51554, n51833, n50981, n63013, n51296, n51832, n51295, 
        n25391, n30079, n6_adj_5865, n51294, n30075, n63011, n60438, 
        n27715, n30072, n51293, n51831, n51830, n71192, n63009, 
        n58928, n51829, n51828, n51827, n51826, n63007, n25508, 
        n27661, n63001, n30062, n58190, n27643, n25515, n19_adj_5866, 
        n71180, n4_adj_5867, n70427, n71174, n4_adj_5868, n18_adj_5869, 
        n20_adj_5870, n31_adj_5871, n71168, n71165, n27635, n62999, 
        n27629, n62997, n30059, n30056, n61707, n62991, n51292, 
        n51825, n20183, n61826, n62985, n344, n71162, n69454, 
        n30053, n51824, n51823, n51291, n62983, n58002, n27585, 
        n271, n51290, n62979, n25522, n60489, n30049, n70773, 
        n51822, n50993, n51289, n71156, n30046, n27561, n62973, 
        n51821, n51820, n51819, n198, n204, n51818, n51817, n51816, 
        n51527, n51526, n15_adj_5872, n71000, n131, n51525, n62963, 
        n51288, n51287, n51524, n51286, n125, n70997, n51815, 
        n51523, n51285, n51522, n51521, n110, n62953, n62951, 
        n51814, n62949, n53, n56, n51813, n51520, n51519, n51518, 
        n62947, n51517, n62945, n38, n62943, n51812, n51811, n51810, 
        n62941, n62939, n51516, n51809, n51515, n62937, n62935, 
        n16_adj_5873, n62929, n62923, n51284, n51514, n51283, n51513, 
        n62917, n70994, n51808, n62911, n70991, n51512, n51282, 
        n62905, n61386, n62899, n51281, n51807, n62893, n62891, 
        n70988, n36881, n3_adj_5874, n70202, n62885, n51511, n62883, 
        n26376, n26372, n69097, n26282, n26210, n62873, n67899, 
        n26143, n59055, n62867, n51806, n52457, n36845, n51805, 
        n67879, n62857, n4_adj_5875, n6_adj_5876, n8_adj_5877, n9_adj_5878, 
        n4_adj_5879, n6_adj_5880, n8_adj_5881, n9_adj_5882, n11_adj_5883, 
        n13_adj_5884, n15_adj_5885, n52456, n51804, n51803, n51802, 
        n51801, n62847, n52455, n51800, n51799, n51798, n69435, 
        n51797, n51280, n51796, n52454, n51795, n51794, n52453, 
        n70760, n51793, n38_adj_5886, n39, n40_adj_5887, n41, n42, 
        n43_adj_5888, n44, n45_adj_5889, n29405, n29403, n55, n11597, 
        n25700, n51792, n69434, n62841, n11566, n11564, n51791, 
        n67852, n51493, n51492, n51491, n51790, n51490, n51789, 
        n58751, n62835, n62831, n62823, n59153, n43547, n62817, 
        n62811, n59359, n51489, n51788, n51488, n29091, n58671, 
        n58670, n58669, n58668, n58667, n58666, n58665, n58664, 
        n58663, n58662, n58661, n58660, n58659, n58507, n58658, 
        n58657, n58656, n58655, n58654, n58653, n58652, n58651, 
        n58650, n58649, n58648, n58647, n58646, n58645, n58644, 
        n62801, n58643, n58642, n58641, n58640, n58639, n58638, 
        n67177, n28385, n28370, n28368, n28366, n61551, n28356, 
        n28814, n60449, n28807, n28313, n28311, n28309, n28307, 
        n52452, n54640, n51787, n51487, n51786, n51486, n51485, 
        n51484, n69291, n51785, n52451, n51784, n51783, n51483, 
        n52450, n51482, n51481, n51480, n67171, n52449, n62795, 
        n52448, n52447, n50992, n51479, n6_adj_5890, n51782, n52446, 
        n51478, n4_adj_5891, n52445, n51781, n51780, n58637, n52444, 
        n51779, n51778, n51777, n51776, n51775, n57800, n51774, 
        n51773, n62787, n29402, n62785, n30043, n52443, n25512, 
        n51772, n51771, n25517, n51770, n51769, n71144, n62779, 
        n61367, n51454, n52442, n20136, n51768, n51453, n52441, 
        n51767, n51452, n51451, n30030, n62773, n60367, n51766, 
        n58636, n51450, n52440, n51449, n51448, n51447, n62767, 
        n60372, n43791, n29976, n29973, n29970, n50991, n52439, 
        n52438, n43779, n29964, n29961, n43775, n29958, n51765, 
        n51764, n52437, n43773, n29955, n51763, n51446, n52436, 
        n43771, n62761, n51762, n52435, n29946, n29943, n29940, 
        n43765, n52434, n51761, n29937, n29934, n51445, n51760, 
        n51759, n52433, n52432, n51444, n29930, n43759, n43737, 
        n29901, n58635, n52431, n52430, n51443, n51758, n51442, 
        n51441, n62755, n52429, n51757, n51756, n51440, n51755, 
        n51754, n62751, n51753, n51752, n51751, n52428, n52427, 
        n69091, n51750, n51749, n62749, n51748, n50990, n51747, 
        n51117, n50980, n51746, n51745, n51744, n51743, n51116, 
        n51742, n51741, n51115, n51740, n51424, n51739, n51114, 
        n51423, n51113, n51738, n51422, n2_adj_5892, n3_adj_5893, 
        n4_adj_5894, n5_adj_5895, n6_adj_5896, n7_adj_5897, n8_adj_5898, 
        n9_adj_5899, n10_adj_5900, n11_adj_5901, n12_adj_5902, n13_adj_5903, 
        n14_adj_5904, n15_adj_5905, n16_adj_5906, n17_adj_5907, n18_adj_5908, 
        n19_adj_5909, n20_adj_5910, n21_adj_5911, n22_adj_5912, n23_adj_5913, 
        n24_adj_5914, n25_adj_5915, n26_adj_5916, n27_adj_5917, n28_adj_5918, 
        n29_adj_5919, n30_adj_5920, n31_adj_5921, n32_adj_5922, n51421, 
        n51737, n51420, n51419, n51736, n51735, n51734, n51418, 
        n51417, n51416, n51415, n51112, n51111, n51414, n51110, 
        n51733, n51413, n51109, n51732, n51412, n51731, n51730, 
        n51729, n51411, n51728, n51727, n52229, n51246, n51726, 
        n51245, n52228, n51725, n51108, n51107, n51244, n51106, 
        n51724, n52227, n51243, n51105, n52226, n51723, n51104, 
        n51722, n51103, n51242, n52225, n52224, n51102, n51980, 
        n51721, n51720, n51719, n51718, n51101, n51717, n51241, 
        n51716, n67140, n51240, n51100, n52223, n51979, n51239, 
        n51099, n51098, n51715, n51978, n50989, n51238, n51714, 
        n51977, n51713, n51237, n51097, n51236, n51976, n51712, 
        n51711, n51975, n51710, n51235, n51709, n62735, n51096, 
        n51234, n51974, n51973, n51095, n51708, n51972, n51707, 
        n51706, n50979, n51971, n51705, n51704, n51970, n51703, 
        n51390, n51233, n51969, n51232, n51702, n51231, n51230, 
        n51008, n51389, n70743, n51968, n51967, n51388, n51387, 
        n51229, n51228, n51966, n51965, n51964, n62725, n51963, 
        n51386, n51385, n51007, n51006, n50978, n51384, n51383, 
        n51227, n51962, n51226, n51961, n51382, n51005, n51225, 
        n51224, n51381, n51960, n51004, n51959, n51958, n67130, 
        n51380, n51379, n51957, n51956, n51955, n64026, n51954, 
        n51378, n51953, n51223, n51222, n51952, n67128, n6_adj_5923, 
        n67125, n51951, n51221, n6_adj_5924, n51950, n51220, n12_adj_5925, 
        n51949, n51219, n51218, n51948, n13_adj_5926, n15_adj_5927, 
        n17_adj_5928, n19_adj_5929, n23_adj_5930, n31_adj_5931, n33_adj_5932, 
        n61_adj_5933, n69105, n51947, n51946, n51945, n51944, n22734, 
        n51943, n51942, n58418, n58634, n20209, n51941, n20877, 
        n20873, n58633, n63449, n70727, n4_adj_5934, n58632, n58631, 
        n33697, n58630, n58629, n51940, n51939, n51938, n51217, 
        n51216, n51937, n58628, n12169, n61345, n25385, n70712, 
        n63447, n53546, n25409, n25499, n20138, n20137, n70367, 
        n25490, n63441, n51215, n51214, n51936, n51213, n71132, 
        n25504, n51935, n51934, n53519, n53515, n22979, n50988, 
        n51933, n51932, n51003, n51931, n51930, n63429, n50987, 
        n50986, n63425, n63423, n51929, n53457, n51928, n54113, 
        n51927, n71126, n63417, n63415, n70337, n71120, n70635, 
        n6_adj_5935, n67092, n67087, n67086, n62525, n69998, n62519, 
        n59508, n62513, n57114, n5_adj_5936, n24_adj_5937, n62509, 
        n17_adj_5938, n25_adj_5939, n62503, n62497, n62493, n62487, 
        n57200, n62481, n62477, n62471, n62465, n62461, n62455, 
        n62449, n62445, n62439, n62433, n62429, n58845, n59274, 
        n58684, n58938, n62423, n59027, n62417, n61638, n59007, 
        n59223, n62413, n62407, n71412, n59452, n59124, n62401, 
        n71114, n57450, n30_adj_5940, n28_adj_5941, n26_adj_5942, 
        n25_adj_5943, n22_adj_5944, n61449, n59299, n70615, n4_adj_5945, 
        n61067, n61064, n59430, n59455, n59406, n8_adj_5946, n6_adj_5947, 
        n15_adj_5948, n14_adj_5949, n14_adj_5950, n13_adj_5951, n70158, 
        n69948, n69942, n71084, n69941, n69937, n59477, n60513, 
        n66991, n58887, n60429, n69936, n60364, n63357, n69772, 
        n70596, n71108, n69991, n69741, n59241, n70304, n61932, 
        n69848, n71102, n60442, n69690, n62163, n60464, n62157, 
        n69740, n60479, n69618, n57834, n57838, n57842, n57846, 
        n57850, n57856, n57860, n57864, n57868, n57872, n57882, 
        n60375, n57886, n57890, n4_adj_5952, n57914, n9_adj_5953, 
        n70578, n57932, n57936, n69760, n57968, n57974, n57980, 
        n57986, n61888, n60467, n8_adj_5954, n12_adj_5955, n69762, 
        n69443, n69442, n58060, n62099, n60380, n62091, n62089, 
        n58106, n7_adj_5956, n62071, n70020, n7_adj_5957, n63793, 
        n64304, n63789, n63783, n71096, n63779, n63773, n70554, 
        n66963, n70273, n62029, n64302, n64301, n64298, n58805, 
        n64180, n59215, n60405, n68630, n4_adj_5958, n70528, n68690, 
        n68664, n7_adj_5959;
    
    VCC i2 (.Y(VCC_net));
    SB_LUT4 i1_4_lut (.I0(n19_adj_5929), .I1(n33_adj_5932), .I2(n62929), 
            .I3(n15_adj_5927), .O(n62935));
    defparam i1_4_lut.LUT_INIT = 16'hfffe;
    SB_IO hall2_input (.PACKAGE_PIN(HALL2), .LATCH_INPUT_VALUE(GND_net), 
          .INPUT_CLK(GND_net), .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_1(GND_net), .D_OUT_0(GND_net), .D_IN_0(hall2)) /* synthesis syn_instantiated=1 */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam hall2_input.PIN_TYPE = 6'b000001;
    defparam hall2_input.PULLUP = 1'b1;
    defparam hall2_input.NEG_TRIGGER = 1'b0;
    defparam hall2_input.IO_STANDARD = "SB_LVCMOS";
    SB_IO hall3_input (.PACKAGE_PIN(HALL3), .LATCH_INPUT_VALUE(GND_net), 
          .INPUT_CLK(GND_net), .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_1(GND_net), .D_OUT_0(GND_net), .D_IN_0(hall3)) /* synthesis syn_instantiated=1 */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam hall3_input.PIN_TYPE = 6'b000001;
    defparam hall3_input.PULLUP = 1'b1;
    defparam hall3_input.NEG_TRIGGER = 1'b0;
    defparam hall3_input.IO_STANDARD = "SB_LVCMOS";
    SB_IO tx_output (.PACKAGE_PIN(TX), .LATCH_INPUT_VALUE(GND_net), .INPUT_CLK(GND_net), 
          .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(tx_enable), .D_OUT_1(GND_net), 
          .D_OUT_0(tx_o)) /* synthesis syn_instantiated=1 */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam tx_output.PIN_TYPE = 6'b101001;
    defparam tx_output.PULLUP = 1'b1;
    defparam tx_output.NEG_TRIGGER = 1'b0;
    defparam tx_output.IO_STANDARD = "SB_LVCMOS";
    SB_CARRY encoder0_position_30__I_0_add_1570_19 (.CI(n51718), .I0(n2317), 
            .I1(VCC_net), .CO(n51719));
    SB_LUT4 encoder0_position_30__I_0_i1582_3_lut (.I0(n2323), .I1(n2390), 
            .I2(n2346), .I3(GND_net), .O(n2422));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1582_3_lut.LUT_INIT = 16'hacac;
    SB_DFF dir_183 (.Q(dir), .C(clk16MHz), .D(pwm_setpoint_23__N_207));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_LUT4 i1_4_lut_adj_1742 (.I0(n3217), .I1(n62935), .I2(n3284), .I3(n3237), 
            .O(n62937));
    defparam i1_4_lut_adj_1742.LUT_INIT = 16'heefc;
    SB_LUT4 encoder0_position_30__I_0_add_2039_24_lut (.I0(GND_net), .I1(n3012), 
            .I2(VCC_net), .I3(n51891), .O(n3079)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2039_24_lut.LUT_INIT = 16'hC33C;
    SB_DFFE dti_185 (.Q(dti), .C(clk16MHz), .E(n27561), .D(dti_N_404));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    SB_LUT4 encoder0_position_30__I_0_i1649_3_lut (.I0(n2422), .I1(n2489), 
            .I2(n2445), .I3(GND_net), .O(n2521));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1649_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1743 (.I0(n3216), .I1(n62937), .I2(n3283), .I3(n3237), 
            .O(n62939));
    defparam i1_4_lut_adj_1743.LUT_INIT = 16'heefc;
    SB_LUT4 i1_4_lut_adj_1744 (.I0(n3215), .I1(n62939), .I2(n3282), .I3(n3237), 
            .O(n62941));
    defparam i1_4_lut_adj_1744.LUT_INIT = 16'heefc;
    SB_DFF encoder0_position_scaled_i0 (.Q(encoder0_position_scaled[0]), .C(clk16MHz), 
           .D(encoder0_position_scaled_23__N_43[0]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_CARRY encoder0_position_30__I_0_add_1838_9 (.CI(n51798), .I0(n2727), 
            .I1(VCC_net), .CO(n51799));
    SB_CARRY encoder0_position_30__I_0_add_2039_24 (.CI(n51891), .I0(n3012), 
            .I1(VCC_net), .CO(n51892));
    SB_LUT4 i1_4_lut_adj_1745 (.I0(n3213), .I1(n62941), .I2(n3280), .I3(n3237), 
            .O(n62943));
    defparam i1_4_lut_adj_1745.LUT_INIT = 16'heefc;
    SB_LUT4 i1_4_lut_adj_1746 (.I0(n3212), .I1(n62943), .I2(n3279), .I3(n3237), 
            .O(n62945));
    defparam i1_4_lut_adj_1746.LUT_INIT = 16'heefc;
    SB_LUT4 i1_4_lut_adj_1747 (.I0(n3211), .I1(n62945), .I2(n3278), .I3(n3237), 
            .O(n62947));
    defparam i1_4_lut_adj_1747.LUT_INIT = 16'heefc;
    SB_CARRY encoder0_position_30__I_0_unary_minus_2_add_3_15 (.CI(n52439), 
            .I0(GND_net), .I1(n20_adj_5910), .CO(n52440));
    SB_DFF pwm_setpoint_i0 (.Q(pwm_setpoint[0]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[0]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_LUT4 encoder0_position_30__I_0_i1716_3_lut (.I0(n2521), .I1(n2588), 
            .I2(n2544), .I3(GND_net), .O(n2620));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1716_3_lut.LUT_INIT = 16'hacac;
    SB_DFF encoder1_position_scaled_i0 (.Q(encoder1_position_scaled[0]), .C(clk16MHz), 
           .D(encoder1_position[2]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_LUT4 i16488_2_lut_2_lut_4_lut (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[13] [0]), 
            .O(n30494));   // verilog/coms.v(130[12] 305[6])
    defparam i16488_2_lut_2_lut_4_lut.LUT_INIT = 16'h5555;
    SB_DFF displacement_i0 (.Q(displacement[0]), .C(clk16MHz), .D(displacement_23__N_67[0]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_IO sda_output (.PACKAGE_PIN(SDA), .LATCH_INPUT_VALUE(GND_net), .INPUT_CLK(GND_net), 
          .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(sda_enable), .D_OUT_1(GND_net), 
          .D_OUT_0(sda_out), .D_IN_0(state_7__N_4126[3])) /* synthesis syn_instantiated=1 */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam sda_output.PIN_TYPE = 6'b101001;
    defparam sda_output.PULLUP = 1'b1;
    defparam sda_output.NEG_TRIGGER = 1'b0;
    defparam sda_output.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 i1_4_lut_adj_1748 (.I0(n3210), .I1(n62947), .I2(n3277), .I3(n3237), 
            .O(n62949));
    defparam i1_4_lut_adj_1748.LUT_INIT = 16'heefc;
    SB_IO INHC_pad (.PACKAGE_PIN(INHC), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INHC_c_0));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INHC_pad.PIN_TYPE = 6'b011001;
    defparam INHC_pad.PULLUP = 1'b0;
    defparam INHC_pad.NEG_TRIGGER = 1'b0;
    defparam INHC_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 i1_4_lut_adj_1749 (.I0(n3209), .I1(n62949), .I2(n3276), .I3(n3237), 
            .O(n62951));
    defparam i1_4_lut_adj_1749.LUT_INIT = 16'heefc;
    SB_IO scl_output (.PACKAGE_PIN(SCL), .LATCH_INPUT_VALUE(GND_net), .INPUT_CLK(GND_net), 
          .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(scl_enable), .D_OUT_1(GND_net), 
          .D_OUT_0(scl)) /* synthesis syn_instantiated=1 */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam scl_output.PIN_TYPE = 6'b101001;
    defparam scl_output.PULLUP = 1'b1;
    defparam scl_output.NEG_TRIGGER = 1'b0;
    defparam scl_output.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 encoder0_position_30__I_0_i2198_3_lut (.I0(n3227), .I1(n3294), 
            .I2(n3237), .I3(GND_net), .O(n17_adj_5928));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2198_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16_4_lut (.I0(n3231), .I1(n67092), .I2(n3237), .I3(n3230), 
            .O(n5_adj_5720));
    defparam i16_4_lut.LUT_INIT = 16'hac0c;
    SB_LUT4 encoder0_position_30__I_0_add_1838_8_lut (.I0(GND_net), .I1(n2728), 
            .I2(VCC_net), .I3(n51797), .O(n2795)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1838_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i51709_3_lut (.I0(n957), .I1(n3232), .I2(n3233), .I3(GND_net), 
            .O(n67086));
    defparam i51709_3_lut.LUT_INIT = 16'hecec;
    SB_CARRY encoder0_position_30__I_0_add_766_2 (.CI(VCC_net), .I0(n522), 
            .I1(GND_net), .CO(n51306));
    SB_IO hall1_input (.PACKAGE_PIN(HALL1), .LATCH_INPUT_VALUE(GND_net), 
          .INPUT_CLK(GND_net), .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_1(GND_net), .D_OUT_0(GND_net), .D_IN_0(hall1)) /* synthesis syn_instantiated=1 */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam hall1_input.PIN_TYPE = 6'b000001;
    defparam hall1_input.PULLUP = 1'b1;
    defparam hall1_input.NEG_TRIGGER = 1'b0;
    defparam hall1_input.IO_STANDARD = "SB_LVCMOS";
    \neopixel(CLOCK_SPEED_HZ=16000000)  nx (.VCC_net(VCC_net), .timer({timer}), 
            .clk16MHz(clk16MHz), .GND_net(GND_net), .state({state}), .\neo_pixel_transmitter.t0 ({\neo_pixel_transmitter.t0 }), 
            .n22979(n22979), .neopxl_color({neopxl_color}), .bit_ctr({Open_0, 
            Open_1, Open_2, Open_3, bit_ctr[0]}), .n29595(n29595), 
            .n27855(n27855), .\bit_ctr[3] (bit_ctr[3]), .\bit_ctr[4] (bit_ctr[4]), 
            .\bit_ctr[1] (bit_ctr[1]), .n43547(n43547), .n30238(n30238), 
            .n30237(n30237), .n30236(n30236), .n30235(n30235), .n30234(n30234), 
            .n30233(n30233), .n30232(n30232), .n30231(n30231), .n30230(n30230), 
            .n30224(n30224), .n30139(n30139), .n57450(n57450), .NEOPXL_c(NEOPXL_c), 
            .n66810(n66810), .LED_c(LED_c), .\color_bit_N_502[1] (color_bit_N_502[1]), 
            .n53519(n53519), .n3157(n3157)) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(51[24] 57[2])
    SB_LUT4 encoder0_position_30__I_0_add_699_10_lut (.I0(GND_net), .I1(n1026), 
            .I2(VCC_net), .I3(n51305), .O(n1093)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_699_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1570_18_lut (.I0(GND_net), .I1(n2318), 
            .I2(VCC_net), .I3(n51717), .O(n2385)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1570_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_i1783_3_lut (.I0(n2620), .I1(n2687), 
            .I2(n2643), .I3(GND_net), .O(n2719));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1783_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_add_3_14_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n21_adj_5911), .I3(n52438), .O(n21_adj_5727)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_unary_minus_2_add_3_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1750 (.I0(n3222), .I1(n23_adj_5930), .I2(n3289), 
            .I3(n3237), .O(n62999));
    defparam i1_4_lut_adj_1750.LUT_INIT = 16'heefc;
    SB_LUT4 i1_4_lut_adj_1751 (.I0(n3223), .I1(n31_adj_5931), .I2(n3290), 
            .I3(n3237), .O(n62997));
    defparam i1_4_lut_adj_1751.LUT_INIT = 16'heefc;
    SB_LUT4 i1_4_lut_adj_1752 (.I0(n67086), .I1(n5_adj_5720), .I2(n67087), 
            .I3(n3237), .O(n55096));
    defparam i1_4_lut_adj_1752.LUT_INIT = 16'h88c0;
    SB_LUT4 i1_4_lut_adj_1753 (.I0(n3225), .I1(n17_adj_5928), .I2(n3292), 
            .I3(n3237), .O(n63001));
    defparam i1_4_lut_adj_1753.LUT_INIT = 16'heefc;
    SB_LUT4 encoder0_position_30__I_0_i1850_3_lut (.I0(n2719), .I1(n2786), 
            .I2(n2742), .I3(GND_net), .O(n2818));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1850_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1754 (.I0(n63001), .I1(n55096), .I2(n62997), 
            .I3(n62999), .O(n63007));
    defparam i1_4_lut_adj_1754.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1755 (.I0(n3218), .I1(n63007), .I2(n3285), .I3(n3237), 
            .O(n63009));
    defparam i1_4_lut_adj_1755.LUT_INIT = 16'heefc;
    SB_LUT4 encoder0_position_30__I_0_i1917_3_lut (.I0(n2818), .I1(n2885), 
            .I2(n2841), .I3(GND_net), .O(n2917));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1917_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1756 (.I0(n3214), .I1(n63009), .I2(n3281), .I3(n3237), 
            .O(n63011));
    defparam i1_4_lut_adj_1756.LUT_INIT = 16'heefc;
    SB_LUT4 encoder0_position_30__I_0_add_2039_23_lut (.I0(GND_net), .I1(n3013), 
            .I2(VCC_net), .I3(n51890), .O(n3080)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2039_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_unary_minus_2_add_3_14 (.CI(n52438), 
            .I0(GND_net), .I1(n21_adj_5911), .CO(n52439));
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_add_3_13_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n22_adj_5912), .I3(n52437), .O(n22_adj_5726)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_unary_minus_2_add_3_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1757 (.I0(n3207), .I1(n63011), .I2(n3274), .I3(n3237), 
            .O(n63013));
    defparam i1_4_lut_adj_1757.LUT_INIT = 16'heefc;
    SB_CARRY encoder0_position_30__I_0_unary_minus_2_add_3_13 (.CI(n52437), 
            .I0(GND_net), .I1(n22_adj_5912), .CO(n52438));
    SB_LUT4 i1_4_lut_adj_1758 (.I0(n3208), .I1(n62951), .I2(n3275), .I3(n3237), 
            .O(n62953));
    defparam i1_4_lut_adj_1758.LUT_INIT = 16'heefc;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_add_3_12_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n23_adj_5913), .I3(n52436), .O(n23_adj_5725)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_unary_minus_2_add_3_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1759 (.I0(n63013), .I1(n3206), .I2(n3273), .I3(n3237), 
            .O(n61638));
    defparam i1_4_lut_adj_1759.LUT_INIT = 16'heefa;
    SB_LUT4 encoder0_position_30__I_0_i2176_3_lut (.I0(n3205), .I1(n3272), 
            .I2(n3237), .I3(GND_net), .O(n61_adj_5933));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2176_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i54473_4_lut (.I0(n61_adj_5933), .I1(n64026), .I2(n61638), 
            .I3(n62953), .O(n43737));
    defparam i54473_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i19_1_lut (.I0(encoder1_position_scaled[18]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n7_adj_5821));   // verilog/TinyFPGA_B.v(323[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_i1984_3_lut (.I0(n2917), .I1(n2984), 
            .I2(n2940), .I3(GND_net), .O(n3016));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1984_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_1582_i21_3_lut (.I0(duty[23]), .I1(duty[20]), .I2(n260), 
            .I3(GND_net), .O(n12173));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1582_i21_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i20_1_lut (.I0(encoder1_position_scaled[19]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n6_adj_5822));   // verilog/TinyFPGA_B.v(323[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_245_i20_4_lut (.I0(encoder1_position_scaled[19]), .I1(displacement[19]), 
            .I2(n15_adj_5722), .I3(n15), .O(motor_state_23__N_91[19]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i20_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 encoder0_position_30__I_0_i2110_3_lut (.I0(n3107), .I1(n3174), 
            .I2(n3138), .I3(GND_net), .O(n3206));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2110_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 RX_I_0_1_lut (.I0(RX_c), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(RX_N_2));   // verilog/TinyFPGA_B.v(262[11:14])
    defparam RX_I_0_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_i2109_3_lut (.I0(n3106), .I1(n3173), 
            .I2(n3138), .I3(GND_net), .O(n3205));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2109_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2112_3_lut (.I0(n3109), .I1(n3176), 
            .I2(n3138), .I3(GND_net), .O(n3208));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2112_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2111_3_lut (.I0(n3108), .I1(n3175), 
            .I2(n3138), .I3(GND_net), .O(n3207));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2111_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1983_3_lut (.I0(n2916), .I1(n2983), 
            .I2(n2940), .I3(GND_net), .O(n3015));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1983_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2132_3_lut (.I0(n3129), .I1(n3196), 
            .I2(n3138), .I3(GND_net), .O(n3228));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2132_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2121_3_lut (.I0(n3118), .I1(n3185), 
            .I2(n3138), .I3(GND_net), .O(n3217));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2121_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2128_3_lut (.I0(n3125), .I1(n3192), 
            .I2(n3138), .I3(GND_net), .O(n3224));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2128_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2119_3_lut (.I0(n3116), .I1(n3183), 
            .I2(n3138), .I3(GND_net), .O(n3215));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2119_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2118_3_lut (.I0(n3115), .I1(n3182), 
            .I2(n3138), .I3(GND_net), .O(n3214));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2118_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2115_3_lut (.I0(n3112), .I1(n3179), 
            .I2(n3138), .I3(GND_net), .O(n3211));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2115_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2114_3_lut (.I0(n3111), .I1(n3178), 
            .I2(n3138), .I3(GND_net), .O(n3210));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2114_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2113_3_lut (.I0(n3110), .I1(n3177), 
            .I2(n3138), .I3(GND_net), .O(n3209));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2113_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2117_3_lut (.I0(n3114), .I1(n3181), 
            .I2(n3138), .I3(GND_net), .O(n3213));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2117_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2120_3_lut (.I0(n3117), .I1(n3184), 
            .I2(n3138), .I3(GND_net), .O(n3216));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2120_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2116_3_lut (.I0(n3113), .I1(n3180), 
            .I2(n3138), .I3(GND_net), .O(n3212));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2116_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2126_3_lut (.I0(n3123), .I1(n3190), 
            .I2(n3138), .I3(GND_net), .O(n3222));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2126_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2127_3_lut (.I0(n3124), .I1(n3191), 
            .I2(n3138), .I3(GND_net), .O(n3223));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2127_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2137_3_lut (.I0(n956), .I1(n3201), 
            .I2(n3138), .I3(GND_net), .O(n3233));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2137_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2136_3_lut (.I0(n3133), .I1(n3200), 
            .I2(n3138), .I3(GND_net), .O(n3232));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2136_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_4297_i1_3_lut (.I0(encoder0_position[0]), .I1(n32), .I2(encoder0_position[30]), 
            .I3(GND_net), .O(n957));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam mux_4297_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_i2135_3_lut (.I0(n3132), .I1(n3199), 
            .I2(n3138), .I3(GND_net), .O(n3231));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2135_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2134_3_lut (.I0(n3131), .I1(n3198), 
            .I2(n3138), .I3(GND_net), .O(n3230));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2134_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2133_3_lut (.I0(n3130), .I1(n3197), 
            .I2(n3138), .I3(GND_net), .O(n3229));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2133_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2122_3_lut (.I0(n3119), .I1(n3186), 
            .I2(n3138), .I3(GND_net), .O(n3218));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2122_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2129_3_lut (.I0(n3126), .I1(n3193), 
            .I2(n3138), .I3(GND_net), .O(n3225));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2129_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2130_3_lut (.I0(n3127), .I1(n3194), 
            .I2(n3138), .I3(GND_net), .O(n3226));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2130_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2123_3_lut (.I0(n3120), .I1(n3187), 
            .I2(n3138), .I3(GND_net), .O(n3219));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2123_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2124_3_lut (.I0(n3121), .I1(n3188), 
            .I2(n3138), .I3(GND_net), .O(n3220));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2124_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2131_3_lut (.I0(n3128), .I1(n3195), 
            .I2(n3138), .I3(GND_net), .O(n3227));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2131_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2125_3_lut (.I0(n3122), .I1(n3189), 
            .I2(n3138), .I3(GND_net), .O(n3221));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2125_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i54464_1_lut (.I0(n3237), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n70158));
    defparam i54464_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_4_lut_adj_1760 (.I0(n3219), .I1(n3226), .I2(n3225), .I3(n3218), 
            .O(n63415));
    defparam i1_4_lut_adj_1760.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_30__I_0_add_699_9_lut (.I0(GND_net), .I1(n1027), 
            .I2(VCC_net), .I3(n51304), .O(n1094)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_699_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i29826_3_lut (.I0(n957), .I1(n3232), .I2(n3233), .I3(GND_net), 
            .O(n43727));
    defparam i29826_3_lut.LUT_INIT = 16'hc8c8;
    SB_CARRY encoder0_position_30__I_0_unary_minus_2_add_3_12 (.CI(n52436), 
            .I0(GND_net), .I1(n23_adj_5913), .CO(n52437));
    SB_LUT4 i1_4_lut_adj_1761 (.I0(n3221), .I1(n63415), .I2(n3227), .I3(n3220), 
            .O(n63417));
    defparam i1_4_lut_adj_1761.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1762 (.I0(n3229), .I1(n43727), .I2(n3230), .I3(n3231), 
            .O(n60513));
    defparam i1_4_lut_adj_1762.LUT_INIT = 16'ha080;
    SB_LUT4 i1_2_lut (.I0(n3223), .I1(n3222), .I2(GND_net), .I3(GND_net), 
            .O(n63449));
    defparam i1_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_1763 (.I0(n3212), .I1(n60513), .I2(n3216), .I3(n63417), 
            .O(n63423));
    defparam i1_4_lut_adj_1763.LUT_INIT = 16'hfffe;
    SB_LUT4 i12_4_lut (.I0(\data_out_frame[21] [1]), .I1(n25764), .I2(\data_out_frame[23] [2]), 
            .I3(n54490), .O(n28_adj_5941));
    defparam i12_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i10_4_lut (.I0(n59455), .I1(\data_out_frame[16] [2]), .I2(\data_out_frame[20] [4]), 
            .I3(\data_out_frame[14] [4]), .O(n26_adj_5942));
    defparam i10_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i14_4_lut (.I0(n59477), .I1(n28_adj_5941), .I2(n22_adj_5944), 
            .I3(n59359), .O(n30_adj_5940));
    defparam i14_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 encoder0_position_30__I_0_i1043_3_lut (.I0(n1528), .I1(n1595), 
            .I2(n1554), .I3(GND_net), .O(n1627));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1043_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1764 (.I0(n3215), .I1(n3224), .I2(n3217), .I3(n3228), 
            .O(n63441));
    defparam i1_4_lut_adj_1764.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_30__I_0_i1110_3_lut (.I0(n1627), .I1(n1694), 
            .I2(n1653), .I3(GND_net), .O(n1726));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1110_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i9_4_lut (.I0(\data_out_frame[22] [7]), .I1(n59274), .I2(n54620), 
            .I3(\data_out_frame[23] [1]), .O(n25_adj_5943));
    defparam i9_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 encoder0_position_30__I_0_i1177_3_lut (.I0(n1726), .I1(n1793), 
            .I2(n1752), .I3(GND_net), .O(n1825));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1177_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i44018_4_lut (.I0(reset), .I1(n161), .I2(n43501), .I3(\FRAME_MATCHER.i [0]), 
            .O(n59656));
    defparam i44018_4_lut.LUT_INIT = 16'hefff;
    SB_LUT4 encoder0_position_30__I_0_i1244_3_lut (.I0(n1825), .I1(n1892), 
            .I2(n1851), .I3(GND_net), .O(n1924));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1244_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15889_3_lut (.I0(\data_in_frame[5] [5]), .I1(rx_data[5]), .I2(n59656), 
            .I3(GND_net), .O(n29895));   // verilog/coms.v(130[12] 305[6])
    defparam i15889_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1311_3_lut (.I0(n1924), .I1(n1991), 
            .I2(n1950), .I3(GND_net), .O(n2023));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1311_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1765 (.I0(n3213), .I1(n63423), .I2(n3209), .I3(n63449), 
            .O(n63425));
    defparam i1_4_lut_adj_1765.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1766 (.I0(n3210), .I1(n3211), .I2(n3214), .I3(n63441), 
            .O(n63447));
    defparam i1_4_lut_adj_1766.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_30__I_0_i1378_3_lut (.I0(n2023), .I1(n2090), 
            .I2(n2049), .I3(GND_net), .O(n2122));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1378_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1767 (.I0(n3207), .I1(n63447), .I2(n63425), .I3(n3208), 
            .O(n63429));
    defparam i1_4_lut_adj_1767.LUT_INIT = 16'hfffe;
    SB_LUT4 i54469_4_lut (.I0(n3205), .I1(n3204), .I2(n3206), .I3(n63429), 
            .O(n3237));
    defparam i54469_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 mux_245_i21_4_lut (.I0(encoder1_position_scaled[20]), .I1(displacement[20]), 
            .I2(n15_adj_5722), .I3(n15), .O(motor_state_23__N_91[20]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i21_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i4_4_lut (.I0(\data_out_frame[21] [0]), .I1(\data_out_frame[18] [6]), 
            .I2(n59359), .I3(n6_adj_5924), .O(n53457));
    defparam i4_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut (.I0(\data_out_frame[22] [7]), .I1(\data_out_frame[20] [6]), 
            .I2(\data_out_frame[22] [6]), .I3(GND_net), .O(n59406));   // verilog/coms.v(100[12:26])
    defparam i2_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1768 (.I0(\data_out_frame[23] [2]), .I1(n53457), 
            .I2(GND_net), .I3(GND_net), .O(n59241));
    defparam i1_2_lut_adj_1768.LUT_INIT = 16'h6666;
    SB_LUT4 mux_1582_i22_3_lut (.I0(duty[23]), .I1(duty[21]), .I2(n260), 
            .I3(GND_net), .O(n12171));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1582_i22_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i21_1_lut (.I0(encoder1_position_scaled[20]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n5_adj_5825));   // verilog/TinyFPGA_B.v(323[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_4_lut_adj_1769 (.I0(n23_adj_5860), .I1(o_Rx_DV_N_3488[12]), 
            .I2(n4935), .I3(o_Rx_DV_N_3488[8]), .O(n62029));
    defparam i1_4_lut_adj_1769.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1770 (.I0(o_Rx_DV_N_3488[24]), .I1(n27_adj_5858), 
            .I2(n29_adj_5857), .I3(n62029), .O(r_SM_Main_2__N_3446[1]));
    defparam i1_4_lut_adj_1770.LUT_INIT = 16'hfffe;
    SB_CARRY encoder0_position_30__I_0_add_2039_23 (.CI(n51890), .I0(n3013), 
            .I1(VCC_net), .CO(n51891));
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_add_3_11_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n24_adj_5914), .I3(n52435), .O(n24_adj_5724)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_unary_minus_2_add_3_11_lut.LUT_INIT = 16'hC33C;
    SB_DFFESR delay_counter__i17 (.Q(delay_counter[17]), .C(clk16MHz), .E(n27635), 
            .D(n1222), .R(n28814));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    SB_DFFESR delay_counter__i18 (.Q(delay_counter[18]), .C(clk16MHz), .E(n27635), 
            .D(n1221), .R(n28814));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    SB_DFFESR delay_counter__i19 (.Q(delay_counter[19]), .C(clk16MHz), .E(n27635), 
            .D(n1220), .R(n28814));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    SB_DFFESR delay_counter__i20 (.Q(delay_counter[20]), .C(clk16MHz), .E(n27635), 
            .D(n1219), .R(n28814));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    SB_DFFESR delay_counter__i21 (.Q(delay_counter[21]), .C(clk16MHz), .E(n27635), 
            .D(n1218), .R(n28814));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    SB_DFFESR delay_counter__i22 (.Q(delay_counter[22]), .C(clk16MHz), .E(n27635), 
            .D(n1217), .R(n28814));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i22_1_lut (.I0(encoder1_position_scaled[21]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n4_adj_5795));   // verilog/TinyFPGA_B.v(323[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_DFFESR delay_counter__i23 (.Q(delay_counter[23]), .C(clk16MHz), .E(n27635), 
            .D(n1216), .R(n28814));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    SB_DFFESR delay_counter__i24 (.Q(delay_counter[24]), .C(clk16MHz), .E(n27635), 
            .D(n1215), .R(n28814));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    SB_DFFESR delay_counter__i25 (.Q(delay_counter[25]), .C(clk16MHz), .E(n27635), 
            .D(n1214), .R(n28814));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    SB_DFFESR delay_counter__i26 (.Q(delay_counter[26]), .C(clk16MHz), .E(n27635), 
            .D(n1213), .R(n28814));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    SB_DFFESR delay_counter__i27 (.Q(delay_counter[27]), .C(clk16MHz), .E(n27635), 
            .D(n1212), .R(n28814));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    SB_DFFESR delay_counter__i28 (.Q(delay_counter[28]), .C(clk16MHz), .E(n27635), 
            .D(n1211), .R(n28814));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    SB_DFFESR delay_counter__i29 (.Q(delay_counter[29]), .C(clk16MHz), .E(n27635), 
            .D(n1210), .R(n28814));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i23_1_lut (.I0(encoder1_position_scaled[22]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n3_adj_5796));   // verilog/TinyFPGA_B.v(323[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_DFFESR delay_counter__i30 (.Q(delay_counter[30]), .C(clk16MHz), .E(n27635), 
            .D(n1209), .R(n28814));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    SB_DFFESR delay_counter__i31 (.Q(delay_counter[31]), .C(clk16MHz), .E(n27635), 
            .D(n1208), .R(n28814));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    SB_LUT4 encoder0_position_30__I_0_i1445_3_lut (.I0(n2122), .I1(n2189), 
            .I2(n2148), .I3(GND_net), .O(n2221));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1445_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 n11566_bdd_4_lut_55427 (.I0(n11566), .I1(current[15]), .I2(duty[20]), 
            .I3(n11564), .O(n71174));
    defparam n11566_bdd_4_lut_55427.LUT_INIT = 16'he4aa;
    SB_LUT4 n71174_bdd_4_lut (.I0(n71174), .I1(duty[17]), .I2(n4909), 
            .I3(n11564), .O(pwm_setpoint_23__N_3[17]));
    defparam n71174_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 unary_minus_15_inv_0_i24_1_lut (.I0(duty[23]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(pwm_setpoint_23__N_207));   // verilog/TinyFPGA_B.v(119[24:29])
    defparam unary_minus_15_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_i1512_3_lut (.I0(n2221), .I1(n2288), 
            .I2(n2247), .I3(GND_net), .O(n2320));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1512_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 n11566_bdd_4_lut_55422 (.I0(n11566), .I1(current[15]), .I2(duty[19]), 
            .I3(n11564), .O(n71168));
    defparam n11566_bdd_4_lut_55422.LUT_INIT = 16'he4aa;
    SB_CARRY encoder0_position_30__I_0_unary_minus_2_add_3_11 (.CI(n52435), 
            .I0(GND_net), .I1(n24_adj_5914), .CO(n52436));
    SB_LUT4 n71168_bdd_4_lut (.I0(n71168), .I1(duty[16]), .I2(n4910), 
            .I3(n11564), .O(pwm_setpoint_23__N_3[16]));
    defparam n71168_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 encoder0_position_30__I_0_i1579_3_lut (.I0(n2320), .I1(n2387), 
            .I2(n2346), .I3(GND_net), .O(n2419));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1579_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_55432 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[18] [4]), .I2(\data_out_frame[19] [4]), 
            .I3(byte_transmit_counter[1]), .O(n71162));
    defparam byte_transmit_counter_0__bdd_4_lut_55432.LUT_INIT = 16'he4aa;
    SB_CARRY encoder0_position_30__I_0_add_1838_8 (.CI(n51797), .I0(n2728), 
            .I1(VCC_net), .CO(n51798));
    SB_LUT4 encoder0_position_30__I_0_i2043_3_lut (.I0(n3008), .I1(n3075), 
            .I2(n3039), .I3(GND_net), .O(n3107));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2043_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2042_3_lut (.I0(n3007), .I1(n3074), 
            .I2(n3039), .I3(GND_net), .O(n3106));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2042_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2049_3_lut (.I0(n3014), .I1(n3081), 
            .I2(n3039), .I3(GND_net), .O(n3113));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2049_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2048_3_lut (.I0(n3013), .I1(n3080), 
            .I2(n3039), .I3(GND_net), .O(n3112));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2048_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_adj_1771 (.I0(\data_out_frame[24] [2]), .I1(\data_out_frame[24] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n58978));
    defparam i1_2_lut_adj_1771.LUT_INIT = 16'h6666;
    SB_LUT4 encoder0_position_30__I_0_i2047_3_lut (.I0(n3012), .I1(n3079), 
            .I2(n3039), .I3(GND_net), .O(n3111));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2047_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2046_3_lut (.I0(n3011), .I1(n3078), 
            .I2(n3039), .I3(GND_net), .O(n3110));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2046_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2045_3_lut (.I0(n3010), .I1(n3077), 
            .I2(n3039), .I3(GND_net), .O(n3109));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2045_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 LessThan_1081_i9_2_lut (.I0(r_Clock_Count[4]), .I1(o_Rx_DV_N_3488[4]), 
            .I2(GND_net), .I3(GND_net), .O(n9_adj_5878));   // verilog/uart_rx.v(119[17:57])
    defparam LessThan_1081_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 encoder0_position_30__I_0_i2044_3_lut (.I0(n3009), .I1(n3076), 
            .I2(n3039), .I3(GND_net), .O(n3108));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2044_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2051_3_lut (.I0(n3016), .I1(n3083), 
            .I2(n3039), .I3(GND_net), .O(n3115));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2051_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 n71162_bdd_4_lut (.I0(n71162), .I1(\data_out_frame[17] [4]), 
            .I2(\data_out_frame[16] [4]), .I3(byte_transmit_counter[1]), 
            .O(n71165));
    defparam n71162_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 encoder0_position_30__I_0_i2050_3_lut (.I0(n3015), .I1(n3082), 
            .I2(n3039), .I3(GND_net), .O(n3114));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2050_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2054_3_lut (.I0(n3019), .I1(n3086), 
            .I2(n3039), .I3(GND_net), .O(n3118));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2054_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2053_3_lut (.I0(n3018), .I1(n3085), 
            .I2(n3039), .I3(GND_net), .O(n3117));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2053_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2052_3_lut (.I0(n3017), .I1(n3084), 
            .I2(n3039), .I3(GND_net), .O(n3116));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2052_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2062_3_lut (.I0(n3027), .I1(n3094), 
            .I2(n3039), .I3(GND_net), .O(n3126));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2062_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2055_3_lut (.I0(n3020), .I1(n3087), 
            .I2(n3039), .I3(GND_net), .O(n3119));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2055_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2060_3_lut (.I0(n3025), .I1(n3092), 
            .I2(n3039), .I3(GND_net), .O(n3124));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2060_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2056_3_lut (.I0(n3021), .I1(n3088), 
            .I2(n3039), .I3(GND_net), .O(n3120));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2056_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 LessThan_1081_i4_4_lut (.I0(r_Clock_Count[0]), .I1(o_Rx_DV_N_3488[1]), 
            .I2(r_Clock_Count[1]), .I3(o_Rx_DV_N_3488[0]), .O(n4_adj_5875));   // verilog/uart_rx.v(119[17:57])
    defparam LessThan_1081_i4_4_lut.LUT_INIT = 16'h4d0c;
    SB_LUT4 encoder0_position_30__I_0_i2063_3_lut (.I0(n3028), .I1(n3095), 
            .I2(n3039), .I3(GND_net), .O(n3127));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2063_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 LessThan_1081_i8_3_lut (.I0(n6_adj_5876), .I1(o_Rx_DV_N_3488[4]), 
            .I2(n9_adj_5878), .I3(GND_net), .O(n8_adj_5877));   // verilog/uart_rx.v(119[17:57])
    defparam LessThan_1081_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i54046_4_lut (.I0(n8_adj_5877), .I1(n4_adj_5875), .I2(n9_adj_5878), 
            .I3(n67828), .O(n69740));   // verilog/uart_rx.v(119[17:57])
    defparam i54046_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i54047_3_lut (.I0(n69740), .I1(o_Rx_DV_N_3488[5]), .I2(r_Clock_Count[5]), 
            .I3(GND_net), .O(n69741));   // verilog/uart_rx.v(119[17:57])
    defparam i54047_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 encoder0_position_30__I_0_i2064_3_lut (.I0(n3029), .I1(n3096), 
            .I2(n3039), .I3(GND_net), .O(n3128));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2064_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2058_3_lut (.I0(n3023), .I1(n3090), 
            .I2(n3039), .I3(GND_net), .O(n3122));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2058_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2061_3_lut (.I0(n3026), .I1(n3093), 
            .I2(n3039), .I3(GND_net), .O(n3125));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2061_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2059_3_lut (.I0(n3024), .I1(n3091), 
            .I2(n3039), .I3(GND_net), .O(n3123));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2059_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i53924_3_lut (.I0(n69741), .I1(o_Rx_DV_N_3488[6]), .I2(r_Clock_Count[6]), 
            .I3(GND_net), .O(n69618));   // verilog/uart_rx.v(119[17:57])
    defparam i53924_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 encoder0_position_30__I_0_i2057_3_lut (.I0(n3022), .I1(n3089), 
            .I2(n3039), .I3(GND_net), .O(n3121));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2057_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_add_2039_22_lut (.I0(GND_net), .I1(n3014), 
            .I2(VCC_net), .I3(n51889), .O(n3081)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2039_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_i2069_3_lut (.I0(n955), .I1(n3101), 
            .I2(n3039), .I3(GND_net), .O(n3133));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2069_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i52643_3_lut (.I0(n69618), .I1(o_Rx_DV_N_3488[7]), .I2(r_Clock_Count[7]), 
            .I3(GND_net), .O(n4935));   // verilog/uart_rx.v(119[17:57])
    defparam i52643_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 encoder0_position_30__I_0_i2068_3_lut (.I0(n3033), .I1(n3100), 
            .I2(n3039), .I3(GND_net), .O(n3132));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2068_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_4297_i2_3_lut (.I0(encoder0_position[1]), .I1(n31), .I2(encoder0_position[30]), 
            .I3(GND_net), .O(n956));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam mux_4297_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_i2067_3_lut (.I0(n3032), .I1(n3099), 
            .I2(n3039), .I3(GND_net), .O(n3131));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2067_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2066_3_lut (.I0(n3031), .I1(n3098), 
            .I2(n3039), .I3(GND_net), .O(n3130));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2066_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2065_3_lut (.I0(n3030), .I1(n3097), 
            .I2(n3039), .I3(GND_net), .O(n3129));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2065_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i54508_1_lut (.I0(n3138), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n70202));
    defparam i54508_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i29824_3_lut (.I0(n956), .I1(n3132), .I2(n3133), .I3(GND_net), 
            .O(n43725));
    defparam i29824_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i1_4_lut_adj_1772 (.I0(n3121), .I1(n3123), .I2(n3125), .I3(n3122), 
            .O(n62749));
    defparam i1_4_lut_adj_1772.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1773 (.I0(o_Rx_DV_N_3488[12]), .I1(n4935), .I2(o_Rx_DV_N_3488[8]), 
            .I3(n61449), .O(n62157));
    defparam i1_4_lut_adj_1773.LUT_INIT = 16'hfeff;
    SB_LUT4 i1_4_lut_adj_1774 (.I0(n3128), .I1(n3127), .I2(n3120), .I3(n3124), 
            .O(n62751));
    defparam i1_4_lut_adj_1774.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1775 (.I0(n62751), .I1(n62749), .I2(n3119), .I3(n3126), 
            .O(n62755));
    defparam i1_4_lut_adj_1775.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_add_3_10_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n25_adj_5915), .I3(n52434), .O(n25_adj_5723)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_unary_minus_2_add_3_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1776 (.I0(n3129), .I1(n43725), .I2(n3130), .I3(n3131), 
            .O(n60467));
    defparam i1_4_lut_adj_1776.LUT_INIT = 16'ha080;
    SB_LUT4 i1_4_lut_adj_1777 (.I0(o_Rx_DV_N_3488[24]), .I1(n29_adj_5857), 
            .I2(n23_adj_5860), .I3(n62157), .O(n62163));
    defparam i1_4_lut_adj_1777.LUT_INIT = 16'hfffe;
    SB_CARRY encoder0_position_30__I_0_unary_minus_2_add_3_10 (.CI(n52434), 
            .I0(GND_net), .I1(n25_adj_5915), .CO(n52435));
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_add_3_9_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n26_adj_5916), .I3(n52433), .O(n26)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_unary_minus_2_add_3_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1778 (.I0(n3116), .I1(n3117), .I2(n62755), .I3(n3118), 
            .O(n62761));
    defparam i1_4_lut_adj_1778.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1779 (.I0(n3114), .I1(n3115), .I2(n62761), .I3(n60467), 
            .O(n62767));
    defparam i1_4_lut_adj_1779.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1780 (.I0(n3111), .I1(n3112), .I2(n3113), .I3(n62767), 
            .O(n62773));
    defparam i1_4_lut_adj_1780.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1781 (.I0(n3108), .I1(n3109), .I2(n3110), .I3(n62773), 
            .O(n62779));
    defparam i1_4_lut_adj_1781.LUT_INIT = 16'hfffe;
    SB_LUT4 i54511_4_lut (.I0(n3106), .I1(n3105), .I2(n3107), .I3(n62779), 
            .O(n3138));
    defparam i54511_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i24_1_lut (.I0(encoder1_position_scaled[23]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n2_adj_5797));   // verilog/TinyFPGA_B.v(323[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_16_inv_0_i1_1_lut (.I0(current[0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_5719));   // verilog/TinyFPGA_B.v(121[16:24])
    defparam unary_minus_16_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_245_i22_4_lut (.I0(encoder1_position_scaled[21]), .I1(displacement[21]), 
            .I2(n15_adj_5722), .I3(n15), .O(motor_state_23__N_91[21]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i22_4_lut.LUT_INIT = 16'h0aca;
    SB_CARRY encoder0_position_30__I_0_unary_minus_2_add_3_9 (.CI(n52433), 
            .I0(GND_net), .I1(n26_adj_5916), .CO(n52434));
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_add_3_8_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n27_adj_5917), .I3(n52432), .O(n27)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_unary_minus_2_add_3_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_adj_1782 (.I0(\data_out_frame[20] [4]), .I1(n59223), 
            .I2(GND_net), .I3(GND_net), .O(n58938));   // verilog/coms.v(100[12:26])
    defparam i1_2_lut_adj_1782.LUT_INIT = 16'h6666;
    SB_LUT4 encoder0_position_30__I_0_i1646_3_lut (.I0(n2419), .I1(n2486), 
            .I2(n2445), .I3(GND_net), .O(n2518));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1646_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_30__I_0_unary_minus_2_add_3_8 (.CI(n52432), 
            .I0(GND_net), .I1(n27_adj_5917), .CO(n52433));
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_add_3_7_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n28_adj_5918), .I3(n52431), .O(n28)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_unary_minus_2_add_3_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_unary_minus_2_add_3_7 (.CI(n52431), 
            .I0(GND_net), .I1(n28_adj_5918), .CO(n52432));
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_add_3_6_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n29_adj_5919), .I3(n52430), .O(n29)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_unary_minus_2_add_3_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_unary_minus_2_add_3_6 (.CI(n52430), 
            .I0(GND_net), .I1(n29_adj_5919), .CO(n52431));
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_add_3_5_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n30_adj_5920), .I3(n52429), .O(n30)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_unary_minus_2_add_3_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_inv_0_i2_1_lut (.I0(current[1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n24_adj_5718));   // verilog/TinyFPGA_B.v(121[16:24])
    defparam unary_minus_16_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_i1975_3_lut (.I0(n2908), .I1(n2975), 
            .I2(n2940), .I3(GND_net), .O(n3007));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1975_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1977_3_lut (.I0(n2910), .I1(n2977), 
            .I2(n2940), .I3(GND_net), .O(n3009));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1977_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1976_3_lut (.I0(n2909), .I1(n2976), 
            .I2(n2940), .I3(GND_net), .O(n3008));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1976_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1979_3_lut (.I0(n2912), .I1(n2979), 
            .I2(n2940), .I3(GND_net), .O(n3011));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1979_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1978_3_lut (.I0(n2911), .I1(n2978), 
            .I2(n2940), .I3(GND_net), .O(n3010));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1978_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i54547_1_lut (.I0(n3039), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n70241));
    defparam i54547_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_4_lut_adj_1783 (.I0(n3027), .I1(n3021), .I2(n3020), .I3(n3023), 
            .O(n63321));
    defparam i1_4_lut_adj_1783.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_3_lut (.I0(n3026), .I1(n3018), .I2(n3019), .I3(GND_net), 
            .O(n63319));
    defparam i1_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i29872_4_lut (.I0(n955), .I1(n3031), .I2(n3032), .I3(n3033), 
            .O(n43773));
    defparam i29872_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 i1_4_lut_adj_1784 (.I0(n3016), .I1(n3017), .I2(n63319), .I3(n63321), 
            .O(n63327));
    defparam i1_4_lut_adj_1784.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1785 (.I0(n3029), .I1(n63327), .I2(n43773), .I3(n3030), 
            .O(n63329));
    defparam i1_4_lut_adj_1785.LUT_INIT = 16'heccc;
    SB_LUT4 i1_4_lut_adj_1786 (.I0(n3022), .I1(n3024), .I2(n3028), .I3(n3025), 
            .O(n63351));
    defparam i1_4_lut_adj_1786.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1787 (.I0(n3010), .I1(n3011), .I2(n3014), .I3(n63329), 
            .O(n63335));
    defparam i1_4_lut_adj_1787.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1788 (.I0(n3012), .I1(n3013), .I2(n3015), .I3(n63351), 
            .O(n63357));
    defparam i1_4_lut_adj_1788.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1789 (.I0(n3008), .I1(n63357), .I2(n63335), .I3(n3009), 
            .O(n63339));
    defparam i1_4_lut_adj_1789.LUT_INIT = 16'hfffe;
    SB_LUT4 i54550_3_lut (.I0(n3007), .I1(n3006), .I2(n63339), .I3(GND_net), 
            .O(n3039));
    defparam i54550_3_lut.LUT_INIT = 16'h0101;
    SB_CARRY encoder0_position_30__I_0_add_2039_22 (.CI(n51889), .I0(n3014), 
            .I1(VCC_net), .CO(n51890));
    SB_CARRY encoder0_position_30__I_0_unary_minus_2_add_3_5 (.CI(n52429), 
            .I0(GND_net), .I1(n30_adj_5920), .CO(n52430));
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_add_3_4_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n31_adj_5921), .I3(n52428), .O(n31)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_unary_minus_2_add_3_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_unary_minus_2_add_3_4 (.CI(n52428), 
            .I0(GND_net), .I1(n31_adj_5921), .CO(n52429));
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_add_3_3_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n32_adj_5922), .I3(n52427), .O(n32)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_unary_minus_2_add_3_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1838_7_lut (.I0(GND_net), .I1(n2729), 
            .I2(GND_net), .I3(n51796), .O(n2796)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1838_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_151_5_lut (.I0(GND_net), .I1(delay_counter[3]), .I2(GND_net), 
            .I3(n50980), .O(n1236)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i11_2_lut (.I0(\data_out_frame[18] [4]), .I1(\data_out_frame[18] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n25764));   // verilog/coms.v(100[12:26])
    defparam i11_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY encoder0_position_30__I_0_unary_minus_2_add_3_3 (.CI(n52427), 
            .I0(GND_net), .I1(n32_adj_5922), .CO(n52428));
    SB_CARRY encoder0_position_30__I_0_unary_minus_2_add_3_2 (.CI(VCC_net), 
            .I0(GND_net), .I1(VCC_net), .CO(n52427));
    SB_DFF pwm_setpoint_i1 (.Q(pwm_setpoint[1]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[1]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_DFF pwm_setpoint_i3 (.Q(pwm_setpoint[3]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[3]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_CARRY encoder0_position_30__I_0_add_1838_7 (.CI(n51796), .I0(n2729), 
            .I1(GND_net), .CO(n51797));
    SB_LUT4 encoder0_position_30__I_0_add_2039_21_lut (.I0(GND_net), .I1(n3015), 
            .I2(VCC_net), .I3(n51888), .O(n3082)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2039_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2039_21 (.CI(n51888), .I0(n3015), 
            .I1(VCC_net), .CO(n51889));
    SB_IO INLC_pad (.PACKAGE_PIN(INLC), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INLC_c_0));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INLC_pad.PIN_TYPE = 6'b011001;
    defparam INLC_pad.PULLUP = 1'b0;
    defparam INLC_pad.NEG_TRIGGER = 1'b0;
    defparam INLC_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 encoder0_position_30__I_0_i1713_3_lut (.I0(n2518), .I1(n2585), 
            .I2(n2544), .I3(GND_net), .O(n2617));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1713_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_1582_i23_3_lut (.I0(duty[23]), .I1(duty[22]), .I2(n260), 
            .I3(GND_net), .O(n12169));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1582_i23_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 n11566_bdd_4_lut_55417 (.I0(n11566), .I1(current[15]), .I2(duty[18]), 
            .I3(n11564), .O(n71156));
    defparam n11566_bdd_4_lut_55417.LUT_INIT = 16'he4aa;
    SB_LUT4 mux_245_i23_4_lut (.I0(encoder1_position_scaled[22]), .I1(displacement[22]), 
            .I2(n15_adj_5722), .I3(n15), .O(motor_state_23__N_91[22]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i23_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 encoder0_position_30__I_0_add_2039_20_lut (.I0(GND_net), .I1(n3016), 
            .I2(VCC_net), .I3(n51887), .O(n3083)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2039_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 n71156_bdd_4_lut (.I0(n71156), .I1(duty[15]), .I2(n4911), 
            .I3(n11564), .O(pwm_setpoint_23__N_3[15]));
    defparam n71156_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_CARRY encoder0_position_30__I_0_add_2039_20 (.CI(n51887), .I0(n3016), 
            .I1(VCC_net), .CO(n51888));
    SB_LUT4 encoder0_position_30__I_0_add_2039_19_lut (.I0(GND_net), .I1(n3017), 
            .I2(VCC_net), .I3(n51886), .O(n3084)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2039_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i54677_1_lut (.I0(n2544), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n70371));
    defparam i54677_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_30__I_0_add_1570_18 (.CI(n51717), .I0(n2318), 
            .I1(VCC_net), .CO(n51718));
    SB_LUT4 unary_minus_16_inv_0_i3_1_lut (.I0(current[2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_5717));   // verilog/TinyFPGA_B.v(121[16:24])
    defparam unary_minus_16_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_30__I_0_add_2039_19 (.CI(n51886), .I0(n3017), 
            .I1(VCC_net), .CO(n51887));
    SB_LUT4 unary_minus_16_inv_0_i4_1_lut (.I0(current[3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n22_adj_5716));   // verilog/TinyFPGA_B.v(121[16:24])
    defparam unary_minus_16_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_GB_IO CLK_pad (.PACKAGE_PIN(CLK), .OUTPUT_ENABLE(VCC_net), .GLOBAL_BUFFER_OUTPUT(clk16MHz));   // verilog/TinyFPGA_B.v(3[9:12])
    defparam CLK_pad.PIN_TYPE = 6'b000001;
    defparam CLK_pad.PULLUP = 1'b0;
    defparam CLK_pad.NEG_TRIGGER = 1'b0;
    defparam CLK_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 encoder0_position_30__I_0_add_2039_18_lut (.I0(GND_net), .I1(n3018), 
            .I2(VCC_net), .I3(n51885), .O(n3085)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2039_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1838_6_lut (.I0(GND_net), .I1(n2730), 
            .I2(GND_net), .I3(n51795), .O(n2797)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1838_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1838_6 (.CI(n51795), .I0(n2730), 
            .I1(GND_net), .CO(n51796));
    SB_LUT4 encoder0_position_30__I_0_add_1570_17_lut (.I0(GND_net), .I1(n2319), 
            .I2(VCC_net), .I3(n51716), .O(n2386)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1570_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_i1780_3_lut (.I0(n2617), .I1(n2684), 
            .I2(n2643), .I3(GND_net), .O(n2716));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1780_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_add_1101_16_lut (.I0(n70615), .I1(n1620), 
            .I2(VCC_net), .I3(n51424), .O(n1719)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1101_16_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_30__I_0_add_1101_15_lut (.I0(GND_net), .I1(n1621), 
            .I2(VCC_net), .I3(n51423), .O(n1688)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1101_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_699_9 (.CI(n51304), .I0(n1027), 
            .I1(VCC_net), .CO(n51305));
    SB_CARRY add_151_14 (.CI(n50989), .I0(delay_counter[12]), .I1(GND_net), 
            .CO(n50990));
    SB_LUT4 encoder0_position_30__I_0_add_699_8_lut (.I0(GND_net), .I1(n1028), 
            .I2(VCC_net), .I3(n51303), .O(n1095)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_699_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1101_15 (.CI(n51423), .I0(n1621), 
            .I1(VCC_net), .CO(n51424));
    SB_CARRY encoder0_position_30__I_0_add_699_8 (.CI(n51303), .I0(n1028), 
            .I1(VCC_net), .CO(n51304));
    SB_LUT4 encoder0_position_30__I_0_add_699_7_lut (.I0(GND_net), .I1(n1029), 
            .I2(GND_net), .I3(n51302), .O(n1096)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_699_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_699_7 (.CI(n51302), .I0(n1029), 
            .I1(GND_net), .CO(n51303));
    SB_LUT4 encoder0_position_30__I_0_add_1101_14_lut (.I0(GND_net), .I1(n1622), 
            .I2(VCC_net), .I3(n51422), .O(n1689)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1101_14_lut.LUT_INIT = 16'hC33C;
    SB_DFF pwm_setpoint_i2 (.Q(pwm_setpoint[2]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[2]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_LUT4 encoder0_position_30__I_0_add_1838_5_lut (.I0(GND_net), .I1(n2731), 
            .I2(VCC_net), .I3(n51794), .O(n2798)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1838_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1101_14 (.CI(n51422), .I0(n1622), 
            .I1(VCC_net), .CO(n51423));
    SB_LUT4 i54579_1_lut (.I0(n2940), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n70273));
    defparam i54579_1_lut.LUT_INIT = 16'h5555;
    SB_DFF encoder0_position_scaled_i23 (.Q(encoder0_position_scaled[23]), 
           .C(clk16MHz), .D(encoder0_position_scaled_23__N_43[23]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_LUT4 encoder0_position_30__I_0_add_699_6_lut (.I0(GND_net), .I1(n1030), 
            .I2(GND_net), .I3(n51301), .O(n1097)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_699_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1101_13_lut (.I0(GND_net), .I1(n1623), 
            .I2(VCC_net), .I3(n51421), .O(n1690)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1101_13_lut.LUT_INIT = 16'hC33C;
    SB_DFF encoder0_position_scaled_i22 (.Q(encoder0_position_scaled[22]), 
           .C(clk16MHz), .D(encoder0_position_scaled_23__N_43[22]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_CARRY encoder0_position_30__I_0_add_699_6 (.CI(n51301), .I0(n1030), 
            .I1(GND_net), .CO(n51302));
    SB_LUT4 mux_4297_i11_3_lut (.I0(encoder0_position[10]), .I1(n22_adj_5726), 
            .I2(encoder0_position[30]), .I3(GND_net), .O(n947));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam mux_4297_i11_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_add_699_5_lut (.I0(GND_net), .I1(n1031), 
            .I2(VCC_net), .I3(n51300), .O(n1098)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_699_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2039_18 (.CI(n51885), .I0(n3018), 
            .I1(VCC_net), .CO(n51886));
    SB_CARRY encoder0_position_30__I_0_add_1570_17 (.CI(n51716), .I0(n2319), 
            .I1(VCC_net), .CO(n51717));
    SB_DFF encoder0_position_scaled_i21 (.Q(encoder0_position_scaled[21]), 
           .C(clk16MHz), .D(encoder0_position_scaled_23__N_43[21]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF encoder0_position_scaled_i20 (.Q(encoder0_position_scaled[20]), 
           .C(clk16MHz), .D(encoder0_position_scaled_23__N_43[20]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF encoder0_position_scaled_i19 (.Q(encoder0_position_scaled[19]), 
           .C(clk16MHz), .D(encoder0_position_scaled_23__N_43[19]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_CARRY encoder0_position_30__I_0_add_699_5 (.CI(n51300), .I0(n1031), 
            .I1(VCC_net), .CO(n51301));
    SB_DFF encoder0_position_scaled_i18 (.Q(encoder0_position_scaled[18]), 
           .C(clk16MHz), .D(encoder0_position_scaled_23__N_43[18]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_LUT4 encoder0_position_30__I_0_i1525_3_lut (.I0(n947), .I1(n2301), 
            .I2(n2247), .I3(GND_net), .O(n2333));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1525_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_30__I_0_add_1101_13 (.CI(n51421), .I0(n1623), 
            .I1(VCC_net), .CO(n51422));
    SB_LUT4 encoder0_position_30__I_0_add_699_4_lut (.I0(GND_net), .I1(n1032), 
            .I2(GND_net), .I3(n51299), .O(n1099)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_699_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_i1592_3_lut (.I0(n2333), .I1(n2400), 
            .I2(n2346), .I3(GND_net), .O(n2432));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1592_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_add_2039_17_lut (.I0(GND_net), .I1(n3019), 
            .I2(VCC_net), .I3(n51884), .O(n3086)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2039_17_lut.LUT_INIT = 16'hC33C;
    SB_DFF encoder0_position_scaled_i17 (.Q(encoder0_position_scaled[17]), 
           .C(clk16MHz), .D(encoder0_position_scaled_23__N_43[17]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF encoder0_position_scaled_i16 (.Q(encoder0_position_scaled[16]), 
           .C(clk16MHz), .D(encoder0_position_scaled_23__N_43[16]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF encoder0_position_scaled_i15 (.Q(encoder0_position_scaled[15]), 
           .C(clk16MHz), .D(encoder0_position_scaled_23__N_43[15]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF encoder0_position_scaled_i14 (.Q(encoder0_position_scaled[14]), 
           .C(clk16MHz), .D(encoder0_position_scaled_23__N_43[14]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF encoder0_position_scaled_i13 (.Q(encoder0_position_scaled[13]), 
           .C(clk16MHz), .D(encoder0_position_scaled_23__N_43[13]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_CARRY encoder0_position_30__I_0_add_699_4 (.CI(n51299), .I0(n1032), 
            .I1(GND_net), .CO(n51300));
    SB_LUT4 encoder0_position_30__I_0_add_1101_12_lut (.I0(GND_net), .I1(n1624), 
            .I2(VCC_net), .I3(n51420), .O(n1691)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1101_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_i1659_3_lut (.I0(n2432), .I1(n2499), 
            .I2(n2445), .I3(GND_net), .O(n2531));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1659_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_30__I_0_add_1838_5 (.CI(n51794), .I0(n2731), 
            .I1(VCC_net), .CO(n51795));
    SB_LUT4 encoder0_position_30__I_0_i1726_3_lut (.I0(n2531), .I1(n2598), 
            .I2(n2544), .I3(GND_net), .O(n2630));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1726_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1793_3_lut (.I0(n2630), .I1(n2697), 
            .I2(n2643), .I3(GND_net), .O(n2729));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1793_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_30__I_0_add_1101_12 (.CI(n51420), .I0(n1624), 
            .I1(VCC_net), .CO(n51421));
    SB_LUT4 encoder0_position_30__I_0_add_699_3_lut (.I0(GND_net), .I1(n1033), 
            .I2(VCC_net), .I3(n51298), .O(n1100)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_699_3_lut.LUT_INIT = 16'hC33C;
    SB_DFF encoder0_position_scaled_i12 (.Q(encoder0_position_scaled[12]), 
           .C(clk16MHz), .D(encoder0_position_scaled_23__N_43[12]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF encoder0_position_scaled_i11 (.Q(encoder0_position_scaled[11]), 
           .C(clk16MHz), .D(encoder0_position_scaled_23__N_43[11]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_CARRY encoder0_position_30__I_0_add_699_3 (.CI(n51298), .I0(n1033), 
            .I1(VCC_net), .CO(n51299));
    SB_DFF encoder0_position_scaled_i10 (.Q(encoder0_position_scaled[10]), 
           .C(clk16MHz), .D(encoder0_position_scaled_23__N_43[10]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF encoder0_position_scaled_i9 (.Q(encoder0_position_scaled[9]), .C(clk16MHz), 
           .D(encoder0_position_scaled_23__N_43[9]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF encoder0_position_scaled_i8 (.Q(encoder0_position_scaled[8]), .C(clk16MHz), 
           .D(encoder0_position_scaled_23__N_43[8]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF encoder0_position_scaled_i7 (.Q(encoder0_position_scaled[7]), .C(clk16MHz), 
           .D(encoder0_position_scaled_23__N_43[7]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_LUT4 encoder0_position_30__I_0_add_1101_11_lut (.I0(GND_net), .I1(n1625), 
            .I2(VCC_net), .I3(n51419), .O(n1692)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1101_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_inv_0_i2_1_lut (.I0(encoder0_position[0]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n32_adj_5922));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_unary_minus_2_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_DFF encoder0_position_scaled_i6 (.Q(encoder0_position_scaled[6]), .C(clk16MHz), 
           .D(encoder0_position_scaled_23__N_43[6]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF encoder0_position_scaled_i5 (.Q(encoder0_position_scaled[5]), .C(clk16MHz), 
           .D(encoder0_position_scaled_23__N_43[5]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF encoder0_position_scaled_i4 (.Q(encoder0_position_scaled[4]), .C(clk16MHz), 
           .D(encoder0_position_scaled_23__N_43[4]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF encoder0_position_scaled_i3 (.Q(encoder0_position_scaled[3]), .C(clk16MHz), 
           .D(encoder0_position_scaled_23__N_43[3]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_inv_0_i3_1_lut (.I0(encoder0_position[1]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n31_adj_5921));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_unary_minus_2_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_DFF encoder0_position_scaled_i2 (.Q(encoder0_position_scaled[2]), .C(clk16MHz), 
           .D(encoder0_position_scaled_23__N_43[2]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF encoder0_position_scaled_i1 (.Q(encoder0_position_scaled[1]), .C(clk16MHz), 
           .D(encoder0_position_scaled_23__N_43[1]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_LUT4 encoder0_position_30__I_0_add_1838_4_lut (.I0(GND_net), .I1(n2732), 
            .I2(GND_net), .I3(n51793), .O(n2799)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1838_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_699_2_lut (.I0(GND_net), .I1(n521), 
            .I2(GND_net), .I3(VCC_net), .O(n1101)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_699_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1101_11 (.CI(n51419), .I0(n1625), 
            .I1(VCC_net), .CO(n51420));
    SB_LUT4 encoder0_position_30__I_0_add_1570_16_lut (.I0(GND_net), .I1(n2320), 
            .I2(VCC_net), .I3(n51715), .O(n2387)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1570_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1101_10_lut (.I0(GND_net), .I1(n1626), 
            .I2(VCC_net), .I3(n51418), .O(n1693)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1101_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_i1847_3_lut (.I0(n2716), .I1(n2783), 
            .I2(n2742), .I3(GND_net), .O(n2815));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1847_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_30__I_0_add_699_2 (.CI(VCC_net), .I0(n521), 
            .I1(GND_net), .CO(n51298));
    SB_LUT4 i1_4_lut_adj_1790 (.I0(control_mode[6]), .I1(control_mode[2]), 
            .I2(control_mode[4]), .I3(control_mode[5]), .O(n63553));   // verilog/TinyFPGA_B.v(286[5:22])
    defparam i1_4_lut_adj_1790.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_inv_0_i4_1_lut (.I0(encoder0_position[2]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n30_adj_5920));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_unary_minus_2_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_3_lut_adj_1791 (.I0(n63553), .I1(control_mode[7]), .I2(control_mode[3]), 
            .I3(GND_net), .O(n42369));   // verilog/TinyFPGA_B.v(286[5:22])
    defparam i1_3_lut_adj_1791.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_2_lut_adj_1792 (.I0(n25385), .I1(control_mode[1]), .I2(GND_net), 
            .I3(GND_net), .O(n15));   // verilog/TinyFPGA_B.v(287[5:22])
    defparam i1_2_lut_adj_1792.LUT_INIT = 16'hbbbb;
    SB_LUT4 i1_3_lut_adj_1793 (.I0(control_mode[0]), .I1(n42369), .I2(control_mode[1]), 
            .I3(GND_net), .O(n15_adj_5722));   // verilog/TinyFPGA_B.v(286[5:22])
    defparam i1_3_lut_adj_1793.LUT_INIT = 16'hfdfd;
    SB_LUT4 i16_4_lut_adj_1794 (.I0(encoder1_position_scaled[23]), .I1(displacement[23]), 
            .I2(n15_adj_5722), .I3(n15), .O(n15_adj_5872));
    defparam i16_4_lut_adj_1794.LUT_INIT = 16'h0aca;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_inv_0_i5_1_lut (.I0(encoder0_position[3]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n29_adj_5919));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_unary_minus_2_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_inv_0_i6_1_lut (.I0(encoder0_position[4]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n28_adj_5918));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_unary_minus_2_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_inv_0_i7_1_lut (.I0(encoder0_position[5]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n27_adj_5917));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_unary_minus_2_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_30__I_0_add_1101_10 (.CI(n51418), .I0(n1626), 
            .I1(VCC_net), .CO(n51419));
    SB_LUT4 encoder0_position_30__I_0_add_1101_9_lut (.I0(GND_net), .I1(n1627), 
            .I2(VCC_net), .I3(n51417), .O(n1694)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1101_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_632_9_lut (.I0(n960), .I1(n927), 
            .I2(VCC_net), .I3(n51297), .O(n1026)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_632_9_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_30__I_0_add_632_8_lut (.I0(GND_net), .I1(n928), 
            .I2(VCC_net), .I3(n51296), .O(n995)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_632_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1570_16 (.CI(n51715), .I0(n2320), 
            .I1(VCC_net), .CO(n51716));
    SB_CARRY encoder0_position_30__I_0_add_2039_17 (.CI(n51884), .I0(n3019), 
            .I1(VCC_net), .CO(n51885));
    SB_LUT4 encoder0_position_30__I_0_add_1570_15_lut (.I0(GND_net), .I1(n2321), 
            .I2(VCC_net), .I3(n51714), .O(n2388)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1570_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_632_8 (.CI(n51296), .I0(n928), 
            .I1(VCC_net), .CO(n51297));
    SB_LUT4 encoder0_position_30__I_0_add_632_7_lut (.I0(GND_net), .I1(n929), 
            .I2(GND_net), .I3(n51295), .O(n996)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_632_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1101_9 (.CI(n51417), .I0(n1627), 
            .I1(VCC_net), .CO(n51418));
    SB_CARRY encoder0_position_30__I_0_add_632_7 (.CI(n51295), .I0(n929), 
            .I1(GND_net), .CO(n51296));
    SB_LUT4 encoder0_position_30__I_0_add_1101_8_lut (.I0(GND_net), .I1(n1628), 
            .I2(VCC_net), .I3(n51416), .O(n1695)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1101_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1570_15 (.CI(n51714), .I0(n2321), 
            .I1(VCC_net), .CO(n51715));
    SB_LUT4 encoder0_position_30__I_0_add_632_6_lut (.I0(GND_net), .I1(n930), 
            .I2(GND_net), .I3(n51294), .O(n997)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_632_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1101_8 (.CI(n51416), .I0(n1628), 
            .I1(VCC_net), .CO(n51417));
    SB_LUT4 encoder0_position_30__I_0_add_1101_7_lut (.I0(GND_net), .I1(n1629), 
            .I2(GND_net), .I3(n51415), .O(n1696)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1101_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1101_7 (.CI(n51415), .I0(n1629), 
            .I1(GND_net), .CO(n51416));
    SB_LUT4 encoder0_position_30__I_0_add_1101_6_lut (.I0(GND_net), .I1(n1630), 
            .I2(GND_net), .I3(n51414), .O(n1697)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1101_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1838_4 (.CI(n51793), .I0(n2732), 
            .I1(GND_net), .CO(n51794));
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_inv_0_i8_1_lut (.I0(encoder0_position[6]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n26_adj_5916));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_unary_minus_2_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_30__I_0_add_632_6 (.CI(n51294), .I0(n930), 
            .I1(GND_net), .CO(n51295));
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_inv_0_i9_1_lut (.I0(encoder0_position[7]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n25_adj_5915));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_unary_minus_2_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_add_632_5_lut (.I0(GND_net), .I1(n931), 
            .I2(VCC_net), .I3(n51293), .O(n998)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_632_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_2039_16_lut (.I0(GND_net), .I1(n3020), 
            .I2(VCC_net), .I3(n51883), .O(n3087)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2039_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_i1982_3_lut (.I0(n2915), .I1(n2982), 
            .I2(n2940), .I3(GND_net), .O(n3014));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1982_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_30__I_0_add_632_5 (.CI(n51293), .I0(n931), 
            .I1(VCC_net), .CO(n51294));
    SB_LUT4 encoder0_position_30__I_0_add_632_4_lut (.I0(GND_net), .I1(n932), 
            .I2(GND_net), .I3(n51292), .O(n999)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_632_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1838_3_lut (.I0(GND_net), .I1(n2733), 
            .I2(VCC_net), .I3(n51792), .O(n2800)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1838_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_632_4 (.CI(n51292), .I0(n932), 
            .I1(GND_net), .CO(n51293));
    SB_CARRY encoder0_position_30__I_0_add_2039_16 (.CI(n51883), .I0(n3020), 
            .I1(VCC_net), .CO(n51884));
    SB_LUT4 i14_2_lut (.I0(\data_out_frame[18] [7]), .I1(\data_out_frame[18] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n2076));   // verilog/coms.v(100[12:26])
    defparam i14_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1795 (.I0(n70020), .I1(n59055), .I2(GND_net), 
            .I3(GND_net), .O(n59027));
    defparam i1_2_lut_adj_1795.LUT_INIT = 16'h9999;
    SB_CARRY encoder0_position_30__I_0_add_1101_6 (.CI(n51414), .I0(n1630), 
            .I1(GND_net), .CO(n51415));
    SB_CARRY encoder0_position_30__I_0_add_1838_3 (.CI(n51792), .I0(n2733), 
            .I1(VCC_net), .CO(n51793));
    SB_LUT4 encoder0_position_30__I_0_add_2039_15_lut (.I0(GND_net), .I1(n3021), 
            .I2(VCC_net), .I3(n51882), .O(n3088)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2039_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1570_14_lut (.I0(GND_net), .I1(n2322), 
            .I2(VCC_net), .I3(n51713), .O(n2389)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1570_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_632_3_lut (.I0(GND_net), .I1(n933), 
            .I2(VCC_net), .I3(n51291), .O(n1000)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_632_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1838_2_lut (.I0(GND_net), .I1(n952), 
            .I2(GND_net), .I3(VCC_net), .O(n2801)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1838_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1101_5_lut (.I0(GND_net), .I1(n1631), 
            .I2(VCC_net), .I3(n51413), .O(n1698)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1101_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_632_3 (.CI(n51291), .I0(n933), 
            .I1(VCC_net), .CO(n51292));
    SB_LUT4 encoder0_position_30__I_0_add_632_2_lut (.I0(GND_net), .I1(n520), 
            .I2(GND_net), .I3(VCC_net), .O(n1001)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_632_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_632_2 (.CI(VCC_net), .I0(n520), 
            .I1(GND_net), .CO(n51291));
    SB_CARRY encoder0_position_30__I_0_add_1101_5 (.CI(n51413), .I0(n1631), 
            .I1(VCC_net), .CO(n51414));
    SB_LUT4 encoder0_position_30__I_0_add_565_8_lut (.I0(n861), .I1(n828), 
            .I2(VCC_net), .I3(n51290), .O(n927)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_565_8_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_30__I_0_add_565_7_lut (.I0(GND_net), .I1(n829), 
            .I2(GND_net), .I3(n51289), .O(n896)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_565_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 n11566_bdd_4_lut_55407 (.I0(n11566), .I1(current[15]), .I2(duty[17]), 
            .I3(n11564), .O(n71144));
    defparam n11566_bdd_4_lut_55407.LUT_INIT = 16'he4aa;
    SB_LUT4 encoder0_position_30__I_0_add_1302_19_lut (.I0(n70454), .I1(n1917), 
            .I2(VCC_net), .I3(n51527), .O(n2016)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1302_19_lut.LUT_INIT = 16'h8228;
    SB_LUT4 n71144_bdd_4_lut (.I0(n71144), .I1(duty[14]), .I2(n4912), 
            .I3(n11564), .O(pwm_setpoint_23__N_3[14]));
    defparam n71144_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_CARRY encoder0_position_30__I_0_add_1570_14 (.CI(n51713), .I0(n2322), 
            .I1(VCC_net), .CO(n51714));
    SB_LUT4 encoder0_position_30__I_0_add_1101_4_lut (.I0(GND_net), .I1(n1632), 
            .I2(GND_net), .I3(n51412), .O(n1699)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1101_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1302_18_lut (.I0(GND_net), .I1(n1918), 
            .I2(VCC_net), .I3(n51526), .O(n1985)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1302_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1101_4 (.CI(n51412), .I0(n1632), 
            .I1(GND_net), .CO(n51413));
    SB_LUT4 encoder0_position_30__I_0_add_1101_3_lut (.I0(GND_net), .I1(n1633), 
            .I2(VCC_net), .I3(n51411), .O(n1700)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1101_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1101_3 (.CI(n51411), .I0(n1633), 
            .I1(VCC_net), .CO(n51412));
    SB_CARRY encoder0_position_30__I_0_add_565_7 (.CI(n51289), .I0(n829), 
            .I1(GND_net), .CO(n51290));
    SB_LUT4 encoder0_position_30__I_0_add_565_6_lut (.I0(GND_net), .I1(n830), 
            .I2(GND_net), .I3(n51288), .O(n897)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_565_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1302_18 (.CI(n51526), .I0(n1918), 
            .I1(VCC_net), .CO(n51527));
    SB_CARRY encoder0_position_30__I_0_add_565_6 (.CI(n51288), .I0(n830), 
            .I1(GND_net), .CO(n51289));
    SB_LUT4 encoder0_position_30__I_0_add_1101_2_lut (.I0(GND_net), .I1(n941), 
            .I2(GND_net), .I3(VCC_net), .O(n1701)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1101_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_565_5_lut (.I0(GND_net), .I1(n831), 
            .I2(VCC_net), .I3(n51287), .O(n898)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_565_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1302_17_lut (.I0(GND_net), .I1(n1919), 
            .I2(VCC_net), .I3(n51525), .O(n1986)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1302_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_565_5 (.CI(n51287), .I0(n831), 
            .I1(VCC_net), .CO(n51288));
    SB_LUT4 encoder0_position_30__I_0_add_1570_13_lut (.I0(GND_net), .I1(n2323), 
            .I2(VCC_net), .I3(n51712), .O(n2390)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1570_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_i1854_3_lut (.I0(n2723), .I1(n2790), 
            .I2(n2742), .I3(GND_net), .O(n2822));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1854_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_add_565_4_lut (.I0(GND_net), .I1(n832), 
            .I2(GND_net), .I3(n51286), .O(n899)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_565_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1302_17 (.CI(n51525), .I0(n1919), 
            .I1(VCC_net), .CO(n51526));
    SB_CARRY encoder0_position_30__I_0_add_1570_13 (.CI(n51712), .I0(n2323), 
            .I1(VCC_net), .CO(n51713));
    SB_CARRY encoder0_position_30__I_0_add_1101_2 (.CI(VCC_net), .I0(n941), 
            .I1(GND_net), .CO(n51411));
    SB_CARRY encoder0_position_30__I_0_add_565_4 (.CI(n51286), .I0(n832), 
            .I1(GND_net), .CO(n51287));
    SB_CARRY encoder0_position_30__I_0_add_1838_2 (.CI(VCC_net), .I0(n952), 
            .I1(GND_net), .CO(n51792));
    SB_LUT4 i13_2_lut (.I0(\data_out_frame[16] [6]), .I1(\data_out_frame[16] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n26372));   // verilog/coms.v(100[12:26])
    defparam i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 encoder0_position_30__I_0_add_565_3_lut (.I0(GND_net), .I1(n833), 
            .I2(VCC_net), .I3(n51285), .O(n900)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_565_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2039_15 (.CI(n51882), .I0(n3021), 
            .I1(VCC_net), .CO(n51883));
    SB_LUT4 encoder0_position_30__I_0_add_2039_14_lut (.I0(GND_net), .I1(n3022), 
            .I2(VCC_net), .I3(n51881), .O(n3089)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2039_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2039_14 (.CI(n51881), .I0(n3022), 
            .I1(VCC_net), .CO(n51882));
    SB_LUT4 add_151_13_lut (.I0(GND_net), .I1(delay_counter[11]), .I2(GND_net), 
            .I3(n50988), .O(n1228)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_13_lut.LUT_INIT = 16'hC33C;
    SB_IO CS_pad (.PACKAGE_PIN(CS), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(CS_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam CS_pad.PIN_TYPE = 6'b011001;
    defparam CS_pad.PULLUP = 1'b0;
    defparam CS_pad.NEG_TRIGGER = 1'b0;
    defparam CS_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 encoder0_position_30__I_0_add_1302_16_lut (.I0(GND_net), .I1(n1920), 
            .I2(VCC_net), .I3(n51524), .O(n1987)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1302_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1570_12_lut (.I0(GND_net), .I1(n2324), 
            .I2(VCC_net), .I3(n51711), .O(n2391)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1570_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1302_16 (.CI(n51524), .I0(n1920), 
            .I1(VCC_net), .CO(n51525));
    SB_CARRY encoder0_position_30__I_0_add_565_3 (.CI(n51285), .I0(n833), 
            .I1(VCC_net), .CO(n51286));
    SB_CARRY encoder0_position_30__I_0_add_1570_12 (.CI(n51711), .I0(n2324), 
            .I1(VCC_net), .CO(n51712));
    SB_LUT4 encoder0_position_30__I_0_add_1771_26_lut (.I0(n70427), .I1(n2610), 
            .I2(VCC_net), .I3(n51791), .O(n2709)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1771_26_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_30__I_0_add_2039_13_lut (.I0(GND_net), .I1(n3023), 
            .I2(VCC_net), .I3(n51880), .O(n3090)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2039_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1771_25_lut (.I0(GND_net), .I1(n2611), 
            .I2(VCC_net), .I3(n51790), .O(n2678)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1771_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1570_11_lut (.I0(GND_net), .I1(n2325), 
            .I2(VCC_net), .I3(n51710), .O(n2392)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1570_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1302_15_lut (.I0(GND_net), .I1(n1921), 
            .I2(VCC_net), .I3(n51523), .O(n1988)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1302_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_565_2_lut (.I0(GND_net), .I1(n519), 
            .I2(GND_net), .I3(VCC_net), .O(n901)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_565_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_11_i23_2_lut (.I0(current[11]), .I1(duty[11]), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_5741));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i23_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY encoder0_position_30__I_0_add_565_2 (.CI(VCC_net), .I0(n519), 
            .I1(GND_net), .CO(n51285));
    SB_LUT4 LessThan_11_i7_2_lut (.I0(current[3]), .I1(duty[3]), .I2(GND_net), 
            .I3(GND_net), .O(n7_adj_5752));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i7_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY encoder0_position_30__I_0_add_1771_25 (.CI(n51790), .I0(n2611), 
            .I1(VCC_net), .CO(n51791));
    SB_CARRY encoder0_position_30__I_0_add_1570_11 (.CI(n51710), .I0(n2325), 
            .I1(VCC_net), .CO(n51711));
    SB_LUT4 LessThan_11_i9_2_lut (.I0(current[4]), .I1(duty[4]), .I2(GND_net), 
            .I3(GND_net), .O(n9_adj_5750));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_11_i17_2_lut (.I0(current[8]), .I1(duty[8]), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_5744));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i17_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY encoder0_position_30__I_0_add_1302_15 (.CI(n51523), .I0(n1921), 
            .I1(VCC_net), .CO(n51524));
    SB_LUT4 encoder0_position_30__I_0_add_1302_14_lut (.I0(GND_net), .I1(n1922), 
            .I2(VCC_net), .I3(n51522), .O(n1989)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1302_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1570_10_lut (.I0(GND_net), .I1(n2326), 
            .I2(VCC_net), .I3(n51709), .O(n2393)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1570_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1302_14 (.CI(n51522), .I0(n1922), 
            .I1(VCC_net), .CO(n51523));
    SB_LUT4 encoder0_position_30__I_0_add_1302_13_lut (.I0(GND_net), .I1(n1923), 
            .I2(VCC_net), .I3(n51521), .O(n1990)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1302_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2452_7_lut (.I0(GND_net), .I1(n402), .I2(GND_net), .I3(n51284), 
            .O(n7442)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2452_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_11_i19_2_lut (.I0(current[9]), .I1(duty[9]), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_5743));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_2452_6_lut (.I0(GND_net), .I1(n403), .I2(GND_net), .I3(n51283), 
            .O(n7443)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2452_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2452_6 (.CI(n51283), .I0(n403), .I1(GND_net), .CO(n51284));
    SB_CARRY encoder0_position_30__I_0_add_1302_13 (.CI(n51521), .I0(n1923), 
            .I1(VCC_net), .CO(n51522));
    SB_LUT4 encoder0_position_30__I_0_add_1302_12_lut (.I0(GND_net), .I1(n1924), 
            .I2(VCC_net), .I3(n51520), .O(n1991)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1302_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1570_10 (.CI(n51709), .I0(n2326), 
            .I1(VCC_net), .CO(n51710));
    SB_LUT4 add_2452_5_lut (.I0(GND_net), .I1(n404), .I2(VCC_net), .I3(n51282), 
            .O(n7444)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2452_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_11_i21_2_lut (.I0(current[10]), .I1(duty[10]), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_5742));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i21_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY encoder0_position_30__I_0_add_1302_12 (.CI(n51520), .I0(n1924), 
            .I1(VCC_net), .CO(n51521));
    SB_LUT4 LessThan_11_i11_2_lut (.I0(current[5]), .I1(duty[5]), .I2(GND_net), 
            .I3(GND_net), .O(n11_adj_5748));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_11_i13_2_lut (.I0(current[6]), .I1(duty[6]), .I2(GND_net), 
            .I3(GND_net), .O(n13_adj_5747));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_11_i15_2_lut (.I0(current[7]), .I1(duty[7]), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_5746));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i15_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY encoder0_position_30__I_0_add_2039_13 (.CI(n51880), .I0(n3023), 
            .I1(VCC_net), .CO(n51881));
    SB_CARRY add_2452_5 (.CI(n51282), .I0(n404), .I1(VCC_net), .CO(n51283));
    SB_LUT4 LessThan_14_i15_2_lut (.I0(current[7]), .I1(current_limit[7]), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_5699));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam LessThan_14_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_14_i13_2_lut (.I0(current[6]), .I1(current_limit[6]), 
            .I2(GND_net), .I3(GND_net), .O(n13_adj_5700));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam LessThan_14_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 unary_minus_16_inv_0_i5_1_lut (.I0(current[4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_5715));   // verilog/TinyFPGA_B.v(121[16:24])
    defparam unary_minus_16_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 LessThan_14_i19_2_lut (.I0(current[9]), .I1(current_limit[9]), 
            .I2(GND_net), .I3(GND_net), .O(n19));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam LessThan_14_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 encoder0_position_30__I_0_add_1771_24_lut (.I0(GND_net), .I1(n2612), 
            .I2(VCC_net), .I3(n51789), .O(n2679)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1771_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_inv_0_i6_1_lut (.I0(current[5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n20_adj_5714));   // verilog/TinyFPGA_B.v(121[16:24])
    defparam unary_minus_16_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_add_2039_12_lut (.I0(GND_net), .I1(n3024), 
            .I2(VCC_net), .I3(n51879), .O(n3091)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2039_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_14_i17_2_lut (.I0(current[8]), .I1(current_limit[8]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_5697));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam LessThan_14_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_14_i7_2_lut (.I0(current[3]), .I1(current_limit[3]), 
            .I2(GND_net), .I3(GND_net), .O(n7_adj_5704));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam LessThan_14_i7_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_14_i9_2_lut (.I0(current[4]), .I1(current_limit[4]), 
            .I2(GND_net), .I3(GND_net), .O(n9_adj_5702));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam LessThan_14_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_2452_4_lut (.I0(GND_net), .I1(n405), .I2(GND_net), .I3(n51281), 
            .O(n7445)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2452_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2039_12 (.CI(n51879), .I0(n3024), 
            .I1(VCC_net), .CO(n51880));
    SB_CARRY encoder0_position_30__I_0_add_1771_24 (.CI(n51789), .I0(n2612), 
            .I1(VCC_net), .CO(n51790));
    SB_LUT4 encoder0_position_30__I_0_add_1302_11_lut (.I0(GND_net), .I1(n1925), 
            .I2(VCC_net), .I3(n51519), .O(n1992)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1302_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2452_4 (.CI(n51281), .I0(n405), .I1(GND_net), .CO(n51282));
    SB_LUT4 encoder0_position_30__I_0_add_2039_11_lut (.I0(GND_net), .I1(n3025), 
            .I2(VCC_net), .I3(n51878), .O(n3092)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2039_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1302_11 (.CI(n51519), .I0(n1925), 
            .I1(VCC_net), .CO(n51520));
    SB_CARRY encoder0_position_30__I_0_add_2039_11 (.CI(n51878), .I0(n3025), 
            .I1(VCC_net), .CO(n51879));
    SB_LUT4 encoder0_position_30__I_0_add_1771_23_lut (.I0(GND_net), .I1(n2613), 
            .I2(VCC_net), .I3(n51788), .O(n2680)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1771_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1771_23 (.CI(n51788), .I0(n2613), 
            .I1(VCC_net), .CO(n51789));
    SB_LUT4 encoder0_position_30__I_0_add_2039_10_lut (.I0(GND_net), .I1(n3026), 
            .I2(VCC_net), .I3(n51877), .O(n3093)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2039_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2039_10 (.CI(n51877), .I0(n3026), 
            .I1(VCC_net), .CO(n51878));
    SB_LUT4 encoder0_position_30__I_0_add_1771_22_lut (.I0(GND_net), .I1(n2614), 
            .I2(VCC_net), .I3(n51787), .O(n2681)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1771_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1302_10_lut (.I0(GND_net), .I1(n1926), 
            .I2(VCC_net), .I3(n51518), .O(n1993)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1302_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1302_10 (.CI(n51518), .I0(n1926), 
            .I1(VCC_net), .CO(n51519));
    SB_LUT4 encoder0_position_30__I_0_add_1570_9_lut (.I0(GND_net), .I1(n2327), 
            .I2(VCC_net), .I3(n51708), .O(n2394)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1570_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_2039_9_lut (.I0(GND_net), .I1(n3027), 
            .I2(VCC_net), .I3(n51876), .O(n3094)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2039_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1771_22 (.CI(n51787), .I0(n2614), 
            .I1(VCC_net), .CO(n51788));
    SB_CARRY encoder0_position_30__I_0_add_2039_9 (.CI(n51876), .I0(n3027), 
            .I1(VCC_net), .CO(n51877));
    SB_LUT4 unary_minus_16_inv_0_i7_1_lut (.I0(current[6]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_5713));   // verilog/TinyFPGA_B.v(121[16:24])
    defparam unary_minus_16_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_inv_0_i13_1_lut (.I0(encoder0_position[11]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n21_adj_5911));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_unary_minus_2_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i54610_1_lut (.I0(n2841), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n70304));
    defparam i54610_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 LessThan_14_i11_2_lut (.I0(current[5]), .I1(current_limit[5]), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_5701));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam LessThan_14_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_14_i5_2_lut (.I0(current[2]), .I1(current_limit[2]), 
            .I2(GND_net), .I3(GND_net), .O(n5_adj_5706));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam LessThan_14_i5_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i52205_4_lut (.I0(n11_adj_5701), .I1(n9_adj_5702), .I2(n7_adj_5704), 
            .I3(n5_adj_5706), .O(n67899));
    defparam i52205_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 encoder0_position_30__I_0_add_1302_9_lut (.I0(GND_net), .I1(n1927), 
            .I2(VCC_net), .I3(n51517), .O(n1994)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1302_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_2039_8_lut (.I0(GND_net), .I1(n3028), 
            .I2(VCC_net), .I3(n51875), .O(n3095)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2039_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1570_9 (.CI(n51708), .I0(n2327), 
            .I1(VCC_net), .CO(n51709));
    SB_LUT4 LessThan_14_i16_3_lut (.I0(n8_adj_5703), .I1(current_limit[9]), 
            .I2(n19), .I3(GND_net), .O(n16_adj_5698));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam LessThan_14_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_14_i4_4_lut (.I0(current_limit[0]), .I1(current_limit[1]), 
            .I2(current[1]), .I3(current[0]), .O(n4_adj_5707));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam LessThan_14_i4_4_lut.LUT_INIT = 16'h0c8e;
    SB_LUT4 i53748_3_lut (.I0(n4_adj_5707), .I1(current_limit[5]), .I2(n11_adj_5701), 
            .I3(GND_net), .O(n69442));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam i53748_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_30__I_0_add_1302_9 (.CI(n51517), .I0(n1927), 
            .I1(VCC_net), .CO(n51518));
    SB_LUT4 i53749_3_lut (.I0(n69442), .I1(current_limit[6]), .I2(n13_adj_5700), 
            .I3(GND_net), .O(n69443));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam i53749_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_16_inv_0_i8_1_lut (.I0(current[7]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n18));   // verilog/TinyFPGA_B.v(121[16:24])
    defparam unary_minus_16_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i52185_4_lut (.I0(n17_adj_5697), .I1(n15_adj_5699), .I2(n13_adj_5700), 
            .I3(n67899), .O(n67879));
    defparam i52185_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 unary_minus_16_inv_0_i9_1_lut (.I0(current[8]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_5712));   // verilog/TinyFPGA_B.v(121[16:24])
    defparam unary_minus_16_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_4297_i22_3_lut (.I0(encoder0_position[21]), .I1(n11_adj_5740), 
            .I2(encoder0_position[30]), .I3(GND_net), .O(n522));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam mux_4297_i22_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i54066_4_lut (.I0(n16_adj_5698), .I1(n6_adj_5705), .I2(n19), 
            .I3(n67852), .O(n69760));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam i54066_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i52500_3_lut (.I0(n69443), .I1(current_limit[7]), .I2(n15_adj_5699), 
            .I3(GND_net), .O(n68194));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam i52500_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_30__I_0_add_2039_8 (.CI(n51875), .I0(n3028), 
            .I1(VCC_net), .CO(n51876));
    SB_LUT4 encoder0_position_30__I_0_add_2039_7_lut (.I0(GND_net), .I1(n3029), 
            .I2(GND_net), .I3(n51874), .O(n3096)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2039_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i54242_4_lut (.I0(n68194), .I1(n69760), .I2(n19), .I3(n67879), 
            .O(n69936));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam i54242_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i54243_3_lut (.I0(n69936), .I1(current_limit[10]), .I2(current[10]), 
            .I3(GND_net), .O(n69937));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam i54243_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 mux_4297_i12_3_lut (.I0(encoder0_position[11]), .I1(n21_adj_5727), 
            .I2(encoder0_position[30]), .I3(GND_net), .O(n946));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam mux_4297_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_i1921_3_lut (.I0(n2822), .I1(n2889), 
            .I2(n2841), .I3(GND_net), .O(n2921));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1921_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_add_1771_21_lut (.I0(GND_net), .I1(n2615), 
            .I2(VCC_net), .I3(n51786), .O(n2682)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1771_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_i1457_3_lut (.I0(n946), .I1(n2201), 
            .I2(n2148), .I3(GND_net), .O(n2233));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1457_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i54168_3_lut (.I0(n69937), .I1(current_limit[11]), .I2(current[11]), 
            .I3(GND_net), .O(n24));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam i54168_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 encoder0_position_30__I_0_add_1570_8_lut (.I0(GND_net), .I1(n2328), 
            .I2(VCC_net), .I3(n51707), .O(n2395)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1570_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1771_21 (.CI(n51786), .I0(n2615), 
            .I1(VCC_net), .CO(n51787));
    SB_LUT4 i1_4_lut_adj_1796 (.I0(current_limit[13]), .I1(n24), .I2(current_limit[14]), 
            .I3(current_limit[12]), .O(n61064));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam i1_4_lut_adj_1796.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1797 (.I0(current_limit[13]), .I1(n24), .I2(current_limit[14]), 
            .I3(current_limit[12]), .O(n61067));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam i1_4_lut_adj_1797.LUT_INIT = 16'h8000;
    SB_CARRY encoder0_position_30__I_0_add_2039_7 (.CI(n51874), .I0(n3029), 
            .I1(GND_net), .CO(n51875));
    SB_LUT4 i1_4_lut_adj_1798 (.I0(current[15]), .I1(current_limit[15]), 
            .I2(n61067), .I3(n61064), .O(n260));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam i1_4_lut_adj_1798.LUT_INIT = 16'hb3a2;
    SB_LUT4 encoder0_position_30__I_0_i1524_3_lut (.I0(n2233), .I1(n2300), 
            .I2(n2247), .I3(GND_net), .O(n2332));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1524_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1591_3_lut (.I0(n2332), .I1(n2399), 
            .I2(n2346), .I3(GND_net), .O(n2431));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1591_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 LessThan_17_i15_2_lut (.I0(duty[7]), .I1(n303), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_5693));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam LessThan_17_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_2452_3_lut (.I0(GND_net), .I1(n625), .I2(VCC_net), .I3(n51280), 
            .O(n7446)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2452_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_2039_6_lut (.I0(GND_net), .I1(n3030), 
            .I2(GND_net), .I3(n51873), .O(n3097)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2039_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_i1658_3_lut (.I0(n2431), .I1(n2498), 
            .I2(n2445), .I3(GND_net), .O(n2530));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1658_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_30__I_0_add_2039_6 (.CI(n51873), .I0(n3030), 
            .I1(GND_net), .CO(n51874));
    SB_CARRY encoder0_position_30__I_0_add_1570_8 (.CI(n51707), .I0(n2328), 
            .I1(VCC_net), .CO(n51708));
    SB_LUT4 LessThan_17_i13_2_lut (.I0(duty[6]), .I1(n304), .I2(GND_net), 
            .I3(GND_net), .O(n13));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam LessThan_17_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 encoder0_position_30__I_0_i1725_3_lut (.I0(n2530), .I1(n2597), 
            .I2(n2544), .I3(GND_net), .O(n2629));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1725_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_add_1302_8_lut (.I0(GND_net), .I1(n1928), 
            .I2(VCC_net), .I3(n51516), .O(n1995)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1302_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_i1792_3_lut (.I0(n2629), .I1(n2696), 
            .I2(n2643), .I3(GND_net), .O(n2728));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1792_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_add_1570_7_lut (.I0(GND_net), .I1(n2329), 
            .I2(GND_net), .I3(n51706), .O(n2396)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1570_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_17_i17_2_lut (.I0(duty[8]), .I1(n302), .I2(GND_net), 
            .I3(GND_net), .O(n17));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam LessThan_17_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_17_i19_2_lut (.I0(duty[9]), .I1(n301), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_5708));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam LessThan_17_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_17_i7_2_lut (.I0(duty[3]), .I1(n307), .I2(GND_net), 
            .I3(GND_net), .O(n7_adj_5694));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam LessThan_17_i7_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_2452_3 (.CI(n51280), .I0(n625), .I1(VCC_net), .CO(n51281));
    SB_CARRY encoder0_position_30__I_0_add_1570_7 (.CI(n51706), .I0(n2329), 
            .I1(GND_net), .CO(n51707));
    SB_CARRY encoder0_position_30__I_0_add_1302_8 (.CI(n51516), .I0(n1928), 
            .I1(VCC_net), .CO(n51517));
    SB_LUT4 LessThan_17_i9_2_lut (.I0(duty[4]), .I1(n306), .I2(GND_net), 
            .I3(GND_net), .O(n9));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam LessThan_17_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 encoder0_position_30__I_0_add_1771_20_lut (.I0(GND_net), .I1(n2616), 
            .I2(VCC_net), .I3(n51785), .O(n2683)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1771_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1302_7_lut (.I0(GND_net), .I1(n1929), 
            .I2(GND_net), .I3(n51515), .O(n1996)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1302_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1570_6_lut (.I0(GND_net), .I1(n2330), 
            .I2(GND_net), .I3(n51705), .O(n2397)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1570_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_17_i11_2_lut (.I0(duty[5]), .I1(n305), .I2(GND_net), 
            .I3(GND_net), .O(n11));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam LessThan_17_i11_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY encoder0_position_30__I_0_add_1570_6 (.CI(n51705), .I0(n2330), 
            .I1(GND_net), .CO(n51706));
    SB_LUT4 LessThan_17_i5_2_lut (.I0(duty[2]), .I1(n308), .I2(GND_net), 
            .I3(GND_net), .O(n5));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam LessThan_17_i5_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY encoder0_position_30__I_0_add_1302_7 (.CI(n51515), .I0(n1929), 
            .I1(GND_net), .CO(n51516));
    SB_LUT4 encoder0_position_30__I_0_add_1302_6_lut (.I0(GND_net), .I1(n1930), 
            .I2(GND_net), .I3(n51514), .O(n1997)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1302_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i52128_4_lut (.I0(n11), .I1(n9), .I2(n7_adj_5694), .I3(n5), 
            .O(n67822));
    defparam i52128_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 LessThan_17_i8_3_lut (.I0(n306), .I1(n302), .I2(n17), .I3(GND_net), 
            .O(n8));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam LessThan_17_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_17_i6_3_lut (.I0(n308), .I1(n307), .I2(n7_adj_5694), 
            .I3(GND_net), .O(n6_adj_5695));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam LessThan_17_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_30__I_0_add_1771_20 (.CI(n51785), .I0(n2616), 
            .I1(VCC_net), .CO(n51786));
    SB_CARRY encoder0_position_30__I_0_add_1302_6 (.CI(n51514), .I0(n1930), 
            .I1(GND_net), .CO(n51515));
    SB_LUT4 encoder0_position_30__I_0_add_1771_19_lut (.I0(GND_net), .I1(n2617), 
            .I2(VCC_net), .I3(n51784), .O(n2684)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1771_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_2039_5_lut (.I0(GND_net), .I1(n3031), 
            .I2(VCC_net), .I3(n51872), .O(n3098)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2039_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2039_5 (.CI(n51872), .I0(n3031), 
            .I1(VCC_net), .CO(n51873));
    SB_CARRY encoder0_position_30__I_0_add_1771_19 (.CI(n51784), .I0(n2617), 
            .I1(VCC_net), .CO(n51785));
    SB_LUT4 encoder0_position_30__I_0_add_2039_4_lut (.I0(GND_net), .I1(n3032), 
            .I2(GND_net), .I3(n51871), .O(n3099)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2039_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_17_i16_3_lut (.I0(n8), .I1(n301), .I2(n19_adj_5708), 
            .I3(GND_net), .O(n16));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam LessThan_17_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_30__I_0_add_2039_4 (.CI(n51871), .I0(n3032), 
            .I1(GND_net), .CO(n51872));
    SB_LUT4 add_151_33_lut (.I0(GND_net), .I1(delay_counter[31]), .I2(GND_net), 
            .I3(n51008), .O(n1208)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_33_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1771_18_lut (.I0(GND_net), .I1(n2618), 
            .I2(VCC_net), .I3(n51783), .O(n2685)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1771_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i2_3_lut_adj_1799 (.I0(duty[15]), .I1(duty[20]), .I2(n294), 
            .I3(GND_net), .O(n12_adj_5842));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam i2_3_lut_adj_1799.LUT_INIT = 16'h7e7e;
    SB_LUT4 i6_4_lut (.I0(duty[13]), .I1(n12_adj_5842), .I2(duty[21]), 
            .I3(n294), .O(n16_adj_5840));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam i6_4_lut.LUT_INIT = 16'hdffe;
    SB_LUT4 i4_3_lut (.I0(duty[19]), .I1(duty[16]), .I2(n294), .I3(GND_net), 
            .O(n14_adj_5841));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam i4_3_lut.LUT_INIT = 16'h7e7e;
    SB_LUT4 encoder0_position_30__I_0_add_2039_3_lut (.I0(GND_net), .I1(n3033), 
            .I2(VCC_net), .I3(n51870), .O(n3100)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2039_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_17_i10_3_lut (.I0(n305), .I1(n304), .I2(n13), .I3(GND_net), 
            .O(n10));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam LessThan_17_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_17_i4_3_lut (.I0(n66963), .I1(n309), .I2(duty[1]), 
            .I3(GND_net), .O(n4_adj_5696));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam LessThan_17_i4_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 LessThan_17_i12_3_lut (.I0(n10), .I1(n303), .I2(n15_adj_5693), 
            .I3(GND_net), .O(n12));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam LessThan_17_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52116_4_lut (.I0(n17), .I1(n15_adj_5693), .I2(n13), .I3(n67822), 
            .O(n67810));
    defparam i52116_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 add_2452_2_lut (.I0(GND_net), .I1(n518), .I2(GND_net), .I3(VCC_net), 
            .O(n7447)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2452_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1771_18 (.CI(n51783), .I0(n2618), 
            .I1(VCC_net), .CO(n51784));
    SB_LUT4 i54068_4_lut (.I0(n16), .I1(n6_adj_5695), .I2(n19_adj_5708), 
            .I3(n67804), .O(n69762));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam i54068_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 encoder0_position_30__I_0_add_1570_5_lut (.I0(GND_net), .I1(n2331), 
            .I2(VCC_net), .I3(n51704), .O(n2398)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1570_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2039_3 (.CI(n51870), .I0(n3033), 
            .I1(VCC_net), .CO(n51871));
    SB_LUT4 encoder0_position_30__I_0_add_1302_5_lut (.I0(GND_net), .I1(n1931), 
            .I2(VCC_net), .I3(n51513), .O(n1998)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1302_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1302_5 (.CI(n51513), .I0(n1931), 
            .I1(VCC_net), .CO(n51514));
    SB_LUT4 add_151_32_lut (.I0(GND_net), .I1(delay_counter[30]), .I2(GND_net), 
            .I3(n51007), .O(n1209)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_32_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1771_17_lut (.I0(GND_net), .I1(n2619), 
            .I2(VCC_net), .I3(n51782), .O(n2686)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1771_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1771_17 (.CI(n51782), .I0(n2619), 
            .I1(VCC_net), .CO(n51783));
    SB_LUT4 encoder0_position_30__I_0_add_1302_4_lut (.I0(GND_net), .I1(n1932), 
            .I2(GND_net), .I3(n51512), .O(n1999)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1302_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i53212_4_lut (.I0(n12), .I1(n4_adj_5696), .I2(n15_adj_5693), 
            .I3(n67816), .O(n68906));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam i53212_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 encoder0_position_30__I_0_add_2039_2_lut (.I0(GND_net), .I1(n955), 
            .I2(GND_net), .I3(VCC_net), .O(n3101)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2039_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i54247_4_lut (.I0(n68906), .I1(n69762), .I2(n19_adj_5708), 
            .I3(n67810), .O(n69941));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam i54247_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i54248_3_lut (.I0(n69941), .I1(n300), .I2(duty[10]), .I3(GND_net), 
            .O(n69942));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam i54248_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i54154_3_lut (.I0(n69942), .I1(n299), .I2(duty[11]), .I3(GND_net), 
            .O(n69848));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam i54154_3_lut.LUT_INIT = 16'h8e8e;
    SB_CARRY encoder0_position_30__I_0_add_1302_4 (.CI(n51512), .I0(n1932), 
            .I1(GND_net), .CO(n51513));
    SB_CARRY add_2452_2 (.CI(VCC_net), .I0(n518), .I1(GND_net), .CO(n51280));
    SB_IO CS_CLK_pad (.PACKAGE_PIN(CS_CLK), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(CS_CLK_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam CS_CLK_pad.PIN_TYPE = 6'b011001;
    defparam CS_CLK_pad.PULLUP = 1'b0;
    defparam CS_CLK_pad.NEG_TRIGGER = 1'b0;
    defparam CS_CLK_pad.IO_STANDARD = "SB_LVCMOS";
    SB_CARRY add_151_13 (.CI(n50988), .I0(delay_counter[11]), .I1(GND_net), 
            .CO(n50989));
    SB_LUT4 n11566_bdd_4_lut_55397 (.I0(n11566), .I1(current[15]), .I2(duty[16]), 
            .I3(n11564), .O(n71132));
    defparam n11566_bdd_4_lut_55397.LUT_INIT = 16'he4aa;
    SB_LUT4 n71132_bdd_4_lut (.I0(n71132), .I1(duty[13]), .I2(n4913), 
            .I3(n11564), .O(pwm_setpoint_23__N_3[13]));
    defparam n71132_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 encoder0_position_30__I_0_i1923_3_lut (.I0(n2824), .I1(n2891), 
            .I2(n2841), .I3(GND_net), .O(n2923));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1923_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 n11566_bdd_4_lut_55387 (.I0(n11566), .I1(current[15]), .I2(duty[15]), 
            .I3(n11564), .O(n71126));
    defparam n11566_bdd_4_lut_55387.LUT_INIT = 16'he4aa;
    SB_LUT4 n71126_bdd_4_lut (.I0(n71126), .I1(duty[12]), .I2(n4914), 
            .I3(n11564), .O(pwm_setpoint_23__N_3[12]));
    defparam n71126_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 encoder0_position_30__I_0_i1912_3_lut (.I0(n2813), .I1(n2880), 
            .I2(n2841), .I3(GND_net), .O(n2912));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1912_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 n11566_bdd_4_lut_55382 (.I0(n11566), .I1(current[11]), .I2(duty[14]), 
            .I3(n11564), .O(n71120));
    defparam n11566_bdd_4_lut_55382.LUT_INIT = 16'he4aa;
    SB_LUT4 n71120_bdd_4_lut (.I0(n71120), .I1(duty[11]), .I2(n4915), 
            .I3(n11564), .O(pwm_setpoint_23__N_3[11]));
    defparam n71120_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 encoder0_position_30__I_0_i1914_3_lut (.I0(n2815), .I1(n2882), 
            .I2(n2841), .I3(GND_net), .O(n2914));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1914_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 n11566_bdd_4_lut_55377 (.I0(n11566), .I1(current[10]), .I2(duty[13]), 
            .I3(n11564), .O(n71114));
    defparam n11566_bdd_4_lut_55377.LUT_INIT = 16'he4aa;
    SB_LUT4 n71114_bdd_4_lut (.I0(n71114), .I1(duty[10]), .I2(n4916), 
            .I3(n11564), .O(pwm_setpoint_23__N_3[10]));
    defparam n71114_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 encoder0_position_30__I_0_i1508_3_lut (.I0(n2217_adj_5853), .I1(n2284), 
            .I2(n2247), .I3(GND_net), .O(n2316));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1508_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 n11566_bdd_4_lut_55372 (.I0(n11566), .I1(current[9]), .I2(duty[12]), 
            .I3(n11564), .O(n71108));
    defparam n11566_bdd_4_lut_55372.LUT_INIT = 16'he4aa;
    SB_LUT4 n71108_bdd_4_lut (.I0(n71108), .I1(duty[9]), .I2(n4917), .I3(n11564), 
            .O(pwm_setpoint_23__N_3[9]));
    defparam n71108_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 encoder0_position_30__I_0_i1575_3_lut (.I0(n2316), .I1(n2383), 
            .I2(n2346), .I3(GND_net), .O(n2415));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1575_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 n11566_bdd_4_lut_55367 (.I0(n11566), .I1(current[8]), .I2(duty[11]), 
            .I3(n11564), .O(n71102));
    defparam n11566_bdd_4_lut_55367.LUT_INIT = 16'he4aa;
    SB_LUT4 n71102_bdd_4_lut (.I0(n71102), .I1(duty[8]), .I2(n4918), .I3(n11564), 
            .O(pwm_setpoint_23__N_3[8]));
    defparam n71102_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 encoder0_position_30__I_0_i1642_3_lut (.I0(n2415), .I1(n2482), 
            .I2(n2445), .I3(GND_net), .O(n2514));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1642_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 n11566_bdd_4_lut_55362 (.I0(n11566), .I1(current[7]), .I2(duty[10]), 
            .I3(n11564), .O(n71096));
    defparam n11566_bdd_4_lut_55362.LUT_INIT = 16'he4aa;
    SB_LUT4 n71096_bdd_4_lut (.I0(n71096), .I1(duty[7]), .I2(n4919), .I3(n11564), 
            .O(pwm_setpoint_23__N_3[7]));
    defparam n71096_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 encoder0_position_30__I_0_i1709_3_lut (.I0(n2514), .I1(n2581), 
            .I2(n2544), .I3(GND_net), .O(n2613));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1709_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 n11566_bdd_4_lut_55357 (.I0(n11566), .I1(current[6]), .I2(duty[9]), 
            .I3(n11564), .O(n71090));
    defparam n11566_bdd_4_lut_55357.LUT_INIT = 16'he4aa;
    SB_LUT4 n71090_bdd_4_lut (.I0(n71090), .I1(duty[6]), .I2(n4920), .I3(n11564), 
            .O(pwm_setpoint_23__N_3[6]));
    defparam n71090_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 encoder0_position_30__I_0_i1776_3_lut (.I0(n2613), .I1(n2680), 
            .I2(n2643), .I3(GND_net), .O(n2712));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1776_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_add_1302_3_lut (.I0(GND_net), .I1(n1933), 
            .I2(VCC_net), .I3(n51511), .O(n2000)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1302_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_151_32 (.CI(n51007), .I0(delay_counter[30]), .I1(GND_net), 
            .CO(n51008));
    SB_LUT4 encoder0_position_30__I_0_add_1771_16_lut (.I0(GND_net), .I1(n2620), 
            .I2(VCC_net), .I3(n51781), .O(n2687)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1771_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i8_4_lut (.I0(duty[14]), .I1(n16_adj_5840), .I2(duty[18]), 
            .I3(n294), .O(n18_adj_5838));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam i8_4_lut.LUT_INIT = 16'hdffe;
    SB_CARRY encoder0_position_30__I_0_add_1570_5 (.CI(n51704), .I0(n2331), 
            .I1(VCC_net), .CO(n51705));
    SB_LUT4 add_151_12_lut (.I0(GND_net), .I1(delay_counter[10]), .I2(GND_net), 
            .I3(n50987), .O(n1229)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1570_4_lut (.I0(GND_net), .I1(n2332), 
            .I2(GND_net), .I3(n51703), .O(n2399)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1570_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2039_2 (.CI(VCC_net), .I0(n955), 
            .I1(GND_net), .CO(n51870));
    SB_LUT4 add_151_31_lut (.I0(GND_net), .I1(delay_counter[29]), .I2(GND_net), 
            .I3(n51006), .O(n1210)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_31_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i7_4_lut (.I0(duty[22]), .I1(n14_adj_5841), .I2(duty[17]), 
            .I3(n294), .O(n17_adj_5839));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam i7_4_lut.LUT_INIT = 16'hdffe;
    SB_LUT4 i53537_3_lut (.I0(n69848), .I1(n298), .I2(duty[12]), .I3(GND_net), 
            .O(n69231));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam i53537_3_lut.LUT_INIT = 16'h8e8e;
    SB_CARRY encoder0_position_30__I_0_add_1302_3 (.CI(n51511), .I0(n1933), 
            .I1(VCC_net), .CO(n51512));
    SB_LUT4 i53538_4_lut (.I0(n69231), .I1(n294), .I2(n17_adj_5839), .I3(n18_adj_5838), 
            .O(n69232));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam i53538_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 encoder0_position_30__I_0_add_1302_2_lut (.I0(GND_net), .I1(n944), 
            .I2(GND_net), .I3(VCC_net), .O(n2001)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1302_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i44113_4_lut (.I0(n260), .I1(duty[23]), .I2(n294), .I3(n69232), 
            .O(n11564));
    defparam i44113_4_lut.LUT_INIT = 16'h1151;
    SB_CARRY add_151_5 (.CI(n50980), .I0(delay_counter[3]), .I1(GND_net), 
            .CO(n50981));
    SB_CARRY add_151_12 (.CI(n50987), .I0(delay_counter[10]), .I1(GND_net), 
            .CO(n50988));
    SB_CARRY encoder0_position_30__I_0_add_1302_2 (.CI(VCC_net), .I0(n944), 
            .I1(GND_net), .CO(n51511));
    SB_CARRY encoder0_position_30__I_0_add_1771_16 (.CI(n51781), .I0(n2620), 
            .I1(VCC_net), .CO(n51782));
    SB_LUT4 encoder0_position_30__I_0_add_1972_29_lut (.I0(n70273), .I1(n2907), 
            .I2(VCC_net), .I3(n51869), .O(n3006)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1972_29_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i52936_3_lut (.I0(n15_adj_5746), .I1(n13_adj_5747), .I2(n11_adj_5748), 
            .I3(GND_net), .O(n68630));
    defparam i52936_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i52896_4_lut (.I0(current[15]), .I1(duty[13]), .I2(duty[14]), 
            .I3(n68630), .O(n68590));
    defparam i52896_4_lut.LUT_INIT = 16'h7eff;
    SB_LUT4 encoder0_position_30__I_0_add_1972_28_lut (.I0(GND_net), .I1(n2908), 
            .I2(VCC_net), .I3(n51868), .O(n2975)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1972_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_151_31 (.CI(n51006), .I0(delay_counter[29]), .I1(GND_net), 
            .CO(n51007));
    SB_LUT4 add_151_4_lut (.I0(GND_net), .I1(delay_counter[2]), .I2(GND_net), 
            .I3(n50979), .O(n1237)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_151_30_lut (.I0(GND_net), .I1(delay_counter[28]), .I2(GND_net), 
            .I3(n51005), .O(n1211)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_30_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_151_11_lut (.I0(GND_net), .I1(delay_counter[9]), .I2(GND_net), 
            .I3(n50986), .O(n1230)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1771_15_lut (.I0(GND_net), .I1(n2621), 
            .I2(VCC_net), .I3(n51780), .O(n2688)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1771_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i2_3_lut_adj_1800 (.I0(n26376), .I1(n36), .I2(\data_out_frame[10] [7]), 
            .I3(GND_net), .O(n58845));   // verilog/coms.v(100[12:26])
    defparam i2_3_lut_adj_1800.LUT_INIT = 16'h9696;
    SB_LUT4 i52027_4_lut (.I0(n21_adj_5742), .I1(n19_adj_5743), .I2(n17_adj_5744), 
            .I3(n9_adj_5750), .O(n67721));
    defparam i52027_4_lut.LUT_INIT = 16'haaab;
    SB_CARRY add_151_30 (.CI(n51005), .I0(delay_counter[28]), .I1(GND_net), 
            .CO(n51006));
    SB_LUT4 add_151_29_lut (.I0(GND_net), .I1(delay_counter[27]), .I2(GND_net), 
            .I3(n51004), .O(n1212)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_29_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_inv_0_i10_1_lut (.I0(current[9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n16_adj_5711));   // verilog/TinyFPGA_B.v(121[16:24])
    defparam unary_minus_16_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 n11566_bdd_4_lut_55352 (.I0(n11566), .I1(current[5]), .I2(duty[8]), 
            .I3(n11564), .O(n71084));
    defparam n11566_bdd_4_lut_55352.LUT_INIT = 16'he4aa;
    SB_LUT4 i52970_4_lut (.I0(n9_adj_5750), .I1(n7_adj_5752), .I2(current[2]), 
            .I3(duty[2]), .O(n68664));
    defparam i52970_4_lut.LUT_INIT = 16'heffe;
    SB_LUT4 i54673_1_lut (.I0(n2742), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n70367));
    defparam i54673_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_151_29 (.CI(n51004), .I0(delay_counter[27]), .I1(GND_net), 
            .CO(n51005));
    SB_LUT4 i54733_1_lut (.I0(n2643), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n70427));
    defparam i54733_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i53411_4_lut (.I0(n15_adj_5746), .I1(n13_adj_5747), .I2(n11_adj_5748), 
            .I3(n68664), .O(n69105));
    defparam i53411_4_lut.LUT_INIT = 16'hfeff;
    SB_CARRY encoder0_position_30__I_0_add_1570_4 (.CI(n51703), .I0(n2332), 
            .I1(GND_net), .CO(n51704));
    SB_CARRY encoder0_position_30__I_0_add_1771_15 (.CI(n51780), .I0(n2621), 
            .I1(VCC_net), .CO(n51781));
    SB_LUT4 i5_4_lut (.I0(\data_out_frame[9] [1]), .I1(n58845), .I2(\data_out_frame[13] [3]), 
            .I3(n26143), .O(n12_adj_5925));   // verilog/coms.v(100[12:26])
    defparam i5_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i53403_4_lut (.I0(n21_adj_5742), .I1(n19_adj_5743), .I2(n17_adj_5744), 
            .I3(n69105), .O(n69097));
    defparam i53403_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i53996_4_lut (.I0(current[15]), .I1(n23_adj_5741), .I2(duty[12]), 
            .I3(n69097), .O(n69690));
    defparam i53996_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 i52902_4_lut (.I0(current[15]), .I1(duty[13]), .I2(duty[14]), 
            .I3(n69690), .O(n68596));
    defparam i52902_4_lut.LUT_INIT = 16'h7eff;
    SB_LUT4 LessThan_11_i4_4_lut (.I0(duty[0]), .I1(duty[1]), .I2(current[1]), 
            .I3(current[0]), .O(n4_adj_5754));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i4_4_lut.LUT_INIT = 16'h0c8e;
    SB_LUT4 i53742_3_lut (.I0(n4_adj_5754), .I1(duty[13]), .I2(current[15]), 
            .I3(GND_net), .O(n69436));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i53742_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 encoder0_position_30__I_0_add_1570_3_lut (.I0(GND_net), .I1(n2333), 
            .I2(VCC_net), .I3(n51702), .O(n2400)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1570_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i28911_2_lut (.I0(pwm_out), .I1(GHC), .I2(GND_net), .I3(GND_net), 
            .O(INHC_c_0));   // verilog/TinyFPGA_B.v(92[16:31])
    defparam i28911_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_inv_0_i14_1_lut (.I0(encoder0_position[12]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n20_adj_5910));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_unary_minus_2_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_4297_i13_3_lut (.I0(encoder0_position[12]), .I1(n20_adj_5728), 
            .I2(encoder0_position[30]), .I3(GND_net), .O(n945));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam mux_4297_i13_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_i1389_3_lut (.I0(n945), .I1(n2101), 
            .I2(n2049), .I3(GND_net), .O(n2133));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1389_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1456_3_lut (.I0(n2133), .I1(n2200), 
            .I2(n2148), .I3(GND_net), .O(n2232));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1456_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1523_3_lut (.I0(n2232), .I1(n2299), 
            .I2(n2247), .I3(GND_net), .O(n2331));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1523_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1590_3_lut (.I0(n2331), .I1(n2398), 
            .I2(n2346), .I3(GND_net), .O(n2430));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1590_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1657_3_lut (.I0(n2430), .I1(n2497), 
            .I2(n2445), .I3(GND_net), .O(n2529));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1657_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 n71084_bdd_4_lut (.I0(n71084), .I1(duty[5]), .I2(n4921), .I3(n11564), 
            .O(pwm_setpoint_23__N_3[5]));
    defparam n71084_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i6_4_lut_adj_1801 (.I0(\data_out_frame[11] [1]), .I1(n12_adj_5925), 
            .I2(n58887), .I3(\data_out_frame[11] [2]), .O(n26210));   // verilog/coms.v(100[12:26])
    defparam i6_4_lut_adj_1801.LUT_INIT = 16'h6996;
    SB_LUT4 i52882_4_lut (.I0(current[15]), .I1(duty[16]), .I2(duty[17]), 
            .I3(n15_adj_5746), .O(n68576));
    defparam i52882_4_lut.LUT_INIT = 16'hff7e;
    SB_LUT4 LessThan_11_i30_4_lut (.I0(duty[7]), .I1(duty[17]), .I2(current[15]), 
            .I3(duty[16]), .O(n30_adj_5736));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i30_4_lut.LUT_INIT = 16'h8f0e;
    SB_LUT4 i51997_4_lut (.I0(current[15]), .I1(duty[15]), .I2(duty[16]), 
            .I3(n68590), .O(n67691));
    defparam i51997_4_lut.LUT_INIT = 16'h5adb;
    SB_LUT4 LessThan_11_i35_rep_170_2_lut (.I0(current[15]), .I1(duty[17]), 
            .I2(GND_net), .I3(GND_net), .O(n71412));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i35_rep_170_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i54078_3_lut (.I0(n30_adj_5736), .I1(n10_adj_5749), .I2(n68576), 
            .I3(GND_net), .O(n69772));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i54078_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i52504_4_lut (.I0(n69436), .I1(duty[15]), .I2(current[15]), 
            .I3(duty[14]), .O(n68198));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i52504_4_lut.LUT_INIT = 16'h8f0e;
    SB_LUT4 i53740_3_lut (.I0(n6_adj_5753), .I1(duty[10]), .I2(n21_adj_5742), 
            .I3(GND_net), .O(n69434));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i53740_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53741_3_lut (.I0(n69434), .I1(duty[11]), .I2(n23_adj_5741), 
            .I3(GND_net), .O(n69435));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i53741_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_i1724_3_lut (.I0(n2529), .I1(n2596), 
            .I2(n2544), .I3(GND_net), .O(n2628));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1724_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_30__I_0_add_1972_28 (.CI(n51868), .I0(n2908), 
            .I1(VCC_net), .CO(n51869));
    SB_LUT4 i53397_4_lut (.I0(current[15]), .I1(n23_adj_5741), .I2(duty[12]), 
            .I3(n67721), .O(n69091));
    defparam i53397_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 encoder0_position_30__I_0_add_1771_14_lut (.I0(GND_net), .I1(n2622), 
            .I2(VCC_net), .I3(n51779), .O(n2689)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1771_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1570_3 (.CI(n51702), .I0(n2333), 
            .I1(VCC_net), .CO(n51703));
    SB_LUT4 encoder0_position_30__I_0_add_1972_27_lut (.I0(GND_net), .I1(n2909), 
            .I2(VCC_net), .I3(n51867), .O(n2976)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1972_27_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_151_28_lut (.I0(GND_net), .I1(delay_counter[26]), .I2(GND_net), 
            .I3(n51003), .O(n1213)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1972_27 (.CI(n51867), .I0(n2909), 
            .I1(VCC_net), .CO(n51868));
    SB_CARRY add_151_28 (.CI(n51003), .I0(delay_counter[26]), .I1(GND_net), 
            .CO(n51004));
    SB_CARRY encoder0_position_30__I_0_add_1771_14 (.CI(n51779), .I0(n2622), 
            .I1(VCC_net), .CO(n51780));
    SB_LUT4 add_151_27_lut (.I0(GND_net), .I1(delay_counter[25]), .I2(GND_net), 
            .I3(n51002), .O(n1214)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_151_27 (.CI(n51002), .I0(delay_counter[25]), .I1(GND_net), 
            .CO(n51003));
    SB_LUT4 LessThan_11_i16_3_lut (.I0(n8_adj_5751), .I1(duty[9]), .I2(n19_adj_5743), 
            .I3(GND_net), .O(n16_adj_5745));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2_3_lut_adj_1802 (.I0(\data_out_frame[18] [7]), .I1(n53515), 
            .I2(\data_out_frame[19] [1]), .I3(GND_net), .O(n59455));
    defparam i2_3_lut_adj_1802.LUT_INIT = 16'h9696;
    SB_LUT4 encoder0_position_30__I_0_add_1972_26_lut (.I0(GND_net), .I1(n2910), 
            .I2(VCC_net), .I3(n51866), .O(n2977)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1972_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1771_13_lut (.I0(GND_net), .I1(n2623), 
            .I2(VCC_net), .I3(n51778), .O(n2690)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1771_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1570_2_lut (.I0(GND_net), .I1(n948), 
            .I2(GND_net), .I3(VCC_net), .O(n2401)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1570_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_151_26_lut (.I0(GND_net), .I1(delay_counter[24]), .I2(GND_net), 
            .I3(n51001), .O(n1215)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_151_26 (.CI(n51001), .I0(delay_counter[24]), .I1(GND_net), 
            .CO(n51002));
    SB_CARRY encoder0_position_30__I_0_add_1570_2 (.CI(VCC_net), .I0(n948), 
            .I1(GND_net), .CO(n51702));
    SB_CARRY encoder0_position_30__I_0_add_1972_26 (.CI(n51866), .I0(n2910), 
            .I1(VCC_net), .CO(n51867));
    SB_LUT4 encoder0_position_30__I_0_i1576_3_lut (.I0(n2317), .I1(n2384), 
            .I2(n2346), .I3(GND_net), .O(n2416));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1576_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_30__I_0_add_1771_13 (.CI(n51778), .I0(n2623), 
            .I1(VCC_net), .CO(n51779));
    SB_LUT4 add_2502_25_lut (.I0(n70773), .I1(n2_adj_5892), .I2(n1059), 
            .I3(n51980), .O(encoder0_position_scaled_23__N_43[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2502_25_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 i52506_3_lut (.I0(n69435), .I1(duty[12]), .I2(current[15]), 
            .I3(GND_net), .O(n68200));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i52506_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 encoder0_position_30__I_0_add_1972_25_lut (.I0(GND_net), .I1(n2911), 
            .I2(VCC_net), .I3(n51865), .O(n2978)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1972_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1771_12_lut (.I0(GND_net), .I1(n2624), 
            .I2(VCC_net), .I3(n51777), .O(n2691)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1771_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1771_12 (.CI(n51777), .I0(n2624), 
            .I1(VCC_net), .CO(n51778));
    SB_CARRY encoder0_position_30__I_0_add_1972_25 (.CI(n51865), .I0(n2911), 
            .I1(VCC_net), .CO(n51866));
    SB_LUT4 encoder0_position_30__I_0_i1791_3_lut (.I0(n2628), .I1(n2695), 
            .I2(n2643), .I3(GND_net), .O(n2727));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1791_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i53760_4_lut (.I0(current[15]), .I1(duty[15]), .I2(duty[16]), 
            .I3(n68596), .O(n69454));
    defparam i53760_4_lut.LUT_INIT = 16'hff7e;
    SB_LUT4 encoder0_position_30__I_0_add_1034_15_lut (.I0(GND_net), .I1(n1521), 
            .I2(VCC_net), .I3(n51390), .O(n1588)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1034_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1771_11_lut (.I0(GND_net), .I1(n2625), 
            .I2(VCC_net), .I3(n51776), .O(n2692)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1771_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2502_24_lut (.I0(n70712), .I1(n2_adj_5892), .I2(n1158), 
            .I3(n51979), .O(encoder0_position_scaled_23__N_43[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2502_24_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 i15886_3_lut (.I0(\data_in_frame[5] [4]), .I1(rx_data[4]), .I2(n59656), 
            .I3(GND_net), .O(n29892));   // verilog/coms.v(130[12] 305[6])
    defparam i15886_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_add_1034_14_lut (.I0(GND_net), .I1(n1522), 
            .I2(VCC_net), .I3(n51389), .O(n1589)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1034_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1771_11 (.CI(n51776), .I0(n2625), 
            .I1(VCC_net), .CO(n51777));
    SB_CARRY encoder0_position_30__I_0_add_1034_14 (.CI(n51389), .I0(n1522), 
            .I1(VCC_net), .CO(n51390));
    SB_LUT4 encoder0_position_30__I_0_add_1034_13_lut (.I0(GND_net), .I1(n1523), 
            .I2(VCC_net), .I3(n51388), .O(n1590)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1034_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1771_10_lut (.I0(GND_net), .I1(n2626), 
            .I2(VCC_net), .I3(n51775), .O(n2693)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1771_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1972_24_lut (.I0(GND_net), .I1(n2912), 
            .I2(VCC_net), .I3(n51864), .O(n2979)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1972_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1972_24 (.CI(n51864), .I0(n2912), 
            .I1(VCC_net), .CO(n51865));
    SB_CARRY add_2502_24 (.CI(n51979), .I0(n2_adj_5892), .I1(n1158), .CO(n51980));
    SB_LUT4 add_2502_23_lut (.I0(n70727), .I1(n2_adj_5892), .I2(n1257), 
            .I3(n51978), .O(encoder0_position_scaled_23__N_43[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2502_23_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2502_23 (.CI(n51978), .I0(n2_adj_5892), .I1(n1257), .CO(n51979));
    SB_CARRY encoder0_position_30__I_0_add_1034_13 (.CI(n51388), .I0(n1523), 
            .I1(VCC_net), .CO(n51389));
    SB_LUT4 encoder0_position_30__I_0_add_1034_12_lut (.I0(GND_net), .I1(n1524), 
            .I2(VCC_net), .I3(n51387), .O(n1591)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1034_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_inv_0_i11_1_lut (.I0(current[10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_5710));   // verilog/TinyFPGA_B.v(121[16:24])
    defparam unary_minus_16_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_30__I_0_add_1034_12 (.CI(n51387), .I0(n1524), 
            .I1(VCC_net), .CO(n51388));
    SB_CARRY encoder0_position_30__I_0_add_1771_10 (.CI(n51775), .I0(n2626), 
            .I1(VCC_net), .CO(n51776));
    SB_LUT4 add_2502_22_lut (.I0(n70743), .I1(n2_adj_5892), .I2(n1356), 
            .I3(n51977), .O(encoder0_position_scaled_23__N_43[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2502_22_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 encoder0_position_30__I_0_add_1771_9_lut (.I0(GND_net), .I1(n2627), 
            .I2(VCC_net), .I3(n51774), .O(n2694)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1771_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1972_23_lut (.I0(GND_net), .I1(n2913), 
            .I2(VCC_net), .I3(n51863), .O(n2980)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1972_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_inv_0_i12_1_lut (.I0(current[11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n14));   // verilog/TinyFPGA_B.v(121[16:24])
    defparam unary_minus_16_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_2502_22 (.CI(n51977), .I0(n2_adj_5892), .I1(n1356), .CO(n51978));
    SB_CARRY encoder0_position_30__I_0_add_1972_23 (.CI(n51863), .I0(n2913), 
            .I1(VCC_net), .CO(n51864));
    SB_LUT4 add_2502_21_lut (.I0(n70760), .I1(n2_adj_5892), .I2(n1455), 
            .I3(n51976), .O(encoder0_position_scaled_23__N_43[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2502_21_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 encoder0_position_30__I_0_add_1034_11_lut (.I0(GND_net), .I1(n1525), 
            .I2(VCC_net), .I3(n51386), .O(n1592)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1034_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2502_21 (.CI(n51976), .I0(n2_adj_5892), .I1(n1455), .CO(n51977));
    SB_LUT4 encoder0_position_30__I_0_add_1972_22_lut (.I0(GND_net), .I1(n2914), 
            .I2(VCC_net), .I3(n51862), .O(n2981)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1972_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1034_11 (.CI(n51386), .I0(n1525), 
            .I1(VCC_net), .CO(n51387));
    SB_LUT4 encoder0_position_30__I_0_add_1034_10_lut (.I0(GND_net), .I1(n1526), 
            .I2(VCC_net), .I3(n51385), .O(n1593)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1034_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1034_10 (.CI(n51385), .I0(n1526), 
            .I1(VCC_net), .CO(n51386));
    SB_LUT4 encoder0_position_30__I_0_add_1034_9_lut (.I0(GND_net), .I1(n1527), 
            .I2(VCC_net), .I3(n51384), .O(n1594)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1034_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2502_20_lut (.I0(n70596), .I1(n2_adj_5892), .I2(n1554), 
            .I3(n51975), .O(encoder0_position_scaled_23__N_43[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2502_20_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY encoder0_position_30__I_0_add_1771_9 (.CI(n51774), .I0(n2627), 
            .I1(VCC_net), .CO(n51775));
    SB_CARRY add_2502_20 (.CI(n51975), .I0(n2_adj_5892), .I1(n1554), .CO(n51976));
    SB_LUT4 add_151_25_lut (.I0(GND_net), .I1(delay_counter[23]), .I2(GND_net), 
            .I3(n51000), .O(n1216)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i54254_4_lut (.I0(n68198), .I1(n69772), .I2(n71412), .I3(n67691), 
            .O(n69948));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i54254_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i53216_3_lut (.I0(n68200), .I1(n16_adj_5745), .I2(n69091), 
            .I3(GND_net), .O(n68910));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i53216_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i54304_4_lut (.I0(n68910), .I1(n69948), .I2(n71412), .I3(n69454), 
            .O(n69998));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i54304_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i54297_4_lut (.I0(n69998), .I1(duty[19]), .I2(current[15]), 
            .I3(duty[18]), .O(n69991));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i54297_4_lut.LUT_INIT = 16'h8f0e;
    SB_LUT4 i2_2_lut (.I0(duty[22]), .I1(current[15]), .I2(GND_net), .I3(GND_net), 
            .O(n6_adj_5760));
    defparam i2_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i53540_4_lut (.I0(n69991), .I1(duty[21]), .I2(current[15]), 
            .I3(duty[20]), .O(n69234));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i53540_4_lut.LUT_INIT = 16'h8f0e;
    SB_LUT4 i7_4_lut_adj_1803 (.I0(n69234), .I1(duty[23]), .I2(n6_adj_5760), 
            .I3(n260), .O(n11566));
    defparam i7_4_lut_adj_1803.LUT_INIT = 16'h3332;
    SB_LUT4 i14_4_lut_adj_1804 (.I0(n58418), .I1(\data_in_frame[4] [4]), 
            .I2(n164), .I3(rx_data[4]), .O(n57918));   // verilog/coms.v(130[12] 305[6])
    defparam i14_4_lut_adj_1804.LUT_INIT = 16'hcac0;
    SB_LUT4 encoder0_position_30__I_0_i1643_3_lut (.I0(n2416), .I1(n2483), 
            .I2(n2445), .I3(GND_net), .O(n2515));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1643_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14_4_lut_adj_1805 (.I0(n58418), .I1(\data_in_frame[4] [5]), 
            .I2(n164), .I3(rx_data[5]), .O(n57916));   // verilog/coms.v(130[12] 305[6])
    defparam i14_4_lut_adj_1805.LUT_INIT = 16'hcac0;
    SB_LUT4 i1_2_lut_adj_1806 (.I0(reset), .I1(n163), .I2(GND_net), .I3(GND_net), 
            .O(n164));
    defparam i1_2_lut_adj_1806.LUT_INIT = 16'heeee;
    SB_CARRY encoder0_position_30__I_0_add_1972_22 (.CI(n51862), .I0(n2914), 
            .I1(VCC_net), .CO(n51863));
    SB_LUT4 i54643_1_lut (.I0(n2445), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n70337));
    defparam i54643_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_add_1972_21_lut (.I0(GND_net), .I1(n2915), 
            .I2(VCC_net), .I3(n51861), .O(n2982)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1972_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_151_25 (.CI(n51000), .I0(delay_counter[23]), .I1(GND_net), 
            .CO(n51001));
    SB_CARRY encoder0_position_30__I_0_add_1972_21 (.CI(n51861), .I0(n2915), 
            .I1(VCC_net), .CO(n51862));
    SB_LUT4 add_2502_19_lut (.I0(n70615), .I1(n2_adj_5892), .I2(n1653), 
            .I3(n51974), .O(encoder0_position_scaled_23__N_43[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2502_19_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2502_19 (.CI(n51974), .I0(n2_adj_5892), .I1(n1653), .CO(n51975));
    SB_LUT4 i54860_1_lut (.I0(n2346), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n70554));
    defparam i54860_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_2502_18_lut (.I0(n70635), .I1(n2_adj_5892), .I2(n1752), 
            .I3(n51973), .O(encoder0_position_scaled_23__N_43[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2502_18_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 unary_minus_16_inv_0_i24_1_lut (.I0(current[15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n2));   // verilog/TinyFPGA_B.v(121[16:24])
    defparam unary_minus_16_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i54834_1_lut (.I0(n2247), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n70528));
    defparam i54834_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i14_4_lut_adj_1807 (.I0(n58418), .I1(\data_in_frame[4] [6]), 
            .I2(n164), .I3(rx_data[6]), .O(n57914));   // verilog/coms.v(130[12] 305[6])
    defparam i14_4_lut_adj_1807.LUT_INIT = 16'hcac0;
    SB_CARRY add_2502_18 (.CI(n51973), .I0(n2_adj_5892), .I1(n1752), .CO(n51974));
    SB_LUT4 i54809_1_lut (.I0(n2148), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n70503));
    defparam i54809_1_lut.LUT_INIT = 16'h5555;
    SB_IO CS_MISO_pad (.PACKAGE_PIN(CS_MISO), .OUTPUT_ENABLE(VCC_net), .D_IN_0(CS_MISO_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam CS_MISO_pad.PIN_TYPE = 6'b000001;
    defparam CS_MISO_pad.PULLUP = 1'b0;
    defparam CS_MISO_pad.NEG_TRIGGER = 1'b0;
    defparam CS_MISO_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 i54783_1_lut (.I0(n2049), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n70477));
    defparam i54783_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_add_1972_20_lut (.I0(GND_net), .I1(n2916), 
            .I2(VCC_net), .I3(n51860), .O(n2983)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1972_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1972_20 (.CI(n51860), .I0(n2916), 
            .I1(VCC_net), .CO(n51861));
    SB_LUT4 add_2502_17_lut (.I0(n70578), .I1(n2_adj_5892), .I2(n1851), 
            .I3(n51972), .O(encoder0_position_scaled_23__N_43[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2502_17_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY encoder0_position_30__I_0_add_1034_9 (.CI(n51384), .I0(n1527), 
            .I1(VCC_net), .CO(n51385));
    SB_LUT4 encoder0_position_30__I_0_add_1034_8_lut (.I0(GND_net), .I1(n1528), 
            .I2(VCC_net), .I3(n51383), .O(n1595)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1034_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1034_8 (.CI(n51383), .I0(n1528), 
            .I1(VCC_net), .CO(n51384));
    SB_LUT4 encoder0_position_30__I_0_add_1034_7_lut (.I0(GND_net), .I1(n1529), 
            .I2(GND_net), .I3(n51382), .O(n1596)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1034_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 n11566_bdd_4_lut_55347 (.I0(n11566), .I1(current[4]), .I2(duty[7]), 
            .I3(n11564), .O(n71072));
    defparam n11566_bdd_4_lut_55347.LUT_INIT = 16'he4aa;
    SB_CARRY add_2502_17 (.CI(n51972), .I0(n2_adj_5892), .I1(n1851), .CO(n51973));
    SB_LUT4 encoder0_position_30__I_0_add_1972_19_lut (.I0(GND_net), .I1(n2917), 
            .I2(VCC_net), .I3(n51859), .O(n2984)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1972_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1972_19 (.CI(n51859), .I0(n2917), 
            .I1(VCC_net), .CO(n51860));
    SB_LUT4 encoder0_position_30__I_0_add_1235_18_lut (.I0(GND_net), .I1(n1818), 
            .I2(VCC_net), .I3(n51493), .O(n1885)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1235_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1034_7 (.CI(n51382), .I0(n1529), 
            .I1(GND_net), .CO(n51383));
    SB_LUT4 add_2502_16_lut (.I0(n70454), .I1(n2_adj_5892), .I2(n1950), 
            .I3(n51971), .O(encoder0_position_scaled_23__N_43[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2502_16_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2502_16 (.CI(n51971), .I0(n2_adj_5892), .I1(n1950), .CO(n51972));
    SB_LUT4 encoder0_position_30__I_0_add_1771_8_lut (.I0(GND_net), .I1(n2628), 
            .I2(VCC_net), .I3(n51773), .O(n2695)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1771_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1034_6_lut (.I0(GND_net), .I1(n1530), 
            .I2(GND_net), .I3(n51381), .O(n1597)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1034_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_151_24_lut (.I0(GND_net), .I1(delay_counter[22]), .I2(GND_net), 
            .I3(n50999), .O(n1217)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i54760_1_lut (.I0(n1950), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n70454));
    defparam i54760_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_30__I_0_add_1771_8 (.CI(n51773), .I0(n2628), 
            .I1(VCC_net), .CO(n51774));
    SB_LUT4 i54884_1_lut (.I0(n1851), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n70578));
    defparam i54884_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i43885_3_lut (.I0(n6_adj_5775), .I1(n7446), .I2(n59507), .I3(GND_net), 
            .O(n59514));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam i43885_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_i1710_3_lut (.I0(n2515), .I1(n2582), 
            .I2(n2544), .I3(GND_net), .O(n2614));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1710_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_add_1771_7_lut (.I0(GND_net), .I1(n2629), 
            .I2(GND_net), .I3(n51772), .O(n2696)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1771_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2502_15_lut (.I0(n70477), .I1(n2_adj_5892), .I2(n2049), 
            .I3(n51970), .O(encoder0_position_scaled_23__N_43[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2502_15_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY encoder0_position_30__I_0_add_1771_7 (.CI(n51772), .I0(n2629), 
            .I1(GND_net), .CO(n51773));
    SB_LUT4 i43886_3_lut (.I0(encoder0_position[26]), .I1(n59514), .I2(encoder0_position[30]), 
            .I3(GND_net), .O(n832));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam i43886_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_add_1972_18_lut (.I0(GND_net), .I1(n2918), 
            .I2(VCC_net), .I3(n51858), .O(n2985)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1972_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1771_6_lut (.I0(GND_net), .I1(n2630), 
            .I2(GND_net), .I3(n51771), .O(n2697)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1771_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2502_15 (.CI(n51970), .I0(n2_adj_5892), .I1(n2049), .CO(n51971));
    SB_CARRY encoder0_position_30__I_0_add_1771_6 (.CI(n51771), .I0(n2630), 
            .I1(GND_net), .CO(n51772));
    SB_CARRY encoder0_position_30__I_0_add_1972_18 (.CI(n51858), .I0(n2918), 
            .I1(VCC_net), .CO(n51859));
    SB_LUT4 encoder0_position_30__I_0_add_1235_17_lut (.I0(GND_net), .I1(n1819), 
            .I2(VCC_net), .I3(n51492), .O(n1886)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1235_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_151_24 (.CI(n50999), .I0(delay_counter[22]), .I1(GND_net), 
            .CO(n51000));
    SB_CARRY encoder0_position_30__I_0_add_1034_6 (.CI(n51381), .I0(n1530), 
            .I1(GND_net), .CO(n51382));
    SB_CARRY encoder0_position_30__I_0_add_1235_17 (.CI(n51492), .I0(n1819), 
            .I1(VCC_net), .CO(n51493));
    SB_LUT4 add_151_23_lut (.I0(GND_net), .I1(delay_counter[21]), .I2(GND_net), 
            .I3(n50998), .O(n1218)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2502_14_lut (.I0(n70503), .I1(n2_adj_5892), .I2(n2148), 
            .I3(n51969), .O(encoder0_position_scaled_23__N_43[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2502_14_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2502_14 (.CI(n51969), .I0(n2_adj_5892), .I1(n2148), .CO(n51970));
    SB_LUT4 encoder0_position_30__I_0_add_1771_5_lut (.I0(GND_net), .I1(n2631), 
            .I2(VCC_net), .I3(n51770), .O(n2698)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1771_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1972_17_lut (.I0(GND_net), .I1(n2919), 
            .I2(VCC_net), .I3(n51857), .O(n2986)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1972_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_i1777_3_lut (.I0(n2614), .I1(n2681), 
            .I2(n2643), .I3(GND_net), .O(n2713));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1777_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1808 (.I0(commutation_state[2]), .I1(commutation_state[1]), 
            .I2(commutation_state_prev[2]), .I3(commutation_state_prev[1]), 
            .O(n4_adj_5845));   // verilog/TinyFPGA_B.v(146[7:48])
    defparam i1_4_lut_adj_1808.LUT_INIT = 16'h7bde;
    SB_LUT4 i15872_3_lut (.I0(\data_in_frame[5] [0]), .I1(rx_data[0]), .I2(n59656), 
            .I3(GND_net), .O(n29878));   // verilog/coms.v(130[12] 305[6])
    defparam i15872_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i2_3_lut_adj_1809 (.I0(commutation_state[0]), .I1(n4_adj_5845), 
            .I2(commutation_state_prev[0]), .I3(GND_net), .O(n15_adj_5755));   // verilog/TinyFPGA_B.v(146[7:48])
    defparam i2_3_lut_adj_1809.LUT_INIT = 16'hdede;
    SB_CARRY encoder0_position_30__I_0_add_1771_5 (.CI(n51770), .I0(n2631), 
            .I1(VCC_net), .CO(n51771));
    SB_LUT4 add_2502_13_lut (.I0(n70528), .I1(n2_adj_5892), .I2(n2247), 
            .I3(n51968), .O(encoder0_position_scaled_23__N_43[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2502_13_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY encoder0_position_30__I_0_add_1972_17 (.CI(n51857), .I0(n2919), 
            .I1(VCC_net), .CO(n51858));
    SB_LUT4 encoder0_position_30__I_0_add_1972_16_lut (.I0(GND_net), .I1(n2920), 
            .I2(VCC_net), .I3(n51856), .O(n2987)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1972_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2502_13 (.CI(n51968), .I0(n2_adj_5892), .I1(n2247), .CO(n51969));
    SB_LUT4 encoder0_position_30__I_0_add_1034_5_lut (.I0(GND_net), .I1(n1531), 
            .I2(VCC_net), .I3(n51380), .O(n1598)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1034_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15875_3_lut (.I0(\data_in_frame[5] [1]), .I1(rx_data[1]), .I2(n59656), 
            .I3(GND_net), .O(n29881));   // verilog/coms.v(130[12] 305[6])
    defparam i15875_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_151_11 (.CI(n50986), .I0(delay_counter[9]), .I1(GND_net), 
            .CO(n50987));
    SB_LUT4 encoder0_position_30__I_0_add_1771_4_lut (.I0(GND_net), .I1(n2632), 
            .I2(GND_net), .I3(n51769), .O(n2699)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1771_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_add_3_15_lut (.I0(GND_net), .I1(GND_net), .I2(n2), 
            .I3(n51246), .O(n294)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_add_3_14_lut (.I0(GND_net), .I1(GND_net), .I2(n2), 
            .I3(n51245), .O(n298)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1972_16 (.CI(n51856), .I0(n2920), 
            .I1(VCC_net), .CO(n51857));
    SB_LUT4 encoder0_position_30__I_0_add_1235_16_lut (.I0(GND_net), .I1(n1820), 
            .I2(VCC_net), .I3(n51491), .O(n1887)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1235_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2502_12_lut (.I0(n70554), .I1(n2_adj_5892), .I2(n2346), 
            .I3(n51967), .O(encoder0_position_scaled_23__N_43[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2502_12_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2502_12 (.CI(n51967), .I0(n2_adj_5892), .I1(n2346), .CO(n51968));
    SB_LUT4 i2_2_lut_adj_1810 (.I0(dti_counter[1]), .I1(dti_counter[2]), 
            .I2(GND_net), .I3(GND_net), .O(n10_adj_5802));   // verilog/TinyFPGA_B.v(171[9:23])
    defparam i2_2_lut_adj_1810.LUT_INIT = 16'heeee;
    SB_LUT4 i54941_1_lut (.I0(n1752), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n70635));
    defparam i54941_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i54921_1_lut (.I0(n1653), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n70615));
    defparam i54921_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i54902_1_lut (.I0(n1554), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n70596));
    defparam i54902_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY unary_minus_16_add_3_14 (.CI(n51245), .I0(GND_net), .I1(n2), 
            .CO(n51246));
    SB_CARRY encoder0_position_30__I_0_add_1235_16 (.CI(n51491), .I0(n1820), 
            .I1(VCC_net), .CO(n51492));
    SB_LUT4 i55066_1_lut (.I0(n1455), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n70760));
    defparam i55066_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_add_1972_15_lut (.I0(GND_net), .I1(n2921), 
            .I2(VCC_net), .I3(n51855), .O(n2988)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1972_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2502_11_lut (.I0(n70337), .I1(n2_adj_5892), .I2(n2445), 
            .I3(n51966), .O(encoder0_position_scaled_23__N_43[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2502_11_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY encoder0_position_30__I_0_add_1972_15 (.CI(n51855), .I0(n2921), 
            .I1(VCC_net), .CO(n51856));
    SB_CARRY add_2502_11 (.CI(n51966), .I0(n2_adj_5892), .I1(n2445), .CO(n51967));
    SB_LUT4 mux_245_i16_4_lut (.I0(encoder1_position_scaled[15]), .I1(displacement[15]), 
            .I2(n15_adj_5722), .I3(n15), .O(motor_state_23__N_91[15]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i16_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i55049_1_lut (.I0(n1356), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n70743));
    defparam i55049_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i55033_1_lut (.I0(n1257), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n70727));
    defparam i55033_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i15750_3_lut (.I0(\data_in_frame[0] [6]), .I1(rx_data[6]), .I2(n7_adj_5957), 
            .I3(GND_net), .O(n29756));   // verilog/coms.v(130[12] 305[6])
    defparam i15750_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i55018_1_lut (.I0(n1158), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n70712));
    defparam i55018_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_30__I_0_add_1034_5 (.CI(n51380), .I0(n1531), 
            .I1(VCC_net), .CO(n51381));
    SB_LUT4 unary_minus_16_add_3_13_lut (.I0(GND_net), .I1(GND_net), .I2(n14), 
            .I3(n51244), .O(n299)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2502_10_lut (.I0(n70371), .I1(n2_adj_5892), .I2(n2544), 
            .I3(n51965), .O(encoder0_position_scaled_23__N_43[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2502_10_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY unary_minus_16_add_3_13 (.CI(n51244), .I0(GND_net), .I1(n14), 
            .CO(n51245));
    SB_CARRY encoder0_position_30__I_0_add_1771_4 (.CI(n51769), .I0(n2632), 
            .I1(GND_net), .CO(n51770));
    SB_LUT4 encoder0_position_30__I_0_add_1972_14_lut (.I0(GND_net), .I1(n2922), 
            .I2(VCC_net), .I3(n51854), .O(n2989)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1972_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1034_4_lut (.I0(GND_net), .I1(n1532), 
            .I2(GND_net), .I3(n51379), .O(n1599)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1034_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1034_4 (.CI(n51379), .I0(n1532), 
            .I1(GND_net), .CO(n51380));
    SB_LUT4 unary_minus_16_add_3_12_lut (.I0(GND_net), .I1(GND_net), .I2(n15_adj_5710), 
            .I3(n51243), .O(n300)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1034_3_lut (.I0(GND_net), .I1(n1533), 
            .I2(VCC_net), .I3(n51378), .O(n1600)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1034_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_151_23 (.CI(n50998), .I0(delay_counter[21]), .I1(GND_net), 
            .CO(n50999));
    SB_CARRY unary_minus_16_add_3_12 (.CI(n51243), .I0(GND_net), .I1(n15_adj_5710), 
            .CO(n51244));
    SB_LUT4 mux_1582_i14_3_lut (.I0(duty[16]), .I1(duty[13]), .I2(n260), 
            .I3(GND_net), .O(n12187));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1582_i14_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i6_4_lut_adj_1811 (.I0(dti_counter[7]), .I1(dti_counter[4]), 
            .I2(dti_counter[5]), .I3(dti_counter[6]), .O(n14_adj_5800));   // verilog/TinyFPGA_B.v(171[9:23])
    defparam i6_4_lut_adj_1811.LUT_INIT = 16'hfffe;
    SB_CARRY add_2502_10 (.CI(n51965), .I0(n2_adj_5892), .I1(n2544), .CO(n51966));
    SB_LUT4 i11_4_lut (.I0(\data_in_frame[23] [2]), .I1(n43503), .I2(n28356), 
            .I3(rx_data[2]), .O(n57968));   // verilog/coms.v(130[12] 305[6])
    defparam i11_4_lut.LUT_INIT = 16'hca0a;
    SB_LUT4 i15879_3_lut (.I0(\data_in_frame[5] [2]), .I1(rx_data[2]), .I2(n59656), 
            .I3(GND_net), .O(n29885));   // verilog/coms.v(130[12] 305[6])
    defparam i15879_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i26923_4_lut (.I0(n61), .I1(n75), .I2(rx_data[1]), .I3(\data_in_frame[23] [1]), 
            .O(n40853));   // verilog/coms.v(94[13:20])
    defparam i26923_4_lut.LUT_INIT = 16'hfac0;
    SB_LUT4 mux_1582_i15_3_lut (.I0(duty[17]), .I1(duty[14]), .I2(n260), 
            .I3(GND_net), .O(n12185));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1582_i15_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 encoder0_position_30__I_0_add_1771_3_lut (.I0(GND_net), .I1(n2633), 
            .I2(VCC_net), .I3(n51768), .O(n2700)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1771_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2502_9_lut (.I0(n70427), .I1(n2_adj_5892), .I2(n2643), 
            .I3(n51964), .O(encoder0_position_scaled_23__N_43[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2502_9_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2502_9 (.CI(n51964), .I0(n2_adj_5892), .I1(n2643), .CO(n51965));
    SB_LUT4 encoder0_position_30__I_0_add_1235_15_lut (.I0(GND_net), .I1(n1821), 
            .I2(VCC_net), .I3(n51490), .O(n1888)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1235_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1034_3 (.CI(n51378), .I0(n1533), 
            .I1(VCC_net), .CO(n51379));
    SB_LUT4 add_2502_8_lut (.I0(n70367), .I1(n2_adj_5892), .I2(n2742), 
            .I3(n51963), .O(encoder0_position_scaled_23__N_43[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2502_8_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 unary_minus_16_add_3_11_lut (.I0(GND_net), .I1(GND_net), .I2(n16_adj_5711), 
            .I3(n51242), .O(n301)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i4880_4_lut (.I0(n25409), .I1(delay_counter[11]), .I2(delay_counter[10]), 
            .I3(delay_counter[9]), .O(n24_adj_5859));
    defparam i4880_4_lut.LUT_INIT = 16'hc8c0;
    SB_CARRY unary_minus_16_add_3_11 (.CI(n51242), .I0(GND_net), .I1(n16_adj_5711), 
            .CO(n51243));
    SB_LUT4 i26924_3_lut (.I0(n40853), .I1(\data_in_frame[23] [1]), .I2(reset), 
            .I3(GND_net), .O(n29764));   // verilog/TinyFPGA_B.v(47[5:10])
    defparam i26924_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7_4_lut_adj_1812 (.I0(dti_counter[0]), .I1(n14_adj_5800), .I2(n10_adj_5802), 
            .I3(dti_counter[3]), .O(n22835));   // verilog/TinyFPGA_B.v(171[9:23])
    defparam i7_4_lut_adj_1812.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_30__I_0_add_1034_2_lut (.I0(GND_net), .I1(n940), 
            .I2(GND_net), .I3(VCC_net), .O(n1601)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1034_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_add_3_10_lut (.I0(GND_net), .I1(GND_net), .I2(n17_adj_5712), 
            .I3(n51241), .O(n302)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i3_4_lut (.I0(\FRAME_MATCHER.i [3]), .I1(n87), .I2(\FRAME_MATCHER.i [4]), 
            .I3(n43501), .O(n61));
    defparam i3_4_lut.LUT_INIT = 16'hefff;
    SB_LUT4 i26908_4_lut (.I0(n61), .I1(n75), .I2(rx_data[0]), .I3(\data_in_frame[23] [0]), 
            .O(n40838));   // verilog/coms.v(94[13:20])
    defparam i26908_4_lut.LUT_INIT = 16'hfac0;
    SB_LUT4 i2_4_lut (.I0(n24_adj_5859), .I1(delay_counter[14]), .I2(delay_counter[12]), 
            .I3(delay_counter[13]), .O(n61386));
    defparam i2_4_lut.LUT_INIT = 16'hc800;
    SB_LUT4 i26909_3_lut (.I0(n40838), .I1(\data_in_frame[23] [0]), .I2(reset), 
            .I3(GND_net), .O(n29765));   // verilog/TinyFPGA_B.v(47[5:10])
    defparam i26909_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2502_8 (.CI(n51963), .I0(n2_adj_5892), .I1(n2742), .CO(n51964));
    SB_CARRY encoder0_position_30__I_0_add_1771_3 (.CI(n51768), .I0(n2633), 
            .I1(VCC_net), .CO(n51769));
    SB_CARRY encoder0_position_30__I_0_add_1235_15 (.CI(n51490), .I0(n1821), 
            .I1(VCC_net), .CO(n51491));
    SB_CARRY encoder0_position_30__I_0_add_1034_2 (.CI(VCC_net), .I0(n940), 
            .I1(GND_net), .CO(n51378));
    SB_CARRY unary_minus_16_add_3_10 (.CI(n51241), .I0(GND_net), .I1(n17_adj_5712), 
            .CO(n51242));
    SB_CARRY add_151_4 (.CI(n50979), .I0(delay_counter[2]), .I1(GND_net), 
            .CO(n50980));
    SB_LUT4 n71072_bdd_4_lut (.I0(n71072), .I1(duty[4]), .I2(n4922), .I3(n11564), 
            .O(pwm_setpoint_23__N_3[4]));
    defparam n71072_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 unary_minus_16_add_3_9_lut (.I0(GND_net), .I1(GND_net), .I2(n18), 
            .I3(n51240), .O(n303)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1235_14_lut (.I0(GND_net), .I1(n1822_adj_5851), 
            .I2(VCC_net), .I3(n51489), .O(n1889)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1235_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_151_10_lut (.I0(GND_net), .I1(delay_counter[8]), .I2(GND_net), 
            .I3(n50985), .O(n1231)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i2_3_lut_adj_1813 (.I0(n61386), .I1(delay_counter[18]), .I2(n25411), 
            .I3(GND_net), .O(n61472));
    defparam i2_3_lut_adj_1813.LUT_INIT = 16'hfefe;
    SB_CARRY unary_minus_16_add_3_9 (.CI(n51240), .I0(GND_net), .I1(n18), 
            .CO(n51241));
    SB_LUT4 i2_4_lut_adj_1814 (.I0(n61472), .I1(delay_counter[23]), .I2(delay_counter[20]), 
            .I3(delay_counter[19]), .O(n7));
    defparam i2_4_lut_adj_1814.LUT_INIT = 16'heccc;
    SB_LUT4 i4_4_lut_adj_1815 (.I0(n7), .I1(delay_counter[21]), .I2(delay_counter[22]), 
            .I3(n25414), .O(n62));
    defparam i4_4_lut_adj_1815.LUT_INIT = 16'hfffe;
    SB_LUT4 i5_4_lut_adj_1816 (.I0(delay_counter[24]), .I1(delay_counter[27]), 
            .I2(delay_counter[28]), .I3(delay_counter[29]), .O(n12_adj_5827));
    defparam i5_4_lut_adj_1816.LUT_INIT = 16'hfffe;
    SB_LUT4 i6_4_lut_adj_1817 (.I0(delay_counter[26]), .I1(n12_adj_5827), 
            .I2(delay_counter[25]), .I3(delay_counter[30]), .O(n25414));
    defparam i6_4_lut_adj_1817.LUT_INIT = 16'hfffe;
    SB_LUT4 i5_3_lut (.I0(delay_counter[3]), .I1(delay_counter[5]), .I2(delay_counter[4]), 
            .I3(GND_net), .O(n14_adj_5949));
    defparam i5_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i6_4_lut_adj_1818 (.I0(delay_counter[1]), .I1(delay_counter[6]), 
            .I2(delay_counter[2]), .I3(delay_counter[8]), .O(n15_adj_5948));
    defparam i6_4_lut_adj_1818.LUT_INIT = 16'hfffe;
    SB_LUT4 i8_4_lut_adj_1819 (.I0(n15_adj_5948), .I1(delay_counter[7]), 
            .I2(n14_adj_5949), .I3(delay_counter[0]), .O(n25409));
    defparam i8_4_lut_adj_1819.LUT_INIT = 16'hfffe;
    SB_LUT4 i15644_3_lut (.I0(\data_in_frame[0] [3]), .I1(rx_data[3]), .I2(n7_adj_5957), 
            .I3(GND_net), .O(n29650));   // verilog/coms.v(130[12] 305[6])
    defparam i15644_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i2_3_lut_adj_1820 (.I0(delay_counter[17]), .I1(delay_counter[16]), 
            .I2(delay_counter[15]), .I3(GND_net), .O(n25411));
    defparam i2_3_lut_adj_1820.LUT_INIT = 16'hfefe;
    SB_LUT4 add_151_22_lut (.I0(GND_net), .I1(delay_counter[20]), .I2(GND_net), 
            .I3(n50997), .O(n1219)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2502_7_lut (.I0(n70304), .I1(n2_adj_5892), .I2(n2841), 
            .I3(n51962), .O(encoder0_position_scaled_23__N_43[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2502_7_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 unary_minus_16_add_3_8_lut (.I0(GND_net), .I1(GND_net), .I2(n19_adj_5713), 
            .I3(n51239), .O(n304)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1235_14 (.CI(n51489), .I0(n1822_adj_5851), 
            .I1(VCC_net), .CO(n51490));
    SB_LUT4 i4885_3_lut (.I0(delay_counter[9]), .I1(delay_counter[10]), 
            .I2(n25409), .I3(GND_net), .O(n22_adj_5861));
    defparam i4885_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i4886_4_lut (.I0(n22_adj_5861), .I1(delay_counter[13]), .I2(delay_counter[12]), 
            .I3(delay_counter[11]), .O(n28_adj_5862));
    defparam i4886_4_lut.LUT_INIT = 16'hccc8;
    SB_CARRY unary_minus_16_add_3_8 (.CI(n51239), .I0(GND_net), .I1(n19_adj_5713), 
            .CO(n51240));
    SB_LUT4 i1_4_lut_adj_1821 (.I0(delay_counter[21]), .I1(delay_counter[20]), 
            .I2(delay_counter[23]), .I3(delay_counter[22]), .O(n4));
    defparam i1_4_lut_adj_1821.LUT_INIT = 16'h8000;
    SB_CARRY add_2502_7 (.CI(n51962), .I0(n2_adj_5892), .I1(n2841), .CO(n51963));
    SB_LUT4 unary_minus_16_add_3_7_lut (.I0(GND_net), .I1(GND_net), .I2(n20_adj_5714), 
            .I3(n51238), .O(n305)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_7 (.CI(n51238), .I0(GND_net), .I1(n20_adj_5714), 
            .CO(n51239));
    SB_LUT4 unary_minus_16_add_3_6_lut (.I0(GND_net), .I1(GND_net), .I2(n21_adj_5715), 
            .I3(n51237), .O(n306)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1235_13_lut (.I0(GND_net), .I1(n1823), 
            .I2(VCC_net), .I3(n51488), .O(n1890)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1235_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1235_13 (.CI(n51488), .I0(n1823), 
            .I1(VCC_net), .CO(n51489));
    SB_CARRY add_151_22 (.CI(n50997), .I0(delay_counter[20]), .I1(GND_net), 
            .CO(n50998));
    SB_LUT4 i2554_4_lut (.I0(n28_adj_5862), .I1(delay_counter[19]), .I2(delay_counter[18]), 
            .I3(n4_adj_5854), .O(n40));
    defparam i2554_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 encoder0_position_30__I_0_add_1771_2_lut (.I0(GND_net), .I1(n951), 
            .I2(GND_net), .I3(VCC_net), .O(n2701)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1771_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i29124_4_lut (.I0(n40), .I1(delay_counter[31]), .I2(n25414), 
            .I3(n4), .O(n1319));   // verilog/TinyFPGA_B.v(379[14:38])
    defparam i29124_4_lut.LUT_INIT = 16'h3230;
    SB_DFF commutation_state_prev_i2 (.Q(commutation_state_prev[2]), .C(clk16MHz), 
           .D(commutation_state[2]));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    SB_LUT4 i15633_3_lut (.I0(\data_in_frame[0] [1]), .I1(rx_data[1]), .I2(n7_adj_5957), 
            .I3(GND_net), .O(n29639));   // verilog/coms.v(130[12] 305[6])
    defparam i15633_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1844_3_lut (.I0(n2713), .I1(n2780), 
            .I2(n2742), .I3(GND_net), .O(n2812));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1844_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i6_4_lut_adj_1822 (.I0(ID[7]), .I1(ID[0]), .I2(ID[5]), .I3(ID[6]), 
            .O(n14_adj_5950));   // verilog/TinyFPGA_B.v(377[12:17])
    defparam i6_4_lut_adj_1822.LUT_INIT = 16'hfffe;
    SB_CARRY unary_minus_16_add_3_6 (.CI(n51237), .I0(GND_net), .I1(n21_adj_5715), 
            .CO(n51238));
    SB_CARRY encoder0_position_30__I_0_add_1771_2 (.CI(VCC_net), .I0(n951), 
            .I1(GND_net), .CO(n51768));
    SB_LUT4 i55007_2_lut (.I0(n22835), .I1(dti), .I2(GND_net), .I3(GND_net), 
            .O(dti_N_404));
    defparam i55007_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 i5_4_lut_adj_1823 (.I0(ID[4]), .I1(ID[1]), .I2(ID[3]), .I3(ID[2]), 
            .O(n13_adj_5951));   // verilog/TinyFPGA_B.v(377[12:17])
    defparam i5_4_lut_adj_1823.LUT_INIT = 16'hfffe;
    SB_LUT4 mux_4297_i25_3_lut (.I0(encoder0_position[24]), .I1(n8_adj_5767), 
            .I2(encoder0_position[30]), .I3(GND_net), .O(n519));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam mux_4297_i25_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i28920_4_lut (.I0(n13_adj_5951), .I1(baudrate[0]), .I2(n14_adj_5950), 
            .I3(n25515), .O(n42812));
    defparam i28920_4_lut.LUT_INIT = 16'hc8fa;
    SB_LUT4 add_2502_6_lut (.I0(n70273), .I1(n2_adj_5892), .I2(n2940), 
            .I3(n51961), .O(encoder0_position_scaled_23__N_43[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2502_6_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 encoder0_position_30__I_0_add_1235_12_lut (.I0(GND_net), .I1(n1824_adj_5852), 
            .I2(VCC_net), .I3(n51487), .O(n1891)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1235_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1235_12 (.CI(n51487), .I0(n1824_adj_5852), 
            .I1(VCC_net), .CO(n51488));
    SB_CARRY add_2502_6 (.CI(n51961), .I0(n2_adj_5892), .I1(n2940), .CO(n51962));
    SB_LUT4 unary_minus_16_add_3_5_lut (.I0(GND_net), .I1(GND_net), .I2(n22_adj_5716), 
            .I3(n51236), .O(n307)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_5 (.CI(n51236), .I0(GND_net), .I1(n22_adj_5716), 
            .CO(n51237));
    SB_LUT4 unary_minus_16_add_3_4_lut (.I0(GND_net), .I1(GND_net), .I2(n23_adj_5717), 
            .I3(n51235), .O(n308)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1704_25_lut (.I0(n70371), .I1(n2511), 
            .I2(VCC_net), .I3(n51767), .O(n2610)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1704_25_lut.LUT_INIT = 16'h8228;
    SB_LUT4 add_1095_25_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_setpoint_23__N_207), 
            .I3(n51117), .O(n4903)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1095_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_1095_24_lut (.I0(GND_net), .I1(GND_net), .I2(n12169), 
            .I3(n51116), .O(n4904)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1095_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1436_21_lut (.I0(GND_net), .I1(n2115), 
            .I2(VCC_net), .I3(n51609), .O(n2182)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1436_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1235_11_lut (.I0(GND_net), .I1(n1825), 
            .I2(VCC_net), .I3(n51486), .O(n1892)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1235_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1972_14 (.CI(n51854), .I0(n2922), 
            .I1(VCC_net), .CO(n51855));
    SB_LUT4 encoder0_position_30__I_0_add_1704_24_lut (.I0(GND_net), .I1(n2512), 
            .I2(VCC_net), .I3(n51766), .O(n2579)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1704_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2502_5_lut (.I0(n70241), .I1(n2_adj_5892), .I2(n3039), 
            .I3(n51960), .O(encoder0_position_scaled_23__N_43[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2502_5_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY unary_minus_16_add_3_4 (.CI(n51235), .I0(GND_net), .I1(n23_adj_5717), 
            .CO(n51236));
    SB_LUT4 unary_minus_16_add_3_3_lut (.I0(GND_net), .I1(GND_net), .I2(n24_adj_5718), 
            .I3(n51234), .O(n309)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15765_3_lut (.I0(\data_in_frame[0] [7]), .I1(rx_data[7]), .I2(n7_adj_5957), 
            .I3(GND_net), .O(n29771));   // verilog/coms.v(130[12] 305[6])
    defparam i15765_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i55079_1_lut (.I0(n1059), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n70773));
    defparam i55079_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_inv_0_i32_1_lut (.I0(encoder0_position[30]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n2_adj_5892));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_unary_minus_2_inv_0_i32_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i29120_2_lut (.I0(n62), .I1(delay_counter[31]), .I2(GND_net), 
            .I3(GND_net), .O(read_N_409));   // verilog/TinyFPGA_B.v(365[12:35])
    defparam i29120_2_lut.LUT_INIT = 16'h2222;
    SB_CARRY encoder0_position_30__I_0_add_1235_11 (.CI(n51486), .I0(n1825), 
            .I1(VCC_net), .CO(n51487));
    SB_LUT4 encoder0_position_30__I_0_add_1235_10_lut (.I0(GND_net), .I1(n1826), 
            .I2(VCC_net), .I3(n51485), .O(n1893)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1235_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1436_20_lut (.I0(GND_net), .I1(n2116), 
            .I2(VCC_net), .I3(n51608), .O(n2183)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1436_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_3 (.CI(n51234), .I0(GND_net), .I1(n24_adj_5718), 
            .CO(n51235));
    SB_CARRY add_1095_24 (.CI(n51116), .I0(GND_net), .I1(n12169), .CO(n51117));
    SB_LUT4 unary_minus_16_add_3_2_lut (.I0(n43055), .I1(GND_net), .I2(n25_adj_5719), 
            .I3(VCC_net), .O(n66963)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY encoder0_position_30__I_0_add_1235_10 (.CI(n51485), .I0(n1826), 
            .I1(VCC_net), .CO(n51486));
    SB_LUT4 encoder0_position_30__I_0_i573_3_lut (.I0(n519), .I1(n901), 
            .I2(n861), .I3(GND_net), .O(n933));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i573_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_add_1235_9_lut (.I0(GND_net), .I1(n1827), 
            .I2(VCC_net), .I3(n51484), .O(n1894)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1235_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2502_5 (.CI(n51960), .I0(n2_adj_5892), .I1(n3039), .CO(n51961));
    SB_CARRY unary_minus_16_add_3_2 (.CI(VCC_net), .I0(GND_net), .I1(n25_adj_5719), 
            .CO(n51234));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_25_lut (.I0(GND_net), .I1(encoder0_position_scaled[23]), 
            .I2(n2_adj_5797), .I3(n51233), .O(displacement_23__N_67[23])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2502_4_lut (.I0(n70202), .I1(n2_adj_5892), .I2(n3138), 
            .I3(n51959), .O(encoder0_position_scaled_23__N_43[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2502_4_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 i14808_4_lut (.I0(n27635), .I1(n1319), .I2(n66991), .I3(n42941), 
            .O(n28814));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i14808_4_lut.LUT_INIT = 16'ha088;
    SB_LUT4 i15396_3_lut (.I0(b_prev_adj_5771), .I1(b_new_adj_5997[1]), 
            .I2(debounce_cnt_N_3833_adj_5772), .I3(GND_net), .O(n29402));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    defparam i15396_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_24_lut (.I0(GND_net), .I1(encoder0_position_scaled[22]), 
            .I2(n3_adj_5796), .I3(n51232), .O(displacement_23__N_67[22])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1436_20 (.CI(n51608), .I0(n2116), 
            .I1(VCC_net), .CO(n51609));
    SB_CARRY add_2502_4 (.CI(n51959), .I0(n2_adj_5892), .I1(n3138), .CO(n51960));
    SB_CARRY encoder0_position_30__I_0_add_1235_9 (.CI(n51484), .I0(n1827), 
            .I1(VCC_net), .CO(n51485));
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_24 (.CI(n51232), .I0(encoder0_position_scaled[22]), 
            .I1(n3_adj_5796), .CO(n51233));
    SB_LUT4 encoder0_position_30__I_0_add_1972_13_lut (.I0(GND_net), .I1(n2923), 
            .I2(VCC_net), .I3(n51853), .O(n2990)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1972_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_23_lut (.I0(GND_net), .I1(encoder0_position_scaled[21]), 
            .I2(n4_adj_5795), .I3(n51231), .O(displacement_23__N_67[21])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i52342_2_lut (.I0(n70919), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n67140));
    defparam i52342_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 encoder0_position_30__I_0_i571_3_lut (.I0(n832), .I1(n899), 
            .I2(n861), .I3(GND_net), .O(n931));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i571_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_30__I_0_add_1704_24 (.CI(n51766), .I0(n2512), 
            .I1(VCC_net), .CO(n51767));
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_inv_0_i10_1_lut (.I0(encoder0_position[8]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n24_adj_5914));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_unary_minus_2_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_30__I_0_add_1972_13 (.CI(n51853), .I0(n2923), 
            .I1(VCC_net), .CO(n51854));
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_23 (.CI(n51231), .I0(encoder0_position_scaled[21]), 
            .I1(n4_adj_5795), .CO(n51232));
    SB_LUT4 i28799_3_lut (.I0(n59656), .I1(rx_data[3]), .I2(\data_in_frame[5] [3]), 
            .I3(GND_net), .O(n29890));   // verilog/coms.v(94[13:20])
    defparam i28799_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_22_lut (.I0(GND_net), .I1(encoder0_position_scaled[20]), 
            .I2(n5_adj_5825), .I3(n51230), .O(displacement_23__N_67[20])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_1095_23_lut (.I0(GND_net), .I1(GND_net), .I2(n12171), 
            .I3(n51115), .O(n4905)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1095_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_22 (.CI(n51230), .I0(encoder0_position_scaled[20]), 
            .I1(n5_adj_5825), .CO(n51231));
    SB_LUT4 encoder0_position_30__I_0_add_1235_8_lut (.I0(GND_net), .I1(n1828), 
            .I2(VCC_net), .I3(n51483), .O(n1895)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1235_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1095_23 (.CI(n51115), .I0(GND_net), .I1(n12171), .CO(n51116));
    SB_CARRY encoder0_position_30__I_0_add_1235_8 (.CI(n51483), .I0(n1828), 
            .I1(VCC_net), .CO(n51484));
    SB_LUT4 encoder0_position_30__I_0_i640_3_lut (.I0(n933), .I1(n1000), 
            .I2(n960), .I3(GND_net), .O(n1032));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i640_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_inv_0_i11_1_lut (.I0(encoder0_position[9]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n23_adj_5913));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_unary_minus_2_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_2502_3_lut (.I0(n70158), .I1(n2_adj_5892), .I2(n3237), 
            .I3(n51958), .O(encoder0_position_scaled_23__N_43[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2502_3_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 encoder0_position_30__I_0_add_1972_12_lut (.I0(GND_net), .I1(n2924), 
            .I2(VCC_net), .I3(n51852), .O(n2991)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1972_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2502_3 (.CI(n51958), .I0(n2_adj_5892), .I1(n3237), .CO(n51959));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_21_lut (.I0(GND_net), .I1(encoder0_position_scaled[19]), 
            .I2(n6_adj_5822), .I3(n51229), .O(displacement_23__N_67[19])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1235_7_lut (.I0(GND_net), .I1(n1829), 
            .I2(GND_net), .I3(n51482), .O(n1896)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1235_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_1095_22_lut (.I0(GND_net), .I1(GND_net), .I2(n12173), 
            .I3(n51114), .O(n4906)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1095_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_21 (.CI(n51229), .I0(encoder0_position_scaled[19]), 
            .I1(n6_adj_5822), .CO(n51230));
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_inv_0_i12_1_lut (.I0(encoder0_position[10]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n22_adj_5912));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_unary_minus_2_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_add_1704_23_lut (.I0(GND_net), .I1(n2513), 
            .I2(VCC_net), .I3(n51765), .O(n2580)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1704_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_i1981_3_lut (.I0(n2914), .I1(n2981), 
            .I2(n2940), .I3(GND_net), .O(n3013));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1981_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_20_lut (.I0(GND_net), .I1(encoder0_position_scaled[18]), 
            .I2(n7_adj_5821), .I3(n51228), .O(displacement_23__N_67[18])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2502_2_lut (.I0(n70164), .I1(n2_adj_5892), .I2(n43737), 
            .I3(VCC_net), .O(encoder0_position_scaled_23__N_43[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2502_2_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 mux_1582_i16_3_lut (.I0(duty[18]), .I1(duty[15]), .I2(n260), 
            .I3(GND_net), .O(n12183));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1582_i16_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 mux_1582_i17_3_lut (.I0(duty[19]), .I1(duty[16]), .I2(n260), 
            .I3(GND_net), .O(n12181));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1582_i17_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 encoder0_position_30__I_0_i707_3_lut (.I0(n1032), .I1(n1099), 
            .I2(n1059), .I3(GND_net), .O(n1131));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i707_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_adj_1824 (.I0(\FRAME_MATCHER.i [5]), .I1(n98), .I2(GND_net), 
            .I3(GND_net), .O(n87));
    defparam i1_2_lut_adj_1824.LUT_INIT = 16'hbbbb;
    SB_LUT4 n11566_bdd_4_lut_55337 (.I0(n11566), .I1(current[3]), .I2(duty[6]), 
            .I3(n11564), .O(n71066));
    defparam n11566_bdd_4_lut_55337.LUT_INIT = 16'he4aa;
    SB_CARRY encoder0_position_30__I_0_add_1972_12 (.CI(n51852), .I0(n2924), 
            .I1(VCC_net), .CO(n51853));
    SB_CARRY add_2502_2 (.CI(VCC_net), .I0(n2_adj_5892), .I1(n43737), 
            .CO(n51958));
    SB_LUT4 encoder0_position_30__I_0_add_1972_11_lut (.I0(GND_net), .I1(n2925), 
            .I2(VCC_net), .I3(n51851), .O(n2992)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1972_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_2173_33_lut (.I0(n70158), .I1(n3204), 
            .I2(VCC_net), .I3(n51957), .O(n64026)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2173_33_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_1095_22 (.CI(n51114), .I0(GND_net), .I1(n12173), .CO(n51115));
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i1_1_lut (.I0(encoder1_position_scaled[0]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n25));   // verilog/TinyFPGA_B.v(323[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_add_2173_32_lut (.I0(GND_net), .I1(n3205), 
            .I2(VCC_net), .I3(n51956), .O(n3272)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2173_32_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_i774_3_lut (.I0(n1131), .I1(n1198), 
            .I2(n1158), .I3(GND_net), .O(n1230_adj_5834));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i774_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i841_3_lut (.I0(n1230_adj_5834), .I1(n1297), 
            .I2(n1257), .I3(GND_net), .O(n1329));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i841_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_30__I_0_add_1972_11 (.CI(n51851), .I0(n2925), 
            .I1(VCC_net), .CO(n51852));
    SB_CARRY encoder0_position_30__I_0_add_1235_7 (.CI(n51482), .I0(n1829), 
            .I1(GND_net), .CO(n51483));
    SB_CARRY encoder0_position_30__I_0_add_2173_32 (.CI(n51956), .I0(n3205), 
            .I1(VCC_net), .CO(n51957));
    SB_LUT4 encoder0_position_30__I_0_add_1972_10_lut (.I0(GND_net), .I1(n2926), 
            .I2(VCC_net), .I3(n51850), .O(n2993)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1972_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_20 (.CI(n51228), .I0(encoder0_position_scaled[18]), 
            .I1(n7_adj_5821), .CO(n51229));
    SB_CARRY encoder0_position_30__I_0_add_1704_23 (.CI(n51765), .I0(n2513), 
            .I1(VCC_net), .CO(n51766));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_19_lut (.I0(GND_net), .I1(encoder0_position_scaled[17]), 
            .I2(n8_adj_5820), .I3(n51227), .O(displacement_23__N_67[17])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_19 (.CI(n51227), .I0(encoder0_position_scaled[17]), 
            .I1(n8_adj_5820), .CO(n51228));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_18_lut (.I0(GND_net), .I1(encoder0_position_scaled[16]), 
            .I2(n9_adj_5819), .I3(n51226), .O(displacement_23__N_67[16])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_18_lut.LUT_INIT = 16'hC33C;
    SB_IO RX_pad (.PACKAGE_PIN(RX), .OUTPUT_ENABLE(VCC_net), .D_IN_0(RX_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam RX_pad.PIN_TYPE = 6'b000001;
    defparam RX_pad.PULLUP = 1'b0;
    defparam RX_pad.NEG_TRIGGER = 1'b0;
    defparam RX_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO ENCODER1_B_pad (.PACKAGE_PIN(ENCODER1_B), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(ENCODER1_B_N));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ENCODER1_B_pad.PIN_TYPE = 6'b000001;
    defparam ENCODER1_B_pad.PULLUP = 1'b0;
    defparam ENCODER1_B_pad.NEG_TRIGGER = 1'b0;
    defparam ENCODER1_B_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO ENCODER1_A_pad (.PACKAGE_PIN(ENCODER1_A), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(ENCODER1_A_N));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ENCODER1_A_pad.PIN_TYPE = 6'b000001;
    defparam ENCODER1_A_pad.PULLUP = 1'b0;
    defparam ENCODER1_A_pad.NEG_TRIGGER = 1'b0;
    defparam ENCODER1_A_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO ENCODER0_B_pad (.PACKAGE_PIN(ENCODER0_B), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(ENCODER0_B_N));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ENCODER0_B_pad.PIN_TYPE = 6'b000001;
    defparam ENCODER0_B_pad.PULLUP = 1'b0;
    defparam ENCODER0_B_pad.NEG_TRIGGER = 1'b0;
    defparam ENCODER0_B_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO ENCODER0_A_pad (.PACKAGE_PIN(ENCODER0_A), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(ENCODER0_A_N));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ENCODER0_A_pad.PIN_TYPE = 6'b000001;
    defparam ENCODER0_A_pad.PULLUP = 1'b0;
    defparam ENCODER0_A_pad.NEG_TRIGGER = 1'b0;
    defparam ENCODER0_A_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO INHA_pad (.PACKAGE_PIN(INHA), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INHA_c_0));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INHA_pad.PIN_TYPE = 6'b011001;
    defparam INHA_pad.PULLUP = 1'b0;
    defparam INHA_pad.NEG_TRIGGER = 1'b0;
    defparam INHA_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO INLB_pad (.PACKAGE_PIN(INLB), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INLB_c_0));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INLB_pad.PIN_TYPE = 6'b011001;
    defparam INLB_pad.PULLUP = 1'b0;
    defparam INLB_pad.NEG_TRIGGER = 1'b0;
    defparam INLB_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO INLA_pad (.PACKAGE_PIN(INLA), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INLA_c_0));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INLA_pad.PIN_TYPE = 6'b011001;
    defparam INLA_pad.PULLUP = 1'b0;
    defparam INLA_pad.NEG_TRIGGER = 1'b0;
    defparam INLA_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO INHB_pad (.PACKAGE_PIN(INHB), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INHB_c_0));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INHB_pad.PIN_TYPE = 6'b011001;
    defparam INHB_pad.PULLUP = 1'b0;
    defparam INHB_pad.NEG_TRIGGER = 1'b0;
    defparam INHB_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DE_pad (.PACKAGE_PIN(DE), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DE_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DE_pad.PIN_TYPE = 6'b011001;
    defparam DE_pad.PULLUP = 1'b0;
    defparam DE_pad.NEG_TRIGGER = 1'b0;
    defparam DE_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 encoder0_position_30__I_0_add_2173_31_lut (.I0(GND_net), .I1(n3206), 
            .I2(VCC_net), .I3(n51955), .O(n3273)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2173_31_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15577_3_lut (.I0(\data_in_frame[21] [7]), .I1(rx_data[7]), 
            .I2(n61932), .I3(GND_net), .O(n29583));   // verilog/coms.v(130[12] 305[6])
    defparam i15577_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i908_3_lut (.I0(n1329), .I1(n1396), 
            .I2(n1356), .I3(GND_net), .O(n1428));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i908_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 n71066_bdd_4_lut (.I0(n71066), .I1(duty[3]), .I2(n4923), .I3(n11564), 
            .O(pwm_setpoint_23__N_3[3]));
    defparam n71066_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 encoder0_position_30__I_0_i1843_3_lut (.I0(n2712), .I1(n2779), 
            .I2(n2742), .I3(GND_net), .O(n2811));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1843_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i2_1_lut (.I0(encoder1_position_scaled[1]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n24_adj_5709));   // verilog/TinyFPGA_B.v(323[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 n11566_bdd_4_lut_55332 (.I0(n11566), .I1(current[2]), .I2(duty[5]), 
            .I3(n11564), .O(n71060));
    defparam n11566_bdd_4_lut_55332.LUT_INIT = 16'he4aa;
    SB_LUT4 encoder0_position_30__I_0_i975_3_lut (.I0(n1428), .I1(n1495), 
            .I2(n1455), .I3(GND_net), .O(n1527));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i975_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 n71060_bdd_4_lut (.I0(n71060), .I1(duty[2]), .I2(n4924), .I3(n11564), 
            .O(pwm_setpoint_23__N_3[2]));
    defparam n71060_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 encoder0_position_30__I_0_i1911_3_lut (.I0(n2812), .I1(n2879), 
            .I2(n2841), .I3(GND_net), .O(n2911));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1911_3_lut.LUT_INIT = 16'hacac;
    SB_DFF dti_counter_1933__i0 (.Q(dti_counter[0]), .C(clk16MHz), .D(n55));   // verilog/TinyFPGA_B.v(174[23:37])
    SB_LUT4 n11566_bdd_4_lut_55327 (.I0(n11566), .I1(current[1]), .I2(duty[4]), 
            .I3(n11564), .O(n71054));
    defparam n11566_bdd_4_lut_55327.LUT_INIT = 16'he4aa;
    SB_LUT4 n71054_bdd_4_lut (.I0(n71054), .I1(duty[1]), .I2(n4925), .I3(n11564), 
            .O(pwm_setpoint_23__N_3[1]));
    defparam n71054_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 encoder0_position_30__I_0_i1910_3_lut (.I0(n2811), .I1(n2878), 
            .I2(n2841), .I3(GND_net), .O(n2910));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1910_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i638_3_lut (.I0(n931), .I1(n998), 
            .I2(n960), .I3(GND_net), .O(n1030));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i638_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_i705_3_lut (.I0(n1030), .I1(n1097), 
            .I2(n1059), .I3(GND_net), .O(n1129));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i705_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_18 (.CI(n51226), .I0(encoder0_position_scaled[16]), 
            .I1(n9_adj_5819), .CO(n51227));
    SB_LUT4 encoder0_position_30__I_0_add_1436_19_lut (.I0(GND_net), .I1(n2117), 
            .I2(VCC_net), .I3(n51607), .O(n2184)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1436_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_4297_i3_3_lut (.I0(encoder0_position[2]), .I1(n30), .I2(encoder0_position[30]), 
            .I3(GND_net), .O(n955));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam mux_4297_i3_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_i1581_3_lut (.I0(n2322), .I1(n2389), 
            .I2(n2346), .I3(GND_net), .O(n2421));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1581_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15572_3_lut (.I0(\data_in_frame[21] [6]), .I1(rx_data[6]), 
            .I2(n61932), .I3(GND_net), .O(n29578));   // verilog/coms.v(130[12] 305[6])
    defparam i15572_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1648_3_lut (.I0(n2421), .I1(n2488), 
            .I2(n2445), .I3(GND_net), .O(n2520));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1648_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1715_3_lut (.I0(n2520), .I1(n2587), 
            .I2(n2544), .I3(GND_net), .O(n2619));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1715_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_add_1235_6_lut (.I0(GND_net), .I1(n1830), 
            .I2(GND_net), .I3(n51481), .O(n1897)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1235_6_lut.LUT_INIT = 16'hC33C;
    SB_DFF commutation_state_prev_i1 (.Q(commutation_state_prev[1]), .C(clk16MHz), 
           .D(commutation_state[1]));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    SB_LUT4 add_1095_21_lut (.I0(GND_net), .I1(GND_net), .I2(n12175), 
            .I3(n51113), .O(n4907)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1095_21_lut.LUT_INIT = 16'hC33C;
    SB_DFF pwm_setpoint_i23 (.Q(pwm_setpoint[23]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[23]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_LUT4 encoder0_position_30__I_0_i772_3_lut (.I0(n1129), .I1(n1196), 
            .I2(n1158), .I3(GND_net), .O(n1228_adj_5832));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i772_3_lut.LUT_INIT = 16'hacac;
    SB_DFF pwm_setpoint_i22 (.Q(pwm_setpoint[22]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[22]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_LUT4 encoder0_position_30__I_0_i839_3_lut (.I0(n1228_adj_5832), .I1(n1295), 
            .I2(n1257), .I3(GND_net), .O(n1327));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i839_3_lut.LUT_INIT = 16'hacac;
    SB_DFF pwm_setpoint_i21 (.Q(pwm_setpoint[21]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[21]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_LUT4 encoder0_position_30__I_0_i906_3_lut (.I0(n1327), .I1(n1394), 
            .I2(n1356), .I3(GND_net), .O(n1426));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i906_3_lut.LUT_INIT = 16'hacac;
    SB_DFF pwm_setpoint_i20 (.Q(pwm_setpoint[20]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[20]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_LUT4 encoder0_position_30__I_0_i973_3_lut (.I0(n1426), .I1(n1493), 
            .I2(n1455), .I3(GND_net), .O(n1525));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i973_3_lut.LUT_INIT = 16'hacac;
    SB_DFF pwm_setpoint_i19 (.Q(pwm_setpoint[19]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[19]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_LUT4 encoder0_position_30__I_0_i1040_3_lut (.I0(n1525), .I1(n1592), 
            .I2(n1554), .I3(GND_net), .O(n1624));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1040_3_lut.LUT_INIT = 16'hacac;
    SB_DFF pwm_setpoint_i18 (.Q(pwm_setpoint[18]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[18]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_LUT4 encoder0_position_30__I_0_i1107_3_lut (.I0(n1624), .I1(n1691), 
            .I2(n1653), .I3(GND_net), .O(n1723));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1107_3_lut.LUT_INIT = 16'hacac;
    SB_DFF pwm_setpoint_i17 (.Q(pwm_setpoint[17]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[17]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_LUT4 encoder0_position_30__I_0_i1174_3_lut (.I0(n1723), .I1(n1790_adj_5847), 
            .I2(n1752), .I3(GND_net), .O(n1822_adj_5851));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1174_3_lut.LUT_INIT = 16'hacac;
    SB_DFF pwm_setpoint_i16 (.Q(pwm_setpoint[16]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[16]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_LUT4 encoder0_position_30__I_0_i1241_3_lut (.I0(n1822_adj_5851), .I1(n1889), 
            .I2(n1851), .I3(GND_net), .O(n1921));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1241_3_lut.LUT_INIT = 16'hacac;
    SB_DFF pwm_setpoint_i15 (.Q(pwm_setpoint[15]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[15]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_LUT4 encoder0_position_30__I_0_i1308_3_lut (.I0(n1921), .I1(n1988), 
            .I2(n1950), .I3(GND_net), .O(n2020));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1308_3_lut.LUT_INIT = 16'hacac;
    SB_DFF pwm_setpoint_i14 (.Q(pwm_setpoint[14]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[14]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_LUT4 encoder0_position_30__I_0_i1375_3_lut (.I0(n2020), .I1(n2087), 
            .I2(n2049), .I3(GND_net), .O(n2119));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1375_3_lut.LUT_INIT = 16'hacac;
    SB_DFF pwm_setpoint_i13 (.Q(pwm_setpoint[13]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[13]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_LUT4 mux_4297_i26_3_lut (.I0(encoder0_position[25]), .I1(n7_adj_5774), 
            .I2(encoder0_position[30]), .I3(GND_net), .O(n518));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam mux_4297_i26_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF pwm_setpoint_i12 (.Q(pwm_setpoint[12]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[12]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_LUT4 i1_4_lut_adj_1825 (.I0(n4_adj_5780), .I1(n5_adj_5779), .I2(n518), 
            .I3(n6_adj_5775), .O(n5_adj_5936));
    defparam i1_4_lut_adj_1825.LUT_INIT = 16'heeea;
    SB_DFF pwm_setpoint_i11 (.Q(pwm_setpoint[11]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[11]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_LUT4 i1_3_lut_adj_1826 (.I0(n3), .I1(n2_adj_5781), .I2(n5_adj_5936), 
            .I3(GND_net), .O(n59507));
    defparam i1_3_lut_adj_1826.LUT_INIT = 16'h8080;
    SB_DFF pwm_setpoint_i10 (.Q(pwm_setpoint[10]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[10]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_LUT4 i43879_3_lut (.I0(n3), .I1(n7443), .I2(n59507), .I3(GND_net), 
            .O(n59508));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam i43879_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF pwm_setpoint_i9 (.Q(pwm_setpoint[9]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[9]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_LUT4 i43880_3_lut (.I0(encoder0_position[29]), .I1(n59508), .I2(encoder0_position[30]), 
            .I3(GND_net), .O(n829));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam i43880_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF pwm_setpoint_i8 (.Q(pwm_setpoint[8]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[8]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_LUT4 encoder0_position_30__I_0_i568_3_lut (.I0(n829), .I1(n896), 
            .I2(n861), .I3(GND_net), .O(n928));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i568_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF pwm_setpoint_i7 (.Q(pwm_setpoint[7]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[7]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_LUT4 encoder0_position_30__I_0_i635_3_lut (.I0(n928), .I1(n995), 
            .I2(n960), .I3(GND_net), .O(n1027));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i635_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF pwm_setpoint_i6 (.Q(pwm_setpoint[6]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[6]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_LUT4 encoder0_position_30__I_0_i702_3_lut (.I0(n1027), .I1(n1094), 
            .I2(n1059), .I3(GND_net), .O(n1126));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i702_3_lut.LUT_INIT = 16'hacac;
    SB_DFF pwm_setpoint_i5 (.Q(pwm_setpoint[5]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[5]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_CARRY encoder0_position_30__I_0_add_1972_10 (.CI(n51850), .I0(n2926), 
            .I1(VCC_net), .CO(n51851));
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_inv_0_i15_1_lut (.I0(encoder0_position[13]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n19_adj_5909));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_unary_minus_2_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_i1042_3_lut (.I0(n1527), .I1(n1594), 
            .I2(n1554), .I3(GND_net), .O(n1626));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1042_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_inv_0_i16_1_lut (.I0(encoder0_position[14]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n18_adj_5908));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_unary_minus_2_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_inv_0_i17_1_lut (.I0(encoder0_position[15]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n17_adj_5907));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_unary_minus_2_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_DFF pwm_setpoint_i4 (.Q(pwm_setpoint[4]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[4]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_CARRY encoder0_position_30__I_0_add_2173_31 (.CI(n51955), .I0(n3206), 
            .I1(VCC_net), .CO(n51956));
    SB_LUT4 encoder0_position_30__I_0_i1507_3_lut (.I0(n2216), .I1(n2283), 
            .I2(n2247), .I3(GND_net), .O(n2315));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1507_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_inv_0_i18_1_lut (.I0(encoder0_position[16]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n16_adj_5906));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_unary_minus_2_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_inv_0_i19_1_lut (.I0(encoder0_position[17]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n15_adj_5905));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_unary_minus_2_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_inv_0_i20_1_lut (.I0(encoder0_position[18]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n14_adj_5904));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_unary_minus_2_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_1095_21 (.CI(n51113), .I0(GND_net), .I1(n12175), .CO(n51114));
    SB_LUT4 encoder0_position_30__I_0_i1109_3_lut (.I0(n1626), .I1(n1693), 
            .I2(n1653), .I3(GND_net), .O(n1725));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1109_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1176_3_lut (.I0(n1725), .I1(n1792_adj_5848), 
            .I2(n1752), .I3(GND_net), .O(n1824_adj_5852));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1176_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_inv_0_i21_1_lut (.I0(encoder0_position[19]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n13_adj_5903));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_unary_minus_2_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_inv_0_i22_1_lut (.I0(encoder0_position[20]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n12_adj_5902));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_unary_minus_2_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_DFF read_197 (.Q(state_7__N_3918[0]), .C(clk16MHz), .D(n61826));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_inv_0_i23_1_lut (.I0(encoder0_position[21]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n11_adj_5901));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_unary_minus_2_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_inv_0_i24_1_lut (.I0(encoder0_position[22]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n10_adj_5900));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_unary_minus_2_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_inv_0_i25_1_lut (.I0(encoder0_position[23]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n9_adj_5899));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_unary_minus_2_inv_0_i25_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_4297_i4_3_lut (.I0(encoder0_position[3]), .I1(n29), .I2(encoder0_position[30]), 
            .I3(GND_net), .O(n954));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam mux_4297_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_i2001_3_lut (.I0(n954), .I1(n3001), 
            .I2(n2940), .I3(GND_net), .O(n3033));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2001_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_inv_0_i26_1_lut (.I0(encoder0_position[24]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n8_adj_5898));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_unary_minus_2_inv_0_i26_1_lut.LUT_INIT = 16'h5555;
    SB_DFFESR delay_counter__i1 (.Q(delay_counter[1]), .C(clk16MHz), .E(n27635), 
            .D(n1238), .R(n28814));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_inv_0_i27_1_lut (.I0(encoder0_position[25]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n7_adj_5897));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_unary_minus_2_inv_0_i27_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_inv_0_i28_1_lut (.I0(encoder0_position[26]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n6_adj_5896));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_unary_minus_2_inv_0_i28_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_inv_0_i29_1_lut (.I0(encoder0_position[27]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n5_adj_5895));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_unary_minus_2_inv_0_i29_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_inv_0_i30_1_lut (.I0(encoder0_position[28]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n4_adj_5894));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_unary_minus_2_inv_0_i30_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_inv_0_i31_1_lut (.I0(encoder0_position[29]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n3_adj_5893));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_unary_minus_2_inv_0_i31_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_4297_i5_3_lut (.I0(encoder0_position[4]), .I1(n28), .I2(encoder0_position[30]), 
            .I3(GND_net), .O(n953));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam mux_4297_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_1827 (.I0(\PID_CONTROLLER.integral_23__N_3715 [12]), 
            .I1(Ki[1]), .I2(GND_net), .I3(GND_net), .O(n110));
    defparam i1_2_lut_adj_1827.LUT_INIT = 16'h8888;
    SB_LUT4 encoder0_position_30__I_0_i1933_3_lut (.I0(n953), .I1(n2901), 
            .I2(n2841), .I3(GND_net), .O(n2933));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1933_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2000_3_lut (.I0(n2933), .I1(n3000), 
            .I2(n2940), .I3(GND_net), .O(n3032));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2000_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1865_3_lut (.I0(n952), .I1(n2801), 
            .I2(n2742), .I3(GND_net), .O(n2833));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1865_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1932_3_lut (.I0(n2833), .I1(n2900), 
            .I2(n2841), .I3(GND_net), .O(n2932));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1932_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1999_3_lut (.I0(n2932), .I1(n2999), 
            .I2(n2940), .I3(GND_net), .O(n3031));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1999_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_adj_1828 (.I0(n60815), .I1(n62089), .I2(GND_net), 
            .I3(GND_net), .O(n62091));
    defparam i1_2_lut_adj_1828.LUT_INIT = 16'heeee;
    SB_LUT4 i22921_3_lut (.I0(n214), .I1(IntegralLimit[17]), .I2(n155), 
            .I3(GND_net), .O(n36881));
    defparam i22921_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFESR delay_counter__i2 (.Q(delay_counter[2]), .C(clk16MHz), .E(n27635), 
            .D(n1237), .R(n28814));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    SB_DFFESR delay_counter__i3 (.Q(delay_counter[3]), .C(clk16MHz), .E(n27635), 
            .D(n1236), .R(n28814));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    SB_DFFESR delay_counter__i4 (.Q(delay_counter[4]), .C(clk16MHz), .E(n27635), 
            .D(n1235), .R(n28814));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    SB_DFFESR delay_counter__i5 (.Q(delay_counter[5]), .C(clk16MHz), .E(n27635), 
            .D(n1234), .R(n28814));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    SB_DFFESR delay_counter__i6 (.Q(delay_counter[6]), .C(clk16MHz), .E(n27635), 
            .D(n1233), .R(n28814));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    SB_DFFESR delay_counter__i7 (.Q(delay_counter[7]), .C(clk16MHz), .E(n27635), 
            .D(n1232), .R(n28814));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    SB_DFFESR delay_counter__i8 (.Q(delay_counter[8]), .C(clk16MHz), .E(n27635), 
            .D(n1231), .R(n28814));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    SB_DFFESR delay_counter__i9 (.Q(delay_counter[9]), .C(clk16MHz), .E(n27635), 
            .D(n1230), .R(n28814));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    SB_DFFESR delay_counter__i10 (.Q(delay_counter[10]), .C(clk16MHz), .E(n27635), 
            .D(n1229), .R(n28814));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    SB_DFFESR delay_counter__i11 (.Q(delay_counter[11]), .C(clk16MHz), .E(n27635), 
            .D(n1228), .R(n28814));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    SB_DFFESR delay_counter__i12 (.Q(delay_counter[12]), .C(clk16MHz), .E(n27635), 
            .D(n1227), .R(n28814));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    SB_DFFESR delay_counter__i13 (.Q(delay_counter[13]), .C(clk16MHz), .E(n27635), 
            .D(n1226), .R(n28814));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    SB_DFFESR delay_counter__i14 (.Q(delay_counter[14]), .C(clk16MHz), .E(n27635), 
            .D(n1225), .R(n28814));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    SB_DFFESR delay_counter__i15 (.Q(delay_counter[15]), .C(clk16MHz), .E(n27635), 
            .D(n1224), .R(n28814));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    SB_DFFESR delay_counter__i16 (.Q(delay_counter[16]), .C(clk16MHz), .E(n27635), 
            .D(n1223), .R(n28814));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    SB_DFF commutation_state_i2 (.Q(commutation_state[2]), .C(clk16MHz), 
           .D(n59505));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    SB_LUT4 i1_2_lut_adj_1829 (.I0(n36881), .I1(Ki[0]), .I2(GND_net), 
            .I3(GND_net), .O(n53));
    defparam i1_2_lut_adj_1829.LUT_INIT = 16'h8888;
    SB_LUT4 encoder0_position_30__I_0_i1243_3_lut (.I0(n1824_adj_5852), .I1(n1891), 
            .I2(n1851), .I3(GND_net), .O(n1923));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1243_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1310_3_lut (.I0(n1923), .I1(n1990), 
            .I2(n1950), .I3(GND_net), .O(n2022));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1310_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1377_3_lut (.I0(n2022), .I1(n2089), 
            .I2(n2049), .I3(GND_net), .O(n2121));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1377_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1864_3_lut (.I0(n2733), .I1(n2800), 
            .I2(n2742), .I3(GND_net), .O(n2832));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1864_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1931_3_lut (.I0(n2832), .I1(n2899), 
            .I2(n2841), .I3(GND_net), .O(n2931));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1931_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1998_3_lut (.I0(n2931), .I1(n2998), 
            .I2(n2940), .I3(GND_net), .O(n3030));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1998_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i769_3_lut (.I0(n1126), .I1(n1193), 
            .I2(n1158), .I3(GND_net), .O(n1225_adj_5829));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i769_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_17_lut (.I0(GND_net), .I1(encoder0_position_scaled[15]), 
            .I2(n10_adj_5818), .I3(n51225), .O(displacement_23__N_67[15])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_17 (.CI(n51225), .I0(encoder0_position_scaled[15]), 
            .I1(n10_adj_5818), .CO(n51226));
    SB_CARRY encoder0_position_30__I_0_add_1436_19 (.CI(n51607), .I0(n2117), 
            .I1(VCC_net), .CO(n51608));
    SB_LUT4 add_1095_20_lut (.I0(GND_net), .I1(GND_net), .I2(n12177), 
            .I3(n51112), .O(n4908)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1095_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1095_20 (.CI(n51112), .I0(GND_net), .I1(n12177), .CO(n51113));
    SB_LUT4 encoder0_position_30__I_0_add_1704_22_lut (.I0(GND_net), .I1(n2514), 
            .I2(VCC_net), .I3(n51764), .O(n2581)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1704_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_16_lut (.I0(GND_net), .I1(encoder0_position_scaled[14]), 
            .I2(n11_adj_5817), .I3(n51224), .O(displacement_23__N_67[14])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_16 (.CI(n51224), .I0(encoder0_position_scaled[14]), 
            .I1(n11_adj_5817), .CO(n51225));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_15_lut (.I0(GND_net), .I1(encoder0_position_scaled[13]), 
            .I2(n12_adj_5806), .I3(n51223), .O(displacement_23__N_67[13])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_i1574_3_lut (.I0(n2315), .I1(n2382), 
            .I2(n2346), .I3(GND_net), .O(n2414));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1574_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1444_3_lut (.I0(n2121), .I1(n2188), 
            .I2(n2148), .I3(GND_net), .O(n2220));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1444_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1511_3_lut (.I0(n2220), .I1(n2287), 
            .I2(n2247), .I3(GND_net), .O(n2319));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1511_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1578_3_lut (.I0(n2319), .I1(n2386), 
            .I2(n2346), .I3(GND_net), .O(n2418));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1578_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_4297_i27_3_lut (.I0(encoder0_position[26]), .I1(n6_adj_5775), 
            .I2(encoder0_position[30]), .I3(GND_net), .O(n625));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam mux_4297_i27_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_i1645_3_lut (.I0(n2418), .I1(n2485), 
            .I2(n2445), .I3(GND_net), .O(n2517));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1645_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i836_3_lut (.I0(n1225_adj_5829), .I1(n1292), 
            .I2(n1257), .I3(GND_net), .O(n1324));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i836_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1712_3_lut (.I0(n2517), .I1(n2584), 
            .I2(n2544), .I3(GND_net), .O(n2616));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1712_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_adj_1830 (.I0(\PID_CONTROLLER.integral_23__N_3715 [12]), 
            .I1(Ki[0]), .I2(GND_net), .I3(GND_net), .O(n38));
    defparam i1_2_lut_adj_1830.LUT_INIT = 16'h8888;
    SB_LUT4 encoder0_position_30__I_0_i1997_3_lut (.I0(n2930), .I1(n2997), 
            .I2(n2940), .I3(GND_net), .O(n3029));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1997_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1779_3_lut (.I0(n2616), .I1(n2683), 
            .I2(n2643), .I3(GND_net), .O(n2715));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1779_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1996_3_lut (.I0(n2929), .I1(n2996), 
            .I2(n2940), .I3(GND_net), .O(n3028));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1996_3_lut.LUT_INIT = 16'hacac;
    SB_IO NEOPXL_pad (.PACKAGE_PIN(NEOPXL), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(NEOPXL_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam NEOPXL_pad.PIN_TYPE = 6'b011001;
    defparam NEOPXL_pad.PULLUP = 1'b0;
    defparam NEOPXL_pad.NEG_TRIGGER = 1'b0;
    defparam NEOPXL_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO USBPU_pad (.PACKAGE_PIN(USBPU), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(GND_net));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam USBPU_pad.PIN_TYPE = 6'b011001;
    defparam USBPU_pad.PULLUP = 1'b0;
    defparam USBPU_pad.NEG_TRIGGER = 1'b0;
    defparam USBPU_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 encoder0_position_30__I_0_i1846_3_lut (.I0(n2715), .I1(n2782), 
            .I2(n2742), .I3(GND_net), .O(n2814));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1846_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1861_3_lut (.I0(n2730), .I1(n2797), 
            .I2(n2742), .I3(GND_net), .O(n2829));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1861_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1928_3_lut (.I0(n2829), .I1(n2896), 
            .I2(n2841), .I3(GND_net), .O(n2928));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1928_3_lut.LUT_INIT = 16'hacac;
    SB_IO LED_pad (.PACKAGE_PIN(LED), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(LED_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam LED_pad.PIN_TYPE = 6'b011001;
    defparam LED_pad.PULLUP = 1'b0;
    defparam LED_pad.NEG_TRIGGER = 1'b0;
    defparam LED_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 encoder0_position_30__I_0_i1995_3_lut (.I0(n2928), .I1(n2995), 
            .I2(n2940), .I3(GND_net), .O(n3027));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1995_3_lut.LUT_INIT = 16'hacac;
    SB_DFFESR dti_counter_1933__i1 (.Q(dti_counter[1]), .C(clk16MHz), .E(n27715), 
            .D(n44), .R(n29091));   // verilog/TinyFPGA_B.v(174[23:37])
    SB_DFFESR dti_counter_1933__i2 (.Q(dti_counter[2]), .C(clk16MHz), .E(n27715), 
            .D(n43_adj_5888), .R(n29091));   // verilog/TinyFPGA_B.v(174[23:37])
    SB_DFFESR dti_counter_1933__i3 (.Q(dti_counter[3]), .C(clk16MHz), .E(n27715), 
            .D(n42), .R(n29091));   // verilog/TinyFPGA_B.v(174[23:37])
    SB_DFFESR dti_counter_1933__i4 (.Q(dti_counter[4]), .C(clk16MHz), .E(n27715), 
            .D(n41), .R(n29091));   // verilog/TinyFPGA_B.v(174[23:37])
    SB_DFFESR dti_counter_1933__i5 (.Q(dti_counter[5]), .C(clk16MHz), .E(n27715), 
            .D(n40_adj_5887), .R(n29091));   // verilog/TinyFPGA_B.v(174[23:37])
    SB_DFFESR dti_counter_1933__i6 (.Q(dti_counter[6]), .C(clk16MHz), .E(n27715), 
            .D(n39), .R(n29091));   // verilog/TinyFPGA_B.v(174[23:37])
    SB_DFFESR dti_counter_1933__i7 (.Q(dti_counter[7]), .C(clk16MHz), .E(n27715), 
            .D(n38_adj_5886), .R(n29091));   // verilog/TinyFPGA_B.v(174[23:37])
    SB_LUT4 encoder0_position_30__I_0_i903_3_lut (.I0(n1324), .I1(n1391), 
            .I2(n1356), .I3(GND_net), .O(n1423));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i903_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15637_3_lut_3_lut (.I0(\FRAME_MATCHER.rx_data_ready_prev ), .I1(rx_data_ready), 
            .I2(reset), .I3(GND_net), .O(n29643));   // verilog/coms.v(130[12] 305[6])
    defparam i15637_3_lut_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_4297_i9_3_lut (.I0(encoder0_position[8]), .I1(n24_adj_5724), 
            .I2(encoder0_position[30]), .I3(GND_net), .O(n949));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam mux_4297_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_add_1972_9_lut (.I0(GND_net), .I1(n2927), 
            .I2(VCC_net), .I3(n51849), .O(n2994)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1972_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1235_6 (.CI(n51481), .I0(n1830), 
            .I1(GND_net), .CO(n51482));
    SB_LUT4 encoder0_position_30__I_0_i1661_3_lut (.I0(n949), .I1(n2501), 
            .I2(n2445), .I3(GND_net), .O(n2533));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1661_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1860_3_lut (.I0(n2729), .I1(n2796), 
            .I2(n2742), .I3(GND_net), .O(n2828));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1860_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1927_3_lut (.I0(n2828), .I1(n2895), 
            .I2(n2841), .I3(GND_net), .O(n2927));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1927_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1994_3_lut (.I0(n2927), .I1(n2994), 
            .I2(n2940), .I3(GND_net), .O(n3026));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1994_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1859_3_lut (.I0(n2728), .I1(n2795), 
            .I2(n2742), .I3(GND_net), .O(n2827));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1859_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 n11566_bdd_4_lut_55322 (.I0(n11566), .I1(current[0]), .I2(duty[3]), 
            .I3(n11564), .O(n71048));
    defparam n11566_bdd_4_lut_55322.LUT_INIT = 16'he4aa;
    SB_LUT4 encoder0_position_30__I_0_i1926_3_lut (.I0(n2827), .I1(n2894), 
            .I2(n2841), .I3(GND_net), .O(n2926));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1926_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1993_3_lut (.I0(n2926), .I1(n2993), 
            .I2(n2940), .I3(GND_net), .O(n3025));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1993_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i970_3_lut (.I0(n1423), .I1(n1490), 
            .I2(n1455), .I3(GND_net), .O(n1522));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i970_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1037_3_lut (.I0(n1522), .I1(n1589), 
            .I2(n1554), .I3(GND_net), .O(n1621));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1037_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_4297_i28_3_lut (.I0(encoder0_position[27]), .I1(n5_adj_5779), 
            .I2(encoder0_position[30]), .I3(GND_net), .O(n405));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam mux_4297_i28_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15622_3_lut_4_lut (.I0(n1742), .I1(b_prev), .I2(a_new[1]), 
            .I3(position_31__N_3836), .O(n29628));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    defparam i15622_3_lut_4_lut.LUT_INIT = 16'h3caa;
    SB_LUT4 encoder0_position_30__I_0_i1858_3_lut (.I0(n2727), .I1(n2794), 
            .I2(n2742), .I3(GND_net), .O(n2826));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1858_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_add_2173_30_lut (.I0(GND_net), .I1(n3207), 
            .I2(VCC_net), .I3(n51954), .O(n3274)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2173_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_15 (.CI(n51223), .I0(encoder0_position_scaled[13]), 
            .I1(n12_adj_5806), .CO(n51224));
    SB_CARRY encoder0_position_30__I_0_add_2173_30 (.CI(n51954), .I0(n3207), 
            .I1(VCC_net), .CO(n51955));
    SB_LUT4 encoder0_position_30__I_0_i1925_3_lut (.I0(n2826), .I1(n2893), 
            .I2(n2841), .I3(GND_net), .O(n2925));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1925_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15608_3_lut_4_lut (.I0(n1784), .I1(b_prev_adj_5771), .I2(a_new_adj_5996[1]), 
            .I3(position_31__N_3836_adj_5773), .O(n29614));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    defparam i15608_3_lut_4_lut.LUT_INIT = 16'h3caa;
    SB_LUT4 encoder0_position_30__I_0_i1992_3_lut (.I0(n2925), .I1(n2992), 
            .I2(n2940), .I3(GND_net), .O(n3024));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1992_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1104_3_lut (.I0(n1621), .I1(n1688), 
            .I2(n1653), .I3(GND_net), .O(n1720));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1104_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1171_3_lut (.I0(n1720), .I1(n1787), 
            .I2(n1752), .I3(GND_net), .O(n1819));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1171_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1238_3_lut (.I0(n1819), .I1(n1886), 
            .I2(n1851), .I3(GND_net), .O(n1918));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1238_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1305_3_lut (.I0(n1918), .I1(n1985), 
            .I2(n1950), .I3(GND_net), .O(n2017));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1305_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1372_3_lut (.I0(n2017), .I1(n2084), 
            .I2(n2049), .I3(GND_net), .O(n2116));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1372_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1440_3_lut (.I0(n2117), .I1(n2184), 
            .I2(n2148), .I3(GND_net), .O(n2216));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1440_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1438_3_lut (.I0(n2115), .I1(n2182), 
            .I2(n2148), .I3(GND_net), .O(n2214));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1438_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1439_3_lut (.I0(n2116), .I1(n2183), 
            .I2(n2148), .I3(GND_net), .O(n2215));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1439_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i29858_4_lut (.I0(n519), .I1(n831), .I2(n832), .I3(n833), 
            .O(n43759));
    defparam i29858_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 i29966_4_lut (.I0(n829), .I1(n828), .I2(n43759), .I3(n830), 
            .O(n861));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam i29966_4_lut.LUT_INIT = 16'heccc;
    SB_LUT4 i43883_3_lut (.I0(n5_adj_5779), .I1(n7445), .I2(n59507), .I3(GND_net), 
            .O(n59512));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam i43883_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_4297_i29_3_lut (.I0(encoder0_position[28]), .I1(n4_adj_5780), 
            .I2(encoder0_position[30]), .I3(GND_net), .O(n404));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam mux_4297_i29_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i43884_3_lut (.I0(encoder0_position[27]), .I1(n59512), .I2(encoder0_position[30]), 
            .I3(GND_net), .O(n831));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam i43884_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_add_1436_18_lut (.I0(GND_net), .I1(n2118), 
            .I2(VCC_net), .I3(n51606), .O(n2185)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1436_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i29788_4_lut (.I0(n520), .I1(n931), .I2(n932), .I3(n933), 
            .O(n43689));
    defparam i29788_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 i1_2_lut_adj_1831 (.I0(n929), .I1(n930), .I2(GND_net), .I3(GND_net), 
            .O(n62963));
    defparam i1_2_lut_adj_1831.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut_adj_1832 (.I0(n927), .I1(n62963), .I2(n928), .I3(n43689), 
            .O(n960));
    defparam i1_4_lut_adj_1832.LUT_INIT = 16'hfefa;
    SB_LUT4 encoder0_position_30__I_0_i570_3_lut (.I0(n831), .I1(n898), 
            .I2(n861), .I3(GND_net), .O(n930));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i570_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29794_3_lut (.I0(n521), .I1(n1032), .I2(n1033), .I3(GND_net), 
            .O(n43695));
    defparam i29794_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 encoder0_position_30__I_0_i1641_3_lut (.I0(n2414), .I1(n2481), 
            .I2(n2445), .I3(GND_net), .O(n2513));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1641_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_add_2173_29_lut (.I0(GND_net), .I1(n3208), 
            .I2(VCC_net), .I3(n51953), .O(n3275)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2173_29_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1833 (.I0(n1029), .I1(n43695), .I2(n1030), .I3(n1031), 
            .O(n60367));
    defparam i1_4_lut_adj_1833.LUT_INIT = 16'ha080;
    SB_LUT4 i55082_4_lut (.I0(n1026), .I1(n60367), .I2(n1027), .I3(n1028), 
            .O(n1059));
    defparam i55082_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_30__I_0_i637_3_lut (.I0(n930), .I1(n997), 
            .I2(n960), .I3(GND_net), .O(n1029));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i637_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_30__I_0_add_1972_9 (.CI(n51849), .I0(n2927), 
            .I1(VCC_net), .CO(n51850));
    SB_LUT4 i29864_4_lut (.I0(n522), .I1(n1131), .I2(n1132), .I3(n1133), 
            .O(n43765));
    defparam i29864_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 i1_3_lut_adj_1834 (.I0(n1126), .I1(n1127), .I2(n1128), .I3(GND_net), 
            .O(n62735));
    defparam i1_3_lut_adj_1834.LUT_INIT = 16'hfefe;
    SB_CARRY encoder0_position_30__I_0_add_1704_22 (.CI(n51764), .I0(n2514), 
            .I1(VCC_net), .CO(n51765));
    SB_LUT4 i1_2_lut_adj_1835 (.I0(n1129), .I1(n1130), .I2(GND_net), .I3(GND_net), 
            .O(n62973));
    defparam i1_2_lut_adj_1835.LUT_INIT = 16'h8888;
    SB_LUT4 i55021_4_lut (.I0(n62973), .I1(n1125), .I2(n62735), .I3(n43765), 
            .O(n1158));
    defparam i55021_4_lut.LUT_INIT = 16'h0103;
    SB_LUT4 encoder0_position_30__I_0_i704_3_lut (.I0(n1029), .I1(n1096), 
            .I2(n1059), .I3(GND_net), .O(n1128));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i704_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i29790_3_lut (.I0(n937), .I1(n1232_adj_5836), .I2(n1233_adj_5837), 
            .I3(GND_net), .O(n43691));
    defparam i29790_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i1_3_lut_adj_1836 (.I0(n1226_adj_5830), .I1(n1227_adj_5831), 
            .I2(n1228_adj_5832), .I3(GND_net), .O(n63021));
    defparam i1_3_lut_adj_1836.LUT_INIT = 16'hfefe;
    SB_LUT4 encoder0_position_30__I_0_i1708_3_lut (.I0(n2513), .I1(n2580), 
            .I2(n2544), .I3(GND_net), .O(n2612));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1708_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1837 (.I0(n1229_adj_5833), .I1(n43691), .I2(n1230_adj_5834), 
            .I3(n1231_adj_5835), .O(n60364));
    defparam i1_4_lut_adj_1837.LUT_INIT = 16'ha080;
    SB_LUT4 i55036_4_lut (.I0(n1225_adj_5829), .I1(n1224_adj_5828), .I2(n60364), 
            .I3(n63021), .O(n1257));
    defparam i55036_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_30__I_0_add_1704_21_lut (.I0(GND_net), .I1(n2515), 
            .I2(VCC_net), .I3(n51763), .O(n2582)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1704_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_i771_3_lut (.I0(n1128), .I1(n1195), 
            .I2(n1158), .I3(GND_net), .O(n1227_adj_5831));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i771_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i29782_3_lut (.I0(n938), .I1(n1332), .I2(n1333), .I3(GND_net), 
            .O(n43683));
    defparam i29782_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i1_4_lut_adj_1838 (.I0(n1325), .I1(n1326), .I2(n1327), .I3(n1328), 
            .O(n62857));
    defparam i1_4_lut_adj_1838.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_30__I_0_add_1972_8_lut (.I0(GND_net), .I1(n2928), 
            .I2(VCC_net), .I3(n51848), .O(n2995)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1972_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1839 (.I0(n1329), .I1(n43683), .I2(n1330), .I3(n1331), 
            .O(n60362));
    defparam i1_4_lut_adj_1839.LUT_INIT = 16'ha080;
    SB_LUT4 i55052_4_lut (.I0(n60362), .I1(n1323), .I2(n1324), .I3(n62857), 
            .O(n1356));
    defparam i55052_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_30__I_0_i838_3_lut (.I0(n1227_adj_5831), .I1(n1294), 
            .I2(n1257), .I3(GND_net), .O(n1326));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i838_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_30__I_0_add_1704_21 (.CI(n51763), .I0(n2515), 
            .I1(VCC_net), .CO(n51764));
    SB_CARRY encoder0_position_30__I_0_add_1972_8 (.CI(n51848), .I0(n2928), 
            .I1(VCC_net), .CO(n51849));
    SB_LUT4 encoder0_position_30__I_0_add_1704_20_lut (.I0(GND_net), .I1(n2516), 
            .I2(VCC_net), .I3(n51762), .O(n2583)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1704_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15575_4_lut_4_lut (.I0(tx_active), .I1(r_SM_Main_adj_6027[1]), 
            .I2(r_SM_Main_adj_6027[2]), .I3(n6_adj_5935), .O(n29581));   // verilog/uart_tx.v(41[10] 144[8])
    defparam i15575_4_lut_4_lut.LUT_INIT = 16'ha3aa;
    SB_LUT4 encoder0_position_30__I_0_i1728_3_lut (.I0(n2533), .I1(n2600), 
            .I2(n2544), .I3(GND_net), .O(n2632));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1728_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_4297_i30_3_lut (.I0(encoder0_position[29]), .I1(n3), .I2(encoder0_position[30]), 
            .I3(GND_net), .O(n403));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam mux_4297_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_30__I_0_add_2173_29 (.CI(n51953), .I0(n3208), 
            .I1(VCC_net), .CO(n51954));
    SB_LUT4 i6041_2_lut (.I0(n2_adj_5781), .I1(encoder0_position[30]), .I2(GND_net), 
            .I3(GND_net), .O(n402));
    defparam i6041_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 encoder0_position_30__I_0_add_1972_7_lut (.I0(GND_net), .I1(n2929), 
            .I2(GND_net), .I3(n51847), .O(n2996)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1972_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1235_5_lut (.I0(GND_net), .I1(n1831), 
            .I2(VCC_net), .I3(n51480), .O(n1898)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1235_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1704_20 (.CI(n51762), .I0(n2516), 
            .I1(VCC_net), .CO(n51763));
    SB_LUT4 encoder0_position_30__I_0_add_2173_28_lut (.I0(GND_net), .I1(n3209), 
            .I2(VCC_net), .I3(n51952), .O(n3276)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2173_28_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1704_19_lut (.I0(GND_net), .I1(n2517), 
            .I2(VCC_net), .I3(n51761), .O(n2584)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1704_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1972_7 (.CI(n51847), .I0(n2929), 
            .I1(GND_net), .CO(n51848));
    SB_CARRY encoder0_position_30__I_0_add_1704_19 (.CI(n51761), .I0(n2517), 
            .I1(VCC_net), .CO(n51762));
    SB_CARRY encoder0_position_30__I_0_add_2173_28 (.CI(n51952), .I0(n3209), 
            .I1(VCC_net), .CO(n51953));
    SB_LUT4 encoder0_position_30__I_0_add_1704_18_lut (.I0(GND_net), .I1(n2518), 
            .I2(VCC_net), .I3(n51760), .O(n2585)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1704_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_4297_i14_3_lut (.I0(encoder0_position[13]), .I1(n19_adj_5729), 
            .I2(encoder0_position[30]), .I3(GND_net), .O(n944));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam mux_4297_i14_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_add_2173_27_lut (.I0(GND_net), .I1(n3210), 
            .I2(VCC_net), .I3(n51951), .O(n3277)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2173_27_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_i1321_3_lut (.I0(n944), .I1(n2001), 
            .I2(n1950), .I3(GND_net), .O(n2033));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1321_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1388_3_lut (.I0(n2033), .I1(n2100), 
            .I2(n2049), .I3(GND_net), .O(n2132));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1388_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_30__I_0_add_1235_5 (.CI(n51480), .I0(n1831), 
            .I1(VCC_net), .CO(n51481));
    SB_LUT4 encoder0_position_30__I_0_add_1972_6_lut (.I0(GND_net), .I1(n2930), 
            .I2(GND_net), .I3(n51846), .O(n2997)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1972_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1704_18 (.CI(n51760), .I0(n2518), 
            .I1(VCC_net), .CO(n51761));
    SB_LUT4 encoder0_position_30__I_0_i1455_3_lut (.I0(n2132), .I1(n2199), 
            .I2(n2148), .I3(GND_net), .O(n2231));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1455_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1522_3_lut (.I0(n2231), .I1(n2298), 
            .I2(n2247), .I3(GND_net), .O(n2330));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1522_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1589_3_lut (.I0(n2330), .I1(n2397), 
            .I2(n2346), .I3(GND_net), .O(n2429));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1589_3_lut.LUT_INIT = 16'hacac;
    SB_DFFE \ID_READOUT_FSM.state__i0  (.Q(\ID_READOUT_FSM.state [0]), .C(clk16MHz), 
            .E(VCC_net), .D(n57114));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    SB_LUT4 encoder0_position_30__I_0_i1656_3_lut (.I0(n2429), .I1(n2496), 
            .I2(n2445), .I3(GND_net), .O(n2528));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1656_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1723_3_lut (.I0(n2528), .I1(n2595), 
            .I2(n2544), .I3(GND_net), .O(n2627));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1723_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1790_3_lut (.I0(n2627), .I1(n2694), 
            .I2(n2643), .I3(GND_net), .O(n2726));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1790_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 n71048_bdd_4_lut (.I0(n71048), .I1(duty[0]), .I2(n4926), .I3(n11564), 
            .O(pwm_setpoint_23__N_3[0]));
    defparam n71048_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFFE commutation_state_i1 (.Q(commutation_state[1]), .C(clk16MHz), 
            .E(VCC_net), .D(n30406));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    SB_LUT4 encoder0_position_30__I_0_i1857_3_lut (.I0(n2726), .I1(n2793), 
            .I2(n2742), .I3(GND_net), .O(n2825));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1857_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_30__I_0_add_1436_18 (.CI(n51606), .I0(n2118), 
            .I1(VCC_net), .CO(n51607));
    SB_CARRY encoder0_position_30__I_0_add_2173_27 (.CI(n51951), .I0(n3210), 
            .I1(VCC_net), .CO(n51952));
    SB_LUT4 encoder0_position_30__I_0_add_1704_17_lut (.I0(GND_net), .I1(n2519), 
            .I2(VCC_net), .I3(n51759), .O(n2586)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1704_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1436_17_lut (.I0(GND_net), .I1(n2119), 
            .I2(VCC_net), .I3(n51605), .O(n2186)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1436_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1972_6 (.CI(n51846), .I0(n2930), 
            .I1(GND_net), .CO(n51847));
    SB_LUT4 encoder0_position_30__I_0_i1924_3_lut (.I0(n2825), .I1(n2892), 
            .I2(n2841), .I3(GND_net), .O(n2924));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1924_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1991_3_lut (.I0(n2924), .I1(n2991), 
            .I2(n2940), .I3(GND_net), .O(n3023));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1991_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_add_1235_4_lut (.I0(GND_net), .I1(n1832), 
            .I2(GND_net), .I3(n51479), .O(n1899)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1235_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_2173_26_lut (.I0(GND_net), .I1(n3211), 
            .I2(VCC_net), .I3(n51950), .O(n3278)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2173_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2173_26 (.CI(n51950), .I0(n3211), 
            .I1(VCC_net), .CO(n51951));
    SB_CARRY encoder0_position_30__I_0_add_1704_17 (.CI(n51759), .I0(n2519), 
            .I1(VCC_net), .CO(n51760));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_14_lut (.I0(GND_net), .I1(encoder0_position_scaled[12]), 
            .I2(n13_adj_5805), .I3(n51222), .O(displacement_23__N_67[12])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1704_16_lut (.I0(GND_net), .I1(n2520), 
            .I2(VCC_net), .I3(n51758), .O(n2587)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1704_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_14 (.CI(n51222), .I0(encoder0_position_scaled[12]), 
            .I1(n13_adj_5805), .CO(n51223));
    SB_LUT4 encoder0_position_30__I_0_add_2173_25_lut (.I0(GND_net), .I1(n3212), 
            .I2(VCC_net), .I3(n51949), .O(n3279)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2173_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2173_25 (.CI(n51949), .I0(n3212), 
            .I1(VCC_net), .CO(n51950));
    SB_LUT4 encoder0_position_30__I_0_add_2173_24_lut (.I0(GND_net), .I1(n3213), 
            .I2(VCC_net), .I3(n51948), .O(n3280)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2173_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1436_17 (.CI(n51605), .I0(n2119), 
            .I1(VCC_net), .CO(n51606));
    SB_LUT4 encoder0_position_30__I_0_add_1436_16_lut (.I0(GND_net), .I1(n2120), 
            .I2(VCC_net), .I3(n51604), .O(n2187)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1436_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2173_24 (.CI(n51948), .I0(n3213), 
            .I1(VCC_net), .CO(n51949));
    SB_LUT4 encoder0_position_30__I_0_add_1972_5_lut (.I0(GND_net), .I1(n2931), 
            .I2(VCC_net), .I3(n51845), .O(n2998)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1972_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1235_4 (.CI(n51479), .I0(n1832), 
            .I1(GND_net), .CO(n51480));
    SB_CARRY encoder0_position_30__I_0_add_1704_16 (.CI(n51758), .I0(n2520), 
            .I1(VCC_net), .CO(n51759));
    SB_LUT4 encoder0_position_30__I_0_i1775_3_lut (.I0(n2612), .I1(n2679), 
            .I2(n2643), .I3(GND_net), .O(n2711));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1775_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_30__I_0_add_1972_5 (.CI(n51845), .I0(n2931), 
            .I1(VCC_net), .CO(n51846));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_13_lut (.I0(GND_net), .I1(encoder0_position_scaled[11]), 
            .I2(n14_adj_5804), .I3(n51221), .O(displacement_23__N_67[11])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_2173_23_lut (.I0(GND_net), .I1(n3214), 
            .I2(VCC_net), .I3(n51947), .O(n3281)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2173_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2173_23 (.CI(n51947), .I0(n3214), 
            .I1(VCC_net), .CO(n51948));
    SB_LUT4 i29778_3_lut (.I0(n939), .I1(n1432), .I2(n1433), .I3(GND_net), 
            .O(n43679));
    defparam i29778_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 encoder0_position_30__I_0_add_1972_4_lut (.I0(GND_net), .I1(n2932), 
            .I2(GND_net), .I3(n51844), .O(n2999)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1972_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_13 (.CI(n51221), .I0(encoder0_position_scaled[11]), 
            .I1(n14_adj_5804), .CO(n51222));
    SB_LUT4 encoder0_position_30__I_0_add_1235_3_lut (.I0(GND_net), .I1(n1833), 
            .I2(VCC_net), .I3(n51478), .O(n1900)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1235_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_2173_22_lut (.I0(GND_net), .I1(n3215), 
            .I2(VCC_net), .I3(n51946), .O(n3282)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2173_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_967_14_lut (.I0(n70760), .I1(n1422), 
            .I2(VCC_net), .I3(n51364), .O(n1521)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_967_14_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_12_lut (.I0(GND_net), .I1(encoder0_position_scaled[10]), 
            .I2(n15_adj_5803), .I3(n51220), .O(displacement_23__N_67[10])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2173_22 (.CI(n51946), .I0(n3215), 
            .I1(VCC_net), .CO(n51947));
    SB_LUT4 encoder0_position_30__I_0_add_967_13_lut (.I0(GND_net), .I1(n1423), 
            .I2(VCC_net), .I3(n51363), .O(n1490)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_967_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_i1990_3_lut (.I0(n2923), .I1(n2990), 
            .I2(n2940), .I3(GND_net), .O(n3022));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1990_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_12 (.CI(n51220), .I0(encoder0_position_scaled[10]), 
            .I1(n15_adj_5803), .CO(n51221));
    SB_CARRY encoder0_position_30__I_0_add_1436_16 (.CI(n51604), .I0(n2120), 
            .I1(VCC_net), .CO(n51605));
    SB_LUT4 i15668_3_lut_4_lut_4_lut (.I0(\data_in_frame[23] [4]), .I1(rx_data[4]), 
            .I2(reset), .I3(n75), .O(n29674));   // verilog/coms.v(130[12] 305[6])
    defparam i15668_3_lut_4_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 encoder0_position_30__I_0_add_1704_15_lut (.I0(GND_net), .I1(n2521), 
            .I2(VCC_net), .I3(n51757), .O(n2588)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1704_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_2173_21_lut (.I0(GND_net), .I1(n3216), 
            .I2(VCC_net), .I3(n51945), .O(n3283)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2173_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1436_15_lut (.I0(GND_net), .I1(n2121), 
            .I2(VCC_net), .I3(n51603), .O(n2188)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1436_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1235_3 (.CI(n51478), .I0(n1833), 
            .I1(VCC_net), .CO(n51479));
    SB_CARRY encoder0_position_30__I_0_add_967_13 (.CI(n51363), .I0(n1423), 
            .I1(VCC_net), .CO(n51364));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_11_lut (.I0(GND_net), .I1(encoder0_position_scaled[9]), 
            .I2(n16_adj_5799), .I3(n51219), .O(displacement_23__N_67[9])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2173_21 (.CI(n51945), .I0(n3216), 
            .I1(VCC_net), .CO(n51946));
    SB_DFF \ID_READOUT_FSM.state__i1  (.Q(\ID_READOUT_FSM.state [1]), .C(clk16MHz), 
           .D(n17_adj_5938));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    SB_LUT4 encoder0_position_30__I_0_add_2173_20_lut (.I0(GND_net), .I1(n3217), 
            .I2(VCC_net), .I3(n51944), .O(n3284)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2173_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_967_12_lut (.I0(GND_net), .I1(n1424), 
            .I2(VCC_net), .I3(n51362), .O(n1491)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_967_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2173_20 (.CI(n51944), .I0(n3217), 
            .I1(VCC_net), .CO(n51945));
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_11 (.CI(n51219), .I0(encoder0_position_scaled[9]), 
            .I1(n16_adj_5799), .CO(n51220));
    SB_CARRY encoder0_position_30__I_0_add_1972_4 (.CI(n51844), .I0(n2932), 
            .I1(GND_net), .CO(n51845));
    SB_LUT4 encoder0_position_30__I_0_add_1235_2_lut (.I0(GND_net), .I1(n943), 
            .I2(GND_net), .I3(VCC_net), .O(n1901)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1235_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_967_12 (.CI(n51362), .I0(n1424), 
            .I1(VCC_net), .CO(n51363));
    SB_LUT4 encoder0_position_30__I_0_i1506_3_lut (.I0(n2215), .I1(n2282), 
            .I2(n2247), .I3(GND_net), .O(n2314));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1506_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_add_2173_19_lut (.I0(GND_net), .I1(n3218), 
            .I2(VCC_net), .I3(n51943), .O(n3285)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2173_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15662_3_lut_4_lut_4_lut (.I0(\data_in_frame[23] [3]), .I1(rx_data[3]), 
            .I2(reset), .I3(n75), .O(n29668));   // verilog/coms.v(130[12] 305[6])
    defparam i15662_3_lut_4_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 encoder0_position_30__I_0_i1573_3_lut (.I0(n2314), .I1(n2381), 
            .I2(n2346), .I3(GND_net), .O(n2413));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1573_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_10_lut (.I0(GND_net), .I1(encoder0_position_scaled[8]), 
            .I2(n17_adj_5794), .I3(n51218), .O(displacement_23__N_67[8])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1972_3_lut (.I0(GND_net), .I1(n2933), 
            .I2(VCC_net), .I3(n51843), .O(n3000)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1972_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1972_3 (.CI(n51843), .I0(n2933), 
            .I1(VCC_net), .CO(n51844));
    SB_LUT4 encoder0_position_30__I_0_add_967_11_lut (.I0(GND_net), .I1(n1425), 
            .I2(VCC_net), .I3(n51361), .O(n1492)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_967_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_10 (.CI(n51218), .I0(encoder0_position_scaled[8]), 
            .I1(n17_adj_5794), .CO(n51219));
    SB_CARRY encoder0_position_30__I_0_add_1436_15 (.CI(n51603), .I0(n2121), 
            .I1(VCC_net), .CO(n51604));
    SB_CARRY encoder0_position_30__I_0_add_2173_19 (.CI(n51943), .I0(n3218), 
            .I1(VCC_net), .CO(n51944));
    SB_LUT4 encoder0_position_30__I_0_add_1972_2_lut (.I0(GND_net), .I1(n954), 
            .I2(GND_net), .I3(VCC_net), .O(n3001)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1972_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1704_15 (.CI(n51757), .I0(n2521), 
            .I1(VCC_net), .CO(n51758));
    SB_LUT4 encoder0_position_30__I_0_add_1436_14_lut (.I0(GND_net), .I1(n2122), 
            .I2(VCC_net), .I3(n51602), .O(n2189)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1436_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1704_14_lut (.I0(GND_net), .I1(n2522), 
            .I2(VCC_net), .I3(n51756), .O(n2589)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1704_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_i1105_3_lut (.I0(n1622), .I1(n1689), 
            .I2(n1653), .I3(GND_net), .O(n1721));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1105_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_add_2173_18_lut (.I0(GND_net), .I1(n3219), 
            .I2(VCC_net), .I3(n51942), .O(n3286)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2173_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1972_2 (.CI(VCC_net), .I0(n954), 
            .I1(GND_net), .CO(n51843));
    SB_CARRY encoder0_position_30__I_0_add_1436_14 (.CI(n51602), .I0(n2122), 
            .I1(VCC_net), .CO(n51603));
    SB_CARRY encoder0_position_30__I_0_add_1704_14 (.CI(n51756), .I0(n2522), 
            .I1(VCC_net), .CO(n51757));
    SB_LUT4 encoder0_position_30__I_0_i1172_3_lut (.I0(n1721), .I1(n1788_adj_5846), 
            .I2(n1752), .I3(GND_net), .O(n1820));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1172_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_add_1905_28_lut (.I0(n70304), .I1(n2808), 
            .I2(VCC_net), .I3(n51842), .O(n2907)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1905_28_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_30__I_0_i1239_3_lut (.I0(n1820), .I1(n1887), 
            .I2(n1851), .I3(GND_net), .O(n1919));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1239_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_add_1704_13_lut (.I0(GND_net), .I1(n2523), 
            .I2(VCC_net), .I3(n51755), .O(n2590)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1704_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1436_13_lut (.I0(GND_net), .I1(n2123), 
            .I2(VCC_net), .I3(n51601), .O(n2190)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1436_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1235_2 (.CI(VCC_net), .I0(n943), 
            .I1(GND_net), .CO(n51478));
    SB_CARRY encoder0_position_30__I_0_add_967_11 (.CI(n51361), .I0(n1425), 
            .I1(VCC_net), .CO(n51362));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_9_lut (.I0(GND_net), .I1(encoder0_position_scaled[7]), 
            .I2(n18_adj_5793), .I3(n51217), .O(displacement_23__N_67[7])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1436_13 (.CI(n51601), .I0(n2123), 
            .I1(VCC_net), .CO(n51602));
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_9 (.CI(n51217), .I0(encoder0_position_scaled[7]), 
            .I1(n18_adj_5793), .CO(n51218));
    SB_LUT4 encoder0_position_30__I_0_i1237_3_lut (.I0(n1818), .I1(n1885), 
            .I2(n1851), .I3(GND_net), .O(n1917));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1237_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_add_967_10_lut (.I0(GND_net), .I1(n1426), 
            .I2(VCC_net), .I3(n51360), .O(n1493)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_967_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_8_lut (.I0(GND_net), .I1(encoder0_position_scaled[6]), 
            .I2(n19_adj_5792), .I3(n51216), .O(displacement_23__N_67[6])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_i1795_3_lut (.I0(n2632), .I1(n2699), 
            .I2(n2643), .I3(GND_net), .O(n2731));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1795_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_151_21_lut (.I0(GND_net), .I1(delay_counter[19]), .I2(GND_net), 
            .I3(n50996), .O(n1220)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1704_13 (.CI(n51755), .I0(n2523), 
            .I1(VCC_net), .CO(n51756));
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_8 (.CI(n51216), .I0(encoder0_position_scaled[6]), 
            .I1(n19_adj_5792), .CO(n51217));
    SB_CARRY encoder0_position_30__I_0_add_2173_18 (.CI(n51942), .I0(n3219), 
            .I1(VCC_net), .CO(n51943));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_7_lut (.I0(GND_net), .I1(encoder0_position_scaled[5]), 
            .I2(n20), .I3(n51215), .O(displacement_23__N_67[5])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_967_10 (.CI(n51360), .I0(n1426), 
            .I1(VCC_net), .CO(n51361));
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_7 (.CI(n51215), .I0(encoder0_position_scaled[5]), 
            .I1(n20), .CO(n51216));
    SB_LUT4 i1_3_lut_adj_1840 (.I0(n5_adj_5936), .I1(n3), .I2(encoder0_position[30]), 
            .I3(GND_net), .O(n63103));
    defparam i1_3_lut_adj_1840.LUT_INIT = 16'h8080;
    SB_LUT4 encoder0_position_30__I_0_add_967_9_lut (.I0(GND_net), .I1(n1427), 
            .I2(VCC_net), .I3(n51359), .O(n1494)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_967_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_i500_4_lut (.I0(n2_adj_5781), .I1(n7442), 
            .I2(n63103), .I3(encoder0_position[30]), .O(n828));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i500_4_lut.LUT_INIT = 16'h8a80;
    SB_LUT4 i1_2_lut_4_lut_4_lut (.I0(\FRAME_MATCHER.state [3]), .I1(reset), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[8] [2]), 
            .O(n58623));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_6_lut (.I0(GND_net), .I1(encoder0_position_scaled[4]), 
            .I2(n21), .I3(n51214), .O(displacement_23__N_67[4])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_4297_i6_3_lut (.I0(encoder0_position[5]), .I1(n27), .I2(encoder0_position[30]), 
            .I3(GND_net), .O(n952));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam mux_4297_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_i1112_3_lut (.I0(n1629), .I1(n1696), 
            .I2(n1653), .I3(GND_net), .O(n1728));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1112_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_add_1436_12_lut (.I0(GND_net), .I1(n2124), 
            .I2(VCC_net), .I3(n51600), .O(n2191)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1436_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_i1179_3_lut (.I0(n1728), .I1(n1795), 
            .I2(n1752), .I3(GND_net), .O(n1827));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1179_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_151_21 (.CI(n50996), .I0(delay_counter[19]), .I1(GND_net), 
            .CO(n50997));
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_6 (.CI(n51214), .I0(encoder0_position_scaled[4]), 
            .I1(n21), .CO(n51215));
    SB_LUT4 encoder0_position_30__I_0_i1246_3_lut (.I0(n1827), .I1(n1894), 
            .I2(n1851), .I3(GND_net), .O(n1926));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1246_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_add_2173_17_lut (.I0(GND_net), .I1(n3220), 
            .I2(VCC_net), .I3(n51941), .O(n3287)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2173_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_5_lut (.I0(GND_net), .I1(encoder0_position_scaled[3]), 
            .I2(n22), .I3(n51213), .O(displacement_23__N_67[3])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1436_12 (.CI(n51600), .I0(n2124), 
            .I1(VCC_net), .CO(n51601));
    SB_LUT4 add_1095_19_lut (.I0(GND_net), .I1(GND_net), .I2(n12179), 
            .I3(n51111), .O(n4909)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1095_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_967_9 (.CI(n51359), .I0(n1427), 
            .I1(VCC_net), .CO(n51360));
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_5 (.CI(n51213), .I0(encoder0_position_scaled[3]), 
            .I1(n22), .CO(n51214));
    SB_LUT4 encoder0_position_30__I_0_i1862_3_lut (.I0(n2731), .I1(n2798), 
            .I2(n2742), .I3(GND_net), .O(n2830));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1862_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_30__I_0_add_2173_17 (.CI(n51941), .I0(n3220), 
            .I1(VCC_net), .CO(n51942));
    SB_LUT4 encoder0_position_30__I_0_add_967_8_lut (.I0(GND_net), .I1(n1428), 
            .I2(VCC_net), .I3(n51358), .O(n1495)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_967_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_967_8 (.CI(n51358), .I0(n1428), 
            .I1(VCC_net), .CO(n51359));
    SB_LUT4 mux_4297_i17_3_lut (.I0(encoder0_position[16]), .I1(n16_adj_5732), 
            .I2(encoder0_position[30]), .I3(GND_net), .O(n941));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam mux_4297_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_4_lut (.I0(GND_net), .I1(encoder0_position_scaled[2]), 
            .I2(n23), .I3(n51212), .O(displacement_23__N_67[2])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_i1313_3_lut (.I0(n1926), .I1(n1993), 
            .I2(n1950), .I3(GND_net), .O(n2025));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1313_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1380_3_lut (.I0(n2025), .I1(n2092), 
            .I2(n2049), .I3(GND_net), .O(n2124));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1380_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1447_3_lut (.I0(n2124), .I1(n2191), 
            .I2(n2148), .I3(GND_net), .O(n2223));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1447_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1514_3_lut (.I0(n2223), .I1(n2290), 
            .I2(n2247), .I3(GND_net), .O(n2322));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1514_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_4297_i16_3_lut (.I0(encoder0_position[15]), .I1(n17_adj_5731), 
            .I2(encoder0_position[30]), .I3(GND_net), .O(n942));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam mux_4297_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_i1185_3_lut (.I0(n942), .I1(n1801), 
            .I2(n1752), .I3(GND_net), .O(n1833));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1185_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1252_3_lut (.I0(n1833), .I1(n1900), 
            .I2(n1851), .I3(GND_net), .O(n1932));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1252_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1841 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[8] [3]), 
            .O(n58622));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1841.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_i1319_3_lut (.I0(n1932), .I1(n1999), 
            .I2(n1950), .I3(GND_net), .O(n2031));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1319_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_4 (.CI(n51212), .I0(encoder0_position_scaled[2]), 
            .I1(n23), .CO(n51213));
    SB_CARRY add_1095_19 (.CI(n51111), .I0(GND_net), .I1(n12179), .CO(n51112));
    SB_LUT4 encoder0_position_30__I_0_i1640_3_lut (.I0(n2413), .I1(n2480), 
            .I2(n2445), .I3(GND_net), .O(n2512));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1640_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1707_3_lut (.I0(n2512), .I1(n2579), 
            .I2(n2544), .I3(GND_net), .O(n2611));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1707_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_add_1436_11_lut (.I0(GND_net), .I1(n2125), 
            .I2(VCC_net), .I3(n51599), .O(n2192)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1436_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i3_1_lut (.I0(encoder1_position_scaled[2]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n23));   // verilog/TinyFPGA_B.v(323[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_i1386_3_lut (.I0(n2031), .I1(n2098), 
            .I2(n2049), .I3(GND_net), .O(n2130));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1386_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1117_3_lut (.I0(n941), .I1(n1701), 
            .I2(n1653), .I3(GND_net), .O(n1733));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1117_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1184_3_lut (.I0(n1733), .I1(n1800), 
            .I2(n1752), .I3(GND_net), .O(n1832));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1184_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1251_3_lut (.I0(n1832), .I1(n1899), 
            .I2(n1851), .I3(GND_net), .O(n1931));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1251_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1318_3_lut (.I0(n1931), .I1(n1998), 
            .I2(n1950), .I3(GND_net), .O(n2030));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1318_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1385_3_lut (.I0(n2030), .I1(n2097), 
            .I2(n2049), .I3(GND_net), .O(n2129));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1385_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1452_3_lut (.I0(n2129), .I1(n2196), 
            .I2(n2148), .I3(GND_net), .O(n2228));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1452_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1519_3_lut (.I0(n2228), .I1(n2295), 
            .I2(n2247), .I3(GND_net), .O(n2327));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1519_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1453_3_lut (.I0(n2130), .I1(n2197), 
            .I2(n2148), .I3(GND_net), .O(n2229));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1453_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1520_3_lut (.I0(n2229), .I1(n2296), 
            .I2(n2247), .I3(GND_net), .O(n2328));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1520_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1587_3_lut (.I0(n2328), .I1(n2395), 
            .I2(n2346), .I3(GND_net), .O(n2427));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1587_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1654_3_lut (.I0(n2427), .I1(n2494), 
            .I2(n2445), .I3(GND_net), .O(n2526));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1654_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15569_3_lut (.I0(\data_in_frame[21] [5]), .I1(rx_data[5]), 
            .I2(n61932), .I3(GND_net), .O(n29575));   // verilog/coms.v(130[12] 305[6])
    defparam i15569_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1721_3_lut (.I0(n2526), .I1(n2593), 
            .I2(n2544), .I3(GND_net), .O(n2625));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1721_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_add_1704_12_lut (.I0(GND_net), .I1(n2524), 
            .I2(VCC_net), .I3(n51754), .O(n2591)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1704_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_i1586_3_lut (.I0(n2327), .I1(n2394), 
            .I2(n2346), .I3(GND_net), .O(n2426));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1586_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1653_3_lut (.I0(n2426), .I1(n2493), 
            .I2(n2445), .I3(GND_net), .O(n2525));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1653_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1720_3_lut (.I0(n2525), .I1(n2592), 
            .I2(n2544), .I3(GND_net), .O(n2624));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1720_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1788_3_lut (.I0(n2625), .I1(n2692), 
            .I2(n2643), .I3(GND_net), .O(n2724));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1788_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1787_3_lut (.I0(n2624), .I1(n2691), 
            .I2(n2643), .I3(GND_net), .O(n2723));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1787_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1855_3_lut (.I0(n2724), .I1(n2791), 
            .I2(n2742), .I3(GND_net), .O(n2823));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1855_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i43887_3_lut (.I0(n7_adj_5774), .I1(n7447), .I2(n59507), .I3(GND_net), 
            .O(n59516));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam i43887_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_i1922_3_lut (.I0(n2823), .I1(n2890), 
            .I2(n2841), .I3(GND_net), .O(n2922));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1922_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1989_3_lut (.I0(n2922), .I1(n2989), 
            .I2(n2940), .I3(GND_net), .O(n3021));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1989_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i43888_3_lut (.I0(encoder0_position[25]), .I1(n59516), .I2(encoder0_position[30]), 
            .I3(GND_net), .O(n833));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam i43888_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1842 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[8] [4]), 
            .O(n58621));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1842.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_i572_3_lut (.I0(n833), .I1(n900), 
            .I2(n861), .I3(GND_net), .O(n932));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i572_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_i639_3_lut (.I0(n932), .I1(n999), 
            .I2(n960), .I3(GND_net), .O(n1031));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i639_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_i706_3_lut (.I0(n1031), .I1(n1098), 
            .I2(n1059), .I3(GND_net), .O(n1130));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i706_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_1582_i18_3_lut (.I0(duty[20]), .I1(duty[17]), .I2(n260), 
            .I3(GND_net), .O(n12179));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1582_i18_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 encoder0_position_30__I_0_i773_3_lut (.I0(n1130), .I1(n1197), 
            .I2(n1158), .I3(GND_net), .O(n1229_adj_5833));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i773_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i840_3_lut (.I0(n1229_adj_5833), .I1(n1296), 
            .I2(n1257), .I3(GND_net), .O(n1328));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i840_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_30__I_0_add_1436_11 (.CI(n51599), .I0(n2125), 
            .I1(VCC_net), .CO(n51600));
    SB_LUT4 encoder0_position_30__I_0_add_1436_10_lut (.I0(GND_net), .I1(n2126), 
            .I2(VCC_net), .I3(n51598), .O(n2193)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1436_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_i907_3_lut (.I0(n1328), .I1(n1395), 
            .I2(n1356), .I3(GND_net), .O(n1427));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i907_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1843 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[8] [5]), 
            .O(n58620));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1843.LUT_INIT = 16'h2300;
    SB_CARRY encoder0_position_30__I_0_add_1436_10 (.CI(n51598), .I0(n2126), 
            .I1(VCC_net), .CO(n51599));
    SB_LUT4 encoder0_position_30__I_0_i974_3_lut (.I0(n1427), .I1(n1494), 
            .I2(n1455), .I3(GND_net), .O(n1526));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i974_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1041_3_lut (.I0(n1526), .I1(n1593), 
            .I2(n1554), .I3(GND_net), .O(n1625));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1041_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1108_3_lut (.I0(n1625), .I1(n1692), 
            .I2(n1653), .I3(GND_net), .O(n1724));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1108_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i4_1_lut (.I0(encoder1_position_scaled[3]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n22));   // verilog/TinyFPGA_B.v(323[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_i1175_3_lut (.I0(n1724), .I1(n1791), 
            .I2(n1752), .I3(GND_net), .O(n1823));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1175_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16585_2_lut_4_lut (.I0(reset), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2873));   // verilog/coms.v(130[12] 305[6])
    defparam i16585_2_lut_4_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_i1242_3_lut (.I0(n1823), .I1(n1890), 
            .I2(n1851), .I3(GND_net), .O(n1922));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1242_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1844 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[8] [6]), 
            .O(n58671));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1844.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_i1309_3_lut (.I0(n1922), .I1(n1989), 
            .I2(n1950), .I3(GND_net), .O(n2021));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1309_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1376_3_lut (.I0(n2021), .I1(n2088), 
            .I2(n2049), .I3(GND_net), .O(n2120));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1376_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_3_lut (.I0(GND_net), .I1(encoder0_position_scaled[1]), 
            .I2(n24_adj_5709), .I3(n51211), .O(displacement_23__N_67[1])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_967_7_lut (.I0(GND_net), .I1(n1429), 
            .I2(GND_net), .I3(n51357), .O(n1496)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_967_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_967_7 (.CI(n51357), .I0(n1429), 
            .I1(GND_net), .CO(n51358));
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1845 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[8] [7]), 
            .O(n58619));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1845.LUT_INIT = 16'h2300;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_3 (.CI(n51211), .I0(encoder0_position_scaled[1]), 
            .I1(n24_adj_5709), .CO(n51212));
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1846 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[9] [0]), 
            .O(n58495));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1846.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1847 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[9] [1]), 
            .O(n58618));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1847.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_i1443_3_lut (.I0(n2120), .I1(n2187), 
            .I2(n2148), .I3(GND_net), .O(n2219));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1443_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_30__I_0_add_1704_12 (.CI(n51754), .I0(n2524), 
            .I1(VCC_net), .CO(n51755));
    SB_LUT4 encoder0_position_30__I_0_add_2173_16_lut (.I0(GND_net), .I1(n3221), 
            .I2(VCC_net), .I3(n51940), .O(n3288)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2173_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1848 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[9] [2]), 
            .O(n58617));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1848.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i5_1_lut (.I0(encoder1_position_scaled[4]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n21));   // verilog/TinyFPGA_B.v(323[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1849 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[9] [3]), 
            .O(n58616));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1849.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1850 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[9] [4]), 
            .O(n58615));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1850.LUT_INIT = 16'h2300;
    SB_CARRY encoder0_position_30__I_0_add_2173_16 (.CI(n51940), .I0(n3221), 
            .I1(VCC_net), .CO(n51941));
    SB_LUT4 encoder0_position_30__I_0_add_2173_15_lut (.I0(GND_net), .I1(n3222), 
            .I2(VCC_net), .I3(n51939), .O(n3289)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2173_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1851 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[9] [5]), 
            .O(n58614));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1851.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1852 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[9] [6]), 
            .O(n58613));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1852.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1853 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[9] [7]), 
            .O(n58612));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1853.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_add_1905_27_lut (.I0(GND_net), .I1(n2809), 
            .I2(VCC_net), .I3(n51841), .O(n2876)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1905_27_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1854 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[10] [0]), 
            .O(n58611));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1854.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_add_1436_9_lut (.I0(GND_net), .I1(n2127), 
            .I2(VCC_net), .I3(n51597), .O(n2194)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1436_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1855 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[10] [1]), 
            .O(n58610));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1855.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_add_1704_11_lut (.I0(GND_net), .I1(n2525), 
            .I2(VCC_net), .I3(n51753), .O(n2592)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1704_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1856 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[10] [2]), 
            .O(n58609));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1856.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1857 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[10] [3]), 
            .O(n58608));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1857.LUT_INIT = 16'h2300;
    SB_CARRY encoder0_position_30__I_0_add_1704_11 (.CI(n51753), .I0(n2525), 
            .I1(VCC_net), .CO(n51754));
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i6_1_lut (.I0(encoder1_position_scaled[5]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n20));   // verilog/TinyFPGA_B.v(323[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i7_1_lut (.I0(encoder1_position_scaled[6]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n19_adj_5792));   // verilog/TinyFPGA_B.v(323[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_30__I_0_add_2173_15 (.CI(n51939), .I0(n3222), 
            .I1(VCC_net), .CO(n51940));
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1858 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[10] [4]), 
            .O(n58607));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1858.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1859 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[10] [5]), 
            .O(n58606));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1859.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_i1510_3_lut (.I0(n2219), .I1(n2286), 
            .I2(n2247), .I3(GND_net), .O(n2318));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1510_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15564_3_lut (.I0(\data_in_frame[21] [4]), .I1(rx_data[4]), 
            .I2(n61932), .I3(GND_net), .O(n29570));   // verilog/coms.v(130[12] 305[6])
    defparam i15564_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_2_lut (.I0(GND_net), .I1(encoder0_position_scaled[0]), 
            .I2(n25), .I3(VCC_net), .O(displacement_23__N_67[0])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_967_6_lut (.I0(GND_net), .I1(n1430), 
            .I2(GND_net), .I3(n51356), .O(n1497)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_967_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i8_1_lut (.I0(encoder1_position_scaled[7]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n18_adj_5793));   // verilog/TinyFPGA_B.v(323[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_2 (.CI(VCC_net), .I0(encoder0_position_scaled[0]), 
            .I1(n25), .CO(n51211));
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1860 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[10] [6]), 
            .O(n58605));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1860.LUT_INIT = 16'h2300;
    SB_LUT4 i15545_3_lut (.I0(\data_in_frame[21] [3]), .I1(rx_data[3]), 
            .I2(n61932), .I3(GND_net), .O(n29551));   // verilog/coms.v(130[12] 305[6])
    defparam i15545_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_4297_i7_3_lut (.I0(encoder0_position[6]), .I1(n26), .I2(encoder0_position[30]), 
            .I3(GND_net), .O(n951));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam mux_4297_i7_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_i1797_3_lut (.I0(n951), .I1(n2701), 
            .I2(n2643), .I3(GND_net), .O(n2733));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1797_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1577_3_lut (.I0(n2318), .I1(n2385), 
            .I2(n2346), .I3(GND_net), .O(n2417));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1577_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_add_2173_14_lut (.I0(GND_net), .I1(n3223), 
            .I2(VCC_net), .I3(n51938), .O(n3290)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2173_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_i1644_3_lut (.I0(n2417), .I1(n2484), 
            .I2(n2445), .I3(GND_net), .O(n2516));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1644_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15536_3_lut (.I0(\data_in_frame[21] [2]), .I1(rx_data[2]), 
            .I2(n61932), .I3(GND_net), .O(n29542));   // verilog/coms.v(130[12] 305[6])
    defparam i15536_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_adj_1861 (.I0(n1427), .I1(n1428), .I2(GND_net), .I3(GND_net), 
            .O(n63047));
    defparam i1_2_lut_adj_1861.LUT_INIT = 16'heeee;
    SB_CARRY encoder0_position_30__I_0_add_1905_27 (.CI(n51841), .I0(n2809), 
            .I1(VCC_net), .CO(n51842));
    SB_LUT4 encoder0_position_30__I_0_i1988_3_lut (.I0(n2921), .I1(n2988), 
            .I2(n2940), .I3(GND_net), .O(n3020));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1988_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i777_3_lut (.I0(n522), .I1(n1201), 
            .I2(n1158), .I3(GND_net), .O(n1233_adj_5837));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i777_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i844_3_lut (.I0(n1233_adj_5837), .I1(n1300), 
            .I2(n1257), .I3(GND_net), .O(n1332));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i844_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i911_3_lut (.I0(n1332), .I1(n1399), 
            .I2(n1356), .I3(GND_net), .O(n1431));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i911_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15533_3_lut (.I0(\data_in_frame[21] [1]), .I1(rx_data[1]), 
            .I2(n61932), .I3(GND_net), .O(n29539));   // verilog/coms.v(130[12] 305[6])
    defparam i15533_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i978_3_lut (.I0(n1431), .I1(n1498), 
            .I2(n1455), .I3(GND_net), .O(n1530));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i978_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1045_3_lut (.I0(n1530), .I1(n1597), 
            .I2(n1554), .I3(GND_net), .O(n1629));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1045_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15529_3_lut (.I0(\data_in_frame[21] [0]), .I1(rx_data[0]), 
            .I2(n61932), .I3(GND_net), .O(n29535));   // verilog/coms.v(130[12] 305[6])
    defparam i15529_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_30__I_0_add_967_6 (.CI(n51356), .I0(n1430), 
            .I1(GND_net), .CO(n51357));
    SB_LUT4 i12_4_lut_adj_1862 (.I0(\data_in_frame[20] [6]), .I1(n28307), 
            .I2(n160), .I3(rx_data[6]), .O(n57974));   // verilog/coms.v(130[12] 305[6])
    defparam i12_4_lut_adj_1862.LUT_INIT = 16'ha3a0;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i9_1_lut (.I0(encoder1_position_scaled[8]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n17_adj_5794));   // verilog/TinyFPGA_B.v(323[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_1095_18_lut (.I0(GND_net), .I1(GND_net), .I2(n12181), 
            .I3(n51110), .O(n4910)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1095_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_967_5_lut (.I0(GND_net), .I1(n1431), 
            .I2(VCC_net), .I3(n51355), .O(n1498)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_967_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1095_18 (.CI(n51110), .I0(GND_net), .I1(n12181), .CO(n51111));
    SB_LUT4 add_1095_17_lut (.I0(GND_net), .I1(GND_net), .I2(n12183), 
            .I3(n51109), .O(n4911)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1095_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1436_9 (.CI(n51597), .I0(n2127), 
            .I1(VCC_net), .CO(n51598));
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1863 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[10] [7]), 
            .O(n58604));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1863.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1864 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[11] [0]), 
            .O(n58603));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1864.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1865 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[11] [1]), 
            .O(n58602));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1865.LUT_INIT = 16'h2300;
    SB_CARRY encoder0_position_30__I_0_add_2173_14 (.CI(n51938), .I0(n3223), 
            .I1(VCC_net), .CO(n51939));
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1866 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[11] [2]), 
            .O(n58601));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1866.LUT_INIT = 16'h2300;
    SB_CARRY encoder0_position_30__I_0_add_967_5 (.CI(n51355), .I0(n1431), 
            .I1(VCC_net), .CO(n51356));
    SB_LUT4 encoder0_position_30__I_0_add_2173_13_lut (.I0(GND_net), .I1(n3224), 
            .I2(VCC_net), .I3(n51937), .O(n3291)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2173_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1704_10_lut (.I0(GND_net), .I1(n2526), 
            .I2(VCC_net), .I3(n51752), .O(n2593)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1704_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1095_17 (.CI(n51109), .I0(GND_net), .I1(n12183), .CO(n51110));
    SB_DFF reset_198 (.Q(reset), .C(clk16MHz), .D(n57200));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    SB_LUT4 i12_4_lut_adj_1867 (.I0(\data_in_frame[20] [2]), .I1(n28307), 
            .I2(n160), .I3(rx_data[2]), .O(n57980));   // verilog/coms.v(130[12] 305[6])
    defparam i12_4_lut_adj_1867.LUT_INIT = 16'ha3a0;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1868 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[11] [3]), 
            .O(n58600));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1868.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1869 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[11] [4]), 
            .O(n58599));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1869.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1870 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[11] [5]), 
            .O(n58598));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1870.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1871 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[11] [6]), 
            .O(n58597));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1871.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_i1711_3_lut (.I0(n2516), .I1(n2583), 
            .I2(n2544), .I3(GND_net), .O(n2615));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1711_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1872 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[11] [7]), 
            .O(n58596));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1872.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1873 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[12] [0]), 
            .O(n58595));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1873.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1874 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[12] [1]), 
            .O(n58594));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1874.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1875 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[12] [2]), 
            .O(n58593));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1875.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_i1774_3_lut (.I0(n2611), .I1(n2678), 
            .I2(n2643), .I3(GND_net), .O(n2710));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1774_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1876 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[12] [3]), 
            .O(n58592));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1876.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1877 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[12] [4]), 
            .O(n58591));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1877.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_3_lut (.I0(n15_adj_5755), .I1(n22835), .I2(dti), 
            .I3(GND_net), .O(n27715));
    defparam i1_2_lut_3_lut.LUT_INIT = 16'heaea;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1878 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[12] [5]), 
            .O(n58590));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1878.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_adj_1879 (.I0(reset), .I1(n159), .I2(GND_net), .I3(GND_net), 
            .O(n160));
    defparam i1_2_lut_adj_1879.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1880 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[12] [6]), 
            .O(n58589));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1880.LUT_INIT = 16'h2300;
    SB_LUT4 i15089_2_lut_3_lut (.I0(n15_adj_5755), .I1(n22835), .I2(dti), 
            .I3(GND_net), .O(n29091));   // verilog/TinyFPGA_B.v(174[23:37])
    defparam i15089_2_lut_3_lut.LUT_INIT = 16'h2a2a;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1881 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[12] [7]), 
            .O(n58588));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1881.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1882 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[13] [0]), 
            .O(n28975));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1882.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_i1778_3_lut (.I0(n2615), .I1(n2682), 
            .I2(n2643), .I3(GND_net), .O(n2714));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1778_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1883 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[13] [1]), 
            .O(n58587));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1883.LUT_INIT = 16'h2300;
    SB_LUT4 i12_4_lut_adj_1884 (.I0(\data_in_frame[20] [0]), .I1(n28307), 
            .I2(n160), .I3(rx_data[0]), .O(n57986));   // verilog/coms.v(130[12] 305[6])
    defparam i12_4_lut_adj_1884.LUT_INIT = 16'ha3a0;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1885 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[13] [2]), 
            .O(n58586));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1885.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1886 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[13] [3]), 
            .O(n58585));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1886.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1887 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[13] [4]), 
            .O(n58584));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1887.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1888 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[13] [5]), 
            .O(n58583));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1888.LUT_INIT = 16'h2300;
    SB_CARRY encoder0_position_30__I_0_add_2173_13 (.CI(n51937), .I0(n3224), 
            .I1(VCC_net), .CO(n51938));
    SB_LUT4 i1_4_lut_adj_1889 (.I0(n1429), .I1(n43679), .I2(n1430), .I3(n1431), 
            .O(n60375));
    defparam i1_4_lut_adj_1889.LUT_INIT = 16'ha080;
    SB_LUT4 encoder0_position_30__I_0_add_1905_26_lut (.I0(GND_net), .I1(n2810), 
            .I2(VCC_net), .I3(n51840), .O(n2877)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1905_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_1095_16_lut (.I0(GND_net), .I1(GND_net), .I2(n12185), 
            .I3(n51108), .O(n4912)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1095_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1905_26 (.CI(n51840), .I0(n2810), 
            .I1(VCC_net), .CO(n51841));
    SB_CARRY encoder0_position_30__I_0_add_1704_10 (.CI(n51752), .I0(n2526), 
            .I1(VCC_net), .CO(n51753));
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1890 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[13] [6]), 
            .O(n58582));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1890.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_add_1704_9_lut (.I0(GND_net), .I1(n2527), 
            .I2(VCC_net), .I3(n51751), .O(n2594)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1704_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1891 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[13] [7]), 
            .O(n58581));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1891.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1892 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[14] [0]), 
            .O(n58580));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1892.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_add_967_4_lut (.I0(GND_net), .I1(n1432), 
            .I2(GND_net), .I3(n51354), .O(n1499)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_967_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_967_4 (.CI(n51354), .I0(n1432), 
            .I1(GND_net), .CO(n51355));
    SB_LUT4 encoder0_position_30__I_0_i1845_3_lut (.I0(n2714), .I1(n2781), 
            .I2(n2742), .I3(GND_net), .O(n2813));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1845_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_1095_16 (.CI(n51108), .I0(GND_net), .I1(n12185), .CO(n51109));
    SB_LUT4 encoder0_position_30__I_0_add_1905_25_lut (.I0(GND_net), .I1(n2811), 
            .I2(VCC_net), .I3(n51839), .O(n2878)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1905_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1704_9 (.CI(n51751), .I0(n2527), 
            .I1(VCC_net), .CO(n51752));
    SB_LUT4 add_1095_15_lut (.I0(GND_net), .I1(GND_net), .I2(n12187), 
            .I3(n51107), .O(n4913)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1095_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1704_8_lut (.I0(GND_net), .I1(n2528), 
            .I2(VCC_net), .I3(n51750), .O(n2595)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1704_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1436_8_lut (.I0(GND_net), .I1(n2128), 
            .I2(VCC_net), .I3(n51596), .O(n2195)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1436_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1704_8 (.CI(n51750), .I0(n2528), 
            .I1(VCC_net), .CO(n51751));
    SB_LUT4 encoder0_position_30__I_0_add_2173_12_lut (.I0(GND_net), .I1(n3225), 
            .I2(VCC_net), .I3(n51936), .O(n3292)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2173_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1905_25 (.CI(n51839), .I0(n2811), 
            .I1(VCC_net), .CO(n51840));
    SB_LUT4 encoder0_position_30__I_0_i1841_3_lut (.I0(n2710), .I1(n2777), 
            .I2(n2742), .I3(GND_net), .O(n2809));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1841_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_add_1905_24_lut (.I0(GND_net), .I1(n2812), 
            .I2(VCC_net), .I3(n51838), .O(n2879)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1905_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_151_10 (.CI(n50985), .I0(delay_counter[8]), .I1(GND_net), 
            .CO(n50986));
    SB_LUT4 encoder0_position_30__I_0_add_967_3_lut (.I0(GND_net), .I1(n1433), 
            .I2(VCC_net), .I3(n51353), .O(n1500)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_967_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1893 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[14] [1]), 
            .O(n58579));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1893.LUT_INIT = 16'h2300;
    SB_LUT4 mux_4297_i15_3_lut (.I0(encoder0_position[14]), .I1(n18_adj_5730), 
            .I2(encoder0_position[30]), .I3(GND_net), .O(n943));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam mux_4297_i15_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1894 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[14] [2]), 
            .O(n58578));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1894.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_i1253_3_lut (.I0(n943), .I1(n1901), 
            .I2(n1851), .I3(GND_net), .O(n1933));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1253_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_30__I_0_add_2173_12 (.CI(n51936), .I0(n3225), 
            .I1(VCC_net), .CO(n51937));
    SB_CARRY encoder0_position_30__I_0_add_1905_24 (.CI(n51838), .I0(n2812), 
            .I1(VCC_net), .CO(n51839));
    SB_LUT4 encoder0_position_30__I_0_add_1704_7_lut (.I0(GND_net), .I1(n2529), 
            .I2(GND_net), .I3(n51749), .O(n2596)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1704_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_4297_i8_3_lut (.I0(encoder0_position[7]), .I1(n25_adj_5723), 
            .I2(encoder0_position[30]), .I3(GND_net), .O(n950));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam mux_4297_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_i1729_3_lut (.I0(n950), .I1(n2601), 
            .I2(n2544), .I3(GND_net), .O(n2633));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1729_3_lut.LUT_INIT = 16'hacac;
    SB_DFFESR delay_counter__i0 (.Q(delay_counter[0]), .C(clk16MHz), .E(n27635), 
            .D(n1239), .R(n28814));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    SB_LUT4 encoder0_position_30__I_0_i1796_3_lut (.I0(n2633), .I1(n2700), 
            .I2(n2643), .I3(GND_net), .O(n2732));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1796_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1895 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[14] [3]), 
            .O(n58577));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1895.LUT_INIT = 16'h2300;
    SB_CARRY encoder0_position_30__I_0_add_1436_8 (.CI(n51596), .I0(n2128), 
            .I1(VCC_net), .CO(n51597));
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1896 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[14] [4]), 
            .O(n58576));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1896.LUT_INIT = 16'h2300;
    SB_LUT4 i1_4_lut_adj_1897 (.I0(n1424), .I1(n1425), .I2(n1426), .I3(n63047), 
            .O(n63053));
    defparam i1_4_lut_adj_1897.LUT_INIT = 16'hfffe;
    SB_LUT4 i55069_4_lut (.I0(n1423), .I1(n1422), .I2(n63053), .I3(n60375), 
            .O(n1455));
    defparam i55069_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_30__I_0_i905_3_lut (.I0(n1326), .I1(n1393), 
            .I2(n1356), .I3(GND_net), .O(n1425));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i905_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i29776_3_lut (.I0(n940), .I1(n1532), .I2(n1533), .I3(GND_net), 
            .O(n43677));
    defparam i29776_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1898 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[14] [5]), 
            .O(n58575));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1898.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_add_1905_23_lut (.I0(GND_net), .I1(n2813), 
            .I2(VCC_net), .I3(n51837), .O(n2880)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1905_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_967_3 (.CI(n51353), .I0(n1433), 
            .I1(VCC_net), .CO(n51354));
    SB_LUT4 encoder0_position_30__I_0_add_1436_7_lut (.I0(GND_net), .I1(n2129), 
            .I2(GND_net), .I3(n51595), .O(n2196)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1436_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_967_2_lut (.I0(GND_net), .I1(n939), 
            .I2(GND_net), .I3(VCC_net), .O(n1501)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_967_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1704_7 (.CI(n51749), .I0(n2529), 
            .I1(GND_net), .CO(n51750));
    SB_LUT4 i1_4_lut_adj_1899 (.I0(o_Rx_DV_N_3488[12]), .I1(n4935), .I2(o_Rx_DV_N_3488[8]), 
            .I3(n62449), .O(n62455));
    defparam i1_4_lut_adj_1899.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1900 (.I0(o_Rx_DV_N_3488[24]), .I1(n29_adj_5857), 
            .I2(n23_adj_5860), .I3(n62455), .O(n62461));
    defparam i1_4_lut_adj_1900.LUT_INIT = 16'hfffe;
    SB_DFFESR GHC_192 (.Q(GHC), .C(clk16MHz), .E(n27585), .D(GHC_N_391), 
            .R(n28807));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    SB_DFFESR GHB_190 (.Q(GHB), .C(clk16MHz), .E(n27585), .D(GHB_N_377), 
            .R(n28807));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    SB_DFF displacement_i23 (.Q(displacement[23]), .C(clk16MHz), .D(displacement_23__N_67[23]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_LUT4 encoder0_position_30__I_0_add_2173_11_lut (.I0(GND_net), .I1(n3226), 
            .I2(VCC_net), .I3(n51935), .O(n3293)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2173_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i16114_4_lut (.I0(r_Rx_Data), .I1(rx_data[1]), .I2(n62461), 
            .I3(n27_adj_5858), .O(n30120));   // verilog/uart_rx.v(50[10] 145[8])
    defparam i16114_4_lut.LUT_INIT = 16'hccca;
    SB_DFFESR GHA_188 (.Q(GHA), .C(clk16MHz), .E(n27585), .D(GHA_N_355), 
            .R(n28807));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    SB_DFFESS commutation_state_i0 (.Q(commutation_state[0]), .C(clk16MHz), 
            .E(n7_adj_5959), .D(commutation_state_7__N_208[0]), .S(commutation_state_7__N_216));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    SB_DFFESR GLA_189 (.Q(INLA_c_0), .C(clk16MHz), .E(n27585), .D(GLA_N_372), 
            .R(n28807));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    SB_DFF displacement_i22 (.Q(displacement[22]), .C(clk16MHz), .D(displacement_23__N_67[22]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1901 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[14] [6]), 
            .O(n58574));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1901.LUT_INIT = 16'h2300;
    SB_DFFESR GLB_191 (.Q(INLB_c_0), .C(clk16MHz), .E(n27585), .D(GLB_N_386), 
            .R(n28807));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    SB_DFF displacement_i21 (.Q(displacement[21]), .C(clk16MHz), .D(displacement_23__N_67[21]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_CARRY encoder0_position_30__I_0_add_1436_7 (.CI(n51595), .I0(n2129), 
            .I1(GND_net), .CO(n51596));
    SB_DFFESR GLC_193 (.Q(INLC_c_0), .C(clk16MHz), .E(n27585), .D(GLC_N_400), 
            .R(n28807));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1902 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[14] [7]), 
            .O(n58573));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1902.LUT_INIT = 16'h2300;
    SB_DFF displacement_i20 (.Q(displacement[20]), .C(clk16MHz), .D(displacement_23__N_67[20]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF displacement_i19 (.Q(displacement[19]), .C(clk16MHz), .D(displacement_23__N_67[19]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF displacement_i18 (.Q(displacement[18]), .C(clk16MHz), .D(displacement_23__N_67[18]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF displacement_i17 (.Q(displacement[17]), .C(clk16MHz), .D(displacement_23__N_67[17]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF displacement_i16 (.Q(displacement[16]), .C(clk16MHz), .D(displacement_23__N_67[16]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF displacement_i15 (.Q(displacement[15]), .C(clk16MHz), .D(displacement_23__N_67[15]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF displacement_i14 (.Q(displacement[14]), .C(clk16MHz), .D(displacement_23__N_67[14]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF displacement_i13 (.Q(displacement[13]), .C(clk16MHz), .D(displacement_23__N_67[13]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF displacement_i12 (.Q(displacement[12]), .C(clk16MHz), .D(displacement_23__N_67[12]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF displacement_i11 (.Q(displacement[11]), .C(clk16MHz), .D(displacement_23__N_67[11]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF displacement_i10 (.Q(displacement[10]), .C(clk16MHz), .D(displacement_23__N_67[10]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF displacement_i9 (.Q(displacement[9]), .C(clk16MHz), .D(displacement_23__N_67[9]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF displacement_i8 (.Q(displacement[8]), .C(clk16MHz), .D(displacement_23__N_67[8]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF displacement_i7 (.Q(displacement[7]), .C(clk16MHz), .D(displacement_23__N_67[7]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF displacement_i6 (.Q(displacement[6]), .C(clk16MHz), .D(displacement_23__N_67[6]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF displacement_i5 (.Q(displacement[5]), .C(clk16MHz), .D(displacement_23__N_67[5]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF displacement_i4 (.Q(displacement[4]), .C(clk16MHz), .D(displacement_23__N_67[4]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF displacement_i3 (.Q(displacement[3]), .C(clk16MHz), .D(displacement_23__N_67[3]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF displacement_i2 (.Q(displacement[2]), .C(clk16MHz), .D(displacement_23__N_67[2]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF displacement_i1 (.Q(displacement[1]), .C(clk16MHz), .D(displacement_23__N_67[1]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF encoder1_position_scaled_i23 (.Q(encoder1_position_scaled[23]), 
           .C(clk16MHz), .D(encoder1_position[25]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF encoder1_position_scaled_i22 (.Q(encoder1_position_scaled[22]), 
           .C(clk16MHz), .D(encoder1_position[24]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF encoder1_position_scaled_i21 (.Q(encoder1_position_scaled[21]), 
           .C(clk16MHz), .D(encoder1_position[23]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF encoder1_position_scaled_i20 (.Q(encoder1_position_scaled[20]), 
           .C(clk16MHz), .D(encoder1_position[22]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF encoder1_position_scaled_i19 (.Q(encoder1_position_scaled[19]), 
           .C(clk16MHz), .D(encoder1_position[21]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF encoder1_position_scaled_i18 (.Q(encoder1_position_scaled[18]), 
           .C(clk16MHz), .D(encoder1_position[20]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF encoder1_position_scaled_i17 (.Q(encoder1_position_scaled[17]), 
           .C(clk16MHz), .D(encoder1_position[19]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF encoder1_position_scaled_i16 (.Q(encoder1_position_scaled[16]), 
           .C(clk16MHz), .D(encoder1_position[18]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF commutation_state_prev_i0 (.Q(commutation_state_prev[0]), .C(clk16MHz), 
           .D(commutation_state[0]));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    SB_DFF encoder1_position_scaled_i15 (.Q(encoder1_position_scaled[15]), 
           .C(clk16MHz), .D(encoder1_position[17]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF encoder1_position_scaled_i14 (.Q(encoder1_position_scaled[14]), 
           .C(clk16MHz), .D(encoder1_position[16]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF encoder1_position_scaled_i13 (.Q(encoder1_position_scaled[13]), 
           .C(clk16MHz), .D(encoder1_position[15]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF encoder1_position_scaled_i12 (.Q(encoder1_position_scaled[12]), 
           .C(clk16MHz), .D(encoder1_position[14]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF encoder1_position_scaled_i11 (.Q(encoder1_position_scaled[11]), 
           .C(clk16MHz), .D(encoder1_position[13]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF encoder1_position_scaled_i10 (.Q(encoder1_position_scaled[10]), 
           .C(clk16MHz), .D(encoder1_position[12]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF encoder1_position_scaled_i9 (.Q(encoder1_position_scaled[9]), .C(clk16MHz), 
           .D(encoder1_position[11]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF encoder1_position_scaled_i8 (.Q(encoder1_position_scaled[8]), .C(clk16MHz), 
           .D(encoder1_position[10]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF encoder1_position_scaled_i7 (.Q(encoder1_position_scaled[7]), .C(clk16MHz), 
           .D(encoder1_position[9]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF encoder1_position_scaled_i6 (.Q(encoder1_position_scaled[6]), .C(clk16MHz), 
           .D(encoder1_position[8]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF encoder1_position_scaled_i5 (.Q(encoder1_position_scaled[5]), .C(clk16MHz), 
           .D(encoder1_position[7]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF encoder1_position_scaled_i4 (.Q(encoder1_position_scaled[4]), .C(clk16MHz), 
           .D(encoder1_position[6]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF encoder1_position_scaled_i3 (.Q(encoder1_position_scaled[3]), .C(clk16MHz), 
           .D(encoder1_position[5]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF encoder1_position_scaled_i2 (.Q(encoder1_position_scaled[2]), .C(clk16MHz), 
           .D(encoder1_position[4]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF encoder1_position_scaled_i1 (.Q(encoder1_position_scaled[1]), .C(clk16MHz), 
           .D(encoder1_position[3]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    GND i1 (.Y(GND_net));
    SB_CARRY encoder0_position_30__I_0_add_1905_23 (.CI(n51837), .I0(n2813), 
            .I1(VCC_net), .CO(n51838));
    SB_CARRY encoder0_position_30__I_0_add_967_2 (.CI(VCC_net), .I0(n939), 
            .I1(GND_net), .CO(n51353));
    SB_CARRY encoder0_position_30__I_0_add_2173_11 (.CI(n51935), .I0(n3226), 
            .I1(VCC_net), .CO(n51936));
    SB_LUT4 encoder0_position_30__I_0_add_1704_6_lut (.I0(GND_net), .I1(n2530), 
            .I2(GND_net), .I3(n51748), .O(n2597)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1704_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1704_6 (.CI(n51748), .I0(n2530), 
            .I1(GND_net), .CO(n51749));
    SB_LUT4 encoder0_position_30__I_0_add_1436_6_lut (.I0(GND_net), .I1(n2130), 
            .I2(GND_net), .I3(n51594), .O(n2197)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1436_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1704_5_lut (.I0(GND_net), .I1(n2531), 
            .I2(VCC_net), .I3(n51747), .O(n2598)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1704_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1095_15 (.CI(n51107), .I0(GND_net), .I1(n12187), .CO(n51108));
    SB_LUT4 encoder0_position_30__I_0_add_1905_22_lut (.I0(GND_net), .I1(n2814), 
            .I2(VCC_net), .I3(n51836), .O(n2881)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1905_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1905_22 (.CI(n51836), .I0(n2814), 
            .I1(VCC_net), .CO(n51837));
    SB_LUT4 add_1095_14_lut (.I0(GND_net), .I1(GND_net), .I2(n12189), 
            .I3(n51106), .O(n4914)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1095_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1905_21_lut (.I0(GND_net), .I1(n2815), 
            .I2(VCC_net), .I3(n51835), .O(n2882)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1905_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1905_21 (.CI(n51835), .I0(n2815), 
            .I1(VCC_net), .CO(n51836));
    SB_CARRY encoder0_position_30__I_0_add_1436_6 (.CI(n51594), .I0(n2130), 
            .I1(GND_net), .CO(n51595));
    SB_LUT4 add_151_20_lut (.I0(GND_net), .I1(delay_counter[18]), .I2(GND_net), 
            .I3(n50995), .O(n1221)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1436_5_lut (.I0(GND_net), .I1(n2131), 
            .I2(VCC_net), .I3(n51593), .O(n2198)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1436_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1436_5 (.CI(n51593), .I0(n2131), 
            .I1(VCC_net), .CO(n51594));
    SB_LUT4 encoder0_position_30__I_0_i1842_3_lut (.I0(n2711), .I1(n2778), 
            .I2(n2742), .I3(GND_net), .O(n2810));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1842_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_1095_14 (.CI(n51106), .I0(GND_net), .I1(n12189), .CO(n51107));
    SB_CARRY encoder0_position_30__I_0_add_1704_5 (.CI(n51747), .I0(n2531), 
            .I1(VCC_net), .CO(n51748));
    SB_LUT4 encoder0_position_30__I_0_add_2173_10_lut (.I0(GND_net), .I1(n3227), 
            .I2(VCC_net), .I3(n51934), .O(n3294)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2173_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1903 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[15] [0]), 
            .O(n28959));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1903.LUT_INIT = 16'h2300;
    SB_LUT4 add_1095_13_lut (.I0(GND_net), .I1(GND_net), .I2(n12191), 
            .I3(n51105), .O(n4915)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1095_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1095_13 (.CI(n51105), .I0(GND_net), .I1(n12191), .CO(n51106));
    SB_CARRY encoder0_position_30__I_0_add_2173_10 (.CI(n51934), .I0(n3227), 
            .I1(VCC_net), .CO(n51935));
    SB_LUT4 encoder0_position_30__I_0_add_1436_4_lut (.I0(GND_net), .I1(n2132), 
            .I2(GND_net), .I3(n51592), .O(n2199)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1436_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1436_4 (.CI(n51592), .I0(n2132), 
            .I1(GND_net), .CO(n51593));
    SB_LUT4 encoder0_position_30__I_0_add_1704_4_lut (.I0(GND_net), .I1(n2532), 
            .I2(GND_net), .I3(n51746), .O(n2599)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1704_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1905_20_lut (.I0(GND_net), .I1(n2816), 
            .I2(VCC_net), .I3(n51834), .O(n2883)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1905_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1905_20 (.CI(n51834), .I0(n2816), 
            .I1(VCC_net), .CO(n51835));
    SB_LUT4 encoder0_position_30__I_0_add_2173_9_lut (.I0(GND_net), .I1(n3228), 
            .I2(VCC_net), .I3(n51933), .O(n3295)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2173_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1704_4 (.CI(n51746), .I0(n2532), 
            .I1(GND_net), .CO(n51747));
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1904 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[15] [1]), 
            .O(n58572));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1904.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_add_1704_3_lut (.I0(GND_net), .I1(n2533), 
            .I2(VCC_net), .I3(n51745), .O(n2600)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1704_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1905_19_lut (.I0(GND_net), .I1(n2817), 
            .I2(VCC_net), .I3(n51833), .O(n2884)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1905_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1905 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[15] [2]), 
            .O(n58571));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1905.LUT_INIT = 16'h2300;
    SB_CARRY add_151_20 (.CI(n50995), .I0(delay_counter[18]), .I1(GND_net), 
            .CO(n50996));
    SB_CARRY encoder0_position_30__I_0_add_2173_9 (.CI(n51933), .I0(n3228), 
            .I1(VCC_net), .CO(n51934));
    SB_CARRY encoder0_position_30__I_0_add_1905_19 (.CI(n51833), .I0(n2817), 
            .I1(VCC_net), .CO(n51834));
    SB_LUT4 encoder0_position_30__I_0_add_1905_18_lut (.I0(GND_net), .I1(n2818), 
            .I2(VCC_net), .I3(n51832), .O(n2885)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1905_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1436_3_lut (.I0(GND_net), .I1(n2133), 
            .I2(VCC_net), .I3(n51591), .O(n2200)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1436_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1704_3 (.CI(n51745), .I0(n2533), 
            .I1(VCC_net), .CO(n51746));
    SB_LUT4 encoder0_position_30__I_0_add_1704_2_lut (.I0(GND_net), .I1(n950), 
            .I2(GND_net), .I3(VCC_net), .O(n2601)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1704_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1436_3 (.CI(n51591), .I0(n2133), 
            .I1(VCC_net), .CO(n51592));
    SB_CARRY encoder0_position_30__I_0_add_1905_18 (.CI(n51832), .I0(n2818), 
            .I1(VCC_net), .CO(n51833));
    SB_LUT4 encoder0_position_30__I_0_add_1905_17_lut (.I0(GND_net), .I1(n2819), 
            .I2(VCC_net), .I3(n51831), .O(n2886)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1905_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1906 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[15] [3]), 
            .O(n58570));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1906.LUT_INIT = 16'h2300;
    SB_LUT4 i1_4_lut_adj_1907 (.I0(o_Rx_DV_N_3488[12]), .I1(n4935), .I2(o_Rx_DV_N_3488[8]), 
            .I3(n62433), .O(n62439));
    defparam i1_4_lut_adj_1907.LUT_INIT = 16'hfffe;
    SB_CARRY encoder0_position_30__I_0_add_1704_2 (.CI(VCC_net), .I0(n950), 
            .I1(GND_net), .CO(n51745));
    SB_LUT4 encoder0_position_30__I_0_add_2173_8_lut (.I0(GND_net), .I1(n3229), 
            .I2(GND_net), .I3(n51932), .O(n3296)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2173_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1905_17 (.CI(n51831), .I0(n2819), 
            .I1(VCC_net), .CO(n51832));
    SB_LUT4 encoder0_position_30__I_0_add_1905_16_lut (.I0(GND_net), .I1(n2820_adj_5856), 
            .I2(VCC_net), .I3(n51830), .O(n2887)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1905_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1637_24_lut (.I0(n70337), .I1(n2412), 
            .I2(VCC_net), .I3(n51744), .O(n2511)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1637_24_lut.LUT_INIT = 16'h8228;
    SB_CARRY encoder0_position_30__I_0_add_2173_8 (.CI(n51932), .I0(n3229), 
            .I1(GND_net), .CO(n51933));
    SB_LUT4 encoder0_position_30__I_0_add_2173_7_lut (.I0(n3298), .I1(n3230), 
            .I2(GND_net), .I3(n51931), .O(n67092)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2173_7_lut.LUT_INIT = 16'h8228;
    SB_CARRY encoder0_position_30__I_0_add_2173_7 (.CI(n51931), .I0(n3230), 
            .I1(GND_net), .CO(n51932));
    SB_LUT4 encoder0_position_30__I_0_add_1637_23_lut (.I0(GND_net), .I1(n2413), 
            .I2(VCC_net), .I3(n51743), .O(n2480)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1637_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1436_2_lut (.I0(GND_net), .I1(n946), 
            .I2(GND_net), .I3(VCC_net), .O(n2201)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1436_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1908 (.I0(o_Rx_DV_N_3488[24]), .I1(n29_adj_5857), 
            .I2(n23_adj_5860), .I3(n62439), .O(n62445));
    defparam i1_4_lut_adj_1908.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_30__I_0_add_2173_6_lut (.I0(GND_net), .I1(n3231), 
            .I2(VCC_net), .I3(n51930), .O(n3298)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2173_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_1095_12_lut (.I0(GND_net), .I1(GND_net), .I2(n12193), 
            .I3(n51104), .O(n4916)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1095_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2173_6 (.CI(n51930), .I0(n3231), 
            .I1(VCC_net), .CO(n51931));
    SB_CARRY encoder0_position_30__I_0_add_1905_16 (.CI(n51830), .I0(n2820_adj_5856), 
            .I1(VCC_net), .CO(n51831));
    SB_LUT4 encoder0_position_30__I_0_add_1905_15_lut (.I0(GND_net), .I1(n2821), 
            .I2(VCC_net), .I3(n51829), .O(n2888)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1905_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1095_12 (.CI(n51104), .I0(GND_net), .I1(n12193), .CO(n51105));
    SB_CARRY encoder0_position_30__I_0_add_1637_23 (.CI(n51743), .I0(n2413), 
            .I1(VCC_net), .CO(n51744));
    SB_LUT4 add_1095_11_lut (.I0(GND_net), .I1(GND_net), .I2(n12195), 
            .I3(n51103), .O(n4917)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1095_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1905_15 (.CI(n51829), .I0(n2821), 
            .I1(VCC_net), .CO(n51830));
    SB_LUT4 encoder0_position_30__I_0_add_1637_22_lut (.I0(GND_net), .I1(n2414), 
            .I2(VCC_net), .I3(n51742), .O(n2481)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1637_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1436_2 (.CI(VCC_net), .I0(n946), 
            .I1(GND_net), .CO(n51591));
    SB_CARRY add_1095_11 (.CI(n51103), .I0(GND_net), .I1(n12195), .CO(n51104));
    SB_LUT4 encoder0_position_30__I_0_add_2173_5_lut (.I0(n6_adj_5923), .I1(n3232), 
            .I2(GND_net), .I3(n51929), .O(n67087)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2173_5_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 i16115_4_lut (.I0(r_Rx_Data), .I1(rx_data[2]), .I2(n62445), 
            .I3(n27_adj_5858), .O(n30121));   // verilog/uart_rx.v(50[10] 145[8])
    defparam i16115_4_lut.LUT_INIT = 16'hccca;
    SB_CARRY encoder0_position_30__I_0_add_1637_22 (.CI(n51742), .I0(n2414), 
            .I1(VCC_net), .CO(n51743));
    SB_LUT4 encoder0_position_30__I_0_add_1637_21_lut (.I0(GND_net), .I1(n2415), 
            .I2(VCC_net), .I3(n51741), .O(n2482)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1637_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2173_5 (.CI(n51929), .I0(n3232), 
            .I1(GND_net), .CO(n51930));
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1909 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[15] [4]), 
            .O(n58569));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1909.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1910 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[15] [5]), 
            .O(n58568));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1910.LUT_INIT = 16'h2300;
    SB_LUT4 add_1095_10_lut (.I0(GND_net), .I1(GND_net), .I2(n12197), 
            .I3(n51102), .O(n4918)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1095_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_2173_4_lut (.I0(n3301), .I1(n3233), 
            .I2(VCC_net), .I3(n51928), .O(n6_adj_5923)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2173_4_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_1095_10 (.CI(n51102), .I0(GND_net), .I1(n12197), .CO(n51103));
    SB_CARRY encoder0_position_30__I_0_add_2173_4 (.CI(n51928), .I0(n3233), 
            .I1(VCC_net), .CO(n51929));
    SB_CARRY encoder0_position_30__I_0_add_1637_21 (.CI(n51741), .I0(n2415), 
            .I1(VCC_net), .CO(n51742));
    SB_LUT4 add_151_19_lut (.I0(GND_net), .I1(delay_counter[17]), .I2(GND_net), 
            .I3(n50994), .O(n1222)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1905_14_lut (.I0(GND_net), .I1(n2822), 
            .I2(VCC_net), .I3(n51828), .O(n2889)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1905_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1911 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[15] [6]), 
            .O(n58567));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1911.LUT_INIT = 16'h2300;
    SB_LUT4 add_1095_9_lut (.I0(GND_net), .I1(GND_net), .I2(n12199), .I3(n51101), 
            .O(n4919)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1095_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1912 (.I0(o_Rx_DV_N_3488[12]), .I1(n4935), .I2(o_Rx_DV_N_3488[8]), 
            .I3(n62481), .O(n62487));
    defparam i1_4_lut_adj_1912.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_30__I_0_add_2173_3_lut (.I0(GND_net), .I1(n957), 
            .I2(GND_net), .I3(n51927), .O(n3301)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2173_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1095_9 (.CI(n51101), .I0(GND_net), .I1(n12199), .CO(n51102));
    SB_LUT4 encoder0_position_30__I_0_add_1637_20_lut (.I0(GND_net), .I1(n2416), 
            .I2(VCC_net), .I3(n51740), .O(n2483)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1637_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_1095_8_lut (.I0(GND_net), .I1(GND_net), .I2(n12201), .I3(n51100), 
            .O(n4920)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1095_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2173_3 (.CI(n51927), .I0(n957), 
            .I1(GND_net), .CO(n51928));
    SB_CARRY encoder0_position_30__I_0_add_1637_20 (.CI(n51740), .I0(n2416), 
            .I1(VCC_net), .CO(n51741));
    SB_CARRY add_1095_8 (.CI(n51100), .I0(GND_net), .I1(n12201), .CO(n51101));
    SB_CARRY encoder0_position_30__I_0_add_2173_2 (.CI(VCC_net), .I0(GND_net), 
            .I1(VCC_net), .CO(n51927));
    SB_CARRY add_151_19 (.CI(n50994), .I0(delay_counter[17]), .I1(GND_net), 
            .CO(n50995));
    SB_LUT4 encoder0_position_30__I_0_add_2106_31_lut (.I0(n70202), .I1(n3105), 
            .I2(VCC_net), .I3(n51926), .O(n3204)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2106_31_lut.LUT_INIT = 16'h8228;
    SB_CARRY encoder0_position_30__I_0_add_1905_14 (.CI(n51828), .I0(n2822), 
            .I1(VCC_net), .CO(n51829));
    SB_LUT4 encoder0_position_30__I_0_add_1637_19_lut (.I0(GND_net), .I1(n2417), 
            .I2(VCC_net), .I3(n51739), .O(n2484)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1637_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1913 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[15] [7]), 
            .O(n58566));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1913.LUT_INIT = 16'h2300;
    SB_CARRY encoder0_position_30__I_0_add_1637_19 (.CI(n51739), .I0(n2417), 
            .I1(VCC_net), .CO(n51740));
    SB_LUT4 encoder0_position_30__I_0_add_2106_30_lut (.I0(GND_net), .I1(n3106), 
            .I2(VCC_net), .I3(n51925), .O(n3173)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2106_30_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1637_18_lut (.I0(GND_net), .I1(n2418), 
            .I2(VCC_net), .I3(n51738), .O(n2485)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1637_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2106_30 (.CI(n51925), .I0(n3106), 
            .I1(VCC_net), .CO(n51926));
    SB_LUT4 encoder0_position_30__I_0_add_1905_13_lut (.I0(GND_net), .I1(n2823), 
            .I2(VCC_net), .I3(n51827), .O(n2890)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1905_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_2106_29_lut (.I0(GND_net), .I1(n3107), 
            .I2(VCC_net), .I3(n51924), .O(n3174)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2106_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1905_13 (.CI(n51827), .I0(n2823), 
            .I1(VCC_net), .CO(n51828));
    SB_LUT4 encoder0_position_30__I_0_add_1905_12_lut (.I0(GND_net), .I1(n2824), 
            .I2(VCC_net), .I3(n51826), .O(n2891)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1905_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2106_29 (.CI(n51924), .I0(n3107), 
            .I1(VCC_net), .CO(n51925));
    SB_CARRY encoder0_position_30__I_0_add_1905_12 (.CI(n51826), .I0(n2824), 
            .I1(VCC_net), .CO(n51827));
    SB_LUT4 encoder0_position_30__I_0_add_2106_28_lut (.I0(GND_net), .I1(n3108), 
            .I2(VCC_net), .I3(n51923), .O(n3175)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2106_28_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_1095_7_lut (.I0(GND_net), .I1(GND_net), .I2(n12203), .I3(n51099), 
            .O(n4921)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1095_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2106_28 (.CI(n51923), .I0(n3108), 
            .I1(VCC_net), .CO(n51924));
    SB_LUT4 encoder0_position_30__I_0_add_1905_11_lut (.I0(GND_net), .I1(n2825), 
            .I2(VCC_net), .I3(n51825), .O(n2892)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1905_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_i1320_3_lut (.I0(n1933), .I1(n2000), 
            .I2(n1950), .I3(GND_net), .O(n2032));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1320_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_1095_7 (.CI(n51099), .I0(GND_net), .I1(n12203), .CO(n51100));
    SB_LUT4 i1_4_lut_adj_1914 (.I0(o_Rx_DV_N_3488[24]), .I1(n29_adj_5857), 
            .I2(n23_adj_5860), .I3(n62487), .O(n62493));
    defparam i1_4_lut_adj_1914.LUT_INIT = 16'hfffe;
    SB_LUT4 add_151_18_lut (.I0(GND_net), .I1(delay_counter[16]), .I2(GND_net), 
            .I3(n50993), .O(n1223)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_1095_6_lut (.I0(GND_net), .I1(GND_net), .I2(n12205), .I3(n51098), 
            .O(n4922)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1095_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_2106_27_lut (.I0(GND_net), .I1(n3109), 
            .I2(VCC_net), .I3(n51922), .O(n3176)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2106_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1905_11 (.CI(n51825), .I0(n2825), 
            .I1(VCC_net), .CO(n51826));
    SB_LUT4 encoder0_position_30__I_0_add_1905_10_lut (.I0(GND_net), .I1(n2826), 
            .I2(VCC_net), .I3(n51824), .O(n2893)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1905_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1095_6 (.CI(n51098), .I0(GND_net), .I1(n12205), .CO(n51099));
    SB_CARRY encoder0_position_30__I_0_add_1637_18 (.CI(n51738), .I0(n2418), 
            .I1(VCC_net), .CO(n51739));
    SB_LUT4 encoder0_position_30__I_0_add_1503_22_lut (.I0(n70528), .I1(n2214), 
            .I2(VCC_net), .I3(n51670), .O(n2313)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1503_22_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_151_18 (.CI(n50993), .I0(delay_counter[16]), .I1(GND_net), 
            .CO(n50994));
    SB_LUT4 add_1095_5_lut (.I0(GND_net), .I1(GND_net), .I2(n12207), .I3(n51097), 
            .O(n4923)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1095_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2106_27 (.CI(n51922), .I0(n3109), 
            .I1(VCC_net), .CO(n51923));
    SB_CARRY encoder0_position_30__I_0_add_1905_10 (.CI(n51824), .I0(n2826), 
            .I1(VCC_net), .CO(n51825));
    SB_LUT4 encoder0_position_30__I_0_add_1905_9_lut (.I0(GND_net), .I1(n2827), 
            .I2(VCC_net), .I3(n51823), .O(n2894)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1905_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_2106_26_lut (.I0(GND_net), .I1(n3110), 
            .I2(VCC_net), .I3(n51921), .O(n3177)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2106_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_900_13_lut (.I0(n70743), .I1(n1323), 
            .I2(VCC_net), .I3(n51335), .O(n1422)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_900_13_lut.LUT_INIT = 16'h8228;
    SB_LUT4 add_151_9_lut (.I0(GND_net), .I1(delay_counter[7]), .I2(GND_net), 
            .I3(n50984), .O(n1232)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1637_17_lut (.I0(GND_net), .I1(n2419), 
            .I2(VCC_net), .I3(n51737), .O(n2486)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1637_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_900_12_lut (.I0(GND_net), .I1(n1324), 
            .I2(VCC_net), .I3(n51334), .O(n1391)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_900_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_900_12 (.CI(n51334), .I0(n1324), 
            .I1(VCC_net), .CO(n51335));
    SB_CARRY encoder0_position_30__I_0_add_1905_9 (.CI(n51823), .I0(n2827), 
            .I1(VCC_net), .CO(n51824));
    SB_CARRY encoder0_position_30__I_0_add_2106_26 (.CI(n51921), .I0(n3110), 
            .I1(VCC_net), .CO(n51922));
    SB_LUT4 encoder0_position_30__I_0_add_2106_25_lut (.I0(GND_net), .I1(n3111), 
            .I2(VCC_net), .I3(n51920), .O(n3178)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2106_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2106_25 (.CI(n51920), .I0(n3111), 
            .I1(VCC_net), .CO(n51921));
    SB_LUT4 encoder0_position_30__I_0_add_900_11_lut (.I0(GND_net), .I1(n1325), 
            .I2(VCC_net), .I3(n51333), .O(n1392)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_900_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_900_11 (.CI(n51333), .I0(n1325), 
            .I1(VCC_net), .CO(n51334));
    SB_LUT4 encoder0_position_30__I_0_add_900_10_lut (.I0(GND_net), .I1(n1326), 
            .I2(VCC_net), .I3(n51332), .O(n1393)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_900_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_900_10 (.CI(n51332), .I0(n1326), 
            .I1(VCC_net), .CO(n51333));
    SB_LUT4 encoder0_position_30__I_0_add_2106_24_lut (.I0(GND_net), .I1(n3112), 
            .I2(VCC_net), .I3(n51919), .O(n3179)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2106_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1905_8_lut (.I0(GND_net), .I1(n2828), 
            .I2(VCC_net), .I3(n51822), .O(n2895)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1905_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i16116_4_lut (.I0(r_Rx_Data), .I1(rx_data[3]), .I2(n62493), 
            .I3(n27_adj_5858), .O(n30122));   // verilog/uart_rx.v(50[10] 145[8])
    defparam i16116_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 add_151_17_lut (.I0(GND_net), .I1(delay_counter[15]), .I2(GND_net), 
            .I3(n50992), .O(n1224)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1095_5 (.CI(n51097), .I0(GND_net), .I1(n12207), .CO(n51098));
    SB_CARRY encoder0_position_30__I_0_add_2106_24 (.CI(n51919), .I0(n3112), 
            .I1(VCC_net), .CO(n51920));
    SB_CARRY encoder0_position_30__I_0_add_1637_17 (.CI(n51737), .I0(n2419), 
            .I1(VCC_net), .CO(n51738));
    SB_LUT4 encoder0_position_30__I_0_add_900_9_lut (.I0(GND_net), .I1(n1327), 
            .I2(VCC_net), .I3(n51331), .O(n1394)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_900_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_2106_23_lut (.I0(GND_net), .I1(n3113), 
            .I2(VCC_net), .I3(n51918), .O(n3180)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2106_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1503_21_lut (.I0(GND_net), .I1(n2215), 
            .I2(VCC_net), .I3(n51669), .O(n2282)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1503_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_1095_4_lut (.I0(GND_net), .I1(GND_net), .I2(n12209), .I3(n51096), 
            .O(n4924)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1095_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1503_21 (.CI(n51669), .I0(n2215), 
            .I1(VCC_net), .CO(n51670));
    SB_CARRY encoder0_position_30__I_0_add_1905_8 (.CI(n51822), .I0(n2828), 
            .I1(VCC_net), .CO(n51823));
    SB_LUT4 encoder0_position_30__I_0_add_1637_16_lut (.I0(GND_net), .I1(n2420), 
            .I2(VCC_net), .I3(n51736), .O(n2487)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1637_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1637_16 (.CI(n51736), .I0(n2420), 
            .I1(VCC_net), .CO(n51737));
    SB_LUT4 encoder0_position_30__I_0_add_1503_20_lut (.I0(GND_net), .I1(n2216), 
            .I2(VCC_net), .I3(n51668), .O(n2283)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1503_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1637_15_lut (.I0(GND_net), .I1(n2421), 
            .I2(VCC_net), .I3(n51735), .O(n2488)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1637_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1095_4 (.CI(n51096), .I0(GND_net), .I1(n12209), .CO(n51097));
    SB_CARRY encoder0_position_30__I_0_add_1503_20 (.CI(n51668), .I0(n2216), 
            .I1(VCC_net), .CO(n51669));
    SB_LUT4 encoder0_position_30__I_0_add_1905_7_lut (.I0(GND_net), .I1(n2829), 
            .I2(GND_net), .I3(n51821), .O(n2896)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1905_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1503_19_lut (.I0(GND_net), .I1(n2217_adj_5853), 
            .I2(VCC_net), .I3(n51667), .O(n2284)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1503_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_1095_3_lut (.I0(GND_net), .I1(GND_net), .I2(n12211), .I3(n51095), 
            .O(n4925)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1095_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_900_9 (.CI(n51331), .I0(n1327), 
            .I1(VCC_net), .CO(n51332));
    SB_LUT4 encoder0_position_30__I_0_add_900_8_lut (.I0(GND_net), .I1(n1328), 
            .I2(VCC_net), .I3(n51330), .O(n1395)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_900_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1637_15 (.CI(n51735), .I0(n2421), 
            .I1(VCC_net), .CO(n51736));
    SB_CARRY encoder0_position_30__I_0_add_900_8 (.CI(n51330), .I0(n1328), 
            .I1(VCC_net), .CO(n51331));
    SB_LUT4 encoder0_position_30__I_0_add_1637_14_lut (.I0(GND_net), .I1(n2422), 
            .I2(VCC_net), .I3(n51734), .O(n2489)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1637_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1503_19 (.CI(n51667), .I0(n2217_adj_5853), 
            .I1(VCC_net), .CO(n51668));
    SB_CARRY encoder0_position_30__I_0_add_1905_7 (.CI(n51821), .I0(n2829), 
            .I1(GND_net), .CO(n51822));
    SB_LUT4 encoder0_position_30__I_0_add_1503_18_lut (.I0(GND_net), .I1(n2218), 
            .I2(VCC_net), .I3(n51666), .O(n2285)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1503_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1503_18 (.CI(n51666), .I0(n2218), 
            .I1(VCC_net), .CO(n51667));
    SB_LUT4 encoder0_position_30__I_0_add_900_7_lut (.I0(GND_net), .I1(n1329), 
            .I2(GND_net), .I3(n51329), .O(n1396)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_900_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1905_6_lut (.I0(GND_net), .I1(n2830), 
            .I2(GND_net), .I3(n51820), .O(n2897)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1905_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1637_14 (.CI(n51734), .I0(n2422), 
            .I1(VCC_net), .CO(n51735));
    SB_LUT4 encoder0_position_30__I_0_add_1637_13_lut (.I0(GND_net), .I1(n2423), 
            .I2(VCC_net), .I3(n51733), .O(n2490)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1637_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1637_13 (.CI(n51733), .I0(n2423), 
            .I1(VCC_net), .CO(n51734));
    SB_CARRY encoder0_position_30__I_0_add_1905_6 (.CI(n51820), .I0(n2830), 
            .I1(GND_net), .CO(n51821));
    SB_LUT4 encoder0_position_30__I_0_add_1905_5_lut (.I0(GND_net), .I1(n2831), 
            .I2(VCC_net), .I3(n51819), .O(n2898)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1905_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1637_12_lut (.I0(GND_net), .I1(n2424), 
            .I2(VCC_net), .I3(n51732), .O(n2491)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1637_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_900_7 (.CI(n51329), .I0(n1329), 
            .I1(GND_net), .CO(n51330));
    SB_LUT4 encoder0_position_30__I_0_add_1503_17_lut (.I0(GND_net), .I1(n2219), 
            .I2(VCC_net), .I3(n51665), .O(n2286)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1503_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1637_12 (.CI(n51732), .I0(n2424), 
            .I1(VCC_net), .CO(n51733));
    SB_LUT4 encoder0_position_30__I_0_add_900_6_lut (.I0(GND_net), .I1(n1330), 
            .I2(GND_net), .I3(n51328), .O(n1397)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_900_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1503_17 (.CI(n51665), .I0(n2219), 
            .I1(VCC_net), .CO(n51666));
    SB_CARRY encoder0_position_30__I_0_add_900_6 (.CI(n51328), .I0(n1330), 
            .I1(GND_net), .CO(n51329));
    SB_LUT4 encoder0_position_30__I_0_add_1168_17_lut (.I0(n70635), .I1(n1719), 
            .I2(VCC_net), .I3(n51454), .O(n1818)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1168_17_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_30__I_0_add_900_5_lut (.I0(GND_net), .I1(n1331), 
            .I2(VCC_net), .I3(n51327), .O(n1398)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_900_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i12_2_lut (.I0(pwm_counter[12]), .I1(pwm_setpoint[12]), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_5864));   // verilog/TinyFPGA_B.v(95[20:32])
    defparam i12_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY encoder0_position_30__I_0_add_900_5 (.CI(n51327), .I0(n1331), 
            .I1(VCC_net), .CO(n51328));
    SB_LUT4 encoder0_position_30__I_0_add_1168_16_lut (.I0(GND_net), .I1(n1720), 
            .I2(VCC_net), .I3(n51453), .O(n1787)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1168_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1168_16 (.CI(n51453), .I0(n1720), 
            .I1(VCC_net), .CO(n51454));
    SB_LUT4 encoder0_position_30__I_0_add_1168_15_lut (.I0(GND_net), .I1(n1721), 
            .I2(VCC_net), .I3(n51452), .O(n1788_adj_5846)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1168_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1503_16_lut (.I0(GND_net), .I1(n2220), 
            .I2(VCC_net), .I3(n51664), .O(n2287)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1503_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1503_16 (.CI(n51664), .I0(n2220), 
            .I1(VCC_net), .CO(n51665));
    SB_LUT4 encoder0_position_30__I_0_add_900_4_lut (.I0(GND_net), .I1(n1332), 
            .I2(GND_net), .I3(n51326), .O(n1399)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_900_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_900_4 (.CI(n51326), .I0(n1332), 
            .I1(GND_net), .CO(n51327));
    SB_LUT4 encoder0_position_30__I_0_add_1503_15_lut (.I0(GND_net), .I1(n2221), 
            .I2(VCC_net), .I3(n51663), .O(n2288)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1503_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1095_3 (.CI(n51095), .I0(GND_net), .I1(n12211), .CO(n51096));
    SB_LUT4 encoder0_position_30__I_0_add_1637_11_lut (.I0(GND_net), .I1(n2425), 
            .I2(VCC_net), .I3(n51731), .O(n2492)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1637_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1637_11 (.CI(n51731), .I0(n2425), 
            .I1(VCC_net), .CO(n51732));
    SB_LUT4 encoder0_position_30__I_0_add_900_3_lut (.I0(GND_net), .I1(n1333), 
            .I2(VCC_net), .I3(n51325), .O(n1400)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_900_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_1095_2_lut (.I0(GND_net), .I1(GND_net), .I2(n7_adj_5826), 
            .I3(VCC_net), .O(n4926)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1095_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1095_2 (.CI(VCC_net), .I0(GND_net), .I1(n7_adj_5826), 
            .CO(n51095));
    SB_CARRY encoder0_position_30__I_0_add_1503_15 (.CI(n51663), .I0(n2221), 
            .I1(VCC_net), .CO(n51664));
    SB_CARRY encoder0_position_30__I_0_add_900_3 (.CI(n51325), .I0(n1333), 
            .I1(VCC_net), .CO(n51326));
    SB_CARRY encoder0_position_30__I_0_add_1168_15 (.CI(n51452), .I0(n1721), 
            .I1(VCC_net), .CO(n51453));
    SB_LUT4 encoder0_position_30__I_0_add_900_2_lut (.I0(GND_net), .I1(n938), 
            .I2(GND_net), .I3(VCC_net), .O(n1401)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_900_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1905_5 (.CI(n51819), .I0(n2831), 
            .I1(VCC_net), .CO(n51820));
    SB_CARRY encoder0_position_30__I_0_add_2106_23 (.CI(n51918), .I0(n3113), 
            .I1(VCC_net), .CO(n51919));
    SB_LUT4 encoder0_position_30__I_0_add_1503_14_lut (.I0(GND_net), .I1(n2222), 
            .I2(VCC_net), .I3(n51662), .O(n2289)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1503_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_151_17 (.CI(n50992), .I0(delay_counter[15]), .I1(GND_net), 
            .CO(n50993));
    SB_LUT4 encoder0_position_30__I_0_add_1168_14_lut (.I0(GND_net), .I1(n1722), 
            .I2(VCC_net), .I3(n51451), .O(n1789)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1168_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1637_10_lut (.I0(GND_net), .I1(n2426), 
            .I2(VCC_net), .I3(n51730), .O(n2493)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1637_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1503_14 (.CI(n51662), .I0(n2222), 
            .I1(VCC_net), .CO(n51663));
    SB_LUT4 encoder0_position_30__I_0_add_2106_22_lut (.I0(GND_net), .I1(n3114), 
            .I2(VCC_net), .I3(n51917), .O(n3181)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2106_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1168_14 (.CI(n51451), .I0(n1722), 
            .I1(VCC_net), .CO(n51452));
    SB_LUT4 encoder0_position_30__I_0_add_1168_13_lut (.I0(GND_net), .I1(n1723), 
            .I2(VCC_net), .I3(n51450), .O(n1790_adj_5847)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1168_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_900_2 (.CI(VCC_net), .I0(n938), 
            .I1(GND_net), .CO(n51325));
    SB_LUT4 encoder0_position_30__I_0_add_1503_13_lut (.I0(GND_net), .I1(n2223), 
            .I2(VCC_net), .I3(n51661), .O(n2290)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1503_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1168_13 (.CI(n51450), .I0(n1723), 
            .I1(VCC_net), .CO(n51451));
    SB_LUT4 encoder0_position_30__I_0_add_1905_4_lut (.I0(GND_net), .I1(n2832), 
            .I2(GND_net), .I3(n51818), .O(n2899)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1905_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2106_22 (.CI(n51917), .I0(n3114), 
            .I1(VCC_net), .CO(n51918));
    SB_LUT4 encoder0_position_30__I_0_add_833_12_lut (.I0(n70727), .I1(n1224_adj_5828), 
            .I2(VCC_net), .I3(n51324), .O(n1323)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_833_12_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_30__I_0_add_833_11_lut (.I0(GND_net), .I1(n1225_adj_5829), 
            .I2(VCC_net), .I3(n51323), .O(n1292)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_833_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1503_13 (.CI(n51661), .I0(n2223), 
            .I1(VCC_net), .CO(n51662));
    SB_CARRY encoder0_position_30__I_0_add_833_11 (.CI(n51323), .I0(n1225_adj_5829), 
            .I1(VCC_net), .CO(n51324));
    SB_LUT4 encoder0_position_30__I_0_add_1168_12_lut (.I0(GND_net), .I1(n1724), 
            .I2(VCC_net), .I3(n51449), .O(n1791)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1168_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1369_20_lut (.I0(n70477), .I1(n2016), 
            .I2(VCC_net), .I3(n51571), .O(n2115)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1369_20_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_30__I_0_add_833_10_lut (.I0(GND_net), .I1(n1226_adj_5830), 
            .I2(VCC_net), .I3(n51322), .O(n1293)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_833_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_833_10 (.CI(n51322), .I0(n1226_adj_5830), 
            .I1(VCC_net), .CO(n51323));
    SB_LUT4 add_151_16_lut (.I0(GND_net), .I1(delay_counter[14]), .I2(GND_net), 
            .I3(n50991), .O(n1225)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1168_12 (.CI(n51449), .I0(n1724), 
            .I1(VCC_net), .CO(n51450));
    SB_LUT4 encoder0_position_30__I_0_add_833_9_lut (.I0(GND_net), .I1(n1227_adj_5831), 
            .I2(VCC_net), .I3(n51321), .O(n1294)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_833_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1503_12_lut (.I0(GND_net), .I1(n2224), 
            .I2(VCC_net), .I3(n51660), .O(n2291)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1503_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1503_12 (.CI(n51660), .I0(n2224), 
            .I1(VCC_net), .CO(n51661));
    SB_LUT4 encoder0_position_30__I_0_add_1369_19_lut (.I0(GND_net), .I1(n2017), 
            .I2(VCC_net), .I3(n51570), .O(n2084)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1369_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_833_9 (.CI(n51321), .I0(n1227_adj_5831), 
            .I1(VCC_net), .CO(n51322));
    SB_CARRY add_151_9 (.CI(n50984), .I0(delay_counter[7]), .I1(GND_net), 
            .CO(n50985));
    SB_CARRY encoder0_position_30__I_0_add_1369_19 (.CI(n51570), .I0(n2017), 
            .I1(VCC_net), .CO(n51571));
    SB_LUT4 encoder0_position_30__I_0_add_1168_11_lut (.I0(GND_net), .I1(n1725), 
            .I2(VCC_net), .I3(n51448), .O(n1792_adj_5848)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1168_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1369_18_lut (.I0(GND_net), .I1(n2018), 
            .I2(VCC_net), .I3(n51569), .O(n2085)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1369_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1637_10 (.CI(n51730), .I0(n2426), 
            .I1(VCC_net), .CO(n51731));
    SB_LUT4 encoder0_position_30__I_0_add_1637_9_lut (.I0(GND_net), .I1(n2427), 
            .I2(VCC_net), .I3(n51729), .O(n2494)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1637_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1168_11 (.CI(n51448), .I0(n1725), 
            .I1(VCC_net), .CO(n51449));
    SB_LUT4 encoder0_position_30__I_0_add_833_8_lut (.I0(GND_net), .I1(n1228_adj_5832), 
            .I2(VCC_net), .I3(n51320), .O(n1295)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_833_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1503_11_lut (.I0(GND_net), .I1(n2225), 
            .I2(VCC_net), .I3(n51659), .O(n2292)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1503_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1637_9 (.CI(n51729), .I0(n2427), 
            .I1(VCC_net), .CO(n51730));
    SB_LUT4 add_151_8_lut (.I0(GND_net), .I1(delay_counter[6]), .I2(GND_net), 
            .I3(n50983), .O(n1233)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1168_10_lut (.I0(GND_net), .I1(n1726), 
            .I2(VCC_net), .I3(n51447), .O(n1793)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1168_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1369_18 (.CI(n51569), .I0(n2018), 
            .I1(VCC_net), .CO(n51570));
    SB_CARRY encoder0_position_30__I_0_add_833_8 (.CI(n51320), .I0(n1228_adj_5832), 
            .I1(VCC_net), .CO(n51321));
    SB_LUT4 encoder0_position_30__I_0_add_833_7_lut (.I0(GND_net), .I1(n1229_adj_5833), 
            .I2(GND_net), .I3(n51319), .O(n1296)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_833_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1369_17_lut (.I0(GND_net), .I1(n2019), 
            .I2(VCC_net), .I3(n51568), .O(n2086)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1369_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1637_8_lut (.I0(GND_net), .I1(n2428), 
            .I2(VCC_net), .I3(n51728), .O(n2495)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1637_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1369_17 (.CI(n51568), .I0(n2019), 
            .I1(VCC_net), .CO(n51569));
    SB_CARRY encoder0_position_30__I_0_add_1503_11 (.CI(n51659), .I0(n2225), 
            .I1(VCC_net), .CO(n51660));
    SB_CARRY encoder0_position_30__I_0_add_833_7 (.CI(n51319), .I0(n1229_adj_5833), 
            .I1(GND_net), .CO(n51320));
    SB_LUT4 encoder0_position_30__I_0_add_1369_16_lut (.I0(GND_net), .I1(n2020), 
            .I2(VCC_net), .I3(n51567), .O(n2087)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1369_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1168_10 (.CI(n51447), .I0(n1726), 
            .I1(VCC_net), .CO(n51448));
    SB_CARRY encoder0_position_30__I_0_add_1369_16 (.CI(n51567), .I0(n2020), 
            .I1(VCC_net), .CO(n51568));
    SB_CARRY encoder0_position_30__I_0_add_1637_8 (.CI(n51728), .I0(n2428), 
            .I1(VCC_net), .CO(n51729));
    SB_CARRY encoder0_position_30__I_0_add_1905_4 (.CI(n51818), .I0(n2832), 
            .I1(GND_net), .CO(n51819));
    SB_LUT4 encoder0_position_30__I_0_add_1637_7_lut (.I0(GND_net), .I1(n2429), 
            .I2(GND_net), .I3(n51727), .O(n2496)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1637_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1637_7 (.CI(n51727), .I0(n2429), 
            .I1(GND_net), .CO(n51728));
    SB_LUT4 encoder0_position_30__I_0_add_833_6_lut (.I0(GND_net), .I1(n1230_adj_5834), 
            .I2(GND_net), .I3(n51318), .O(n1297)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_833_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_833_6 (.CI(n51318), .I0(n1230_adj_5834), 
            .I1(GND_net), .CO(n51319));
    SB_LUT4 encoder0_position_30__I_0_add_2106_21_lut (.I0(GND_net), .I1(n3115), 
            .I2(VCC_net), .I3(n51916), .O(n3182)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2106_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1503_10_lut (.I0(GND_net), .I1(n2226), 
            .I2(VCC_net), .I3(n51658), .O(n2293)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1503_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1369_15_lut (.I0(GND_net), .I1(n2021), 
            .I2(VCC_net), .I3(n51566), .O(n2088)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1369_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1168_9_lut (.I0(GND_net), .I1(n1727), 
            .I2(VCC_net), .I3(n51446), .O(n1794_adj_5849)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1168_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1905_3_lut (.I0(GND_net), .I1(n2833), 
            .I2(VCC_net), .I3(n51817), .O(n2900)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1905_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1637_6_lut (.I0(GND_net), .I1(n2430), 
            .I2(GND_net), .I3(n51726), .O(n2497)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1637_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1503_10 (.CI(n51658), .I0(n2226), 
            .I1(VCC_net), .CO(n51659));
    SB_LUT4 add_151_3_lut (.I0(GND_net), .I1(delay_counter[1]), .I2(GND_net), 
            .I3(n50978), .O(n1238)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_833_5_lut (.I0(GND_net), .I1(n1231_adj_5835), 
            .I2(VCC_net), .I3(n51317), .O(n1298)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_833_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1503_9_lut (.I0(GND_net), .I1(n2227), 
            .I2(VCC_net), .I3(n51657), .O(n2294)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1503_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1915 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[16] [0]), 
            .O(n58565));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1915.LUT_INIT = 16'h2300;
    SB_CARRY encoder0_position_30__I_0_add_1905_3 (.CI(n51817), .I0(n2833), 
            .I1(VCC_net), .CO(n51818));
    SB_CARRY encoder0_position_30__I_0_add_1369_15 (.CI(n51566), .I0(n2021), 
            .I1(VCC_net), .CO(n51567));
    SB_CARRY encoder0_position_30__I_0_add_2106_21 (.CI(n51916), .I0(n3115), 
            .I1(VCC_net), .CO(n51917));
    SB_CARRY encoder0_position_30__I_0_add_1637_6 (.CI(n51726), .I0(n2430), 
            .I1(GND_net), .CO(n51727));
    SB_LUT4 encoder0_position_30__I_0_add_1369_14_lut (.I0(GND_net), .I1(n2022), 
            .I2(VCC_net), .I3(n51565), .O(n2089)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1369_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1637_5_lut (.I0(GND_net), .I1(n2431), 
            .I2(VCC_net), .I3(n51725), .O(n2498)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1637_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1369_14 (.CI(n51565), .I0(n2022), 
            .I1(VCC_net), .CO(n51566));
    SB_CARRY encoder0_position_30__I_0_add_1168_9 (.CI(n51446), .I0(n1727), 
            .I1(VCC_net), .CO(n51447));
    SB_CARRY encoder0_position_30__I_0_add_1637_5 (.CI(n51725), .I0(n2431), 
            .I1(VCC_net), .CO(n51726));
    SB_CARRY encoder0_position_30__I_0_add_1503_9 (.CI(n51657), .I0(n2227), 
            .I1(VCC_net), .CO(n51658));
    SB_LUT4 encoder0_position_30__I_0_add_1369_13_lut (.I0(GND_net), .I1(n2023), 
            .I2(VCC_net), .I3(n51564), .O(n2090)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1369_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1503_8_lut (.I0(GND_net), .I1(n2228), 
            .I2(VCC_net), .I3(n51656), .O(n2295)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1503_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_833_5 (.CI(n51317), .I0(n1231_adj_5835), 
            .I1(VCC_net), .CO(n51318));
    SB_CARRY encoder0_position_30__I_0_add_1503_8 (.CI(n51656), .I0(n2228), 
            .I1(VCC_net), .CO(n51657));
    SB_CARRY encoder0_position_30__I_0_add_1369_13 (.CI(n51564), .I0(n2023), 
            .I1(VCC_net), .CO(n51565));
    SB_LUT4 encoder0_position_30__I_0_add_1369_12_lut (.I0(GND_net), .I1(n2024), 
            .I2(VCC_net), .I3(n51563), .O(n2091)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1369_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1369_12 (.CI(n51563), .I0(n2024), 
            .I1(VCC_net), .CO(n51564));
    SB_CARRY add_151_8 (.CI(n50983), .I0(delay_counter[6]), .I1(GND_net), 
            .CO(n50984));
    SB_LUT4 encoder0_position_30__I_0_add_1637_4_lut (.I0(GND_net), .I1(n2432), 
            .I2(GND_net), .I3(n51724), .O(n2499)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1637_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_2106_20_lut (.I0(GND_net), .I1(n3116), 
            .I2(VCC_net), .I3(n51915), .O(n3183)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2106_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1369_11_lut (.I0(GND_net), .I1(n2025), 
            .I2(VCC_net), .I3(n51562), .O(n2092)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1369_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1503_7_lut (.I0(GND_net), .I1(n2229), 
            .I2(GND_net), .I3(n51655), .O(n2296)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1503_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1916 (.I0(o_Rx_DV_N_3488[12]), .I1(n4935), .I2(o_Rx_DV_N_3488[8]), 
            .I3(n62401), .O(n62407));
    defparam i1_4_lut_adj_1916.LUT_INIT = 16'hfffe;
    SB_CARRY encoder0_position_30__I_0_add_1369_11 (.CI(n51562), .I0(n2025), 
            .I1(VCC_net), .CO(n51563));
    SB_LUT4 encoder0_position_30__I_0_add_1905_2_lut (.I0(GND_net), .I1(n953), 
            .I2(GND_net), .I3(VCC_net), .O(n2901)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1905_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1168_8_lut (.I0(GND_net), .I1(n1728), 
            .I2(VCC_net), .I3(n51445), .O(n1795)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1168_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1369_10_lut (.I0(GND_net), .I1(n2026), 
            .I2(VCC_net), .I3(n51561), .O(n2093)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1369_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1905_2 (.CI(VCC_net), .I0(n953), 
            .I1(GND_net), .CO(n51817));
    SB_CARRY encoder0_position_30__I_0_add_2106_20 (.CI(n51915), .I0(n3116), 
            .I1(VCC_net), .CO(n51916));
    SB_CARRY encoder0_position_30__I_0_add_1168_8 (.CI(n51445), .I0(n1728), 
            .I1(VCC_net), .CO(n51446));
    SB_LUT4 encoder0_position_30__I_0_add_1838_27_lut (.I0(n70367), .I1(n2709), 
            .I2(VCC_net), .I3(n51816), .O(n2808)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1838_27_lut.LUT_INIT = 16'h8228;
    SB_CARRY encoder0_position_30__I_0_add_1369_10 (.CI(n51561), .I0(n2026), 
            .I1(VCC_net), .CO(n51562));
    SB_LUT4 i1_4_lut_adj_1917 (.I0(o_Rx_DV_N_3488[24]), .I1(n29_adj_5857), 
            .I2(n23_adj_5860), .I3(n62407), .O(n62413));
    defparam i1_4_lut_adj_1917.LUT_INIT = 16'hfffe;
    SB_CARRY add_151_16 (.CI(n50991), .I0(delay_counter[14]), .I1(GND_net), 
            .CO(n50992));
    SB_CARRY encoder0_position_30__I_0_add_1637_4 (.CI(n51724), .I0(n2432), 
            .I1(GND_net), .CO(n51725));
    SB_LUT4 encoder0_position_30__I_0_add_833_4_lut (.I0(GND_net), .I1(n1232_adj_5836), 
            .I2(GND_net), .I3(n51316), .O(n1299)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_833_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_833_4 (.CI(n51316), .I0(n1232_adj_5836), 
            .I1(GND_net), .CO(n51317));
    SB_CARRY encoder0_position_30__I_0_add_1503_7 (.CI(n51655), .I0(n2229), 
            .I1(GND_net), .CO(n51656));
    SB_LUT4 encoder0_position_30__I_0_add_2106_19_lut (.I0(GND_net), .I1(n3117), 
            .I2(VCC_net), .I3(n51914), .O(n3184)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2106_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1503_6_lut (.I0(GND_net), .I1(n2230), 
            .I2(GND_net), .I3(n51654), .O(n2297)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1503_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1369_9_lut (.I0(GND_net), .I1(n2027), 
            .I2(VCC_net), .I3(n51560), .O(n2094)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1369_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1168_7_lut (.I0(GND_net), .I1(n1729), 
            .I2(GND_net), .I3(n51444), .O(n1796_adj_5850)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1168_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1369_9 (.CI(n51560), .I0(n2027), 
            .I1(VCC_net), .CO(n51561));
    SB_LUT4 encoder0_position_30__I_0_add_1838_26_lut (.I0(GND_net), .I1(n2710), 
            .I2(VCC_net), .I3(n51815), .O(n2777)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1838_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1838_26 (.CI(n51815), .I0(n2710), 
            .I1(VCC_net), .CO(n51816));
    SB_CARRY add_151_3 (.CI(n50978), .I0(delay_counter[1]), .I1(GND_net), 
            .CO(n50979));
    SB_LUT4 encoder0_position_30__I_0_add_1369_8_lut (.I0(GND_net), .I1(n2028), 
            .I2(VCC_net), .I3(n51559), .O(n2095)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1369_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1637_3_lut (.I0(GND_net), .I1(n2433), 
            .I2(VCC_net), .I3(n51723), .O(n2500)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1637_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_833_3_lut (.I0(GND_net), .I1(n1233_adj_5837), 
            .I2(VCC_net), .I3(n51315), .O(n1300)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_833_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1503_6 (.CI(n51654), .I0(n2230), 
            .I1(GND_net), .CO(n51655));
    SB_CARRY encoder0_position_30__I_0_add_2106_19 (.CI(n51914), .I0(n3117), 
            .I1(VCC_net), .CO(n51915));
    SB_CARRY encoder0_position_30__I_0_add_1369_8 (.CI(n51559), .I0(n2028), 
            .I1(VCC_net), .CO(n51560));
    SB_LUT4 add_151_2_lut (.I0(GND_net), .I1(delay_counter[0]), .I2(GND_net), 
            .I3(VCC_net), .O(n1239)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1168_7 (.CI(n51444), .I0(n1729), 
            .I1(GND_net), .CO(n51445));
    SB_LUT4 encoder0_position_30__I_0_add_1369_7_lut (.I0(GND_net), .I1(n2029), 
            .I2(GND_net), .I3(n51558), .O(n2096)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1369_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1369_7 (.CI(n51558), .I0(n2029), 
            .I1(GND_net), .CO(n51559));
    SB_LUT4 encoder0_position_30__I_0_add_1838_25_lut (.I0(GND_net), .I1(n2711), 
            .I2(VCC_net), .I3(n51814), .O(n2778)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1838_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_2106_18_lut (.I0(GND_net), .I1(n3118), 
            .I2(VCC_net), .I3(n51913), .O(n3185)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2106_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1918 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[16] [1]), 
            .O(n58564));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1918.LUT_INIT = 16'h2300;
    SB_CARRY encoder0_position_30__I_0_add_833_3 (.CI(n51315), .I0(n1233_adj_5837), 
            .I1(VCC_net), .CO(n51316));
    SB_LUT4 encoder0_position_30__I_0_add_1168_6_lut (.I0(GND_net), .I1(n1730), 
            .I2(GND_net), .I3(n51443), .O(n1797)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1168_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1503_5_lut (.I0(GND_net), .I1(n2231), 
            .I2(VCC_net), .I3(n51653), .O(n2298)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1503_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_833_2_lut (.I0(GND_net), .I1(n937), 
            .I2(GND_net), .I3(VCC_net), .O(n1301)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_833_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2106_18 (.CI(n51913), .I0(n3118), 
            .I1(VCC_net), .CO(n51914));
    SB_CARRY encoder0_position_30__I_0_add_833_2 (.CI(VCC_net), .I0(n937), 
            .I1(GND_net), .CO(n51315));
    SB_LUT4 encoder0_position_30__I_0_add_1369_6_lut (.I0(GND_net), .I1(n2030), 
            .I2(GND_net), .I3(n51557), .O(n2097)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1369_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1168_6 (.CI(n51443), .I0(n1730), 
            .I1(GND_net), .CO(n51444));
    SB_CARRY encoder0_position_30__I_0_add_1369_6 (.CI(n51557), .I0(n2030), 
            .I1(GND_net), .CO(n51558));
    SB_LUT4 encoder0_position_30__I_0_add_2106_17_lut (.I0(GND_net), .I1(n3119), 
            .I2(VCC_net), .I3(n51912), .O(n3186)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2106_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1838_25 (.CI(n51814), .I0(n2711), 
            .I1(VCC_net), .CO(n51815));
    SB_LUT4 encoder0_position_30__I_0_add_1168_5_lut (.I0(GND_net), .I1(n1731), 
            .I2(VCC_net), .I3(n51442), .O(n1798)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1168_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_766_11_lut (.I0(n70712), .I1(n1125), 
            .I2(VCC_net), .I3(n51314), .O(n1224_adj_5828)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_766_11_lut.LUT_INIT = 16'h8228;
    SB_CARRY encoder0_position_30__I_0_add_1637_3 (.CI(n51723), .I0(n2433), 
            .I1(VCC_net), .CO(n51724));
    SB_CARRY encoder0_position_30__I_0_add_2106_17 (.CI(n51912), .I0(n3119), 
            .I1(VCC_net), .CO(n51913));
    SB_LUT4 i16117_4_lut (.I0(r_Rx_Data), .I1(rx_data[4]), .I2(n62413), 
            .I3(n27_adj_5858), .O(n30123));   // verilog/uart_rx.v(50[10] 145[8])
    defparam i16117_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 encoder0_position_30__I_0_add_766_10_lut (.I0(GND_net), .I1(n1126), 
            .I2(VCC_net), .I3(n51313), .O(n1193)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_766_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_151_7_lut (.I0(GND_net), .I1(delay_counter[5]), .I2(GND_net), 
            .I3(n50982), .O(n1234)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1503_5 (.CI(n51653), .I0(n2231), 
            .I1(VCC_net), .CO(n51654));
    SB_LUT4 encoder0_position_30__I_0_add_1838_24_lut (.I0(GND_net), .I1(n2712), 
            .I2(VCC_net), .I3(n51813), .O(n2779)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1838_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1503_4_lut (.I0(GND_net), .I1(n2232), 
            .I2(GND_net), .I3(n51652), .O(n2299)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1503_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1369_5_lut (.I0(GND_net), .I1(n2031), 
            .I2(VCC_net), .I3(n51556), .O(n2098)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1369_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1369_5 (.CI(n51556), .I0(n2031), 
            .I1(VCC_net), .CO(n51557));
    SB_LUT4 encoder0_position_30__I_0_add_1369_4_lut (.I0(GND_net), .I1(n2032), 
            .I2(GND_net), .I3(n51555), .O(n2099)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1369_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_2106_16_lut (.I0(GND_net), .I1(n3120), 
            .I2(VCC_net), .I3(n51911), .O(n3187)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2106_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1168_5 (.CI(n51442), .I0(n1731), 
            .I1(VCC_net), .CO(n51443));
    SB_LUT4 encoder0_position_30__I_0_add_1168_4_lut (.I0(GND_net), .I1(n1732), 
            .I2(GND_net), .I3(n51441), .O(n1799)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1168_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_766_10 (.CI(n51313), .I0(n1126), 
            .I1(VCC_net), .CO(n51314));
    SB_LUT4 encoder0_position_30__I_0_add_766_9_lut (.I0(GND_net), .I1(n1127), 
            .I2(VCC_net), .I3(n51312), .O(n1194)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_766_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1503_4 (.CI(n51652), .I0(n2232), 
            .I1(GND_net), .CO(n51653));
    SB_CARRY encoder0_position_30__I_0_add_2106_16 (.CI(n51911), .I0(n3120), 
            .I1(VCC_net), .CO(n51912));
    SB_CARRY encoder0_position_30__I_0_add_1369_4 (.CI(n51555), .I0(n2032), 
            .I1(GND_net), .CO(n51556));
    SB_LUT4 encoder0_position_30__I_0_add_2106_15_lut (.I0(GND_net), .I1(n3121), 
            .I2(VCC_net), .I3(n51910), .O(n3188)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2106_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2106_15 (.CI(n51910), .I0(n3121), 
            .I1(VCC_net), .CO(n51911));
    SB_LUT4 add_151_15_lut (.I0(GND_net), .I1(delay_counter[13]), .I2(GND_net), 
            .I3(n50990), .O(n1226)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_766_9 (.CI(n51312), .I0(n1127), 
            .I1(VCC_net), .CO(n51313));
    SB_CARRY encoder0_position_30__I_0_add_1168_4 (.CI(n51441), .I0(n1732), 
            .I1(GND_net), .CO(n51442));
    SB_LUT4 encoder0_position_30__I_0_add_2106_14_lut (.I0(GND_net), .I1(n3122), 
            .I2(VCC_net), .I3(n51909), .O(n3189)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2106_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1838_24 (.CI(n51813), .I0(n2712), 
            .I1(VCC_net), .CO(n51814));
    SB_CARRY add_151_7 (.CI(n50982), .I0(delay_counter[5]), .I1(GND_net), 
            .CO(n50983));
    SB_LUT4 encoder0_position_30__I_0_add_766_8_lut (.I0(GND_net), .I1(n1128), 
            .I2(VCC_net), .I3(n51311), .O(n1195)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_766_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_766_8 (.CI(n51311), .I0(n1128), 
            .I1(VCC_net), .CO(n51312));
    SB_LUT4 encoder0_position_30__I_0_add_1369_3_lut (.I0(GND_net), .I1(n2033), 
            .I2(VCC_net), .I3(n51554), .O(n2100)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1369_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1838_23_lut (.I0(GND_net), .I1(n2713), 
            .I2(VCC_net), .I3(n51812), .O(n2780)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1838_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2106_14 (.CI(n51909), .I0(n3122), 
            .I1(VCC_net), .CO(n51910));
    SB_CARRY encoder0_position_30__I_0_add_1838_23 (.CI(n51812), .I0(n2713), 
            .I1(VCC_net), .CO(n51813));
    SB_CARRY encoder0_position_30__I_0_add_1369_3 (.CI(n51554), .I0(n2033), 
            .I1(VCC_net), .CO(n51555));
    SB_LUT4 encoder0_position_30__I_0_add_2106_13_lut (.I0(GND_net), .I1(n3123), 
            .I2(VCC_net), .I3(n51908), .O(n3190)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2106_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1637_2_lut (.I0(GND_net), .I1(n949), 
            .I2(GND_net), .I3(VCC_net), .O(n2501)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1637_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2106_13 (.CI(n51908), .I0(n3123), 
            .I1(VCC_net), .CO(n51909));
    SB_LUT4 encoder0_position_30__I_0_add_2106_12_lut (.I0(GND_net), .I1(n3124), 
            .I2(VCC_net), .I3(n51907), .O(n3191)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2106_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1168_3_lut (.I0(GND_net), .I1(n1733), 
            .I2(VCC_net), .I3(n51440), .O(n1800)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1168_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1838_22_lut (.I0(GND_net), .I1(n2714), 
            .I2(VCC_net), .I3(n51811), .O(n2781)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1838_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_766_7_lut (.I0(GND_net), .I1(n1129), 
            .I2(GND_net), .I3(n51310), .O(n1196)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_766_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1637_2 (.CI(VCC_net), .I0(n949), 
            .I1(GND_net), .CO(n51723));
    SB_CARRY add_151_15 (.CI(n50990), .I0(delay_counter[13]), .I1(GND_net), 
            .CO(n50991));
    SB_LUT4 add_151_14_lut (.I0(GND_net), .I1(delay_counter[12]), .I2(GND_net), 
            .I3(n50989), .O(n1227)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1168_3 (.CI(n51440), .I0(n1733), 
            .I1(VCC_net), .CO(n51441));
    SB_LUT4 encoder0_position_30__I_0_add_1503_3_lut (.I0(GND_net), .I1(n2233), 
            .I2(VCC_net), .I3(n51651), .O(n2300)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1503_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1919 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[16] [2]), 
            .O(n58496));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1919.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1920 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[16] [3]), 
            .O(n58499));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1920.LUT_INIT = 16'h2300;
    SB_LUT4 i1_4_lut_adj_1921 (.I0(o_Rx_DV_N_3488[12]), .I1(n4935), .I2(o_Rx_DV_N_3488[8]), 
            .I3(n62465), .O(n62471));
    defparam i1_4_lut_adj_1921.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1922 (.I0(o_Rx_DV_N_3488[24]), .I1(n29_adj_5857), 
            .I2(n23_adj_5860), .I3(n62471), .O(n62477));
    defparam i1_4_lut_adj_1922.LUT_INIT = 16'hfffe;
    SB_LUT4 i16118_4_lut (.I0(r_Rx_Data), .I1(rx_data[5]), .I2(n62477), 
            .I3(n27_adj_5858), .O(n30124));   // verilog/uart_rx.v(50[10] 145[8])
    defparam i16118_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1923 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[16] [4]), 
            .O(n28947));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1923.LUT_INIT = 16'h2300;
    SB_CARRY encoder0_position_30__I_0_add_1838_22 (.CI(n51811), .I0(n2714), 
            .I1(VCC_net), .CO(n51812));
    SB_LUT4 encoder0_position_30__I_0_add_1369_2_lut (.I0(GND_net), .I1(n945), 
            .I2(GND_net), .I3(VCC_net), .O(n2101)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1369_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1168_2_lut (.I0(GND_net), .I1(n942), 
            .I2(GND_net), .I3(VCC_net), .O(n1801)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1168_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_766_7 (.CI(n51310), .I0(n1129), 
            .I1(GND_net), .CO(n51311));
    SB_CARRY encoder0_position_30__I_0_add_2106_12 (.CI(n51907), .I0(n3124), 
            .I1(VCC_net), .CO(n51908));
    SB_LUT4 encoder0_position_30__I_0_add_1570_23_lut (.I0(n70554), .I1(n2313), 
            .I2(VCC_net), .I3(n51722), .O(n2412)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1570_23_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_30__I_0_add_1838_21_lut (.I0(GND_net), .I1(n2715), 
            .I2(VCC_net), .I3(n51810), .O(n2782)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1838_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1168_2 (.CI(VCC_net), .I0(n942), 
            .I1(GND_net), .CO(n51440));
    SB_CARRY add_151_2 (.CI(VCC_net), .I0(delay_counter[0]), .I1(GND_net), 
            .CO(n50978));
    SB_LUT4 encoder0_position_30__I_0_add_2106_11_lut (.I0(GND_net), .I1(n3125), 
            .I2(VCC_net), .I3(n51906), .O(n3192)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2106_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1503_3 (.CI(n51651), .I0(n2233), 
            .I1(VCC_net), .CO(n51652));
    SB_CARRY encoder0_position_30__I_0_add_2106_11 (.CI(n51906), .I0(n3125), 
            .I1(VCC_net), .CO(n51907));
    SB_LUT4 encoder0_position_30__I_0_add_2106_10_lut (.I0(GND_net), .I1(n3126), 
            .I2(VCC_net), .I3(n51905), .O(n3193)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2106_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1924 (.I0(o_Rx_DV_N_3488[12]), .I1(n4935), .I2(o_Rx_DV_N_3488[8]), 
            .I3(n62513), .O(n62519));
    defparam i1_4_lut_adj_1924.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1925 (.I0(o_Rx_DV_N_3488[24]), .I1(n29_adj_5857), 
            .I2(n23_adj_5860), .I3(n62519), .O(n62525));
    defparam i1_4_lut_adj_1925.LUT_INIT = 16'hfffe;
    SB_CARRY encoder0_position_30__I_0_add_1369_2 (.CI(VCC_net), .I0(n945), 
            .I1(GND_net), .CO(n51554));
    SB_CARRY encoder0_position_30__I_0_add_1838_21 (.CI(n51810), .I0(n2715), 
            .I1(VCC_net), .CO(n51811));
    SB_LUT4 encoder0_position_30__I_0_add_1503_2_lut (.I0(GND_net), .I1(n947), 
            .I2(GND_net), .I3(VCC_net), .O(n2301)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1503_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1838_20_lut (.I0(GND_net), .I1(n2716), 
            .I2(VCC_net), .I3(n51809), .O(n2783)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1838_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1838_20 (.CI(n51809), .I0(n2716), 
            .I1(VCC_net), .CO(n51810));
    SB_LUT4 encoder0_position_30__I_0_i1387_3_lut (.I0(n2032), .I1(n2099), 
            .I2(n2049), .I3(GND_net), .O(n2131));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1387_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1926 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[16] [5]), 
            .O(n58500));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1926.LUT_INIT = 16'h2300;
    SB_LUT4 i1_3_lut_adj_1927 (.I0(n1525), .I1(n1528), .I2(n1527), .I3(GND_net), 
            .O(n62725));
    defparam i1_3_lut_adj_1927.LUT_INIT = 16'hfefe;
    SB_LUT4 encoder0_position_30__I_0_i1454_3_lut (.I0(n2131), .I1(n2198), 
            .I2(n2148), .I3(GND_net), .O(n2230));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1454_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16119_4_lut (.I0(r_Rx_Data), .I1(rx_data[6]), .I2(n62525), 
            .I3(n27_adj_5858), .O(n30125));   // verilog/uart_rx.v(50[10] 145[8])
    defparam i16119_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1928 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[16] [6]), 
            .O(n28945));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1928.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1929 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[16] [7]), 
            .O(n58501));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1929.LUT_INIT = 16'h2300;
    SB_LUT4 i1_4_lut_adj_1930 (.I0(o_Rx_DV_N_3488[12]), .I1(n4935), .I2(o_Rx_DV_N_3488[8]), 
            .I3(n62417), .O(n62423));
    defparam i1_4_lut_adj_1930.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1931 (.I0(o_Rx_DV_N_3488[24]), .I1(n29_adj_5857), 
            .I2(n23_adj_5860), .I3(n62423), .O(n62429));
    defparam i1_4_lut_adj_1931.LUT_INIT = 16'hfffe;
    SB_LUT4 i16120_4_lut (.I0(r_Rx_Data), .I1(rx_data[7]), .I2(n62429), 
            .I3(n27_adj_5858), .O(n30126));   // verilog/uart_rx.v(50[10] 145[8])
    defparam i16120_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 encoder0_position_30__I_0_add_1838_19_lut (.I0(GND_net), .I1(n2717), 
            .I2(VCC_net), .I3(n51808), .O(n2784)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1838_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1932 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[17] [0]), 
            .O(n58503));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1932.LUT_INIT = 16'h2300;
    SB_CARRY encoder0_position_30__I_0_add_2106_10 (.CI(n51905), .I0(n3126), 
            .I1(VCC_net), .CO(n51906));
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1933 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[17] [1]), 
            .O(n58505));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1933.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1934 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[17] [2]), 
            .O(n58507));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1934.LUT_INIT = 16'h2300;
    SB_LUT4 i16122_4_lut (.I0(state_7__N_4126[3]), .I1(data_adj_6007[1]), 
            .I2(n10_adj_5761), .I3(n25517), .O(n30128));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i16122_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i16123_4_lut (.I0(state_7__N_4126[3]), .I1(data_adj_6007[2]), 
            .I2(n4_adj_5756), .I3(n25522), .O(n30129));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i16123_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i16124_4_lut (.I0(state_7__N_4126[3]), .I1(data_adj_6007[3]), 
            .I2(n4_adj_5756), .I3(n25517), .O(n30130));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i16124_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i16125_4_lut (.I0(state_7__N_4126[3]), .I1(data_adj_6007[4]), 
            .I2(n4_adj_5757), .I3(n25522), .O(n30131));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i16125_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i16126_4_lut (.I0(state_7__N_4126[3]), .I1(data_adj_6007[5]), 
            .I2(n4_adj_5757), .I3(n25517), .O(n30132));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i16126_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i16127_4_lut (.I0(state_7__N_4126[3]), .I1(data_adj_6007[6]), 
            .I2(n42994), .I3(n25522), .O(n30133));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i16127_4_lut.LUT_INIT = 16'hccac;
    SB_LUT4 mux_4297_i18_3_lut (.I0(encoder0_position[17]), .I1(n15_adj_5735), 
            .I2(encoder0_position[30]), .I3(GND_net), .O(n940));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam mux_4297_i18_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_i1049_3_lut (.I0(n940), .I1(n1601), 
            .I2(n1554), .I3(GND_net), .O(n1633));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1049_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1116_3_lut (.I0(n1633), .I1(n1700), 
            .I2(n1653), .I3(GND_net), .O(n1732));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1116_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1183_3_lut (.I0(n1732), .I1(n1799), 
            .I2(n1752), .I3(GND_net), .O(n1831));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1183_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1250_3_lut (.I0(n1831), .I1(n1898), 
            .I2(n1851), .I3(GND_net), .O(n1930));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1250_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1317_3_lut (.I0(n1930), .I1(n1997), 
            .I2(n1950), .I3(GND_net), .O(n2029));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1317_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1935 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[17] [3]), 
            .O(n58508));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1935.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_i1384_3_lut (.I0(n2029), .I1(n2096), 
            .I2(n2049), .I3(GND_net), .O(n2128));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1384_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1451_3_lut (.I0(n2128), .I1(n2195), 
            .I2(n2148), .I3(GND_net), .O(n2227));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1451_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1518_3_lut (.I0(n2227), .I1(n2294), 
            .I2(n2247), .I3(GND_net), .O(n2326));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1518_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1936 (.I0(n1522), .I1(n1521), .I2(n1524), .I3(n1526), 
            .O(n61345));
    defparam i1_4_lut_adj_1936.LUT_INIT = 16'hfffe;
    SB_LUT4 i16128_4_lut (.I0(state_7__N_4126[3]), .I1(data_adj_6007[7]), 
            .I2(n42994), .I3(n25517), .O(n30134));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i16128_4_lut.LUT_INIT = 16'hccac;
    SB_LUT4 encoder0_position_30__I_0_i1585_3_lut (.I0(n2326), .I1(n2393), 
            .I2(n2346), .I3(GND_net), .O(n2425));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1585_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_add_766_6_lut (.I0(GND_net), .I1(n1130), 
            .I2(GND_net), .I3(n51309), .O(n1197)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_766_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1503_2 (.CI(VCC_net), .I0(n947), 
            .I1(GND_net), .CO(n51651));
    SB_CARRY encoder0_position_30__I_0_add_1838_19 (.CI(n51808), .I0(n2717), 
            .I1(VCC_net), .CO(n51809));
    SB_LUT4 dti_counter_1933_add_4_9_lut (.I0(GND_net), .I1(VCC_net), .I2(dti_counter[7]), 
            .I3(n52229), .O(n38_adj_5886)) /* synthesis syn_instantiated=1 */ ;
    defparam dti_counter_1933_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_2106_9_lut (.I0(GND_net), .I1(n3127), 
            .I2(VCC_net), .I3(n51904), .O(n3194)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2106_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1838_18_lut (.I0(GND_net), .I1(n2718), 
            .I2(VCC_net), .I3(n51807), .O(n2785)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1838_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 dti_counter_1933_add_4_8_lut (.I0(GND_net), .I1(VCC_net), .I2(dti_counter[6]), 
            .I3(n52228), .O(n39)) /* synthesis syn_instantiated=1 */ ;
    defparam dti_counter_1933_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY dti_counter_1933_add_4_8 (.CI(n52228), .I0(VCC_net), .I1(dti_counter[6]), 
            .CO(n52229));
    SB_CARRY encoder0_position_30__I_0_add_1838_18 (.CI(n51807), .I0(n2718), 
            .I1(VCC_net), .CO(n51808));
    SB_LUT4 dti_counter_1933_add_4_7_lut (.I0(GND_net), .I1(VCC_net), .I2(dti_counter[5]), 
            .I3(n52227), .O(n40_adj_5887)) /* synthesis syn_instantiated=1 */ ;
    defparam dti_counter_1933_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i51591_4_lut (.I0(bit_ctr[0]), .I1(n66810), .I2(n53519), .I3(color_bit_N_502[1]), 
            .O(n67130));   // verilog/neopixel.v(34[12] 116[6])
    defparam i51591_4_lut.LUT_INIT = 16'h0040;
    SB_LUT4 i26_4_lut (.I0(n22979), .I1(n67130), .I2(state[1]), .I3(n4_adj_5945), 
            .O(n57450));   // verilog/neopixel.v(34[12] 116[6])
    defparam i26_4_lut.LUT_INIT = 16'hf5c5;
    SB_CARRY encoder0_position_30__I_0_add_766_6 (.CI(n51309), .I0(n1130), 
            .I1(GND_net), .CO(n51310));
    SB_CARRY dti_counter_1933_add_4_7 (.CI(n52227), .I0(VCC_net), .I1(dti_counter[5]), 
            .CO(n52228));
    SB_LUT4 encoder0_position_30__I_0_add_1838_17_lut (.I0(GND_net), .I1(n2719), 
            .I2(VCC_net), .I3(n51806), .O(n2786)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1838_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 dti_counter_1933_add_4_6_lut (.I0(GND_net), .I1(VCC_net), .I2(dti_counter[4]), 
            .I3(n52226), .O(n41)) /* synthesis syn_instantiated=1 */ ;
    defparam dti_counter_1933_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2106_9 (.CI(n51904), .I0(n3127), 
            .I1(VCC_net), .CO(n51905));
    SB_LUT4 encoder0_position_30__I_0_add_2106_8_lut (.I0(GND_net), .I1(n3128), 
            .I2(VCC_net), .I3(n51903), .O(n3195)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2106_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY dti_counter_1933_add_4_6 (.CI(n52226), .I0(VCC_net), .I1(dti_counter[4]), 
            .CO(n52227));
    SB_LUT4 dti_counter_1933_add_4_5_lut (.I0(GND_net), .I1(VCC_net), .I2(dti_counter[3]), 
            .I3(n52225), .O(n42)) /* synthesis syn_instantiated=1 */ ;
    defparam dti_counter_1933_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_766_5_lut (.I0(GND_net), .I1(n1131), 
            .I2(VCC_net), .I3(n51308), .O(n1198)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_766_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2106_8 (.CI(n51903), .I0(n3128), 
            .I1(VCC_net), .CO(n51904));
    SB_CARRY encoder0_position_30__I_0_add_1838_17 (.CI(n51806), .I0(n2719), 
            .I1(VCC_net), .CO(n51807));
    SB_LUT4 encoder0_position_30__I_0_add_2106_7_lut (.I0(GND_net), .I1(n3129), 
            .I2(GND_net), .I3(n51902), .O(n3196)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2106_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY dti_counter_1933_add_4_5 (.CI(n52225), .I0(VCC_net), .I1(dti_counter[3]), 
            .CO(n52226));
    SB_LUT4 encoder0_position_30__I_0_i1652_3_lut (.I0(n2425), .I1(n2492), 
            .I2(n2445), .I3(GND_net), .O(n2524));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1652_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_30__I_0_add_766_5 (.CI(n51308), .I0(n1131), 
            .I1(VCC_net), .CO(n51309));
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1937 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[17] [4]), 
            .O(n58509));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1937.LUT_INIT = 16'h2300;
    SB_LUT4 dti_counter_1933_add_4_4_lut (.I0(GND_net), .I1(VCC_net), .I2(dti_counter[2]), 
            .I3(n52224), .O(n43_adj_5888)) /* synthesis syn_instantiated=1 */ ;
    defparam dti_counter_1933_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_i1719_3_lut (.I0(n2524), .I1(n2591), 
            .I2(n2544), .I3(GND_net), .O(n2623));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1719_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_add_766_4_lut (.I0(GND_net), .I1(n1132), 
            .I2(GND_net), .I3(n51307), .O(n1199)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_766_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1570_22_lut (.I0(GND_net), .I1(n2314), 
            .I2(VCC_net), .I3(n51721), .O(n2381)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1570_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1838_16_lut (.I0(GND_net), .I1(n2720), 
            .I2(VCC_net), .I3(n51805), .O(n2787)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1838_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2106_7 (.CI(n51902), .I0(n3129), 
            .I1(GND_net), .CO(n51903));
    SB_LUT4 encoder0_position_30__I_0_i1786_3_lut (.I0(n2623), .I1(n2690), 
            .I2(n2643), .I3(GND_net), .O(n2722));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1786_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_30__I_0_add_1838_16 (.CI(n51805), .I0(n2720), 
            .I1(VCC_net), .CO(n51806));
    SB_CARRY dti_counter_1933_add_4_4 (.CI(n52224), .I0(VCC_net), .I1(dti_counter[2]), 
            .CO(n52225));
    SB_LUT4 encoder0_position_30__I_0_i1853_3_lut (.I0(n2722), .I1(n2789), 
            .I2(n2742), .I3(GND_net), .O(n2821));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1853_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 dti_counter_1933_add_4_3_lut (.I0(GND_net), .I1(VCC_net), .I2(dti_counter[1]), 
            .I3(n52223), .O(n44)) /* synthesis syn_instantiated=1 */ ;
    defparam dti_counter_1933_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_i1920_3_lut (.I0(n2821), .I1(n2888), 
            .I2(n2841), .I3(GND_net), .O(n2920));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1920_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY dti_counter_1933_add_4_3 (.CI(n52223), .I0(VCC_net), .I1(dti_counter[1]), 
            .CO(n52224));
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1938 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[17] [5]), 
            .O(n58510));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1938.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_add_1838_15_lut (.I0(GND_net), .I1(n2721), 
            .I2(VCC_net), .I3(n51804), .O(n2788)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1838_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 dti_counter_1933_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(dti_counter[0]), 
            .I3(VCC_net), .O(n45_adj_5889)) /* synthesis syn_instantiated=1 */ ;
    defparam dti_counter_1933_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_i1987_3_lut (.I0(n2920), .I1(n2987), 
            .I2(n2940), .I3(GND_net), .O(n3019));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1987_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1939 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[17] [6]), 
            .O(n58511));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1939.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1940 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[17] [7]), 
            .O(n58512));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1940.LUT_INIT = 16'h2300;
    SB_CARRY dti_counter_1933_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(dti_counter[0]), 
            .CO(n52223));
    SB_LUT4 encoder0_position_30__I_0_add_2106_6_lut (.I0(GND_net), .I1(n3130), 
            .I2(GND_net), .I3(n51901), .O(n3197)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2106_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2106_6 (.CI(n51901), .I0(n3130), 
            .I1(GND_net), .CO(n51902));
    SB_LUT4 encoder0_position_30__I_0_i1521_3_lut (.I0(n2230), .I1(n2297), 
            .I2(n2247), .I3(GND_net), .O(n2329));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1521_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12_4_lut_adj_1941 (.I0(\data_in_frame[18] [7]), .I1(n28309), 
            .I2(n28366), .I3(rx_data[7]), .O(n57834));   // verilog/coms.v(130[12] 305[6])
    defparam i12_4_lut_adj_1941.LUT_INIT = 16'h3a0a;
    SB_LUT4 i12_4_lut_adj_1942 (.I0(\data_in_frame[18] [6]), .I1(n28309), 
            .I2(n28366), .I3(rx_data[6]), .O(n57838));   // verilog/coms.v(130[12] 305[6])
    defparam i12_4_lut_adj_1942.LUT_INIT = 16'h3a0a;
    SB_LUT4 i12_4_lut_adj_1943 (.I0(\data_in_frame[18] [4]), .I1(n28309), 
            .I2(n28366), .I3(rx_data[4]), .O(n57842));   // verilog/coms.v(130[12] 305[6])
    defparam i12_4_lut_adj_1943.LUT_INIT = 16'h3a0a;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1944 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[18] [0]), 
            .O(n58513));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1944.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_i703_3_lut (.I0(n1028), .I1(n1095), 
            .I2(n1059), .I3(GND_net), .O(n1127));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i703_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i770_3_lut (.I0(n1127), .I1(n1194), 
            .I2(n1158), .I3(GND_net), .O(n1226_adj_5830));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i770_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i837_3_lut (.I0(n1226_adj_5830), .I1(n1293), 
            .I2(n1257), .I3(GND_net), .O(n1325));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i837_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i904_3_lut (.I0(n1325), .I1(n1392), 
            .I2(n1356), .I3(GND_net), .O(n1424));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i904_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_add_2106_5_lut (.I0(GND_net), .I1(n3131), 
            .I2(VCC_net), .I3(n51900), .O(n3198)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2106_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_i971_3_lut (.I0(n1424), .I1(n1491), 
            .I2(n1455), .I3(GND_net), .O(n1523));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i971_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16148_3_lut (.I0(current_limit[6]), .I1(\data_in_frame[21] [6]), 
            .I2(n22734), .I3(GND_net), .O(n30154));   // verilog/coms.v(130[12] 305[6])
    defparam i16148_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1945 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[18] [1]), 
            .O(n58514));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1945.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1946 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[18] [2]), 
            .O(n58515));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1946.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_i1038_3_lut (.I0(n1523), .I1(n1590), 
            .I2(n1554), .I3(GND_net), .O(n1622));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1038_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i43881_3_lut (.I0(n4_adj_5780), .I1(n7444), .I2(n59507), .I3(GND_net), 
            .O(n59510));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam i43881_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48495_2_lut (.I0(data_ready), .I1(\ID_READOUT_FSM.state [0]), 
            .I2(GND_net), .I3(GND_net), .O(n64180));
    defparam i48495_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1947 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[18] [3]), 
            .O(n58493));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1947.LUT_INIT = 16'h2300;
    SB_CARRY encoder0_position_30__I_0_add_2106_5 (.CI(n51900), .I0(n3131), 
            .I1(VCC_net), .CO(n51901));
    SB_LUT4 i55103_4_lut (.I0(\ID_READOUT_FSM.state [1]), .I1(n6615), .I2(n64180), 
            .I3(n25_adj_5939), .O(n17_adj_5938));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i55103_4_lut.LUT_INIT = 16'h88ba;
    SB_LUT4 encoder0_position_30__I_0_i701_3_lut (.I0(n1026), .I1(n1093), 
            .I2(n1059), .I3(GND_net), .O(n1125));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i701_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i43882_3_lut (.I0(encoder0_position[28]), .I1(n59510), .I2(encoder0_position[30]), 
            .I3(GND_net), .O(n830));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam i43882_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_i569_3_lut (.I0(n830), .I1(n897), 
            .I2(n861), .I3(GND_net), .O(n929));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i569_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_i636_3_lut (.I0(n929), .I1(n996), 
            .I2(n960), .I3(GND_net), .O(n1028));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i636_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_i1036_3_lut (.I0(n1521), .I1(n1588), 
            .I2(n1554), .I3(GND_net), .O(n1620));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1036_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i11_4_lut_adj_1948 (.I0(\data_in_frame[23] [6]), .I1(n43503), 
            .I2(n28356), .I3(rx_data[6]), .O(n57996));   // verilog/coms.v(130[12] 305[6])
    defparam i11_4_lut_adj_1948.LUT_INIT = 16'hca0a;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1949 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[18] [4]), 
            .O(n58516));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1949.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i10_1_lut (.I0(encoder1_position_scaled[9]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n16_adj_5799));   // verilog/TinyFPGA_B.v(323[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1950 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[18] [5]), 
            .O(n58517));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1950.LUT_INIT = 16'h2300;
    SB_LUT4 i1_4_lut_adj_1951 (.I0(n1529), .I1(n43677), .I2(n1530), .I3(n1531), 
            .O(n60372));
    defparam i1_4_lut_adj_1951.LUT_INIT = 16'ha080;
    SB_LUT4 i54905_4_lut (.I0(n60372), .I1(n61345), .I2(n1523), .I3(n62725), 
            .O(n1554));
    defparam i54905_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_30__I_0_i1588_3_lut (.I0(n2329), .I1(n2396), 
            .I2(n2346), .I3(GND_net), .O(n2428));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1588_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_30__I_0_add_766_4 (.CI(n51307), .I0(n1132), 
            .I1(GND_net), .CO(n51308));
    SB_CARRY encoder0_position_30__I_0_add_1570_22 (.CI(n51721), .I0(n2314), 
            .I1(VCC_net), .CO(n51722));
    SB_LUT4 add_151_6_lut (.I0(GND_net), .I1(delay_counter[4]), .I2(GND_net), 
            .I3(n50981), .O(n1235)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_766_3_lut (.I0(GND_net), .I1(n1133), 
            .I2(VCC_net), .I3(n51306), .O(n1200)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_766_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_2106_4_lut (.I0(GND_net), .I1(n3132), 
            .I2(GND_net), .I3(n51899), .O(n3199)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2106_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_151_6 (.CI(n50981), .I0(delay_counter[4]), .I1(GND_net), 
            .CO(n50982));
    SB_CARRY encoder0_position_30__I_0_add_2106_4 (.CI(n51899), .I0(n3132), 
            .I1(GND_net), .CO(n51900));
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1952 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[18] [6]), 
            .O(n28929));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1952.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_add_2106_3_lut (.I0(GND_net), .I1(n3133), 
            .I2(VCC_net), .I3(n51898), .O(n3200)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2106_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1838_15 (.CI(n51804), .I0(n2721), 
            .I1(VCC_net), .CO(n51805));
    SB_LUT4 encoder0_position_30__I_0_add_1570_21_lut (.I0(GND_net), .I1(n2315), 
            .I2(VCC_net), .I3(n51720), .O(n2382)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1570_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1953 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[18] [7]), 
            .O(n28928));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1953.LUT_INIT = 16'h2300;
    SB_CARRY encoder0_position_30__I_0_add_2106_3 (.CI(n51898), .I0(n3133), 
            .I1(VCC_net), .CO(n51899));
    SB_LUT4 mux_4297_i10_3_lut (.I0(encoder0_position[9]), .I1(n23_adj_5725), 
            .I2(encoder0_position[30]), .I3(GND_net), .O(n948));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam mux_4297_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_i1593_3_lut (.I0(n948), .I1(n2401), 
            .I2(n2346), .I3(GND_net), .O(n2433));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1593_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_add_1838_14_lut (.I0(GND_net), .I1(n2722), 
            .I2(VCC_net), .I3(n51803), .O(n2789)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1838_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1954 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[19] [0]), 
            .O(n58518));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1954.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_i1660_3_lut (.I0(n2433), .I1(n2500), 
            .I2(n2445), .I3(GND_net), .O(n2532));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1660_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_30__I_0_add_1570_21 (.CI(n51720), .I0(n2315), 
            .I1(VCC_net), .CO(n51721));
    SB_LUT4 encoder0_position_30__I_0_add_2106_2_lut (.I0(GND_net), .I1(n956), 
            .I2(GND_net), .I3(VCC_net), .O(n3201)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2106_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2106_2 (.CI(VCC_net), .I0(n956), 
            .I1(GND_net), .CO(n51898));
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1955 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[19] [1]), 
            .O(n58519));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1955.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_add_2039_30_lut (.I0(n70241), .I1(n3006), 
            .I2(VCC_net), .I3(n51897), .O(n3105)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2039_30_lut.LUT_INIT = 16'h8228;
    SB_CARRY encoder0_position_30__I_0_add_1838_14 (.CI(n51803), .I0(n2722), 
            .I1(VCC_net), .CO(n51804));
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1956 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[19] [2]), 
            .O(n58520));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1956.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1957 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[19] [3]), 
            .O(n58521));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1957.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_i1655_3_lut (.I0(n2428), .I1(n2495), 
            .I2(n2445), .I3(GND_net), .O(n2527));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1655_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16073_3_lut (.I0(\data_in_frame[12] [7]), .I1(rx_data[7]), 
            .I2(n59644), .I3(GND_net), .O(n30079));   // verilog/coms.v(130[12] 305[6])
    defparam i16073_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16069_3_lut (.I0(\data_in_frame[12] [6]), .I1(rx_data[6]), 
            .I2(n59644), .I3(GND_net), .O(n30075));   // verilog/coms.v(130[12] 305[6])
    defparam i16069_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i972_3_lut (.I0(n1425), .I1(n1492), 
            .I2(n1455), .I3(GND_net), .O(n1524));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i972_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1727_3_lut (.I0(n2532), .I1(n2599), 
            .I2(n2544), .I3(GND_net), .O(n2631));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1727_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16163_3_lut (.I0(current_limit[5]), .I1(\data_in_frame[21] [5]), 
            .I2(n22734), .I3(GND_net), .O(n30169));   // verilog/coms.v(130[12] 305[6])
    defparam i16163_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16066_3_lut (.I0(\data_in_frame[12] [5]), .I1(rx_data[5]), 
            .I2(n59644), .I3(GND_net), .O(n30072));   // verilog/coms.v(130[12] 305[6])
    defparam i16066_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1794_3_lut (.I0(n2631), .I1(n2698), 
            .I2(n2643), .I3(GND_net), .O(n2730));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1794_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_add_1838_13_lut (.I0(GND_net), .I1(n2723), 
            .I2(VCC_net), .I3(n51802), .O(n2790)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1838_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_2039_29_lut (.I0(GND_net), .I1(n3007), 
            .I2(VCC_net), .I3(n51896), .O(n3074)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2039_29_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1570_20_lut (.I0(GND_net), .I1(n2316), 
            .I2(VCC_net), .I3(n51719), .O(n2383)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1570_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1838_13 (.CI(n51802), .I0(n2723), 
            .I1(VCC_net), .CO(n51803));
    SB_CARRY encoder0_position_30__I_0_add_2039_29 (.CI(n51896), .I0(n3007), 
            .I1(VCC_net), .CO(n51897));
    SB_LUT4 encoder0_position_30__I_0_add_2039_28_lut (.I0(GND_net), .I1(n3008), 
            .I2(VCC_net), .I3(n51895), .O(n3075)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2039_28_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1838_12_lut (.I0(GND_net), .I1(n2724), 
            .I2(VCC_net), .I3(n51801), .O(n2791)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1838_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2039_28 (.CI(n51895), .I0(n3008), 
            .I1(VCC_net), .CO(n51896));
    SB_LUT4 encoder0_position_30__I_0_add_2039_27_lut (.I0(GND_net), .I1(n3009), 
            .I2(VCC_net), .I3(n51894), .O(n3076)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2039_27_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i54309_3_lut (.I0(rx_data[4]), .I1(\data_in_frame[12] [4]), 
            .I2(n59644), .I3(GND_net), .O(n57936));   // verilog/coms.v(94[13:20])
    defparam i54309_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1958 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[19] [4]), 
            .O(n58522));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1958.LUT_INIT = 16'h2300;
    SB_CARRY encoder0_position_30__I_0_add_2039_27 (.CI(n51894), .I0(n3009), 
            .I1(VCC_net), .CO(n51895));
    SB_LUT4 i54308_3_lut (.I0(rx_data[3]), .I1(\data_in_frame[12] [3]), 
            .I2(n59644), .I3(GND_net), .O(n57932));   // verilog/coms.v(94[13:20])
    defparam i54308_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16056_3_lut (.I0(\data_in_frame[12] [2]), .I1(rx_data[2]), 
            .I2(n59644), .I3(GND_net), .O(n30062));   // verilog/coms.v(130[12] 305[6])
    defparam i16056_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_4297_i19_3_lut (.I0(encoder0_position[18]), .I1(n14_adj_5737), 
            .I2(encoder0_position[30]), .I3(GND_net), .O(n939));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam mux_4297_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_i981_3_lut (.I0(n939), .I1(n1501), 
            .I2(n1455), .I3(GND_net), .O(n1533));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i981_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1048_3_lut (.I0(n1533), .I1(n1600), 
            .I2(n1554), .I3(GND_net), .O(n1632));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1048_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1115_3_lut (.I0(n1632), .I1(n1699), 
            .I2(n1653), .I3(GND_net), .O(n1731));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1115_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1182_3_lut (.I0(n1731), .I1(n1798), 
            .I2(n1752), .I3(GND_net), .O(n1830));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1182_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1249_3_lut (.I0(n1830), .I1(n1897), 
            .I2(n1851), .I3(GND_net), .O(n1929));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1249_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16053_3_lut (.I0(\data_in_frame[12] [1]), .I1(rx_data[1]), 
            .I2(n59644), .I3(GND_net), .O(n30059));   // verilog/coms.v(130[12] 305[6])
    defparam i16053_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1959 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[19] [5]), 
            .O(n58523));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1959.LUT_INIT = 16'h2300;
    SB_LUT4 i16050_3_lut (.I0(\data_in_frame[12] [0]), .I1(rx_data[0]), 
            .I2(n59644), .I3(GND_net), .O(n30056));   // verilog/coms.v(130[12] 305[6])
    defparam i16050_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1316_3_lut (.I0(n1929), .I1(n1996), 
            .I2(n1950), .I3(GND_net), .O(n2028));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1316_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1383_3_lut (.I0(n2028), .I1(n2095), 
            .I2(n2049), .I3(GND_net), .O(n2127));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1383_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1450_3_lut (.I0(n2127), .I1(n2194), 
            .I2(n2148), .I3(GND_net), .O(n2226));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1450_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1517_3_lut (.I0(n2226), .I1(n2293), 
            .I2(n2247), .I3(GND_net), .O(n2325));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1517_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1584_3_lut (.I0(n2325), .I1(n2392), 
            .I2(n2346), .I3(GND_net), .O(n2424));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1584_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1909_3_lut (.I0(n2810), .I1(n2877), 
            .I2(n2841), .I3(GND_net), .O(n2909));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1909_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1651_3_lut (.I0(n2424), .I1(n2491), 
            .I2(n2445), .I3(GND_net), .O(n2523));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1651_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1718_3_lut (.I0(n2523), .I1(n2590), 
            .I2(n2544), .I3(GND_net), .O(n2622));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1718_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1908_3_lut (.I0(n2809), .I1(n2876), 
            .I2(n2841), .I3(GND_net), .O(n2908));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1908_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1785_3_lut (.I0(n2622), .I1(n2689), 
            .I2(n2643), .I3(GND_net), .O(n2721));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1785_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16047_3_lut (.I0(\data_in_frame[11] [7]), .I1(rx_data[7]), 
            .I2(n7_adj_5956), .I3(GND_net), .O(n30053));   // verilog/coms.v(130[12] 305[6])
    defparam i16047_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1852_3_lut (.I0(n2721), .I1(n2788), 
            .I2(n2742), .I3(GND_net), .O(n2820_adj_5856));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1852_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_add_3_33_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n2_adj_5892), .I3(n52457), .O(n2_adj_5781)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_unary_minus_2_add_3_33_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_add_3_32_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n3_adj_5893), .I3(n52456), .O(n3)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_unary_minus_2_add_3_32_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_unary_minus_2_add_3_32 (.CI(n52456), 
            .I0(GND_net), .I1(n3_adj_5893), .CO(n52457));
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_add_3_31_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n4_adj_5894), .I3(n52455), .O(n4_adj_5780)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_unary_minus_2_add_3_31_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_unary_minus_2_add_3_31 (.CI(n52455), 
            .I0(GND_net), .I1(n4_adj_5894), .CO(n52456));
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_add_3_30_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n5_adj_5895), .I3(n52454), .O(n5_adj_5779)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_unary_minus_2_add_3_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_unary_minus_2_add_3_30 (.CI(n52454), 
            .I0(GND_net), .I1(n5_adj_5895), .CO(n52455));
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_add_3_29_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n6_adj_5896), .I3(n52453), .O(n6_adj_5775)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_unary_minus_2_add_3_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_unary_minus_2_add_3_29 (.CI(n52453), 
            .I0(GND_net), .I1(n6_adj_5896), .CO(n52454));
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_add_3_28_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n7_adj_5897), .I3(n52452), .O(n7_adj_5774)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_unary_minus_2_add_3_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_unary_minus_2_add_3_28 (.CI(n52452), 
            .I0(GND_net), .I1(n7_adj_5897), .CO(n52453));
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_add_3_27_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n8_adj_5898), .I3(n52451), .O(n8_adj_5767)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_unary_minus_2_add_3_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_unary_minus_2_add_3_27 (.CI(n52451), 
            .I0(GND_net), .I1(n8_adj_5898), .CO(n52452));
    SB_CARRY encoder0_position_30__I_0_add_766_3 (.CI(n51306), .I0(n1133), 
            .I1(VCC_net), .CO(n51307));
    SB_LUT4 encoder0_position_30__I_0_add_2039_26_lut (.I0(GND_net), .I1(n3010), 
            .I2(VCC_net), .I3(n51893), .O(n3077)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2039_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_add_3_26_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n9_adj_5899), .I3(n52450), .O(n9_adj_5766)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_unary_minus_2_add_3_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i16043_3_lut (.I0(\data_in_frame[11] [6]), .I1(rx_data[6]), 
            .I2(n7_adj_5956), .I3(GND_net), .O(n30049));   // verilog/coms.v(130[12] 305[6])
    defparam i16043_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_30__I_0_unary_minus_2_add_3_26 (.CI(n52450), 
            .I0(GND_net), .I1(n9_adj_5899), .CO(n52451));
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_add_3_25_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n10_adj_5900), .I3(n52449), .O(n10_adj_5765)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_unary_minus_2_add_3_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_unary_minus_2_add_3_25 (.CI(n52449), 
            .I0(GND_net), .I1(n10_adj_5900), .CO(n52450));
    SB_LUT4 i16040_3_lut (.I0(\data_in_frame[11] [5]), .I1(rx_data[5]), 
            .I2(n7_adj_5956), .I3(GND_net), .O(n30046));   // verilog/coms.v(130[12] 305[6])
    defparam i16040_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1919_3_lut (.I0(n2820_adj_5856), .I1(n2887), 
            .I2(n2841), .I3(GND_net), .O(n2919));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1919_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1986_3_lut (.I0(n2919), .I1(n2986), 
            .I2(n2940), .I3(GND_net), .O(n3018));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1986_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_add_3_24_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n11_adj_5901), .I3(n52448), .O(n11_adj_5740)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_unary_minus_2_add_3_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i16037_3_lut (.I0(\data_in_frame[11] [4]), .I1(rx_data[4]), 
            .I2(n7_adj_5956), .I3(GND_net), .O(n30043));   // verilog/coms.v(130[12] 305[6])
    defparam i16037_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_30__I_0_unary_minus_2_add_3_24 (.CI(n52448), 
            .I0(GND_net), .I1(n11_adj_5901), .CO(n52449));
    SB_CARRY encoder0_position_30__I_0_add_1838_12 (.CI(n51801), .I0(n2724), 
            .I1(VCC_net), .CO(n51802));
    SB_CARRY encoder0_position_30__I_0_add_1570_20 (.CI(n51719), .I0(n2316), 
            .I1(VCC_net), .CO(n51720));
    SB_LUT4 encoder0_position_30__I_0_add_1838_11_lut (.I0(GND_net), .I1(n2725), 
            .I2(VCC_net), .I3(n51800), .O(n2792)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1838_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2039_26 (.CI(n51893), .I0(n3010), 
            .I1(VCC_net), .CO(n51894));
    SB_LUT4 encoder0_position_30__I_0_add_766_2_lut (.I0(GND_net), .I1(n522), 
            .I2(GND_net), .I3(VCC_net), .O(n1201)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_766_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_add_3_23_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n12_adj_5902), .I3(n52447), .O(n12_adj_5739)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_unary_minus_2_add_3_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_unary_minus_2_add_3_23 (.CI(n52447), 
            .I0(GND_net), .I1(n12_adj_5902), .CO(n52448));
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_add_3_22_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n13_adj_5903), .I3(n52446), .O(n13_adj_5738)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_unary_minus_2_add_3_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1960 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[19] [6]), 
            .O(n28921));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1960.LUT_INIT = 16'h2300;
    SB_CARRY encoder0_position_30__I_0_add_1838_11 (.CI(n51800), .I0(n2725), 
            .I1(VCC_net), .CO(n51801));
    SB_LUT4 i54310_3_lut (.I0(rx_data[3]), .I1(\data_in_frame[11] [3]), 
            .I2(n7_adj_5956), .I3(GND_net), .O(n58060));   // verilog/coms.v(94[13:20])
    defparam i54310_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i54314_3_lut (.I0(rx_data[2]), .I1(\data_in_frame[11] [2]), 
            .I2(n7_adj_5956), .I3(GND_net), .O(n58108));   // verilog/coms.v(94[13:20])
    defparam i54314_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_i1722_3_lut (.I0(n2527), .I1(n2594), 
            .I2(n2544), .I3(GND_net), .O(n2626));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1722_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_30__I_0_unary_minus_2_add_3_22 (.CI(n52446), 
            .I0(GND_net), .I1(n13_adj_5903), .CO(n52447));
    SB_LUT4 i54313_3_lut (.I0(rx_data[1]), .I1(\data_in_frame[11] [1]), 
            .I2(n7_adj_5956), .I3(GND_net), .O(n58106));   // verilog/coms.v(94[13:20])
    defparam i54313_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1961 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[19] [7]), 
            .O(n58524));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1961.LUT_INIT = 16'h2300;
    SB_LUT4 i2_3_lut_4_lut (.I0(n62), .I1(delay_counter[31]), .I2(data_ready), 
            .I3(\ID_READOUT_FSM.state [0]), .O(n6_adj_5947));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h2022;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1962 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[20] [0]), 
            .O(n58525));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1962.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_add_1570_19_lut (.I0(GND_net), .I1(n2317), 
            .I2(VCC_net), .I3(n51718), .O(n2384)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1570_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_add_3_21_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n14_adj_5904), .I3(n52445), .O(n14_adj_5737)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_unary_minus_2_add_3_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_unary_minus_2_add_3_21 (.CI(n52445), 
            .I0(GND_net), .I1(n14_adj_5904), .CO(n52446));
    SB_LUT4 encoder0_position_30__I_0_add_1838_10_lut (.I0(GND_net), .I1(n2726), 
            .I2(VCC_net), .I3(n51799), .O(n2793)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1838_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_add_3_20_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n15_adj_5905), .I3(n52444), .O(n15_adj_5735)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_unary_minus_2_add_3_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_unary_minus_2_add_3_20 (.CI(n52444), 
            .I0(GND_net), .I1(n15_adj_5905), .CO(n52445));
    SB_LUT4 encoder0_position_30__I_0_add_2039_25_lut (.I0(GND_net), .I1(n3011), 
            .I2(VCC_net), .I3(n51892), .O(n3078)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2039_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2039_25 (.CI(n51892), .I0(n3011), 
            .I1(VCC_net), .CO(n51893));
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_add_3_19_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n16_adj_5906), .I3(n52443), .O(n16_adj_5732)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_unary_minus_2_add_3_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_unary_minus_2_add_3_19 (.CI(n52443), 
            .I0(GND_net), .I1(n16_adj_5906), .CO(n52444));
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_add_3_18_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n17_adj_5907), .I3(n52442), .O(n17_adj_5731)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_unary_minus_2_add_3_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1853_4_lut_4_lut (.I0(\ID_READOUT_FSM.state [0]), .I1(\ID_READOUT_FSM.state [1]), 
            .I2(n1319), .I3(n42812), .O(n6615));   // verilog/TinyFPGA_B.v(361[5] 387[12])
    defparam i1853_4_lut_4_lut.LUT_INIT = 16'hcc8c;
    SB_LUT4 i16024_3_lut (.I0(\data_in_frame[11] [0]), .I1(rx_data[0]), 
            .I2(n7_adj_5956), .I3(GND_net), .O(n30030));   // verilog/coms.v(130[12] 305[6])
    defparam i16024_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_30__I_0_unary_minus_2_add_3_18 (.CI(n52442), 
            .I0(GND_net), .I1(n17_adj_5907), .CO(n52443));
    SB_CARRY encoder0_position_30__I_0_add_1838_10 (.CI(n51799), .I0(n2726), 
            .I1(VCC_net), .CO(n51800));
    SB_LUT4 encoder0_position_30__I_0_add_1838_9_lut (.I0(GND_net), .I1(n2727), 
            .I2(VCC_net), .I3(n51798), .O(n2794)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1838_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_add_3_17_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n18_adj_5908), .I3(n52441), .O(n18_adj_5730)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_unary_minus_2_add_3_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_unary_minus_2_add_3_17 (.CI(n52441), 
            .I0(GND_net), .I1(n18_adj_5908), .CO(n52442));
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_add_3_16_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n19_adj_5909), .I3(n52440), .O(n19_adj_5729)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_unary_minus_2_add_3_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_4_lut (.I0(\ID_READOUT_FSM.state [0]), .I1(\ID_READOUT_FSM.state [1]), 
            .I2(n1319), .I3(n42812), .O(n24_adj_5937));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut.LUT_INIT = 16'hffbf;
    SB_LUT4 i1_4_lut_adj_1963 (.I0(n1625), .I1(n1627), .I2(n1628), .I3(n1626), 
            .O(n63079));
    defparam i1_4_lut_adj_1963.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1964 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[20] [1]), 
            .O(n58526));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1964.LUT_INIT = 16'h2300;
    SB_CARRY encoder0_position_30__I_0_unary_minus_2_add_3_16 (.CI(n52440), 
            .I0(GND_net), .I1(n19_adj_5909), .CO(n52441));
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_add_3_15_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n20_adj_5910), .I3(n52439), .O(n20_adj_5728)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_unary_minus_2_add_3_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1965 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[20] [2]), 
            .O(n58527));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1965.LUT_INIT = 16'h2300;
    SB_LUT4 i52327_2_lut_3_lut (.I0(enable_slow_N_4213), .I1(ready_prev), 
            .I2(state_adj_6008[1]), .I3(GND_net), .O(n67177));   // verilog/eeprom.v(35[8] 81[4])
    defparam i52327_2_lut_3_lut.LUT_INIT = 16'hd0d0;
    SB_LUT4 i1_2_lut_3_lut_adj_1966 (.I0(hall1), .I1(hall2), .I2(n20873), 
            .I3(GND_net), .O(n4_adj_5958));   // verilog/TinyFPGA_B.v(151[7:22])
    defparam i1_2_lut_3_lut_adj_1966.LUT_INIT = 16'hf2f2;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1967 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[20] [3]), 
            .O(n58528));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1967.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1968 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[20] [4]), 
            .O(n58529));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1968.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1969 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[20] [5]), 
            .O(n58530));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1969.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1970 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[20] [6]), 
            .O(n58531));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1970.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1971 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[20] [7]), 
            .O(n58532));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1971.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1972 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[21] [0]), 
            .O(n58533));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1972.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1973 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[21] [1]), 
            .O(n58534));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1973.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1974 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[21] [2]), 
            .O(n58535));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1974.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1975 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[21] [3]), 
            .O(n58536));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1975.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1976 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[21] [4]), 
            .O(n58492));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1976.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1977 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[21] [5]), 
            .O(n58537));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1977.LUT_INIT = 16'h2300;
    SB_LUT4 mux_4297_i23_3_lut (.I0(encoder0_position[22]), .I1(n10_adj_5765), 
            .I2(encoder0_position[30]), .I3(GND_net), .O(n521));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam mux_4297_i23_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16192_3_lut (.I0(current_limit[4]), .I1(\data_in_frame[21] [4]), 
            .I2(n22734), .I3(GND_net), .O(n30198));   // verilog/coms.v(130[12] 305[6])
    defparam i16192_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16193_3_lut (.I0(current_limit[3]), .I1(\data_in_frame[21] [3]), 
            .I2(n22734), .I3(GND_net), .O(n30199));   // verilog/coms.v(130[12] 305[6])
    defparam i16193_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1978 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[21] [6]), 
            .O(n58538));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1978.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_i1789_3_lut (.I0(n2626), .I1(n2693), 
            .I2(n2643), .I3(GND_net), .O(n2725));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1789_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1979 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[21] [7]), 
            .O(n58539));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1979.LUT_INIT = 16'h2300;
    SB_LUT4 i12_3_lut_4_lut (.I0(rx_data_ready), .I1(r_SM_Main[1]), .I2(r_SM_Main[2]), 
            .I3(n27661), .O(n54640));   // verilog/uart_rx.v(50[10] 145[8])
    defparam i12_3_lut_4_lut.LUT_INIT = 16'h0caa;
    SB_LUT4 i15970_3_lut (.I0(\data_in_frame[8] [7]), .I1(rx_data[7]), .I2(n28385), 
            .I3(GND_net), .O(n29976));   // verilog/coms.v(130[12] 305[6])
    defparam i15970_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15967_3_lut (.I0(\data_in_frame[8] [6]), .I1(rx_data[6]), .I2(n28385), 
            .I3(GND_net), .O(n29973));   // verilog/coms.v(130[12] 305[6])
    defparam i15967_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15964_3_lut (.I0(\data_in_frame[8] [5]), .I1(rx_data[5]), .I2(n28385), 
            .I3(GND_net), .O(n29970));   // verilog/coms.v(130[12] 305[6])
    defparam i15964_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i23886_3_lut (.I0(n28385), .I1(rx_data[4]), .I2(\data_in_frame[8] [4]), 
            .I3(GND_net), .O(n30205));   // verilog/coms.v(94[13:20])
    defparam i23886_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1980 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[22] [0]), 
            .O(n28903));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1980.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1981 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[22] [1]), 
            .O(n58540));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1981.LUT_INIT = 16'h2300;
    SB_LUT4 i15958_3_lut (.I0(\data_in_frame[8] [3]), .I1(rx_data[3]), .I2(n28385), 
            .I3(GND_net), .O(n29964));   // verilog/coms.v(130[12] 305[6])
    defparam i15958_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1982 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[22] [2]), 
            .O(n58541));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1982.LUT_INIT = 16'h2300;
    SB_LUT4 i15955_3_lut (.I0(\data_in_frame[8] [2]), .I1(rx_data[2]), .I2(n28385), 
            .I3(GND_net), .O(n29961));   // verilog/coms.v(130[12] 305[6])
    defparam i15955_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15952_3_lut (.I0(\data_in_frame[8] [1]), .I1(rx_data[1]), .I2(n28385), 
            .I3(GND_net), .O(n29958));   // verilog/coms.v(130[12] 305[6])
    defparam i15952_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1983 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[22] [3]), 
            .O(n58494));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1983.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1984 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[22] [4]), 
            .O(n58542));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1984.LUT_INIT = 16'h2300;
    SB_LUT4 i51698_3_lut_4_lut (.I0(state_7__N_4110[0]), .I1(n10_adj_5758), 
            .I2(state_adj_6041[0]), .I3(enable_slow_N_4213), .O(n67171));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i51698_3_lut_4_lut.LUT_INIT = 16'h54fc;
    SB_LUT4 mux_245_i1_4_lut (.I0(encoder1_position_scaled[0]), .I1(displacement[0]), 
            .I2(n15_adj_5722), .I3(n15), .O(motor_state_23__N_91[0]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i1_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1985 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[22] [5]), 
            .O(n58543));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1985.LUT_INIT = 16'h2300;
    SB_LUT4 i15949_3_lut (.I0(\data_in_frame[8] [0]), .I1(rx_data[0]), .I2(n28385), 
            .I3(GND_net), .O(n29955));   // verilog/coms.v(130[12] 305[6])
    defparam i15949_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12_4_lut_adj_1986 (.I0(\data_in_frame[18] [2]), .I1(n28309), 
            .I2(n28366), .I3(rx_data[2]), .O(n57846));   // verilog/coms.v(130[12] 305[6])
    defparam i12_4_lut_adj_1986.LUT_INIT = 16'h3a0a;
    SB_LUT4 i15940_3_lut (.I0(\data_in_frame[7] [5]), .I1(rx_data[5]), .I2(n59638), 
            .I3(GND_net), .O(n29946));   // verilog/coms.v(130[12] 305[6])
    defparam i15940_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15937_3_lut (.I0(\data_in_frame[7] [4]), .I1(rx_data[4]), .I2(n59638), 
            .I3(GND_net), .O(n29943));   // verilog/coms.v(130[12] 305[6])
    defparam i15937_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1987 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[22] [6]), 
            .O(n58544));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1987.LUT_INIT = 16'h2300;
    SB_LUT4 mux_245_i2_4_lut (.I0(encoder1_position_scaled[1]), .I1(displacement[1]), 
            .I2(n15_adj_5722), .I3(n15), .O(motor_state_23__N_91[1]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i2_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1988 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[22] [7]), 
            .O(n58545));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1988.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1989 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[23] [0]), 
            .O(n28895));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1989.LUT_INIT = 16'h2300;
    SB_LUT4 i15934_3_lut (.I0(\data_in_frame[7] [3]), .I1(rx_data[3]), .I2(n59638), 
            .I3(GND_net), .O(n29940));   // verilog/coms.v(130[12] 305[6])
    defparam i15934_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15931_3_lut (.I0(\data_in_frame[7] [2]), .I1(rx_data[2]), .I2(n59638), 
            .I3(GND_net), .O(n29937));   // verilog/coms.v(130[12] 305[6])
    defparam i15931_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_245_i3_4_lut (.I0(encoder1_position_scaled[2]), .I1(displacement[2]), 
            .I2(n15_adj_5722), .I3(n15), .O(motor_state_23__N_91[2]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i3_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1990 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[23] [1]), 
            .O(n28894));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1990.LUT_INIT = 16'h2300;
    SB_LUT4 i15928_3_lut (.I0(\data_in_frame[7] [1]), .I1(rx_data[1]), .I2(n59638), 
            .I3(GND_net), .O(n29934));   // verilog/coms.v(130[12] 305[6])
    defparam i15928_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16212_3_lut (.I0(current_limit[2]), .I1(\data_in_frame[21] [2]), 
            .I2(n22734), .I3(GND_net), .O(n30218));   // verilog/coms.v(130[12] 305[6])
    defparam i16212_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1991 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[23] [2]), 
            .O(n58546));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1991.LUT_INIT = 16'h2300;
    SB_LUT4 i15924_3_lut (.I0(\data_in_frame[7] [0]), .I1(rx_data[0]), .I2(n59638), 
            .I3(GND_net), .O(n29930));   // verilog/coms.v(130[12] 305[6])
    defparam i15924_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1992 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[0] [2]), 
            .O(n58670));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1992.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1993 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[0] [3]), 
            .O(n58669));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1993.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1994 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[0] [4]), 
            .O(n58668));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1994.LUT_INIT = 16'h2300;
    SB_LUT4 mux_245_i4_4_lut (.I0(encoder1_position_scaled[3]), .I1(displacement[3]), 
            .I2(n15_adj_5722), .I3(n15), .O(motor_state_23__N_91[3]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i4_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1995 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[1] [0]), 
            .O(n58667));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1995.LUT_INIT = 16'h2300;
    SB_LUT4 i12_4_lut_adj_1996 (.I0(\data_in_frame[18] [1]), .I1(n28309), 
            .I2(n28366), .I3(rx_data[1]), .O(n57850));   // verilog/coms.v(130[12] 305[6])
    defparam i12_4_lut_adj_1996.LUT_INIT = 16'h3a0a;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1997 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[1] [1]), 
            .O(n58666));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1997.LUT_INIT = 16'h2300;
    SB_LUT4 i16218_3_lut (.I0(\neo_pixel_transmitter.t0 [10]), .I1(timer[10]), 
            .I2(n3157), .I3(GND_net), .O(n30224));   // verilog/neopixel.v(34[12] 116[6])
    defparam i16218_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_1998 (.I0(n40820), .I1(n8_adj_5778), .I2(GND_net), 
            .I3(GND_net), .O(n28366));
    defparam i1_2_lut_adj_1998.LUT_INIT = 16'h2222;
    SB_LUT4 i12_4_lut_adj_1999 (.I0(\data_in_frame[18] [0]), .I1(n28309), 
            .I2(n28366), .I3(rx_data[0]), .O(n57852));   // verilog/coms.v(130[12] 305[6])
    defparam i12_4_lut_adj_1999.LUT_INIT = 16'h3a0a;
    SB_LUT4 i12_4_lut_adj_2000 (.I0(\data_in_frame[17] [7]), .I1(n28311), 
            .I2(n28368), .I3(rx_data[7]), .O(n57856));   // verilog/coms.v(130[12] 305[6])
    defparam i12_4_lut_adj_2000.LUT_INIT = 16'h3a0a;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i11_1_lut (.I0(encoder1_position_scaled[10]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n15_adj_5803));   // verilog/TinyFPGA_B.v(323[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_i1863_3_lut (.I0(n2732), .I1(n2799), 
            .I2(n2742), .I3(GND_net), .O(n2831));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1863_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16224_3_lut (.I0(\neo_pixel_transmitter.t0 [9]), .I1(timer[9]), 
            .I2(n3157), .I3(GND_net), .O(n30230));   // verilog/neopixel.v(34[12] 116[6])
    defparam i16224_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16225_3_lut (.I0(\neo_pixel_transmitter.t0 [8]), .I1(timer[8]), 
            .I2(n3157), .I3(GND_net), .O(n30231));   // verilog/neopixel.v(34[12] 116[6])
    defparam i16225_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16226_3_lut (.I0(\neo_pixel_transmitter.t0 [7]), .I1(timer[7]), 
            .I2(n3157), .I3(GND_net), .O(n30232));   // verilog/neopixel.v(34[12] 116[6])
    defparam i16226_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16227_3_lut (.I0(\neo_pixel_transmitter.t0 [6]), .I1(timer[6]), 
            .I2(n3157), .I3(GND_net), .O(n30233));   // verilog/neopixel.v(34[12] 116[6])
    defparam i16227_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16228_3_lut (.I0(\neo_pixel_transmitter.t0 [5]), .I1(timer[5]), 
            .I2(n3157), .I3(GND_net), .O(n30234));   // verilog/neopixel.v(34[12] 116[6])
    defparam i16228_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_i1856_3_lut (.I0(n2725), .I1(n2792), 
            .I2(n2742), .I3(GND_net), .O(n2824));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1856_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16229_3_lut (.I0(\neo_pixel_transmitter.t0 [4]), .I1(timer[4]), 
            .I2(n3157), .I3(GND_net), .O(n30235));   // verilog/neopixel.v(34[12] 116[6])
    defparam i16229_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16230_3_lut (.I0(\neo_pixel_transmitter.t0 [3]), .I1(timer[3]), 
            .I2(n3157), .I3(GND_net), .O(n30236));   // verilog/neopixel.v(34[12] 116[6])
    defparam i16230_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16231_3_lut (.I0(\neo_pixel_transmitter.t0 [2]), .I1(timer[2]), 
            .I2(n3157), .I3(GND_net), .O(n30237));   // verilog/neopixel.v(34[12] 116[6])
    defparam i16231_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_245_i5_4_lut (.I0(encoder1_position_scaled[4]), .I1(displacement[4]), 
            .I2(n15_adj_5722), .I3(n15), .O(motor_state_23__N_91[4]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i5_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i6559_3_lut_4_lut (.I0(commutation_state[2]), .I1(commutation_state[1]), 
            .I2(commutation_state[0]), .I3(dir), .O(GLC_N_400));   // verilog/TinyFPGA_B.v(200[7] 219[14])
    defparam i6559_3_lut_4_lut.LUT_INIT = 16'hcc21;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2001 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[1] [3]), 
            .O(n58665));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2001.LUT_INIT = 16'h2300;
    SB_LUT4 i6557_3_lut_4_lut (.I0(commutation_state[2]), .I1(commutation_state[1]), 
            .I2(commutation_state[0]), .I3(dir), .O(GHC_N_391));   // verilog/TinyFPGA_B.v(200[7] 219[14])
    defparam i6557_3_lut_4_lut.LUT_INIT = 16'h21cc;
    SB_LUT4 i16232_3_lut (.I0(\neo_pixel_transmitter.t0 [1]), .I1(timer[1]), 
            .I2(n3157), .I3(GND_net), .O(n30238));   // verilog/neopixel.v(34[12] 116[6])
    defparam i16232_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2002 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[1] [5]), 
            .O(n58664));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2002.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2003 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[1] [6]), 
            .O(n58663));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2003.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2004 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[1] [7]), 
            .O(n58662));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2004.LUT_INIT = 16'h2300;
    SB_LUT4 mux_1582_i2_3_lut (.I0(duty[4]), .I1(duty[1]), .I2(n260), 
            .I3(GND_net), .O(n12211));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1582_i2_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2005 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[3] [1]), 
            .O(n58661));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2005.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2006 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[3] [3]), 
            .O(n58660));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2006.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2007 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[3] [4]), 
            .O(n58659));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2007.LUT_INIT = 16'h2300;
    SB_LUT4 i12_4_lut_adj_2008 (.I0(\data_in_frame[17] [6]), .I1(n28311), 
            .I2(n28368), .I3(rx_data[6]), .O(n57860));   // verilog/coms.v(130[12] 305[6])
    defparam i12_4_lut_adj_2008.LUT_INIT = 16'h3a0a;
    SB_LUT4 LessThan_1081_i6_3_lut_3_lut (.I0(r_Clock_Count[3]), .I1(o_Rx_DV_N_3488[3]), 
            .I2(o_Rx_DV_N_3488[2]), .I3(GND_net), .O(n6_adj_5876));   // verilog/uart_rx.v(119[17:57])
    defparam LessThan_1081_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 i12_4_lut_adj_2009 (.I0(\data_in_frame[17] [5]), .I1(n28311), 
            .I2(n28368), .I3(rx_data[5]), .O(n57864));   // verilog/coms.v(130[12] 305[6])
    defparam i12_4_lut_adj_2009.LUT_INIT = 16'h3a0a;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2010 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[3] [6]), 
            .O(n58658));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2010.LUT_INIT = 16'h2300;
    SB_LUT4 i12_4_lut_adj_2011 (.I0(\data_in_frame[17] [4]), .I1(n28311), 
            .I2(n28368), .I3(rx_data[4]), .O(n57868));   // verilog/coms.v(130[12] 305[6])
    defparam i12_4_lut_adj_2011.LUT_INIT = 16'h3a0a;
    SB_LUT4 i52134_3_lut_4_lut (.I0(r_Clock_Count[3]), .I1(o_Rx_DV_N_3488[3]), 
            .I2(o_Rx_DV_N_3488[2]), .I3(r_Clock_Count[2]), .O(n67828));   // verilog/uart_rx.v(119[17:57])
    defparam i52134_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i12_4_lut_adj_2012 (.I0(\data_in_frame[17] [3]), .I1(n28311), 
            .I2(n28368), .I3(rx_data[3]), .O(n57872));   // verilog/coms.v(130[12] 305[6])
    defparam i12_4_lut_adj_2012.LUT_INIT = 16'h3a0a;
    SB_LUT4 i12_4_lut_adj_2013 (.I0(\data_in_frame[17] [2]), .I1(n28311), 
            .I2(n28368), .I3(rx_data[2]), .O(n57874));   // verilog/coms.v(130[12] 305[6])
    defparam i12_4_lut_adj_2013.LUT_INIT = 16'h3a0a;
    SB_LUT4 i12_4_lut_adj_2014 (.I0(\data_in_frame[17] [1]), .I1(n28311), 
            .I2(n28368), .I3(rx_data[1]), .O(n57876));   // verilog/coms.v(130[12] 305[6])
    defparam i12_4_lut_adj_2014.LUT_INIT = 16'h3a0a;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2015 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[3] [7]), 
            .O(n58657));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2015.LUT_INIT = 16'h2300;
    SB_LUT4 mux_1582_i3_3_lut (.I0(duty[5]), .I1(duty[2]), .I2(n260), 
            .I3(GND_net), .O(n12209));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1582_i3_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i1_2_lut_adj_2016 (.I0(n40820), .I1(n8_adj_5798), .I2(GND_net), 
            .I3(GND_net), .O(n28368));
    defparam i1_2_lut_adj_2016.LUT_INIT = 16'h2222;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2017 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[4] [0]), 
            .O(n58506));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2017.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2018 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[4] [1]), 
            .O(n58656));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2018.LUT_INIT = 16'h2300;
    SB_LUT4 i12_4_lut_adj_2019 (.I0(\data_in_frame[17] [0]), .I1(n28311), 
            .I2(n28368), .I3(rx_data[0]), .O(n57878));   // verilog/coms.v(130[12] 305[6])
    defparam i12_4_lut_adj_2019.LUT_INIT = 16'h3a0a;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2020 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[4] [2]), 
            .O(n58655));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2020.LUT_INIT = 16'h2300;
    SB_LUT4 i12_4_lut_adj_2021 (.I0(\data_in_frame[16] [6]), .I1(n28313), 
            .I2(n28370), .I3(rx_data[6]), .O(n57882));   // verilog/coms.v(130[12] 305[6])
    defparam i12_4_lut_adj_2021.LUT_INIT = 16'h3a0a;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2022 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[4] [3]), 
            .O(n58654));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2022.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2023 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[4] [4]), 
            .O(n58653));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2023.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2024 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[4] [5]), 
            .O(n58652));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2024.LUT_INIT = 16'h2300;
    SB_LUT4 i16249_3_lut (.I0(current_limit[1]), .I1(\data_in_frame[21] [1]), 
            .I2(n22734), .I3(GND_net), .O(n30255));   // verilog/coms.v(130[12] 305[6])
    defparam i16249_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12_4_lut_adj_2025 (.I0(\data_in_frame[16] [1]), .I1(n28313), 
            .I2(n28370), .I3(rx_data[1]), .O(n57886));   // verilog/coms.v(130[12] 305[6])
    defparam i12_4_lut_adj_2025.LUT_INIT = 16'h3a0a;
    SB_LUT4 mux_245_i6_4_lut (.I0(encoder1_position_scaled[5]), .I1(displacement[5]), 
            .I2(n15_adj_5722), .I3(n15), .O(motor_state_23__N_91[5]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i6_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2026 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[4] [6]), 
            .O(n58651));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2026.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2027 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[4] [7]), 
            .O(n58650));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2027.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2028 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[5] [0]), 
            .O(n58649));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2028.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2029 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[5] [1]), 
            .O(n58648));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2029.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2030 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[5] [2]), 
            .O(n58647));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2030.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2031 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[5] [3]), 
            .O(n58646));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2031.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2032 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[5] [4]), 
            .O(n58645));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2032.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2033 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[5] [5]), 
            .O(n58644));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2033.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_i709_3_lut (.I0(n521), .I1(n1101), 
            .I2(n1059), .I3(GND_net), .O(n1133));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i709_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2034 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[5] [6]), 
            .O(n58643));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2034.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_adj_2035 (.I0(n40820), .I1(n8_adj_5801), .I2(GND_net), 
            .I3(GND_net), .O(n28370));
    defparam i1_2_lut_adj_2035.LUT_INIT = 16'h2222;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2036 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[5] [7]), 
            .O(n58642));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2036.LUT_INIT = 16'h2300;
    SB_LUT4 i12_4_lut_adj_2037 (.I0(\data_in_frame[16] [0]), .I1(n28313), 
            .I2(n28370), .I3(rx_data[0]), .O(n57890));   // verilog/coms.v(130[12] 305[6])
    defparam i12_4_lut_adj_2037.LUT_INIT = 16'h3a0a;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2038 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[6] [0]), 
            .O(n58641));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2038.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2039 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[6] [1]), 
            .O(n58640));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2039.LUT_INIT = 16'h2300;
    SB_LUT4 i29846_4_lut (.I0(n941), .I1(n1631), .I2(n1632), .I3(n1633), 
            .O(n43747));
    defparam i29846_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2040 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[6] [2]), 
            .O(n58639));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2040.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2041 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[6] [3]), 
            .O(n58638));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2041.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2042 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[6] [4]), 
            .O(n58637));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2042.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_i776_3_lut (.I0(n1133), .I1(n1200), 
            .I2(n1158), .I3(GND_net), .O(n1232_adj_5836));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i776_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2043 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[6] [5]), 
            .O(n58636));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2043.LUT_INIT = 16'h2300;
    SB_LUT4 i15895_3_lut (.I0(\data_in_frame[5] [7]), .I1(rx_data[7]), .I2(n59656), 
            .I3(GND_net), .O(n29901));   // verilog/coms.v(130[12] 305[6])
    defparam i15895_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2044 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[6] [6]), 
            .O(n58635));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2044.LUT_INIT = 16'h2300;
    SB_LUT4 i36842_3_lut_4_lut (.I0(n36845), .I1(Ki[3]), .I2(n4_adj_5863), 
            .I3(n20182), .O(n6_adj_5865));
    defparam i36842_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2045 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[6] [7]), 
            .O(n58634));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2045.LUT_INIT = 16'h2300;
    SB_LUT4 i15892_3_lut (.I0(\data_in_frame[5] [6]), .I1(rx_data[6]), .I2(n59656), 
            .I3(GND_net), .O(n29898));   // verilog/coms.v(130[12] 305[6])
    defparam i15892_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_4297_i24_3_lut (.I0(encoder0_position[23]), .I1(n9_adj_5766), 
            .I2(encoder0_position[30]), .I3(GND_net), .O(n520));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam mux_4297_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2046 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[7] [0]), 
            .O(n58633));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2046.LUT_INIT = 16'h2300;
    SB_LUT4 i1_3_lut_4_lut (.I0(n36845), .I1(Ki[3]), .I2(n4_adj_5863), 
            .I3(n20182), .O(n20136));
    defparam i1_3_lut_4_lut.LUT_INIT = 16'h8778;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2047 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[7] [1]), 
            .O(n58632));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2047.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2048 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[23] [3]), 
            .O(n58547));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2048.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2049 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[23] [4]), 
            .O(n58548));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2049.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2050 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[23] [5]), 
            .O(n58549));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2050.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i12_1_lut (.I0(encoder1_position_scaled[11]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n14_adj_5804));   // verilog/TinyFPGA_B.v(323[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2051 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[23] [6]), 
            .O(n58550));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2051.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2052 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[23] [7]), 
            .O(n58551));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2052.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2053 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[24] [0]), 
            .O(n58552));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2053.LUT_INIT = 16'h2300;
    SB_LUT4 i1_3_lut_4_lut_adj_2054 (.I0(n36845), .I1(Ki[2]), .I2(n50687), 
            .I3(n20183), .O(n20137));
    defparam i1_3_lut_4_lut_adj_2054.LUT_INIT = 16'h8778;
    SB_LUT4 i16267_3_lut (.I0(control_mode[7]), .I1(\data_in_frame[1] [7]), 
            .I2(n22734), .I3(GND_net), .O(n30273));   // verilog/coms.v(130[12] 305[6])
    defparam i16267_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2055 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[24] [1]), 
            .O(n58553));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2055.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2056 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[24] [2]), 
            .O(n58504));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2056.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2057 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[24] [3]), 
            .O(n58498));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2057.LUT_INIT = 16'h2300;
    SB_LUT4 i36834_3_lut_4_lut (.I0(n36845), .I1(Ki[2]), .I2(n50687), 
            .I3(n20183), .O(n4_adj_5863));
    defparam i36834_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2058 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[24] [4]), 
            .O(n58554));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2058.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2059 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[24] [5]), 
            .O(n58555));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2059.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2060 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[24] [6]), 
            .O(n58556));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2060.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2061 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[24] [7]), 
            .O(n58557));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2061.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_i641_3_lut (.I0(n520), .I1(n1001), 
            .I2(n960), .I3(GND_net), .O(n1033));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i641_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2062 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[25] [0]), 
            .O(n58558));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2062.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2063 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[25] [1]), 
            .O(n58497));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2063.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2064 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[25] [2]), 
            .O(n58502));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2064.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2065 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[25] [3]), 
            .O(n58559));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2065.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2066 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[7] [2]), 
            .O(n58631));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2066.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2067 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[7] [3]), 
            .O(n58630));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2067.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2068 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[7] [4]), 
            .O(n58629));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2068.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2069 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[7] [5]), 
            .O(n58628));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2069.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2070 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[25] [4]), 
            .O(n58560));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2070.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2071 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[25] [5]), 
            .O(n58561));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2071.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2072 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[25] [6]), 
            .O(n58562));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2072.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2073 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[25] [7]), 
            .O(n58563));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2073.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_i708_3_lut (.I0(n1033), .I1(n1100), 
            .I2(n1059), .I3(GND_net), .O(n1132));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i708_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2074 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[7] [6]), 
            .O(n58627));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2074.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2075 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[7] [7]), 
            .O(n58626));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2075.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2076 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[8] [0]), 
            .O(n58625));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2076.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2077 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[8] [1]), 
            .O(n58624));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2077.LUT_INIT = 16'h2300;
    SB_LUT4 mux_245_i8_4_lut (.I0(encoder1_position_scaled[7]), .I1(displacement[7]), 
            .I2(n15_adj_5722), .I3(n15), .O(motor_state_23__N_91[7]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i8_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i36821_2_lut_3_lut_4_lut (.I0(n36816), .I1(Ki[0]), .I2(Ki[1]), 
            .I3(n36845), .O(n20138));
    defparam i36821_2_lut_3_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 i36823_2_lut_3_lut_4_lut (.I0(n36816), .I1(Ki[0]), .I2(Ki[1]), 
            .I3(n36845), .O(n50687));
    defparam i36823_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i13_1_lut (.I0(encoder1_position_scaled[12]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n13_adj_5805));   // verilog/TinyFPGA_B.v(323[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_1582_i4_3_lut (.I0(duty[6]), .I1(duty[3]), .I2(n260), 
            .I3(GND_net), .O(n12207));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1582_i4_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i16299_3_lut (.I0(control_mode[6]), .I1(\data_in_frame[1] [6]), 
            .I2(n22734), .I3(GND_net), .O(n30305));   // verilog/coms.v(130[12] 305[6])
    defparam i16299_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16302_3_lut (.I0(current[11]), .I1(data_adj_6015[11]), .I2(n27643), 
            .I3(GND_net), .O(n30308));   // verilog/tli4970.v(35[10] 68[6])
    defparam i16302_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16303_3_lut (.I0(current[10]), .I1(data_adj_6015[10]), .I2(n27643), 
            .I3(GND_net), .O(n30309));   // verilog/tli4970.v(35[10] 68[6])
    defparam i16303_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16304_3_lut (.I0(current[9]), .I1(data_adj_6015[9]), .I2(n27643), 
            .I3(GND_net), .O(n30310));   // verilog/tli4970.v(35[10] 68[6])
    defparam i16304_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16305_3_lut (.I0(current[8]), .I1(data_adj_6015[8]), .I2(n27643), 
            .I3(GND_net), .O(n30311));   // verilog/tli4970.v(35[10] 68[6])
    defparam i16305_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1582_i5_3_lut (.I0(duty[7]), .I1(duty[4]), .I2(n260), 
            .I3(GND_net), .O(n12205));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1582_i5_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i16306_3_lut (.I0(current[7]), .I1(data_adj_6015[7]), .I2(n27643), 
            .I3(GND_net), .O(n30312));   // verilog/tli4970.v(35[10] 68[6])
    defparam i16306_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16307_3_lut (.I0(current[6]), .I1(data_adj_6015[6]), .I2(n27643), 
            .I3(GND_net), .O(n30313));   // verilog/tli4970.v(35[10] 68[6])
    defparam i16307_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_245_i9_4_lut (.I0(encoder1_position_scaled[8]), .I1(displacement[8]), 
            .I2(n15_adj_5722), .I3(n15), .O(motor_state_23__N_91[8]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i9_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i16309_3_lut (.I0(current[5]), .I1(data_adj_6015[5]), .I2(n27643), 
            .I3(GND_net), .O(n30315));   // verilog/tli4970.v(35[10] 68[6])
    defparam i16309_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i28311_3_lut (.I0(current[4]), .I1(data_adj_6015[4]), .I2(n27643), 
            .I3(GND_net), .O(n30316));
    defparam i28311_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16311_3_lut (.I0(current[3]), .I1(data_adj_6015[3]), .I2(n27643), 
            .I3(GND_net), .O(n30317));   // verilog/tli4970.v(35[10] 68[6])
    defparam i16311_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1582_i6_3_lut (.I0(duty[8]), .I1(duty[5]), .I2(n260), 
            .I3(GND_net), .O(n12203));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1582_i6_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i16312_3_lut (.I0(current[2]), .I1(data_adj_6015[2]), .I2(n27643), 
            .I3(GND_net), .O(n30318));   // verilog/tli4970.v(35[10] 68[6])
    defparam i16312_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16313_3_lut (.I0(current[1]), .I1(data_adj_6015[1]), .I2(n27643), 
            .I3(GND_net), .O(n30319));   // verilog/tli4970.v(35[10] 68[6])
    defparam i16313_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_i843_3_lut (.I0(n1232_adj_5836), .I1(n1299), 
            .I2(n1257), .I3(GND_net), .O(n1331));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i843_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_3_lut_4_lut_adj_2078 (.I0(n36816), .I1(Ki[3]), .I2(n4_adj_5891), 
            .I3(n20209), .O(n20181));
    defparam i1_3_lut_4_lut_adj_2078.LUT_INIT = 16'h8778;
    SB_LUT4 i16317_3_lut (.I0(baudrate[31]), .I1(data_adj_6007[7]), .I2(n61888), 
            .I3(GND_net), .O(n30323));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16317_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16318_3_lut (.I0(baudrate[30]), .I1(data_adj_6007[6]), .I2(n61888), 
            .I3(GND_net), .O(n30324));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16318_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i37049_3_lut_4_lut (.I0(n36816), .I1(Ki[3]), .I2(n4_adj_5891), 
            .I3(n20209), .O(n6_adj_5890));
    defparam i37049_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 i16319_3_lut (.I0(baudrate[29]), .I1(data_adj_6007[5]), .I2(n61888), 
            .I3(GND_net), .O(n30325));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16319_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16320_3_lut (.I0(baudrate[28]), .I1(data_adj_6007[4]), .I2(n61888), 
            .I3(GND_net), .O(n30326));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16320_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i910_3_lut (.I0(n1331), .I1(n1398), 
            .I2(n1356), .I3(GND_net), .O(n1430));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i910_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16321_3_lut (.I0(baudrate[27]), .I1(data_adj_6007[3]), .I2(n61888), 
            .I3(GND_net), .O(n30327));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16321_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16322_3_lut (.I0(baudrate[26]), .I1(data_adj_6007[2]), .I2(n61888), 
            .I3(GND_net), .O(n30328));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16322_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_3_lut_adj_2079 (.I0(n1623), .I1(n1624), .I2(n63079), .I3(GND_net), 
            .O(n63083));
    defparam i1_3_lut_adj_2079.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_4_lut_adj_2080 (.I0(n1629), .I1(n63083), .I2(n43747), .I3(n1630), 
            .O(n63085));
    defparam i1_4_lut_adj_2080.LUT_INIT = 16'heccc;
    SB_LUT4 i54924_4_lut (.I0(n1621), .I1(n1620), .I2(n63085), .I3(n1622), 
            .O(n1653));
    defparam i54924_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i16323_3_lut (.I0(baudrate[25]), .I1(data_adj_6007[1]), .I2(n61888), 
            .I3(GND_net), .O(n30329));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16323_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_adj_2081 (.I0(\data_in_frame[5] [6]), .I1(\data_in_frame[5] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n59430));   // verilog/coms.v(99[12:25])
    defparam i1_2_lut_adj_2081.LUT_INIT = 16'h6666;
    SB_LUT4 encoder0_position_30__I_0_i977_3_lut (.I0(n1430), .I1(n1497), 
            .I2(n1455), .I3(GND_net), .O(n1529));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i977_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1039_3_lut (.I0(n1524), .I1(n1591), 
            .I2(n1554), .I3(GND_net), .O(n1623));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1039_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_adj_2082 (.I0(n1728), .I1(n1727), .I2(GND_net), .I3(GND_net), 
            .O(n62911));
    defparam i1_2_lut_adj_2082.LUT_INIT = 16'heeee;
    SB_LUT4 i29698_3_lut (.I0(n942), .I1(n1732), .I2(n1733), .I3(GND_net), 
            .O(n43595));
    defparam i29698_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i16324_3_lut (.I0(baudrate[24]), .I1(data_adj_6007[0]), .I2(n61888), 
            .I3(GND_net), .O(n30330));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16324_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1044_3_lut (.I0(n1529), .I1(n1596), 
            .I2(n1554), .I3(GND_net), .O(n1628));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1044_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i27714_4_lut_4_lut (.I0(encoder1_position_scaled[6]), .I1(displacement[6]), 
            .I2(n15_adj_5722), .I3(n15), .O(n41634));
    defparam i27714_4_lut_4_lut.LUT_INIT = 16'hf535;
    SB_LUT4 i1_4_lut_adj_2083 (.I0(n1724), .I1(n1725), .I2(n62911), .I3(n1726), 
            .O(n62917));
    defparam i1_4_lut_adj_2083.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_30__I_0_i1111_3_lut (.I0(n1628), .I1(n1695), 
            .I2(n1653), .I3(GND_net), .O(n1727));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1111_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1178_3_lut (.I0(n1727), .I1(n1794_adj_5849), 
            .I2(n1752), .I3(GND_net), .O(n1826));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1178_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_2084 (.I0(n1729), .I1(n43595), .I2(n1730), .I3(n1731), 
            .O(n60380));
    defparam i1_4_lut_adj_2084.LUT_INIT = 16'ha080;
    SB_LUT4 encoder0_position_30__I_0_i1245_3_lut (.I0(n1826), .I1(n1893), 
            .I2(n1851), .I3(GND_net), .O(n1925));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1245_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_2085 (.I0(n1722), .I1(n1723), .I2(n60380), .I3(n62917), 
            .O(n62923));
    defparam i1_4_lut_adj_2085.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_30__I_0_i1312_3_lut (.I0(n1925), .I1(n1992), 
            .I2(n1950), .I3(GND_net), .O(n2024));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1312_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i54944_4_lut (.I0(n1720), .I1(n1719), .I2(n1721), .I3(n62923), 
            .O(n1752));
    defparam i54944_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_30__I_0_i1379_3_lut (.I0(n2024), .I1(n2091), 
            .I2(n2049), .I3(GND_net), .O(n2123));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1379_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1106_3_lut (.I0(n1623), .I1(n1690), 
            .I2(n1653), .I3(GND_net), .O(n1722));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1106_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_245_i10_4_lut (.I0(encoder1_position_scaled[9]), .I1(displacement[9]), 
            .I2(n15_adj_5722), .I3(n15), .O(motor_state_23__N_91[9]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i10_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i1_3_lut_adj_2086 (.I0(\data_in_frame[3] [5]), .I1(\data_in_frame[4] [7]), 
            .I2(\data_in_frame[4] [0]), .I3(GND_net), .O(n63773));   // verilog/coms.v(99[12:25])
    defparam i1_3_lut_adj_2086.LUT_INIT = 16'h9696;
    SB_LUT4 i1_4_lut_adj_2087 (.I0(n63773), .I1(n58928), .I2(\data_in_frame[3] [6]), 
            .I3(\data_in_frame[5] [3]), .O(n63779));   // verilog/coms.v(99[12:25])
    defparam i1_4_lut_adj_2087.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_2088 (.I0(n59430), .I1(n63779), .I2(n58805), 
            .I3(n59215), .O(n63783));   // verilog/coms.v(99[12:25])
    defparam i1_4_lut_adj_2088.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_2089 (.I0(n25700), .I1(n59153), .I2(Kp_23__N_748), 
            .I3(n63783), .O(n63789));   // verilog/coms.v(99[12:25])
    defparam i1_4_lut_adj_2089.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_2090 (.I0(n59299), .I1(n59007), .I2(n26282), 
            .I3(n63793), .O(n54113));   // verilog/coms.v(99[12:25])
    defparam i1_4_lut_adj_2090.LUT_INIT = 16'h6996;
    SB_LUT4 i15411_3_lut_4_lut (.I0(\data_in_frame[16] [2]), .I1(rx_data[2]), 
            .I2(n40820), .I3(n8_adj_5801), .O(n29417));   // verilog/coms.v(130[12] 305[6])
    defparam i15411_3_lut_4_lut.LUT_INIT = 16'haaca;
    SB_LUT4 i15414_3_lut_4_lut (.I0(\data_in_frame[16] [3]), .I1(rx_data[3]), 
            .I2(n40820), .I3(n8_adj_5801), .O(n29420));   // verilog/coms.v(130[12] 305[6])
    defparam i15414_3_lut_4_lut.LUT_INIT = 16'haaca;
    SB_LUT4 i15417_3_lut_4_lut (.I0(\data_in_frame[16] [4]), .I1(rx_data[4]), 
            .I2(n40820), .I3(n8_adj_5801), .O(n29423));   // verilog/coms.v(130[12] 305[6])
    defparam i15417_3_lut_4_lut.LUT_INIT = 16'haaca;
    SB_LUT4 i15420_3_lut_4_lut (.I0(\data_in_frame[16] [5]), .I1(rx_data[5]), 
            .I2(n40820), .I3(n8_adj_5801), .O(n29426));   // verilog/coms.v(130[12] 305[6])
    defparam i15420_3_lut_4_lut.LUT_INIT = 16'haaca;
    SB_LUT4 i15426_3_lut_4_lut (.I0(\data_in_frame[16] [7]), .I1(rx_data[7]), 
            .I2(n40820), .I3(n8_adj_5801), .O(n29432));   // verilog/coms.v(130[12] 305[6])
    defparam i15426_3_lut_4_lut.LUT_INIT = 16'haaca;
    SB_LUT4 mux_245_i11_4_lut (.I0(encoder1_position_scaled[10]), .I1(displacement[10]), 
            .I2(n15_adj_5722), .I3(n15), .O(motor_state_23__N_91[10]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i11_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 encoder0_position_30__I_0_i1446_3_lut (.I0(n2123), .I1(n2190), 
            .I2(n2148), .I3(GND_net), .O(n2222));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1446_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i775_3_lut (.I0(n1132), .I1(n1199), 
            .I2(n1158), .I3(GND_net), .O(n1231_adj_5835));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i775_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i6549_3_lut_4_lut_4_lut (.I0(commutation_state[2]), .I1(commutation_state[1]), 
            .I2(dir), .I3(commutation_state[0]), .O(GHA_N_355));   // verilog/TinyFPGA_B.v(179[7] 198[15])
    defparam i6549_3_lut_4_lut_4_lut.LUT_INIT = 16'h12c2;
    SB_LUT4 mux_4297_i20_3_lut (.I0(encoder0_position[19]), .I1(n13_adj_5738), 
            .I2(encoder0_position[30]), .I3(GND_net), .O(n938));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam mux_4297_i20_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_i913_3_lut (.I0(n938), .I1(n1401), 
            .I2(n1356), .I3(GND_net), .O(n1433));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i913_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i980_3_lut (.I0(n1433), .I1(n1500), 
            .I2(n1455), .I3(GND_net), .O(n1532));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i980_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1047_3_lut (.I0(n1532), .I1(n1599), 
            .I2(n1554), .I3(GND_net), .O(n1631));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1047_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i6551_3_lut_4_lut_4_lut (.I0(commutation_state[2]), .I1(commutation_state[1]), 
            .I2(dir), .I3(commutation_state[0]), .O(GLA_N_372));   // verilog/TinyFPGA_B.v(179[7] 198[15])
    defparam i6551_3_lut_4_lut_4_lut.LUT_INIT = 16'h212c;
    SB_LUT4 i6553_3_lut_4_lut_4_lut (.I0(commutation_state[2]), .I1(commutation_state[1]), 
            .I2(dir), .I3(commutation_state[0]), .O(GHB_N_377));
    defparam i6553_3_lut_4_lut_4_lut.LUT_INIT = 16'hc121;
    SB_LUT4 i1_3_lut_adj_2091 (.I0(n1825), .I1(n1824_adj_5852), .I2(n1828), 
            .I3(GND_net), .O(n63109));
    defparam i1_3_lut_adj_2091.LUT_INIT = 16'hfefe;
    SB_LUT4 encoder0_position_30__I_0_i1114_3_lut (.I0(n1631), .I1(n1698), 
            .I2(n1653), .I3(GND_net), .O(n1730));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1114_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1181_3_lut (.I0(n1730), .I1(n1797), 
            .I2(n1752), .I3(GND_net), .O(n1829));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1181_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1248_3_lut (.I0(n1829), .I1(n1896), 
            .I2(n1851), .I3(GND_net), .O(n1928));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1248_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i6555_3_lut_4_lut_4_lut (.I0(commutation_state[2]), .I1(commutation_state[1]), 
            .I2(dir), .I3(commutation_state[0]), .O(GLB_N_386));
    defparam i6555_3_lut_4_lut_4_lut.LUT_INIT = 16'h1c12;
    SB_LUT4 encoder0_position_30__I_0_i1315_3_lut (.I0(n1928), .I1(n1995), 
            .I2(n1950), .I3(GND_net), .O(n2027));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1315_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1382_3_lut (.I0(n2027), .I1(n2094), 
            .I2(n2049), .I3(GND_net), .O(n2126));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1382_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1449_3_lut (.I0(n2126), .I1(n2193), 
            .I2(n2148), .I3(GND_net), .O(n2225));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1449_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1516_3_lut (.I0(n2225), .I1(n2292), 
            .I2(n2247), .I3(GND_net), .O(n2324));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1516_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1583_3_lut (.I0(n2324), .I1(n2391), 
            .I2(n2346), .I3(GND_net), .O(n2423));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1583_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1650_3_lut (.I0(n2423), .I1(n2490), 
            .I2(n2445), .I3(GND_net), .O(n2522));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1650_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1717_3_lut (.I0(n2522), .I1(n2589), 
            .I2(n2544), .I3(GND_net), .O(n2621));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1717_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1784_3_lut (.I0(n2621), .I1(n2688), 
            .I2(n2643), .I3(GND_net), .O(n2720));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1784_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1851_3_lut (.I0(n2720), .I1(n2787), 
            .I2(n2742), .I3(GND_net), .O(n2819));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1851_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1918_3_lut (.I0(n2819), .I1(n2886), 
            .I2(n2841), .I3(GND_net), .O(n2918));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1918_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1985_3_lut (.I0(n2918), .I1(n2985), 
            .I2(n2940), .I3(GND_net), .O(n3017));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1985_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_3_lut_adj_2092 (.I0(n23_adj_5860), .I1(o_Rx_DV_N_3488[12]), 
            .I2(n4938), .I3(GND_net), .O(n62071));
    defparam i1_3_lut_adj_2092.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_4_lut_adj_2093 (.I0(o_Rx_DV_N_3488[24]), .I1(n27_adj_5858), 
            .I2(n29_adj_5857), .I3(n62071), .O(r_SM_Main_2__N_3536[1]));
    defparam i1_4_lut_adj_2093.LUT_INIT = 16'hfffe;
    SB_LUT4 LessThan_1084_i15_2_lut (.I0(r_Clock_Count_adj_6028[7]), .I1(o_Rx_DV_N_3488[7]), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_5885));   // verilog/uart_tx.v(117[17:57])
    defparam LessThan_1084_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_1084_i9_2_lut (.I0(r_Clock_Count_adj_6028[4]), .I1(o_Rx_DV_N_3488[4]), 
            .I2(GND_net), .I3(GND_net), .O(n9_adj_5882));   // verilog/uart_tx.v(117[17:57])
    defparam LessThan_1084_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mux_1582_i7_3_lut (.I0(duty[9]), .I1(duty[6]), .I2(n260), 
            .I3(GND_net), .O(n12201));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1582_i7_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 LessThan_1084_i13_2_lut (.I0(r_Clock_Count_adj_6028[6]), .I1(o_Rx_DV_N_3488[6]), 
            .I2(GND_net), .I3(GND_net), .O(n13_adj_5884));   // verilog/uart_tx.v(117[17:57])
    defparam LessThan_1084_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_1084_i11_2_lut (.I0(r_Clock_Count_adj_6028[5]), .I1(o_Rx_DV_N_3488[5]), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_5883));   // verilog/uart_tx.v(117[17:57])
    defparam LessThan_1084_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i52124_3_lut_4_lut (.I0(r_Clock_Count_adj_6028[3]), .I1(o_Rx_DV_N_3488[3]), 
            .I2(o_Rx_DV_N_3488[2]), .I3(r_Clock_Count_adj_6028[2]), .O(n67818));   // verilog/uart_tx.v(117[17:57])
    defparam i52124_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 LessThan_1084_i4_4_lut (.I0(r_Clock_Count_adj_6028[0]), .I1(o_Rx_DV_N_3488[1]), 
            .I2(r_Clock_Count_adj_6028[1]), .I3(o_Rx_DV_N_3488[0]), .O(n4_adj_5879));   // verilog/uart_tx.v(117[17:57])
    defparam LessThan_1084_i4_4_lut.LUT_INIT = 16'h4d0c;
    SB_LUT4 i53613_3_lut (.I0(n4_adj_5879), .I1(o_Rx_DV_N_3488[5]), .I2(n11_adj_5883), 
            .I3(GND_net), .O(n69307));   // verilog/uart_tx.v(117[17:57])
    defparam i53613_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53614_3_lut (.I0(n69307), .I1(o_Rx_DV_N_3488[6]), .I2(n13_adj_5884), 
            .I3(GND_net), .O(n69308));   // verilog/uart_tx.v(117[17:57])
    defparam i53614_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52996_4_lut (.I0(n13_adj_5884), .I1(n11_adj_5883), .I2(n9_adj_5882), 
            .I3(n67818), .O(n68690));
    defparam i52996_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 LessThan_1084_i8_3_lut (.I0(n6_adj_5880), .I1(o_Rx_DV_N_3488[4]), 
            .I2(n9_adj_5882), .I3(GND_net), .O(n8_adj_5881));   // verilog/uart_tx.v(117[17:57])
    defparam LessThan_1084_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52647_3_lut (.I0(n69308), .I1(o_Rx_DV_N_3488[7]), .I2(n15_adj_5885), 
            .I3(GND_net), .O(n68341));   // verilog/uart_tx.v(117[17:57])
    defparam i52647_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_1084_i6_3_lut_3_lut (.I0(r_Clock_Count_adj_6028[3]), 
            .I1(o_Rx_DV_N_3488[3]), .I2(o_Rx_DV_N_3488[2]), .I3(GND_net), 
            .O(n6_adj_5880));   // verilog/uart_tx.v(117[17:57])
    defparam LessThan_1084_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 i53597_4_lut (.I0(n68341), .I1(n8_adj_5881), .I2(n15_adj_5885), 
            .I3(n68690), .O(n69291));   // verilog/uart_tx.v(117[17:57])
    defparam i53597_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i53598_3_lut (.I0(n69291), .I1(o_Rx_DV_N_3488[8]), .I2(r_Clock_Count_adj_6028[8]), 
            .I3(GND_net), .O(n4938));   // verilog/uart_tx.v(117[17:57])
    defparam i53598_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 encoder0_position_30__I_0_i842_3_lut (.I0(n1231_adj_5835), .I1(n1298), 
            .I2(n1257), .I3(GND_net), .O(n1330));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i842_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_adj_2094 (.I0(n2327), .I1(n2328), .I2(GND_net), .I3(GND_net), 
            .O(n62831));
    defparam i1_2_lut_adj_2094.LUT_INIT = 16'heeee;
    SB_LUT4 i44010_2_lut (.I0(r_SM_Main_adj_6027[2]), .I1(r_SM_Main_adj_6027[0]), 
            .I2(GND_net), .I3(GND_net), .O(n59648));
    defparam i44010_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 encoder0_position_30__I_0_i909_3_lut (.I0(n1330), .I1(n1397), 
            .I2(n1356), .I3(GND_net), .O(n1429));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i909_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_1582_i8_3_lut (.I0(duty[10]), .I1(duty[7]), .I2(n260), 
            .I3(GND_net), .O(n12199));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1582_i8_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 mux_4297_i21_3_lut (.I0(encoder0_position[20]), .I1(n12_adj_5739), 
            .I2(encoder0_position[30]), .I3(GND_net), .O(n937));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam mux_4297_i21_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16357_3_lut (.I0(\PID_CONTROLLER.integral [23]), .I1(\PID_CONTROLLER.integral_23__N_3715 [23]), 
            .I2(control_update), .I3(GND_net), .O(n30363));   // verilog/motorControl.v(41[14] 62[8])
    defparam i16357_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_i845_3_lut (.I0(n937), .I1(n1301), 
            .I2(n1257), .I3(GND_net), .O(n1333));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i845_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16358_3_lut (.I0(\PID_CONTROLLER.integral [22]), .I1(\PID_CONTROLLER.integral_23__N_3715 [22]), 
            .I2(control_update), .I3(GND_net), .O(n30364));   // verilog/motorControl.v(41[14] 62[8])
    defparam i16358_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_i912_3_lut (.I0(n1333), .I1(n1400), 
            .I2(n1356), .I3(GND_net), .O(n1432));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i912_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i979_3_lut (.I0(n1432), .I1(n1499), 
            .I2(n1455), .I3(GND_net), .O(n1531));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i979_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1046_3_lut (.I0(n1531), .I1(n1598), 
            .I2(n1554), .I3(GND_net), .O(n1630));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1046_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1113_3_lut (.I0(n1630), .I1(n1697), 
            .I2(n1653), .I3(GND_net), .O(n1729));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1113_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1180_3_lut (.I0(n1729), .I1(n1796_adj_5850), 
            .I2(n1752), .I3(GND_net), .O(n1828));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1180_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1247_3_lut (.I0(n1828), .I1(n1895), 
            .I2(n1851), .I3(GND_net), .O(n1927));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1247_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1314_3_lut (.I0(n1927), .I1(n1994), 
            .I2(n1950), .I3(GND_net), .O(n2026));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1314_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1381_3_lut (.I0(n2026), .I1(n2093), 
            .I2(n2049), .I3(GND_net), .O(n2125));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1381_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1448_3_lut (.I0(n2125), .I1(n2192), 
            .I2(n2148), .I3(GND_net), .O(n2224));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1448_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1515_3_lut (.I0(n2224), .I1(n2291), 
            .I2(n2247), .I3(GND_net), .O(n2323));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1515_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i29818_3_lut (.I0(n948), .I1(n2332), .I2(n2333), .I3(GND_net), 
            .O(n43719));
    defparam i29818_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i16359_3_lut (.I0(\PID_CONTROLLER.integral [21]), .I1(\PID_CONTROLLER.integral_23__N_3715 [21]), 
            .I2(control_update), .I3(GND_net), .O(n30365));   // verilog/motorControl.v(41[14] 62[8])
    defparam i16359_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16360_3_lut (.I0(\PID_CONTROLLER.integral [20]), .I1(\PID_CONTROLLER.integral_23__N_3715 [20]), 
            .I2(control_update), .I3(GND_net), .O(n30366));   // verilog/motorControl.v(41[14] 62[8])
    defparam i16360_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i22854_3_lut (.I0(n212), .I1(IntegralLimit[19]), .I2(n155), 
            .I3(GND_net), .O(n36816));
    defparam i22854_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i22855_3_lut (.I0(\PID_CONTROLLER.integral [19]), .I1(n36816), 
            .I2(control_update), .I3(GND_net), .O(n30367));   // verilog/motorControl.v(20[7:21])
    defparam i22855_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i22884_3_lut (.I0(n213), .I1(IntegralLimit[18]), .I2(n155), 
            .I3(GND_net), .O(n36845));
    defparam i22884_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i22885_3_lut (.I0(\PID_CONTROLLER.integral [18]), .I1(n36845), 
            .I2(control_update), .I3(GND_net), .O(n30368));   // verilog/motorControl.v(20[7:21])
    defparam i22885_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i22922_3_lut (.I0(\PID_CONTROLLER.integral [17]), .I1(n36881), 
            .I2(control_update), .I3(GND_net), .O(n30369));   // verilog/motorControl.v(20[7:21])
    defparam i22922_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16364_3_lut (.I0(\PID_CONTROLLER.integral [16]), .I1(\PID_CONTROLLER.integral_23__N_3715 [16]), 
            .I2(control_update), .I3(GND_net), .O(n30370));   // verilog/motorControl.v(41[14] 62[8])
    defparam i16364_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16365_3_lut (.I0(\PID_CONTROLLER.integral [15]), .I1(\PID_CONTROLLER.integral_23__N_3715 [15]), 
            .I2(control_update), .I3(GND_net), .O(n30371));   // verilog/motorControl.v(41[14] 62[8])
    defparam i16365_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16366_3_lut (.I0(\PID_CONTROLLER.integral [14]), .I1(\PID_CONTROLLER.integral_23__N_3715 [14]), 
            .I2(control_update), .I3(GND_net), .O(n30372));   // verilog/motorControl.v(41[14] 62[8])
    defparam i16366_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16368_3_lut (.I0(\PID_CONTROLLER.integral [13]), .I1(\PID_CONTROLLER.integral_23__N_3715 [13]), 
            .I2(control_update), .I3(GND_net), .O(n30374));   // verilog/motorControl.v(41[14] 62[8])
    defparam i16368_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i22559_3_lut (.I0(n219), .I1(IntegralLimit[12]), .I2(n155), 
            .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3715 [12]));
    defparam i22559_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i22560_3_lut (.I0(\PID_CONTROLLER.integral [12]), .I1(\PID_CONTROLLER.integral_23__N_3715 [12]), 
            .I2(control_update), .I3(GND_net), .O(n30376));   // verilog/motorControl.v(20[7:21])
    defparam i22560_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16371_3_lut (.I0(\PID_CONTROLLER.integral [11]), .I1(\PID_CONTROLLER.integral_23__N_3715 [11]), 
            .I2(control_update), .I3(GND_net), .O(n30377));   // verilog/motorControl.v(41[14] 62[8])
    defparam i16371_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_245_i12_4_lut (.I0(encoder1_position_scaled[11]), .I1(displacement[11]), 
            .I2(n15_adj_5722), .I3(n15), .O(motor_state_23__N_91[11]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i12_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i16372_3_lut (.I0(\PID_CONTROLLER.integral [10]), .I1(\PID_CONTROLLER.integral_23__N_3715 [10]), 
            .I2(control_update), .I3(GND_net), .O(n30378));   // verilog/motorControl.v(41[14] 62[8])
    defparam i16372_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16373_3_lut (.I0(\PID_CONTROLLER.integral [9]), .I1(\PID_CONTROLLER.integral_23__N_3715 [9]), 
            .I2(control_update), .I3(GND_net), .O(n30379));   // verilog/motorControl.v(41[14] 62[8])
    defparam i16373_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16374_3_lut (.I0(\PID_CONTROLLER.integral [8]), .I1(\PID_CONTROLLER.integral_23__N_3715 [8]), 
            .I2(control_update), .I3(GND_net), .O(n30380));   // verilog/motorControl.v(41[14] 62[8])
    defparam i16374_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16375_3_lut (.I0(\PID_CONTROLLER.integral [7]), .I1(\PID_CONTROLLER.integral_23__N_3715 [7]), 
            .I2(control_update), .I3(GND_net), .O(n30381));   // verilog/motorControl.v(41[14] 62[8])
    defparam i16375_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16376_3_lut (.I0(\PID_CONTROLLER.integral [6]), .I1(\PID_CONTROLLER.integral_23__N_3715 [6]), 
            .I2(control_update), .I3(GND_net), .O(n30382));   // verilog/motorControl.v(41[14] 62[8])
    defparam i16376_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16377_3_lut (.I0(\PID_CONTROLLER.integral [5]), .I1(\PID_CONTROLLER.integral_23__N_3715 [5]), 
            .I2(control_update), .I3(GND_net), .O(n30383));   // verilog/motorControl.v(41[14] 62[8])
    defparam i16377_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1582_i9_3_lut (.I0(duty[11]), .I1(duty[8]), .I2(n260), 
            .I3(GND_net), .O(n12197));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1582_i9_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i16378_3_lut (.I0(\PID_CONTROLLER.integral [4]), .I1(\PID_CONTROLLER.integral_23__N_3715 [4]), 
            .I2(control_update), .I3(GND_net), .O(n30384));   // verilog/motorControl.v(41[14] 62[8])
    defparam i16378_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16379_3_lut (.I0(\PID_CONTROLLER.integral [3]), .I1(\PID_CONTROLLER.integral_23__N_3715 [3]), 
            .I2(control_update), .I3(GND_net), .O(n30385));   // verilog/motorControl.v(41[14] 62[8])
    defparam i16379_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16380_3_lut (.I0(\PID_CONTROLLER.integral [2]), .I1(\PID_CONTROLLER.integral_23__N_3715 [2]), 
            .I2(control_update), .I3(GND_net), .O(n30386));   // verilog/motorControl.v(41[14] 62[8])
    defparam i16380_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16381_3_lut (.I0(\PID_CONTROLLER.integral [1]), .I1(\PID_CONTROLLER.integral_23__N_3715 [1]), 
            .I2(control_update), .I3(GND_net), .O(n30387));   // verilog/motorControl.v(41[14] 62[8])
    defparam i16381_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16385_3_lut (.I0(control_mode[5]), .I1(\data_in_frame[1] [5]), 
            .I2(n22734), .I3(GND_net), .O(n30391));   // verilog/coms.v(130[12] 305[6])
    defparam i16385_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29870_4_lut (.I0(n943), .I1(n1831), .I2(n1832), .I3(n1833), 
            .O(n43771));
    defparam i29870_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 i1_4_lut_adj_2095 (.I0(n2323), .I1(n2325), .I2(n62831), .I3(n2326), 
            .O(n62835));
    defparam i1_4_lut_adj_2095.LUT_INIT = 16'hfffe;
    SB_LUT4 i16400_4_lut (.I0(commutation_state_7__N_27[2]), .I1(commutation_state[1]), 
            .I2(n20873), .I3(n4_adj_5958), .O(n30406));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    defparam i16400_4_lut.LUT_INIT = 16'h5044;
    SB_LUT4 mux_1582_i10_3_lut (.I0(duty[12]), .I1(duty[9]), .I2(n260), 
            .I3(GND_net), .O(n12195));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1582_i10_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i16_4_lut_adj_2096 (.I0(state_adj_6041[0]), .I1(n67171), .I2(n6426), 
            .I3(n6_adj_5721), .O(n8_adj_5954));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i16_4_lut_adj_2096.LUT_INIT = 16'h3afa;
    SB_LUT4 i16404_4_lut (.I0(state_7__N_4126[3]), .I1(data_adj_6007[0]), 
            .I2(n10_adj_5761), .I3(n25522), .O(n30410));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i16404_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i16410_3_lut (.I0(n59702), .I1(r_Bit_Index[0]), .I2(n27901), 
            .I3(GND_net), .O(n30416));   // verilog/uart_rx.v(50[10] 145[8])
    defparam i16410_3_lut.LUT_INIT = 16'h1414;
    SB_LUT4 i1_2_lut_adj_2097 (.I0(r_SM_Main[1]), .I1(r_SM_Main[2]), .I2(GND_net), 
            .I3(GND_net), .O(n58684));   // verilog/uart_rx.v(50[10] 145[8])
    defparam i1_2_lut_adj_2097.LUT_INIT = 16'h2222;
    SB_LUT4 mux_1582_i11_3_lut (.I0(duty[13]), .I1(duty[10]), .I2(n260), 
            .I3(GND_net), .O(n12193));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1582_i11_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i1_4_lut_adj_2098 (.I0(n2329), .I1(n43719), .I2(n2330), .I3(n2331), 
            .O(n60429));
    defparam i1_4_lut_adj_2098.LUT_INIT = 16'ha080;
    SB_LUT4 i1_4_lut_adj_2099 (.I0(n2319), .I1(n2320), .I2(n60429), .I3(n62835), 
            .O(n62841));
    defparam i1_4_lut_adj_2099.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_2100 (.I0(o_Rx_DV_N_3488[12]), .I1(n4935), .I2(o_Rx_DV_N_3488[8]), 
            .I3(n62497), .O(n62503));
    defparam i1_4_lut_adj_2100.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_2101 (.I0(o_Rx_DV_N_3488[24]), .I1(n29_adj_5857), 
            .I2(n23_adj_5860), .I3(n62503), .O(n62509));
    defparam i1_4_lut_adj_2101.LUT_INIT = 16'hfffe;
    SB_LUT4 i16414_4_lut (.I0(r_Rx_Data), .I1(rx_data[0]), .I2(n62509), 
            .I3(n27_adj_5858), .O(n30420));   // verilog/uart_rx.v(50[10] 145[8])
    defparam i16414_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i1_2_lut_adj_2102 (.I0(n36881), .I1(Ki[1]), .I2(GND_net), 
            .I3(GND_net), .O(n125));
    defparam i1_2_lut_adj_2102.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_2103 (.I0(n36845), .I1(Ki[0]), .I2(GND_net), 
            .I3(GND_net), .O(n56));
    defparam i1_2_lut_adj_2103.LUT_INIT = 16'h8888;
    SB_LUT4 i16415_3_lut (.I0(\data_in_frame[0] [0]), .I1(rx_data[0]), .I2(n7_adj_5957), 
            .I3(GND_net), .O(n30421));   // verilog/coms.v(130[12] 305[6])
    defparam i16415_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16418_4_lut (.I0(CS_MISO_c), .I1(data_adj_6015[0]), .I2(n11_adj_5764), 
            .I3(state_7__N_4319), .O(n30424));   // verilog/tli4970.v(35[10] 68[6])
    defparam i16418_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 mux_245_i13_4_lut (.I0(encoder1_position_scaled[12]), .I1(displacement[12]), 
            .I2(n15_adj_5722), .I3(n15), .O(motor_state_23__N_91[12]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i13_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i30_4_lut (.I0(state_7__N_3918[0]), .I1(n25391), .I2(state_adj_6008[1]), 
            .I3(n4_adj_5952), .O(n12_adj_5955));   // verilog/eeprom.v(35[8] 81[4])
    defparam i30_4_lut.LUT_INIT = 16'h0a3a;
    SB_LUT4 i29_4_lut (.I0(n12_adj_5955), .I1(n67177), .I2(state_adj_6008[0]), 
            .I3(state_adj_6008[2]), .O(n58002));   // verilog/eeprom.v(35[8] 81[4])
    defparam i29_4_lut.LUT_INIT = 16'hf0ca;
    SB_LUT4 i1_4_lut_adj_2104 (.I0(n2321), .I1(n2318), .I2(n2322), .I3(n2324), 
            .O(n61551));
    defparam i1_4_lut_adj_2104.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_2105 (.I0(n2316), .I1(n61551), .I2(n2317), .I3(n62841), 
            .O(n62847));
    defparam i1_4_lut_adj_2105.LUT_INIT = 16'hfffe;
    SB_LUT4 i584_2_lut (.I0(n1319), .I1(n42812), .I2(GND_net), .I3(GND_net), 
            .O(n2820));   // verilog/TinyFPGA_B.v(383[18] 385[12])
    defparam i584_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i51595_4_lut (.I0(data_ready), .I1(n6615), .I2(n24_adj_5937), 
            .I3(\ID_READOUT_FSM.state [0]), .O(n67125));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i51595_4_lut.LUT_INIT = 16'hdccc;
    SB_LUT4 i54863_4_lut (.I0(n2314), .I1(n2313), .I2(n2315), .I3(n62847), 
            .O(n2346));
    defparam i54863_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i52271_2_lut (.I0(n24_adj_5937), .I1(n6615), .I2(GND_net), 
            .I3(GND_net), .O(n67128));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i52271_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i49_4_lut (.I0(n67128), .I1(n67125), .I2(\ID_READOUT_FSM.state [0]), 
            .I3(n6_adj_5947), .O(n57114));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i49_4_lut.LUT_INIT = 16'hcac0;
    SB_LUT4 i1_2_lut_adj_2106 (.I0(n36881), .I1(Ki[2]), .I2(GND_net), 
            .I3(GND_net), .O(n198));
    defparam i1_2_lut_adj_2106.LUT_INIT = 16'h8888;
    SB_LUT4 i15602_3_lut_4_lut_4_lut (.I0(reset), .I1(n33697), .I2(\data_in_frame[6] [5]), 
            .I3(neopxl_color[5]), .O(n29608));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i15602_3_lut_4_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i15397_3_lut_4_lut_4_lut (.I0(reset), .I1(n33697), .I2(\data_in_frame[5] [5]), 
            .I3(neopxl_color[13]), .O(n29403));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i15397_3_lut_4_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i15576_3_lut_4_lut_4_lut (.I0(reset), .I1(n33697), .I2(\data_in_frame[5] [2]), 
            .I3(neopxl_color[10]), .O(n29582));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i15576_3_lut_4_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i1_2_lut_adj_2107 (.I0(n36881), .I1(Ki[3]), .I2(GND_net), 
            .I3(GND_net), .O(n271));
    defparam i1_2_lut_adj_2107.LUT_INIT = 16'h8888;
    SB_LUT4 i15600_3_lut_4_lut_4_lut (.I0(reset), .I1(n33697), .I2(\data_in_frame[6] [7]), 
            .I3(neopxl_color[7]), .O(n29606));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i15600_3_lut_4_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i15550_3_lut_4_lut_4_lut (.I0(reset), .I1(n33697), .I2(\data_in_frame[6] [0]), 
            .I3(neopxl_color[0]), .O(n29556));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i15550_3_lut_4_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i16431_3_lut (.I0(current_limit[15]), .I1(\data_in_frame[20] [7]), 
            .I2(n22734), .I3(GND_net), .O(n30437));   // verilog/coms.v(130[12] 305[6])
    defparam i16431_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_i1782_3_lut (.I0(n2619), .I1(n2686), 
            .I2(n2643), .I3(GND_net), .O(n2718));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1782_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16432_3_lut (.I0(current_limit[14]), .I1(\data_in_frame[20] [6]), 
            .I2(n22734), .I3(GND_net), .O(n30438));   // verilog/coms.v(130[12] 305[6])
    defparam i16432_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16433_3_lut (.I0(current_limit[13]), .I1(\data_in_frame[20] [5]), 
            .I2(n22734), .I3(GND_net), .O(n30439));   // verilog/coms.v(130[12] 305[6])
    defparam i16433_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_i1849_3_lut (.I0(n2718), .I1(n2785), 
            .I2(n2742), .I3(GND_net), .O(n2817));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1849_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_245_i14_4_lut (.I0(encoder1_position_scaled[13]), .I1(displacement[13]), 
            .I2(n15_adj_5722), .I3(n15), .O(motor_state_23__N_91[13]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i14_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i1_4_lut_adj_2108 (.I0(n1823), .I1(n63109), .I2(n1827), .I3(n1826), 
            .O(n63113));
    defparam i1_4_lut_adj_2108.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_30__I_0_i1513_3_lut (.I0(n2222), .I1(n2289), 
            .I2(n2247), .I3(GND_net), .O(n2321));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1513_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_2109 (.I0(n2426), .I1(n2425), .I2(n2428), .I3(n2427), 
            .O(n63207));
    defparam i1_4_lut_adj_2109.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_3_lut_adj_2110 (.I0(n1820), .I1(n1821), .I2(n1822_adj_5851), 
            .I3(GND_net), .O(n63119));
    defparam i1_3_lut_adj_2110.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_2_lut_adj_2111 (.I0(n36881), .I1(Ki[4]), .I2(GND_net), 
            .I3(GND_net), .O(n344));
    defparam i1_2_lut_adj_2111.LUT_INIT = 16'h8888;
    SB_LUT4 i28800_3_lut_4_lut_4_lut (.I0(reset), .I1(n33697), .I2(\data_in_frame[5] [3]), 
            .I3(neopxl_color[11]), .O(n29410));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i28800_3_lut_4_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 mux_1582_i12_3_lut (.I0(duty[14]), .I1(duty[11]), .I2(n260), 
            .I3(GND_net), .O(n12191));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1582_i12_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i15399_3_lut_4_lut_4_lut (.I0(reset), .I1(n33697), .I2(\data_in_frame[5] [4]), 
            .I3(neopxl_color[12]), .O(n29405));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i15399_3_lut_4_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i15599_3_lut_4_lut_4_lut (.I0(reset), .I1(n33697), .I2(\data_in_frame[5] [0]), 
            .I3(neopxl_color[8]), .O(n29605));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i15599_3_lut_4_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_55294 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[22] [4]), .I2(\data_out_frame[23] [4]), 
            .I3(byte_transmit_counter[1]), .O(n71000));
    defparam byte_transmit_counter_0__bdd_4_lut_55294.LUT_INIT = 16'he4aa;
    SB_LUT4 i29816_3_lut (.I0(n949), .I1(n2432), .I2(n2433), .I3(GND_net), 
            .O(n43717));
    defparam i29816_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 mux_245_i18_4_lut (.I0(encoder1_position_scaled[17]), .I1(displacement[17]), 
            .I2(n15_adj_5722), .I3(n15), .O(motor_state_23__N_91[17]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i18_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i15598_3_lut_4_lut_4_lut (.I0(reset), .I1(n33697), .I2(\data_in_frame[5] [1]), 
            .I3(neopxl_color[9]), .O(n29604));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i15598_3_lut_4_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i1_4_lut_adj_2112 (.I0(n63207), .I1(n2423), .I2(n2424), .I3(n2421), 
            .O(n63209));
    defparam i1_4_lut_adj_2112.LUT_INIT = 16'hfffe;
    SB_LUT4 mux_1582_i13_3_lut (.I0(duty[15]), .I1(duty[12]), .I2(n260), 
            .I3(GND_net), .O(n12189));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1582_i13_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i1_4_lut_adj_2113 (.I0(n1829), .I1(n63113), .I2(n43771), .I3(n1830), 
            .O(n63115));
    defparam i1_4_lut_adj_2113.LUT_INIT = 16'heccc;
    SB_LUT4 i1_4_lut_adj_2114 (.I0(n2429), .I1(n43717), .I2(n2430), .I3(n2431), 
            .O(n60464));
    defparam i1_4_lut_adj_2114.LUT_INIT = 16'ha080;
    SB_LUT4 i54887_4_lut (.I0(n1818), .I1(n63115), .I2(n63119), .I3(n1819), 
            .O(n1851));
    defparam i54887_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i1_4_lut_adj_2115 (.I0(n2417), .I1(n60464), .I2(n63209), .I3(n2420), 
            .O(n63215));
    defparam i1_4_lut_adj_2115.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_30__I_0_i1173_3_lut (.I0(n1722), .I1(n1789), 
            .I2(n1752), .I3(GND_net), .O(n1821));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1173_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_3_lut_adj_2116 (.I0(n2418), .I1(n2419), .I2(n2422), .I3(GND_net), 
            .O(n63311));
    defparam i1_3_lut_adj_2116.LUT_INIT = 16'hfefe;
    SB_LUT4 n71000_bdd_4_lut (.I0(n71000), .I1(\data_out_frame[21] [4]), 
            .I2(\data_out_frame[20] [4]), .I3(byte_transmit_counter[1]), 
            .O(n71003));
    defparam n71000_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_4_lut_adj_2117 (.I0(n63311), .I1(n2415), .I2(n63215), .I3(n2416), 
            .O(n63219));
    defparam i1_4_lut_adj_2117.LUT_INIT = 16'hfffe;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_55482 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[18] [3]), .I2(\data_out_frame[19] [3]), 
            .I3(byte_transmit_counter[1]), .O(n71222));
    defparam byte_transmit_counter_0__bdd_4_lut_55482.LUT_INIT = 16'he4aa;
    SB_LUT4 i54646_4_lut (.I0(n2413), .I1(n2412), .I2(n2414), .I3(n63219), 
            .O(n2445));
    defparam i54646_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i15601_3_lut_4_lut_4_lut (.I0(reset), .I1(n33697), .I2(\data_in_frame[6] [6]), 
            .I3(neopxl_color[6]), .O(n29607));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i15601_3_lut_4_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i15606_3_lut_4_lut_4_lut (.I0(reset), .I1(n33697), .I2(\data_in_frame[6] [4]), 
            .I3(neopxl_color[4]), .O(n29612));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i15606_3_lut_4_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i23887_3_lut_4_lut_4_lut (.I0(reset), .I1(n33697), .I2(\data_in_frame[6] [3]), 
            .I3(neopxl_color[3]), .O(n29613));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i23887_3_lut_4_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i15625_3_lut_4_lut_4_lut (.I0(reset), .I1(n33697), .I2(\data_in_frame[4] [6]), 
            .I3(neopxl_color[22]), .O(n29631));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i15625_3_lut_4_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i1_2_lut_adj_2118 (.I0(n36881), .I1(Ki[5]), .I2(GND_net), 
            .I3(GND_net), .O(n417));
    defparam i1_2_lut_adj_2118.LUT_INIT = 16'h8888;
    SB_LUT4 i15632_3_lut_4_lut_4_lut (.I0(reset), .I1(n33697), .I2(\data_in_frame[5] [6]), 
            .I3(neopxl_color[14]), .O(n29638));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i15632_3_lut_4_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i15636_3_lut_4_lut_4_lut (.I0(reset), .I1(n33697), .I2(\data_in_frame[6] [1]), 
            .I3(neopxl_color[1]), .O(n29642));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i15636_3_lut_4_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i16104_3_lut_4_lut (.I0(\data_in_frame[23] [7]), .I1(rx_data[7]), 
            .I2(reset), .I3(n75), .O(n30110));   // verilog/coms.v(130[12] 305[6])
    defparam i16104_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i16133_4_lut_4_lut (.I0(n27855), .I1(state[1]), .I2(bit_ctr[1]), 
            .I3(bit_ctr[0]), .O(n30139));   // verilog/neopixel.v(34[12] 116[6])
    defparam i16133_4_lut_4_lut.LUT_INIT = 16'h5270;
    SB_LUT4 i1_2_lut_adj_2119 (.I0(n36816), .I1(Ki[2]), .I2(GND_net), 
            .I3(GND_net), .O(n204));
    defparam i1_2_lut_adj_2119.LUT_INIT = 16'h8888;
    SB_LUT4 i15626_3_lut_4_lut_4_lut (.I0(reset), .I1(n33697), .I2(\data_in_frame[4] [7]), 
            .I3(neopxl_color[23]), .O(n29632));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i15626_3_lut_4_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i15619_3_lut_4_lut_4_lut (.I0(reset), .I1(n33697), .I2(\data_in_frame[4] [1]), 
            .I3(neopxl_color[17]), .O(n29625));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i15619_3_lut_4_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i15462_3_lut_4_lut (.I0(\data_in_frame[18] [3]), .I1(rx_data[3]), 
            .I2(n40820), .I3(n8_adj_5778), .O(n29468));   // verilog/coms.v(130[12] 305[6])
    defparam i15462_3_lut_4_lut.LUT_INIT = 16'haaca;
    SB_LUT4 i15620_3_lut_4_lut_4_lut (.I0(reset), .I1(n33697), .I2(\data_in_frame[4] [2]), 
            .I3(neopxl_color[18]), .O(n29626));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i15620_3_lut_4_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i15621_3_lut_4_lut_4_lut (.I0(reset), .I1(n33697), .I2(\data_in_frame[4] [3]), 
            .I3(neopxl_color[19]), .O(n29627));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i15621_3_lut_4_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i15623_3_lut_4_lut_4_lut (.I0(reset), .I1(n33697), .I2(\data_in_frame[4] [4]), 
            .I3(neopxl_color[20]), .O(n29629));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i15623_3_lut_4_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i15468_3_lut_4_lut (.I0(\data_in_frame[18] [5]), .I1(rx_data[5]), 
            .I2(n40820), .I3(n8_adj_5778), .O(n29474));   // verilog/coms.v(130[12] 305[6])
    defparam i15468_3_lut_4_lut.LUT_INIT = 16'haaca;
    SB_LUT4 i15624_3_lut_4_lut_4_lut (.I0(reset), .I1(n33697), .I2(\data_in_frame[4] [5]), 
            .I3(neopxl_color[21]), .O(n29630));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i15624_3_lut_4_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i15615_3_lut_4_lut_4_lut (.I0(reset), .I1(n33697), .I2(\data_in_frame[6] [2]), 
            .I3(neopxl_color[2]), .O(n29621));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i15615_3_lut_4_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i15617_3_lut_4_lut_4_lut (.I0(reset), .I1(n33697), .I2(\data_in_frame[5] [7]), 
            .I3(neopxl_color[15]), .O(n29623));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i15617_3_lut_4_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i1_2_lut_4_lut_adj_2120 (.I0(state[0]), .I1(bit_ctr[3]), .I2(n43547), 
            .I3(bit_ctr[4]), .O(n4_adj_5945));   // verilog/neopixel.v(34[12] 116[6])
    defparam i1_2_lut_4_lut_adj_2120.LUT_INIT = 16'hd555;
    SB_LUT4 i15618_3_lut_4_lut_4_lut (.I0(reset), .I1(n33697), .I2(\data_in_frame[4] [0]), 
            .I3(neopxl_color[16]), .O(n29624));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i15618_3_lut_4_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i1_2_lut_adj_2121 (.I0(n36816), .I1(Ki[1]), .I2(GND_net), 
            .I3(GND_net), .O(n131));
    defparam i1_2_lut_adj_2121.LUT_INIT = 16'h8888;
    SB_LUT4 i29704_3_lut (.I0(n944), .I1(n1932), .I2(n1933), .I3(GND_net), 
            .O(n43601));
    defparam i29704_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i15514_3_lut_4_lut (.I0(\data_in_frame[20] [4]), .I1(rx_data[4]), 
            .I2(reset), .I3(n159), .O(n29520));   // verilog/coms.v(130[12] 305[6])
    defparam i15514_3_lut_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i15517_3_lut_4_lut (.I0(\data_in_frame[20] [5]), .I1(rx_data[5]), 
            .I2(reset), .I3(n159), .O(n29523));   // verilog/coms.v(130[12] 305[6])
    defparam i15517_3_lut_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i1_2_lut_adj_2122 (.I0(n36881), .I1(Ki[6]), .I2(GND_net), 
            .I3(GND_net), .O(n490));
    defparam i1_2_lut_adj_2122.LUT_INIT = 16'h8888;
    SB_LUT4 encoder0_position_30__I_0_i1580_3_lut (.I0(n2321), .I1(n2388), 
            .I2(n2346), .I3(GND_net), .O(n2420));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1580_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_2123 (.I0(n1925), .I1(n1926), .I2(n1927), .I3(n1928), 
            .O(n62811));
    defparam i1_4_lut_adj_2123.LUT_INIT = 16'hfffe;
    SB_LUT4 i29814_3_lut (.I0(n950), .I1(n2532), .I2(n2533), .I3(GND_net), 
            .O(n43715));
    defparam i29814_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i1_4_lut_adj_2124 (.I0(n1929), .I1(n43601), .I2(n1930), .I3(n1931), 
            .O(n60405));
    defparam i1_4_lut_adj_2124.LUT_INIT = 16'ha080;
    SB_LUT4 i1_4_lut_adj_2125 (.I0(n1922), .I1(n1923), .I2(n1924), .I3(n62811), 
            .O(n62817));
    defparam i1_4_lut_adj_2125.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_3_lut_adj_2126 (.I0(n2527), .I1(n2528), .I2(n2526), .I3(GND_net), 
            .O(n63131));
    defparam i1_3_lut_adj_2126.LUT_INIT = 16'hfefe;
    SB_LUT4 n71222_bdd_4_lut (.I0(n71222), .I1(\data_out_frame[17] [3]), 
            .I2(\data_out_frame[16] [3]), .I3(byte_transmit_counter[1]), 
            .O(n71225));
    defparam n71222_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_4_lut_adj_2127 (.I0(n2520), .I1(n63131), .I2(n2523), .I3(n2524), 
            .O(n63135));
    defparam i1_4_lut_adj_2127.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_adj_2128 (.I0(n2521), .I1(n2525), .I2(GND_net), .I3(GND_net), 
            .O(n62785));
    defparam i1_2_lut_adj_2128.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_2129 (.I0(n2529), .I1(n43715), .I2(n2530), .I3(n2531), 
            .O(n60438));
    defparam i1_4_lut_adj_2129.LUT_INIT = 16'ha080;
    SB_LUT4 i1_4_lut_adj_2130 (.I0(n1920), .I1(n1921), .I2(n62817), .I3(n60405), 
            .O(n62823));
    defparam i1_4_lut_adj_2130.LUT_INIT = 16'hfffe;
    SB_LUT4 i54763_4_lut (.I0(n1918), .I1(n1917), .I2(n1919), .I3(n62823), 
            .O(n1950));
    defparam i54763_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i14_1_lut (.I0(encoder1_position_scaled[13]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n12_adj_5806));   // verilog/TinyFPGA_B.v(323[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_4_lut_adj_2131 (.I0(state_adj_6008[2]), .I1(state_adj_6008[1]), 
            .I2(state_adj_6008[0]), .I3(n42885), .O(n57800));   // verilog/eeprom.v(35[8] 81[4])
    defparam i1_4_lut_adj_2131.LUT_INIT = 16'ha8e8;
    SB_LUT4 encoder0_position_30__I_0_i1240_3_lut (.I0(n1821), .I1(n1888), 
            .I2(n1851), .I3(GND_net), .O(n1920));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1240_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_2132 (.I0(n2516), .I1(n2515), .I2(n2518), .I3(n2522), 
            .O(n61367));
    defparam i1_4_lut_adj_2132.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_adj_2133 (.I0(n2023), .I1(n2026), .I2(GND_net), .I3(GND_net), 
            .O(n63145));
    defparam i1_2_lut_adj_2133.LUT_INIT = 16'heeee;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i15_1_lut (.I0(encoder1_position_scaled[14]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n11_adj_5817));   // verilog/TinyFPGA_B.v(323[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_55279 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [2]), .I2(\data_out_frame[27] [2]), 
            .I3(byte_transmit_counter[1]), .O(n70994));
    defparam byte_transmit_counter_0__bdd_4_lut_55279.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_4_lut_adj_2134 (.I0(n2519), .I1(n62785), .I2(n2517), .I3(n63135), 
            .O(n62787));
    defparam i1_4_lut_adj_2134.LUT_INIT = 16'hfffe;
    SB_LUT4 mux_1582_i19_3_lut (.I0(duty[21]), .I1(duty[18]), .I2(n260), 
            .I3(GND_net), .O(n12177));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1582_i19_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i1_4_lut_adj_2135 (.I0(n2025), .I1(n2027), .I2(n2028), .I3(n2024), 
            .O(n63147));
    defparam i1_4_lut_adj_2135.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_2136 (.I0(n61367), .I1(n2513), .I2(n2514), .I3(n60438), 
            .O(n61361));
    defparam i1_4_lut_adj_2136.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i16_1_lut (.I0(encoder1_position_scaled[15]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n10_adj_5818));   // verilog/TinyFPGA_B.v(323[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i54704_4_lut (.I0(n61361), .I1(n2511), .I2(n2512), .I3(n62787), 
            .O(n2544));
    defparam i54704_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i29708_3_lut (.I0(n945), .I1(n2032), .I2(n2033), .I3(GND_net), 
            .O(n43605));
    defparam i29708_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i1_4_lut_adj_2137 (.I0(n2021), .I1(n2022), .I2(n63147), .I3(n63145), 
            .O(n63153));
    defparam i1_4_lut_adj_2137.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_30__I_0_i1647_3_lut (.I0(n2420), .I1(n2487), 
            .I2(n2445), .I3(GND_net), .O(n2519));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1647_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_2138 (.I0(n2029), .I1(n43605), .I2(n2030), .I3(n2031), 
            .O(n60442));
    defparam i1_4_lut_adj_2138.LUT_INIT = 16'ha080;
    SB_LUT4 n70994_bdd_4_lut (.I0(n70994), .I1(\data_out_frame[25] [2]), 
            .I2(\data_out_frame[24] [2]), .I3(byte_transmit_counter[1]), 
            .O(n70997));
    defparam n70994_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_adj_2139 (.I0(n2626), .I1(n2628), .I2(GND_net), .I3(GND_net), 
            .O(n63229));
    defparam i1_2_lut_adj_2139.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_2140 (.I0(n2625), .I1(n2621), .I2(n2624), .I3(n2627), 
            .O(n63237));
    defparam i1_4_lut_adj_2140.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_2141 (.I0(n2622), .I1(n63229), .I2(n2620), .I3(n2623), 
            .O(n63239));
    defparam i1_4_lut_adj_2141.LUT_INIT = 16'hfffe;
    SB_LUT4 i29812_3_lut (.I0(n951), .I1(n2632), .I2(n2633), .I3(GND_net), 
            .O(n43713));
    defparam i29812_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i1_4_lut_adj_2142 (.I0(n2019), .I1(n60442), .I2(n2020), .I3(n63153), 
            .O(n63159));
    defparam i1_4_lut_adj_2142.LUT_INIT = 16'hfffe;
    SB_LUT4 i54786_4_lut (.I0(n2017), .I1(n2016), .I2(n2018), .I3(n63159), 
            .O(n2049));
    defparam i54786_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i1_4_lut_adj_2143 (.I0(n2618), .I1(n2619), .I2(n63239), .I3(n63237), 
            .O(n63245));
    defparam i1_4_lut_adj_2143.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_30__I_0_i1307_3_lut (.I0(n1920), .I1(n1987), 
            .I2(n1950), .I3(GND_net), .O(n2019));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1307_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_2144 (.I0(n2629), .I1(n43713), .I2(n2630), .I3(n2631), 
            .O(n60479));
    defparam i1_4_lut_adj_2144.LUT_INIT = 16'ha080;
    SB_LUT4 i1_4_lut_adj_2145 (.I0(n2120), .I1(n2121), .I2(n2123), .I3(n2124), 
            .O(n62867));
    defparam i1_4_lut_adj_2145.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_adj_2146 (.I0(n2127), .I1(n2126), .I2(GND_net), .I3(GND_net), 
            .O(n63039));
    defparam i1_2_lut_adj_2146.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_2147 (.I0(n2616), .I1(n60479), .I2(n2617), .I3(n63245), 
            .O(n63251));
    defparam i1_4_lut_adj_2147.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_2148 (.I0(n2613), .I1(n2614), .I2(n2615), .I3(n63251), 
            .O(n63257));
    defparam i1_4_lut_adj_2148.LUT_INIT = 16'hfffe;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_55274 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[22] [3]), .I2(\data_out_frame[23] [3]), 
            .I3(byte_transmit_counter[1]), .O(n70988));
    defparam byte_transmit_counter_0__bdd_4_lut_55274.LUT_INIT = 16'he4aa;
    SB_LUT4 i54736_4_lut (.I0(n2611), .I1(n2610), .I2(n2612), .I3(n63257), 
            .O(n2643));
    defparam i54736_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i15780_3_lut_4_lut (.I0(\data_in_frame[23] [5]), .I1(rx_data[5]), 
            .I2(reset), .I3(n75), .O(n29786));   // verilog/coms.v(130[12] 305[6])
    defparam i15780_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i1_2_lut_2_lut (.I0(reset), .I1(n75), .I2(GND_net), .I3(GND_net), 
            .O(n28356));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i1_4_lut_4_lut (.I0(\ID_READOUT_FSM.state [0]), .I1(\ID_READOUT_FSM.state [1]), 
            .I2(reset), .I3(n42812), .O(n57200));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_4_lut_4_lut.LUT_INIT = 16'hb1f1;
    SB_LUT4 encoder0_position_30__I_0_i1714_3_lut (.I0(n2519), .I1(n2586), 
            .I2(n2544), .I3(GND_net), .O(n2618));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1714_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i54369_3_lut_3_lut (.I0(\ID_READOUT_FSM.state [0]), .I1(\ID_READOUT_FSM.state [1]), 
            .I2(n42812), .I3(GND_net), .O(n27635));
    defparam i54369_3_lut_3_lut.LUT_INIT = 16'h1515;
    SB_LUT4 i51619_2_lut_3_lut (.I0(n62), .I1(delay_counter[31]), .I2(\ID_READOUT_FSM.state [0]), 
            .I3(GND_net), .O(n66991));
    defparam i51619_2_lut_3_lut.LUT_INIT = 16'hf2f2;
    SB_LUT4 n70988_bdd_4_lut (.I0(n70988), .I1(\data_out_frame[21] [3]), 
            .I2(\data_out_frame[20] [3]), .I3(byte_transmit_counter[1]), 
            .O(n70991));
    defparam n70988_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_3_lut_adj_2149 (.I0(n2721), .I1(n2723), .I2(n2727), .I3(GND_net), 
            .O(n62795));
    defparam i1_3_lut_adj_2149.LUT_INIT = 16'hfefe;
    SB_LUT4 i29049_2_lut_3_lut (.I0(\ID_READOUT_FSM.state [0]), .I1(\ID_READOUT_FSM.state [1]), 
            .I2(n42812), .I3(GND_net), .O(n42941));
    defparam i29049_2_lut_3_lut.LUT_INIT = 16'hfbfb;
    SB_LUT4 i1_2_lut_3_lut_adj_2150 (.I0(n15_adj_5755), .I1(n22835), .I2(dti), 
            .I3(GND_net), .O(n27561));
    defparam i1_2_lut_3_lut_adj_2150.LUT_INIT = 16'hbaba;
    SB_LUT4 i1_2_lut_4_lut_adj_2151 (.I0(delay_counter[17]), .I1(delay_counter[16]), 
            .I2(delay_counter[15]), .I3(delay_counter[14]), .O(n4_adj_5854));
    defparam i1_2_lut_4_lut_adj_2151.LUT_INIT = 16'hfffe;
    SB_LUT4 i15523_4_lut (.I0(CS_MISO_c), .I1(data_adj_6015[1]), .I2(n5_adj_5734), 
            .I3(n25512), .O(n29529));   // verilog/tli4970.v(35[10] 68[6])
    defparam i15523_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i15524_4_lut (.I0(CS_MISO_c), .I1(data_adj_6015[2]), .I2(n5_adj_5824), 
            .I3(n25512), .O(n29530));   // verilog/tli4970.v(35[10] 68[6])
    defparam i15524_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i15532_4_lut (.I0(CS_MISO_c), .I1(data_adj_6015[3]), .I2(n6), 
            .I3(n25499), .O(n29538));   // verilog/tli4970.v(35[10] 68[6])
    defparam i15532_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i15539_4_lut (.I0(CS_MISO_c), .I1(data_adj_6015[4]), .I2(n5_adj_5733), 
            .I3(n25504), .O(n29545));   // verilog/tli4970.v(35[10] 68[6])
    defparam i15539_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i1_3_lut_adj_2152 (.I0(n2722), .I1(n2725), .I2(n2728), .I3(GND_net), 
            .O(n62979));
    defparam i1_3_lut_adj_2152.LUT_INIT = 16'hfefe;
    SB_LUT4 i15540_4_lut (.I0(CS_MISO_c), .I1(data_adj_6015[5]), .I2(n5_adj_5734), 
            .I3(n25504), .O(n29546));   // verilog/tli4970.v(35[10] 68[6])
    defparam i15540_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i29878_4_lut (.I0(n952), .I1(n2731), .I2(n2732), .I3(n2733), 
            .O(n43779));
    defparam i29878_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 i15541_4_lut (.I0(CS_MISO_c), .I1(data_adj_6015[6]), .I2(n5_adj_5824), 
            .I3(n25504), .O(n29547));   // verilog/tli4970.v(35[10] 68[6])
    defparam i15541_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i1_4_lut_adj_2153 (.I0(n2720), .I1(n62979), .I2(n2726), .I3(n2724), 
            .O(n62983));
    defparam i1_4_lut_adj_2153.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_2154 (.I0(n2729), .I1(n62983), .I2(n43779), .I3(n2730), 
            .O(n62985));
    defparam i1_4_lut_adj_2154.LUT_INIT = 16'heccc;
    SB_LUT4 i15542_4_lut (.I0(CS_MISO_c), .I1(data_adj_6015[7]), .I2(n6_adj_5762), 
            .I3(n25499), .O(n29548));   // verilog/tli4970.v(35[10] 68[6])
    defparam i15542_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i15543_4_lut (.I0(CS_MISO_c), .I1(data_adj_6015[8]), .I2(n5_adj_5733), 
            .I3(n25508), .O(n29549));   // verilog/tli4970.v(35[10] 68[6])
    defparam i15543_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i2_2_lut_adj_2155 (.I0(hall2), .I1(commutation_state_7__N_27[2]), 
            .I2(GND_net), .I3(GND_net), .O(commutation_state_7__N_216));   // verilog/TinyFPGA_B.v(166[7:32])
    defparam i2_2_lut_adj_2155.LUT_INIT = 16'h4444;
    SB_LUT4 i15544_4_lut (.I0(CS_MISO_c), .I1(data_adj_6015[9]), .I2(n5_adj_5734), 
            .I3(n25508), .O(n29550));   // verilog/tli4970.v(35[10] 68[6])
    defparam i15544_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i29890_4_lut (.I0(n946), .I1(n2131), .I2(n2132), .I3(n2133), 
            .O(n43791));
    defparam i29890_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 i1_3_lut_adj_2156 (.I0(hall3), .I1(hall2), .I2(hall1), .I3(GND_net), 
            .O(commutation_state_7__N_208[0]));   // verilog/TinyFPGA_B.v(163[4] 165[7])
    defparam i1_3_lut_adj_2156.LUT_INIT = 16'h1414;
    SB_LUT4 i1_4_lut_adj_2157 (.I0(n2122), .I1(n2125), .I2(n63039), .I3(n2128), 
            .O(n63043));
    defparam i1_4_lut_adj_2157.LUT_INIT = 16'hfffe;
    SB_LUT4 i55160_4_lut_4_lut_4_lut (.I0(hall3), .I1(hall1), .I2(commutation_state_7__N_27[2]), 
            .I3(hall2), .O(n7_adj_5959));
    defparam i55160_4_lut_4_lut_4_lut.LUT_INIT = 16'h77fc;
    SB_LUT4 i15551_3_lut (.I0(control_mode[0]), .I1(\data_in_frame[1] [0]), 
            .I2(n22734), .I3(GND_net), .O(n29557));   // verilog/coms.v(130[12] 305[6])
    defparam i15551_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15552_3_lut (.I0(current_limit[0]), .I1(\data_in_frame[21] [0]), 
            .I2(n22734), .I3(GND_net), .O(n29558));   // verilog/coms.v(130[12] 305[6])
    defparam i15552_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_2158 (.I0(n2716), .I1(n2717), .I2(n62985), .I3(n2718), 
            .O(n62991));
    defparam i1_4_lut_adj_2158.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_2159 (.I0(n2712), .I1(n2714), .I2(n2719), .I3(n62795), 
            .O(n62801));
    defparam i1_4_lut_adj_2159.LUT_INIT = 16'hfffe;
    SB_LUT4 i15554_3_lut (.I0(\PID_CONTROLLER.integral [0]), .I1(\PID_CONTROLLER.integral_23__N_3715 [0]), 
            .I2(control_update), .I3(GND_net), .O(n29560));   // verilog/motorControl.v(41[14] 62[8])
    defparam i15554_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_2160 (.I0(n2713), .I1(n2711), .I2(n2715), .I3(n62991), 
            .O(n61707));
    defparam i1_4_lut_adj_2160.LUT_INIT = 16'hfffe;
    SB_LUT4 i15556_4_lut (.I0(CS_MISO_c), .I1(data_adj_6015[10]), .I2(n5_adj_5824), 
            .I3(n25508), .O(n29562));   // verilog/tli4970.v(35[10] 68[6])
    defparam i15556_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i1_4_lut_4_lut_adj_2161 (.I0(\ID_READOUT_FSM.state [0]), .I1(\ID_READOUT_FSM.state [1]), 
            .I2(read_N_409), .I3(n2820), .O(n25_adj_5939));   // verilog/TinyFPGA_B.v(376[7:11])
    defparam i1_4_lut_4_lut_adj_2161.LUT_INIT = 16'h5450;
    SB_LUT4 i15557_4_lut (.I0(CS_MISO_c), .I1(data_adj_6015[11]), .I2(n6_adj_5759), 
            .I3(n25499), .O(n29563));   // verilog/tli4970.v(35[10] 68[6])
    defparam i15557_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i1_4_lut_adj_2162 (.I0(state_adj_6008[2]), .I1(data_ready), 
            .I2(n43543), .I3(n25490), .O(n58190));   // verilog/eeprom.v(35[8] 81[4])
    defparam i1_4_lut_adj_2162.LUT_INIT = 16'hcca8;
    SB_LUT4 i15559_3_lut (.I0(current[0]), .I1(data_adj_6015[0]), .I2(n27643), 
            .I3(GND_net), .O(n29565));   // verilog/tli4970.v(35[10] 68[6])
    defparam i15559_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i54676_4_lut (.I0(n2710), .I1(n2709), .I2(n61707), .I3(n62801), 
            .O(n2742));
    defparam i54676_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i15560_4_lut (.I0(rw), .I1(state_adj_6008[1]), .I2(state_adj_6008[2]), 
            .I3(n5772), .O(n29566));   // verilog/eeprom.v(35[8] 81[4])
    defparam i15560_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 LessThan_11_i6_3_lut_3_lut (.I0(duty[2]), .I1(duty[3]), .I2(current[3]), 
            .I3(GND_net), .O(n6_adj_5753));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i6_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i15561_3_lut (.I0(CS_c), .I1(state_adj_6017[0]), .I2(state_adj_6017[1]), 
            .I3(GND_net), .O(n29567));   // verilog/tli4970.v(35[10] 68[6])
    defparam i15561_3_lut.LUT_INIT = 16'ha3a3;
    SB_LUT4 i55142_4_lut (.I0(n15_adj_5763), .I1(clk_out), .I2(state_adj_6017[0]), 
            .I3(state_adj_6017[1]), .O(n9_adj_5953));   // verilog/tli4970.v(35[10] 68[6])
    defparam i55142_4_lut.LUT_INIT = 16'hc8fc;
    SB_LUT4 LessThan_11_i10_3_lut_3_lut (.I0(duty[5]), .I1(duty[6]), .I2(current[6]), 
            .I3(GND_net), .O(n10_adj_5749));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i10_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 LessThan_11_i8_3_lut_3_lut (.I0(duty[4]), .I1(duty[8]), .I2(current[8]), 
            .I3(GND_net), .O(n8_adj_5751));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i8_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i14795_2_lut (.I0(n27585), .I1(dti), .I2(GND_net), .I3(GND_net), 
            .O(n28807));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    defparam i14795_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i15567_4_lut (.I0(saved_addr[0]), .I1(rw), .I2(n58751), .I3(state_7__N_4110[0]), 
            .O(n29573));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i15567_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i54306_4_lut (.I0(commutation_state[1]), .I1(n22835), .I2(dti), 
            .I3(commutation_state[2]), .O(n27585));
    defparam i54306_4_lut.LUT_INIT = 16'hc5cf;
    SB_LUT4 i15568_3_lut (.I0(current_limit[12]), .I1(\data_in_frame[20] [4]), 
            .I2(n22734), .I3(GND_net), .O(n29574));   // verilog/coms.v(130[12] 305[6])
    defparam i15568_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_2163 (.I0(n23_adj_5860), .I1(o_Rx_DV_N_3488[12]), 
            .I2(n4938), .I3(r_SM_Main_adj_6027[0]), .O(n62099));
    defparam i1_4_lut_adj_2163.LUT_INIT = 16'hfeff;
    SB_LUT4 i1_4_lut_adj_2164 (.I0(o_Rx_DV_N_3488[24]), .I1(n27_adj_5858), 
            .I2(n29_adj_5857), .I3(n62099), .O(n60274));
    defparam i1_4_lut_adj_2164.LUT_INIT = 16'hfffe;
    SB_LUT4 mux_243_i1_3_lut_4_lut (.I0(n25385), .I1(control_mode[1]), .I2(motor_state_23__N_91[0]), 
            .I3(encoder0_position_scaled[0]), .O(motor_state[0]));   // verilog/TinyFPGA_B.v(285[5:22])
    defparam mux_243_i1_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 encoder0_position_30__I_0_i1781_3_lut (.I0(n2618), .I1(n2685), 
            .I2(n2643), .I3(GND_net), .O(n2717));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1781_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_243_i2_3_lut_4_lut (.I0(n25385), .I1(control_mode[1]), .I2(motor_state_23__N_91[1]), 
            .I3(encoder0_position_scaled[1]), .O(motor_state[1]));   // verilog/TinyFPGA_B.v(285[5:22])
    defparam mux_243_i2_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 mux_243_i3_3_lut_4_lut (.I0(n25385), .I1(control_mode[1]), .I2(motor_state_23__N_91[2]), 
            .I3(encoder0_position_scaled[2]), .O(motor_state[2]));   // verilog/TinyFPGA_B.v(285[5:22])
    defparam mux_243_i3_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 i29808_3_lut (.I0(n953), .I1(n2832), .I2(n2833), .I3(GND_net), 
            .O(n43709));
    defparam i29808_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 mux_243_i4_3_lut_4_lut (.I0(n25385), .I1(control_mode[1]), .I2(motor_state_23__N_91[3]), 
            .I3(encoder0_position_scaled[3]), .O(motor_state[3]));   // verilog/TinyFPGA_B.v(285[5:22])
    defparam mux_243_i4_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 n11566_bdd_4_lut (.I0(n11566), .I1(current[15]), .I2(duty[22]), 
            .I3(n11564), .O(n71192));
    defparam n11566_bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n71192_bdd_4_lut (.I0(n71192), .I1(duty[19]), .I2(n4907), 
            .I3(n11564), .O(pwm_setpoint_23__N_3[19]));
    defparam n71192_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_4_lut_adj_2165 (.I0(n2116), .I1(n2117), .I2(n2119), .I3(n62867), 
            .O(n62873));
    defparam i1_4_lut_adj_2165.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_2166 (.I0(n2822), .I1(n2827), .I2(n2824), .I3(n2820_adj_5856), 
            .O(n63277));
    defparam i1_4_lut_adj_2166.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_2167 (.I0(n2821), .I1(n2823), .I2(n2826), .I3(n2825), 
            .O(n63279));
    defparam i1_4_lut_adj_2167.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_2168 (.I0(n63279), .I1(n63277), .I2(n2819), .I3(n2828), 
            .O(n63283));
    defparam i1_4_lut_adj_2168.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_2169 (.I0(n2829), .I1(n43709), .I2(n2830), .I3(n2831), 
            .O(n60489));
    defparam i1_4_lut_adj_2169.LUT_INIT = 16'ha080;
    SB_LUT4 mux_243_i5_3_lut_4_lut (.I0(n25385), .I1(control_mode[1]), .I2(motor_state_23__N_91[4]), 
            .I3(encoder0_position_scaled[4]), .O(motor_state[4]));   // verilog/TinyFPGA_B.v(285[5:22])
    defparam mux_243_i5_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 i1_4_lut_adj_2170 (.I0(n2129), .I1(n63043), .I2(n43791), .I3(n2130), 
            .O(n63045));
    defparam i1_4_lut_adj_2170.LUT_INIT = 16'heccc;
    SB_LUT4 i1_4_lut_adj_2171 (.I0(n2816), .I1(n2817), .I2(n63283), .I3(n2818), 
            .O(n63289));
    defparam i1_4_lut_adj_2171.LUT_INIT = 16'hfffe;
    SB_LUT4 i54812_4_lut (.I0(n63045), .I1(n62873), .I2(n2118), .I3(n2115), 
            .O(n2148));
    defparam i54812_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_30__I_0_i1374_3_lut (.I0(n2019), .I1(n2086), 
            .I2(n2049), .I3(GND_net), .O(n2118));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1374_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_2172 (.I0(n2814), .I1(n2815), .I2(n63289), .I3(n60489), 
            .O(n63295));
    defparam i1_4_lut_adj_2172.LUT_INIT = 16'hfffe;
    SB_LUT4 mux_243_i6_3_lut_4_lut (.I0(n25385), .I1(control_mode[1]), .I2(motor_state_23__N_91[5]), 
            .I3(encoder0_position_scaled[5]), .O(motor_state[5]));   // verilog/TinyFPGA_B.v(285[5:22])
    defparam mux_243_i6_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 encoder0_position_30__I_0_i1441_3_lut (.I0(n2118), .I1(n2185), 
            .I2(n2148), .I3(GND_net), .O(n2217_adj_5853));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1441_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_2173 (.I0(n2811), .I1(n2812), .I2(n2813), .I3(n63295), 
            .O(n63301));
    defparam i1_4_lut_adj_2173.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_2174 (.I0(n2223), .I1(n2225), .I2(n2224), .I3(n2222), 
            .O(n63177));
    defparam i1_4_lut_adj_2174.LUT_INIT = 16'hfffe;
    SB_LUT4 i27715_3_lut_4_lut (.I0(n25385), .I1(control_mode[1]), .I2(n41634), 
            .I3(encoder0_position_scaled[6]), .O(n41635));   // verilog/TinyFPGA_B.v(285[5:22])
    defparam i27715_3_lut_4_lut.LUT_INIT = 16'he0f1;
    SB_LUT4 i15589_3_lut (.I0(\neo_pixel_transmitter.t0 [0]), .I1(timer[0]), 
            .I2(n3157), .I3(GND_net), .O(n29595));   // verilog/neopixel.v(34[12] 116[6])
    defparam i15589_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_243_i8_3_lut_4_lut (.I0(n25385), .I1(control_mode[1]), .I2(motor_state_23__N_91[7]), 
            .I3(encoder0_position_scaled[7]), .O(motor_state[7]));   // verilog/TinyFPGA_B.v(285[5:22])
    defparam mux_243_i8_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 i15596_4_lut (.I0(CS_MISO_c), .I1(data_adj_6015[12]), .I2(n5_adj_5733), 
            .I3(n4_adj_5934), .O(n29602));   // verilog/tli4970.v(35[10] 68[6])
    defparam i15596_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i7470_2_lut (.I0(hall3), .I1(hall2), .I2(GND_net), .I3(GND_net), 
            .O(n20873));   // verilog/TinyFPGA_B.v(160[4] 162[7])
    defparam i7470_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i52122_2_lut_4_lut (.I0(duty[6]), .I1(n304), .I2(duty[5]), 
            .I3(n305), .O(n67816));
    defparam i52122_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i8758_2_lut (.I0(hall3), .I1(hall1), .I2(GND_net), .I3(GND_net), 
            .O(commutation_state_7__N_27[2]));   // verilog/TinyFPGA_B.v(166[4] 168[7])
    defparam i8758_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i43877_3_lut (.I0(n4_adj_5958), .I1(commutation_state_7__N_27[2]), 
            .I2(commutation_state[2]), .I3(GND_net), .O(n59505));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    defparam i43877_3_lut.LUT_INIT = 16'hdcdc;
    SB_LUT4 i54613_4_lut (.I0(n2809), .I1(n2808), .I2(n2810), .I3(n63301), 
            .O(n2841));
    defparam i54613_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i1_4_lut_adj_2175 (.I0(n2226), .I1(n63177), .I2(n2227), .I3(n2228), 
            .O(n63179));
    defparam i1_4_lut_adj_2175.LUT_INIT = 16'hfffe;
    motorControl control (.GND_net(GND_net), .control_update(control_update), 
            .duty({duty}), .clk16MHz(clk16MHz), .reset(reset), .\Ki[11] (Ki[11]), 
            .\PID_CONTROLLER.integral_23__N_3715[0] (\PID_CONTROLLER.integral_23__N_3715 [0]), 
            .\Kp[7] (Kp[7]), .\Kp[1] (Kp[1]), .\Kp[0] (Kp[0]), .\Kp[8] (Kp[8]), 
            .\Kp[9] (Kp[9]), .n43055(n43055), .\Kp[10] (Kp[10]), .\Kp[13] (Kp[13]), 
            .\Kp[2] (Kp[2]), .IntegralLimit({IntegralLimit}), .\Kp[11] (Kp[11]), 
            .n155(n155), .\PID_CONTROLLER.integral_23__N_3715[15] (\PID_CONTROLLER.integral_23__N_3715 [15]), 
            .\Ki[1] (Ki[1]), .\PID_CONTROLLER.integral_23__N_3715[14] (\PID_CONTROLLER.integral_23__N_3715 [14]), 
            .\Ki[0] (Ki[0]), .n367(n367), .VCC_net(VCC_net), .n375(n375), 
            .n376(n376), .\Kp[12] (Kp[12]), .\PID_CONTROLLER.integral ({\PID_CONTROLLER.integral }), 
            .\Ki[2] (Ki[2]), .\Kp[3] (Kp[3]), .\Kp[14] (Kp[14]), .n53(n53), 
            .\Kp[4] (Kp[4]), .\Kp[15] (Kp[15]), .\Kp[5] (Kp[5]), .\Kp[6] (Kp[6]), 
            .\Ki[12] (Ki[12]), .\Ki[13] (Ki[13]), .PWMLimit({PWMLimit}), 
            .\Ki[14] (Ki[14]), .\Ki[15] (Ki[15]), .\Ki[4] (Ki[4]), .n4(n4_adj_5868), 
            .setpoint({setpoint}), .n16(n16_adj_5873), .n3(n3_adj_5874), 
            .n18(n18_adj_5869), .\motor_state[21] (motor_state[21]), .\motor_state[20] (motor_state[20]), 
            .\motor_state[19] (motor_state[19]), .\Ki[5] (Ki[5]), .\motor_state[18] (motor_state[18]), 
            .n28(n28_adj_5855), .\PID_CONTROLLER.integral_23__N_3715[13] (\PID_CONTROLLER.integral_23__N_3715 [13]), 
            .\PID_CONTROLLER.integral_23__N_3715[12] (\PID_CONTROLLER.integral_23__N_3715 [12]), 
            .\Ki[3] (Ki[3]), .n214(n214), .\PID_CONTROLLER.integral_23__N_3715[16] (\PID_CONTROLLER.integral_23__N_3715 [16]), 
            .n29560(n29560), .\Ki[6] (Ki[6]), .\Ki[7] (Ki[7]), .\Ki[8] (Ki[8]), 
            .\Ki[9] (Ki[9]), .\Ki[10] (Ki[10]), .\PID_CONTROLLER.integral_23__N_3715[11] (\PID_CONTROLLER.integral_23__N_3715 [11]), 
            .\motor_state[17] (motor_state[17]), .\PID_CONTROLLER.integral_23__N_3715[10] (\PID_CONTROLLER.integral_23__N_3715 [10]), 
            .n30387(n30387), .n30386(n30386), .n30385(n30385), .n30384(n30384), 
            .n30383(n30383), .n30382(n30382), .n30381(n30381), .n30380(n30380), 
            .n30379(n30379), .n30378(n30378), .n30377(n30377), .n30376(n30376), 
            .n30374(n30374), .n30372(n30372), .n30371(n30371), .n30370(n30370), 
            .n30369(n30369), .n30368(n30368), .n30367(n30367), .n30366(n30366), 
            .n30365(n30365), .n30364(n30364), .n30363(n30363), .\PID_CONTROLLER.integral_23__N_3715[9] (\PID_CONTROLLER.integral_23__N_3715 [9]), 
            .\PID_CONTROLLER.integral_23__N_3715[20] (\PID_CONTROLLER.integral_23__N_3715 [20]), 
            .n36816(n36816), .n20183(n20183), .\PID_CONTROLLER.integral_23__N_3715[8] (\PID_CONTROLLER.integral_23__N_3715 [8]), 
            .\PID_CONTROLLER.integral_23__N_3715[23] (\PID_CONTROLLER.integral_23__N_3715 [23]), 
            .n20(n20_adj_5844), .\motor_state[15] (motor_state[15]), .\motor_state[14] (motor_state[14]), 
            .n490(n490), .n417(n417), .n20136(n20136), .n344(n344), 
            .\motor_state[13] (motor_state[13]), .n20137(n20137), .n271(n271), 
            .n20138(n20138), .n198(n198), .\PID_CONTROLLER.integral_23__N_3715[7] (\PID_CONTROLLER.integral_23__N_3715 [7]), 
            .\motor_state[12] (motor_state[12]), .n56(n56), .n125(n125), 
            .\motor_state[11] (motor_state[11]), .n455(n455), .n456(n456), 
            .\motor_state[10] (motor_state[10]), .\motor_state[9] (motor_state[9]), 
            .\motor_state[8] (motor_state[8]), .\motor_state[7] (motor_state[7]), 
            .n41635(n41635), .\motor_state[5] (motor_state[5]), .\motor_state[4] (motor_state[4]), 
            .\motor_state[3] (motor_state[3]), .\motor_state[2] (motor_state[2]), 
            .\motor_state[1] (motor_state[1]), .\motor_state[0] (motor_state[0]), 
            .n401(n401), .n33(n33), .n361(n361), .\PID_CONTROLLER.integral_23__N_3715[6] (\PID_CONTROLLER.integral_23__N_3715 [6]), 
            .\PID_CONTROLLER.integral_23__N_3715[5] (\PID_CONTROLLER.integral_23__N_3715 [5]), 
            .deadband({deadband}), .n38(n38), .n110(n110), .\PID_CONTROLLER.integral_23__N_3715[4] (\PID_CONTROLLER.integral_23__N_3715 [4]), 
            .\PID_CONTROLLER.integral_23__N_3715[3] (\PID_CONTROLLER.integral_23__N_3715 [3]), 
            .\PID_CONTROLLER.integral_23__N_3715[21] (\PID_CONTROLLER.integral_23__N_3715 [21]), 
            .n37330(n37330), .n11597(n11597), .n131(n131), .n204(n204), 
            .n4_adj_30(n4_adj_5891), .n20182(n20182), .n31(n31_adj_5871), 
            .\PID_CONTROLLER.integral_23__N_3715[22] (\PID_CONTROLLER.integral_23__N_3715 [22]), 
            .n20_adj_31(n20_adj_5870), .n212(n212), .n213(n213), .\PID_CONTROLLER.integral_23__N_3715[2] (\PID_CONTROLLER.integral_23__N_3715 [2]), 
            .n219(n219), .n230(n230), .n19(n19_adj_5866), .\PID_CONTROLLER.integral_23__N_3715[1] (\PID_CONTROLLER.integral_23__N_3715 [1]), 
            .n4_adj_32(n4_adj_5867), .n20181(n20181), .n6(n6_adj_5865), 
            .n36845(n36845), .n20209(n20209), .n6_adj_33(n6_adj_5890), 
            .n27629(n27629)) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(290[16] 302[4])
    SB_LUT4 i52110_2_lut_4_lut (.I0(duty[8]), .I1(n302), .I2(duty[4]), 
            .I3(n306), .O(n67804));
    defparam i52110_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 mux_243_i9_3_lut_4_lut (.I0(n25385), .I1(control_mode[1]), .I2(motor_state_23__N_91[8]), 
            .I3(encoder0_position_scaled[8]), .O(motor_state[8]));   // verilog/TinyFPGA_B.v(285[5:22])
    defparam mux_243_i9_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 LessThan_14_i6_3_lut_3_lut (.I0(current_limit[2]), .I1(current_limit[3]), 
            .I2(current[3]), .I3(GND_net), .O(n6_adj_5705));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam LessThan_14_i6_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 encoder0_position_30__I_0_i1848_3_lut (.I0(n2717), .I1(n2784), 
            .I2(n2742), .I3(GND_net), .O(n2816));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1848_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_243_i10_3_lut_4_lut (.I0(n25385), .I1(control_mode[1]), 
            .I2(motor_state_23__N_91[9]), .I3(encoder0_position_scaled[9]), 
            .O(motor_state[9]));   // verilog/TinyFPGA_B.v(285[5:22])
    defparam mux_243_i10_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 i52158_2_lut_4_lut (.I0(current[8]), .I1(current_limit[8]), 
            .I2(current[4]), .I3(current_limit[4]), .O(n67852));
    defparam i52158_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 LessThan_14_i8_3_lut_3_lut (.I0(current_limit[4]), .I1(current_limit[8]), 
            .I2(current[8]), .I3(GND_net), .O(n8_adj_5703));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam LessThan_14_i8_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i15855_3_lut_4_lut (.I0(\data_in_frame[4] [3]), .I1(rx_data[3]), 
            .I2(reset), .I3(n163), .O(n29861));   // verilog/coms.v(130[12] 305[6])
    defparam i15855_3_lut_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i15609_3_lut (.I0(current_limit[11]), .I1(\data_in_frame[20] [3]), 
            .I2(n22734), .I3(GND_net), .O(n29615));   // verilog/coms.v(130[12] 305[6])
    defparam i15609_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_243_i11_3_lut_4_lut (.I0(n25385), .I1(control_mode[1]), 
            .I2(motor_state_23__N_91[10]), .I3(encoder0_position_scaled[10]), 
            .O(motor_state[10]));   // verilog/TinyFPGA_B.v(285[5:22])
    defparam mux_243_i11_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 mux_243_i12_3_lut_4_lut (.I0(n25385), .I1(control_mode[1]), 
            .I2(motor_state_23__N_91[11]), .I3(encoder0_position_scaled[11]), 
            .O(motor_state[11]));   // verilog/TinyFPGA_B.v(285[5:22])
    defparam mux_243_i12_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 i15610_3_lut (.I0(current_limit[10]), .I1(\data_in_frame[20] [2]), 
            .I2(n22734), .I3(GND_net), .O(n29616));   // verilog/coms.v(130[12] 305[6])
    defparam i15610_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15611_3_lut (.I0(current_limit[9]), .I1(\data_in_frame[20] [1]), 
            .I2(n22734), .I3(GND_net), .O(n29617));   // verilog/coms.v(130[12] 305[6])
    defparam i15611_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15612_3_lut (.I0(current_limit[8]), .I1(\data_in_frame[20] [0]), 
            .I2(n22734), .I3(GND_net), .O(n29618));   // verilog/coms.v(130[12] 305[6])
    defparam i15612_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_i1916_3_lut (.I0(n2817), .I1(n2884), 
            .I2(n2841), .I3(GND_net), .O(n2916));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1916_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_245_i15_4_lut (.I0(encoder1_position_scaled[14]), .I1(displacement[14]), 
            .I2(n15_adj_5722), .I3(n15), .O(motor_state_23__N_91[14]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i15_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i3_4_lut_adj_2176 (.I0(\ID_READOUT_FSM.state [1]), .I1(n62), 
            .I2(delay_counter[31]), .I3(\ID_READOUT_FSM.state [0]), .O(n61826));
    defparam i3_4_lut_adj_2176.LUT_INIT = 16'h0004;
    SB_LUT4 i48610_3_lut (.I0(n4906), .I1(duty[20]), .I2(n11566), .I3(GND_net), 
            .O(n64304));
    defparam i48610_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15852_3_lut_4_lut (.I0(\data_in_frame[4] [2]), .I1(rx_data[2]), 
            .I2(reset), .I3(n163), .O(n29858));   // verilog/coms.v(130[12] 305[6])
    defparam i15852_3_lut_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i48612_3_lut (.I0(n64304), .I1(n64302), .I2(n11564), .I3(GND_net), 
            .O(pwm_setpoint_23__N_3[20]));
    defparam i48612_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48607_3_lut (.I0(n4905), .I1(duty[21]), .I2(n11566), .I3(GND_net), 
            .O(n64301));
    defparam i48607_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48609_3_lut (.I0(n64301), .I1(n64302), .I2(n11564), .I3(GND_net), 
            .O(pwm_setpoint_23__N_3[21]));
    defparam i48609_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48608_3_lut (.I0(current[15]), .I1(duty[23]), .I2(n11566), 
            .I3(GND_net), .O(n64302));
    defparam i48608_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48604_3_lut (.I0(n4904), .I1(duty[22]), .I2(n11566), .I3(GND_net), 
            .O(n64298));
    defparam i48604_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48606_3_lut (.I0(n64298), .I1(n64302), .I2(n11564), .I3(GND_net), 
            .O(pwm_setpoint_23__N_3[22]));
    defparam i48606_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7194_3_lut (.I0(n4903), .I1(current[15]), .I2(n11564), .I3(GND_net), 
            .O(n20877));
    defparam i7194_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7195_3_lut (.I0(n20877), .I1(duty[23]), .I2(n11566), .I3(GND_net), 
            .O(pwm_setpoint_23__N_3[23]));
    defparam i7195_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1582_i20_3_lut (.I0(duty[22]), .I1(duty[19]), .I2(n260), 
            .I3(GND_net), .O(n12175));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1582_i20_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 mux_245_i19_4_lut (.I0(encoder1_position_scaled[18]), .I1(displacement[18]), 
            .I2(n15_adj_5722), .I3(n15), .O(motor_state_23__N_91[18]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i19_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 n11566_bdd_4_lut_55437 (.I0(n11566), .I1(current[15]), .I2(duty[21]), 
            .I3(n11564), .O(n71180));
    defparam n11566_bdd_4_lut_55437.LUT_INIT = 16'he4aa;
    SB_LUT4 mux_243_i21_3_lut_4_lut (.I0(n25385), .I1(control_mode[1]), 
            .I2(motor_state_23__N_91[20]), .I3(encoder0_position_scaled[20]), 
            .O(motor_state[20]));   // verilog/TinyFPGA_B.v(285[5:22])
    defparam mux_243_i21_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 i15849_3_lut_4_lut (.I0(\data_in_frame[4] [1]), .I1(rx_data[1]), 
            .I2(reset), .I3(n163), .O(n29855));   // verilog/coms.v(130[12] 305[6])
    defparam i15849_3_lut_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i15845_3_lut_4_lut (.I0(\data_in_frame[4] [0]), .I1(rx_data[0]), 
            .I2(reset), .I3(n163), .O(n29851));   // verilog/coms.v(130[12] 305[6])
    defparam i15845_3_lut_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 mux_243_i19_3_lut_4_lut (.I0(n25385), .I1(control_mode[1]), 
            .I2(motor_state_23__N_91[18]), .I3(encoder0_position_scaled[18]), 
            .O(motor_state[18]));   // verilog/TinyFPGA_B.v(285[5:22])
    defparam mux_243_i19_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 encoder0_position_30__I_0_i1915_3_lut (.I0(n2816), .I1(n2883), 
            .I2(n2841), .I3(GND_net), .O(n2915));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1915_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i28707_3_lut_4_lut (.I0(n25385), .I1(control_mode[1]), .I2(motor_state_23__N_91[22]), 
            .I3(encoder0_position_scaled[22]), .O(n3_adj_5874));   // verilog/TinyFPGA_B.v(285[5:22])
    defparam i28707_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 n71180_bdd_4_lut (.I0(n71180), .I1(duty[18]), .I2(n4908), 
            .I3(n11564), .O(pwm_setpoint_23__N_3[18]));
    defparam n71180_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i17_3_lut_4_lut (.I0(n25385), .I1(control_mode[1]), .I2(n15_adj_5872), 
            .I3(encoder0_position_scaled[23]), .O(n16_adj_5873));   // verilog/TinyFPGA_B.v(285[5:22])
    defparam i17_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 encoder0_position_30__I_0_i1306_3_lut (.I0(n1919), .I1(n1986), 
            .I2(n1950), .I3(GND_net), .O(n2018));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1306_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1930_3_lut (.I0(n2831), .I1(n2898), 
            .I2(n2841), .I3(GND_net), .O(n2930));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1930_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1373_3_lut (.I0(n2018), .I1(n2085), 
            .I2(n2049), .I3(GND_net), .O(n2117));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1373_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_243_i22_3_lut_4_lut (.I0(n25385), .I1(control_mode[1]), 
            .I2(motor_state_23__N_91[21]), .I3(encoder0_position_scaled[21]), 
            .O(motor_state[21]));   // verilog/TinyFPGA_B.v(285[5:22])
    defparam mux_243_i22_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 i29021_2_lut (.I0(n22835), .I1(dti), .I2(GND_net), .I3(GND_net), 
            .O(n42913));
    defparam i29021_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 dti_counter_1933_mux_6_i1_4_lut (.I0(n45_adj_5889), .I1(n15_adj_5755), 
            .I2(n42913), .I3(dti_counter[0]), .O(n55));   // verilog/TinyFPGA_B.v(174[23:37])
    defparam dti_counter_1933_mux_6_i1_4_lut.LUT_INIT = 16'ha3a0;
    SB_LUT4 mux_243_i20_3_lut_4_lut (.I0(n25385), .I1(control_mode[1]), 
            .I2(motor_state_23__N_91[19]), .I3(encoder0_position_scaled[19]), 
            .O(motor_state[19]));   // verilog/TinyFPGA_B.v(285[5:22])
    defparam mux_243_i20_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 encoder0_position_30__I_0_i1929_3_lut (.I0(n2830), .I1(n2897), 
            .I2(n2841), .I3(GND_net), .O(n2929));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1929_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_243_i18_3_lut_4_lut (.I0(n25385), .I1(control_mode[1]), 
            .I2(motor_state_23__N_91[17]), .I3(encoder0_position_scaled[17]), 
            .O(motor_state[17]));   // verilog/TinyFPGA_B.v(285[5:22])
    defparam mux_243_i18_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 i15616_4_lut (.I0(CS_MISO_c), .I1(data_adj_6015[15]), .I2(n42981), 
            .I3(n25499), .O(n29622));   // verilog/tli4970.v(35[10] 68[6])
    defparam i15616_4_lut.LUT_INIT = 16'hccac;
    SB_LUT4 i1_4_lut_adj_2177 (.I0(n2926), .I1(n2925), .I2(n2928), .I3(n2924), 
            .O(n62883));
    defparam i1_4_lut_adj_2177.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_4_lut_adj_2178 (.I0(control_mode[0]), .I1(n63553), 
            .I2(control_mode[7]), .I3(control_mode[3]), .O(n25385));   // verilog/TinyFPGA_B.v(286[5:22])
    defparam i1_2_lut_4_lut_adj_2178.LUT_INIT = 16'hfffe;
    SB_LUT4 mux_243_i13_3_lut_4_lut (.I0(n25385), .I1(control_mode[1]), 
            .I2(motor_state_23__N_91[12]), .I3(encoder0_position_scaled[12]), 
            .O(motor_state[12]));   // verilog/TinyFPGA_B.v(285[5:22])
    defparam mux_243_i13_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 i1_4_lut_adj_2179 (.I0(n62883), .I1(n2927), .I2(n2920), .I3(n2922), 
            .O(n62885));
    defparam i1_4_lut_adj_2179.LUT_INIT = 16'hfffe;
    SB_LUT4 i29822_3_lut (.I0(n947), .I1(n2232), .I2(n2233), .I3(GND_net), 
            .O(n43723));
    defparam i29822_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i29874_4_lut (.I0(n954), .I1(n2931), .I2(n2932), .I3(n2933), 
            .O(n43775));
    defparam i29874_4_lut.LUT_INIT = 16'hfcec;
    \quadrature_decoder(0)  quad_counter1 (.ENCODER1_B_N_keep(ENCODER1_B_N), 
            .n1779(clk16MHz), .ENCODER1_A_N_keep(ENCODER1_A_N), .n1786(n1786), 
            .GND_net(GND_net), .n1788(n1788), .n1790(n1790), .n1792(n1792), 
            .n1794(n1794), .n1796(n1796), .\encoder1_position[25] (encoder1_position[25]), 
            .\encoder1_position[24] (encoder1_position[24]), .\encoder1_position[23] (encoder1_position[23]), 
            .\encoder1_position[22] (encoder1_position[22]), .\encoder1_position[21] (encoder1_position[21]), 
            .\encoder1_position[20] (encoder1_position[20]), .b_prev(b_prev_adj_5771), 
            .\a_new[1] (a_new_adj_5996[1]), .\encoder1_position[19] (encoder1_position[19]), 
            .\encoder1_position[18] (encoder1_position[18]), .\encoder1_position[17] (encoder1_position[17]), 
            .\encoder1_position[16] (encoder1_position[16]), .\encoder1_position[15] (encoder1_position[15]), 
            .\encoder1_position[14] (encoder1_position[14]), .\encoder1_position[13] (encoder1_position[13]), 
            .\encoder1_position[12] (encoder1_position[12]), .\encoder1_position[11] (encoder1_position[11]), 
            .\encoder1_position[10] (encoder1_position[10]), .\encoder1_position[9] (encoder1_position[9]), 
            .\encoder1_position[8] (encoder1_position[8]), .\encoder1_position[7] (encoder1_position[7]), 
            .\encoder1_position[6] (encoder1_position[6]), .\encoder1_position[5] (encoder1_position[5]), 
            .\encoder1_position[4] (encoder1_position[4]), .\encoder1_position[3] (encoder1_position[3]), 
            .\encoder1_position[2] (encoder1_position[2]), .n1822(n1822), 
            .n1824(n1824), .VCC_net(VCC_net), .n29649(n29649), .a_prev(a_prev_adj_5770), 
            .n29614(n29614), .n1784(n1784), .position_31__N_3836(position_31__N_3836_adj_5773), 
            .\b_new[1] (b_new_adj_5997[1]), .n29402(n29402), .debounce_cnt_N_3833(debounce_cnt_N_3833_adj_5772)) /* synthesis lattice_noprune=1 */ ;   // verilog/TinyFPGA_B.v(312[27] 318[6])
    SB_LUT4 i1_4_lut_adj_2180 (.I0(n2219), .I1(n2220), .I2(n63179), .I3(n2221), 
            .O(n63185));
    defparam i1_4_lut_adj_2180.LUT_INIT = 16'hfffe;
    SB_LUT4 mux_243_i15_3_lut_4_lut (.I0(n25385), .I1(control_mode[1]), 
            .I2(motor_state_23__N_91[14]), .I3(encoder0_position_scaled[14]), 
            .O(motor_state[14]));   // verilog/TinyFPGA_B.v(285[5:22])
    defparam mux_243_i15_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 i1_4_lut_adj_2181 (.I0(n2229), .I1(n43723), .I2(n2230), .I3(n2231), 
            .O(n60449));
    defparam i1_4_lut_adj_2181.LUT_INIT = 16'ha080;
    SB_LUT4 i1_2_lut_4_lut_adj_2182 (.I0(\data_out_frame[20] [6]), .I1(\data_out_frame[20] [7]), 
            .I2(\data_out_frame[20] [4]), .I3(n59223), .O(n2217));   // verilog/coms.v(100[12:26])
    defparam i1_2_lut_4_lut_adj_2182.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_2183 (.I0(n2217_adj_5853), .I1(n2218), .I2(n60449), 
            .I3(n63185), .O(n63191));
    defparam i1_4_lut_adj_2183.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_2184 (.I0(n2917), .I1(n2918), .I2(n2919), .I3(n62885), 
            .O(n62891));
    defparam i1_4_lut_adj_2184.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_2185 (.I0(n62891), .I1(n2929), .I2(n43775), .I3(n2930), 
            .O(n62893));
    defparam i1_4_lut_adj_2185.LUT_INIT = 16'heaaa;
    SB_LUT4 i54837_4_lut (.I0(n2215), .I1(n2214), .I2(n2216), .I3(n63191), 
            .O(n2247));
    defparam i54837_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i1_4_lut_adj_2186 (.I0(n2913), .I1(n2915), .I2(n2916), .I3(n62893), 
            .O(n62899));
    defparam i1_4_lut_adj_2186.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_30__I_0_i1442_3_lut (.I0(n2119), .I1(n2186), 
            .I2(n2148), .I3(GND_net), .O(n2218));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1442_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15627_3_lut (.I0(control_mode[1]), .I1(\data_in_frame[1] [1]), 
            .I2(n22734), .I3(GND_net), .O(n29633));   // verilog/coms.v(130[12] 305[6])
    defparam i15627_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15628_3_lut (.I0(control_mode[2]), .I1(\data_in_frame[1] [2]), 
            .I2(n22734), .I3(GND_net), .O(n29634));   // verilog/coms.v(130[12] 305[6])
    defparam i15628_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_2187 (.I0(n2914), .I1(n2912), .I2(n2923), .I3(n2921), 
            .O(n61577));
    defparam i1_4_lut_adj_2187.LUT_INIT = 16'hfffe;
    SB_LUT4 mux_243_i16_3_lut_4_lut (.I0(n25385), .I1(control_mode[1]), 
            .I2(motor_state_23__N_91[15]), .I3(encoder0_position_scaled[15]), 
            .O(motor_state[15]));   // verilog/TinyFPGA_B.v(285[5:22])
    defparam mux_243_i16_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 i21_3_lut_4_lut (.I0(n25385), .I1(control_mode[1]), .I2(n19_adj_5843), 
            .I3(encoder0_position_scaled[16]), .O(n20_adj_5844));   // verilog/TinyFPGA_B.v(285[5:22])
    defparam i21_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 i1_4_lut_adj_2188 (.I0(n2910), .I1(n61577), .I2(n2911), .I3(n62899), 
            .O(n62905));
    defparam i1_4_lut_adj_2188.LUT_INIT = 16'hfffe;
    SB_LUT4 mux_243_i14_3_lut_4_lut (.I0(n25385), .I1(control_mode[1]), 
            .I2(motor_state_23__N_91[13]), .I3(encoder0_position_scaled[13]), 
            .O(motor_state[13]));   // verilog/TinyFPGA_B.v(285[5:22])
    defparam mux_243_i14_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 encoder0_position_30__I_0_i976_3_lut (.I0(n1429), .I1(n1496), 
            .I2(n1455), .I3(GND_net), .O(n1528));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i976_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i54582_4_lut (.I0(n2908), .I1(n2907), .I2(n2909), .I3(n62905), 
            .O(n2940));
    defparam i54582_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_30__I_0_i1509_3_lut (.I0(n2218), .I1(n2285), 
            .I2(n2247), .I3(GND_net), .O(n2317));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1509_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15629_3_lut (.I0(control_mode[3]), .I1(\data_in_frame[1] [3]), 
            .I2(n22734), .I3(GND_net), .O(n29635));   // verilog/coms.v(130[12] 305[6])
    defparam i15629_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15630_3_lut (.I0(control_mode[4]), .I1(\data_in_frame[1] [4]), 
            .I2(n22734), .I3(GND_net), .O(n29636));   // verilog/coms.v(130[12] 305[6])
    defparam i15630_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_i1913_3_lut (.I0(n2814), .I1(n2881), 
            .I2(n2841), .I3(GND_net), .O(n2913));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1913_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1980_3_lut (.I0(n2913), .I1(n2980), 
            .I2(n2940), .I3(GND_net), .O(n3012));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1980_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15631_3_lut (.I0(current_limit[7]), .I1(\data_in_frame[21] [7]), 
            .I2(n22734), .I3(GND_net), .O(n29637));   // verilog/coms.v(130[12] 305[6])
    defparam i15631_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i28910_2_lut (.I0(pwm_out), .I1(GHB), .I2(GND_net), .I3(GND_net), 
            .O(INHB_c_0));   // verilog/TinyFPGA_B.v(90[16:31])
    defparam i28910_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i29039_2_lut (.I0(pwm_out), .I1(GHA), .I2(GND_net), .I3(GND_net), 
            .O(INHA_c_0));   // verilog/TinyFPGA_B.v(88[16:31])
    defparam i29039_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i17_1_lut (.I0(encoder1_position_scaled[16]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n9_adj_5819));   // verilog/TinyFPGA_B.v(323[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i18_1_lut (.I0(encoder1_position_scaled[17]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n8_adj_5820));   // verilog/TinyFPGA_B.v(323[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    coms neopxl_color_23__I_0 (.n29895(n29895), .VCC_net(VCC_net), .\data_in_frame[5] ({\data_in_frame[5] }), 
         .clk16MHz(clk16MHz), .GND_net(GND_net), .n29892(n29892), .\data_out_frame[6] ({\data_out_frame[6] }), 
         .\data_out_frame[5] ({\data_out_frame[5] }), .\data_out_frame[4] ({\data_out_frame[4] }), 
         .\Ki[7] (Ki[7]), .n2873(n2873), .\data_out_frame[8] ({\data_out_frame[8] }), 
         .n58623(n58623), .n58622(n58622), .n29583(n29583), .\data_in_frame[21] ({\data_in_frame[21] }), 
         .\data_out_frame[18] ({\data_out_frame[18] }), .\FRAME_MATCHER.i_31__N_2509 (\FRAME_MATCHER.i_31__N_2509 ), 
         .displacement({displacement}), .\Ki[6] (Ki[6]), .\FRAME_MATCHER.state[3] (\FRAME_MATCHER.state [3]), 
         .\data_out_frame[25] ({\data_out_frame[25] }), .n8(n8_adj_5946), 
         .\data_out_frame[22] ({\data_out_frame[22] }), .\Ki[5] (Ki[5]), 
         .\data_out_frame[23] ({\data_out_frame[23] }), .n59477(n59477), 
         .\data_out_frame[19] ({\data_out_frame[19] }), .n53457(n53457), 
         .n58957(n58957), .\Ki[4] (Ki[4]), .n59223(n59223), .\data_out_frame[16] ({\data_out_frame[16] }), 
         .\data_out_frame[24] ({\data_out_frame[24] }), .n59452(n59452), 
         .n59455(n59455), .n58938(n58938), .n29890(n29890), .n25(n25_adj_5943), 
         .n30(n30_adj_5940), .n26(n26_adj_5942), .n54456(n54456), .n53546(n53546), 
         .\data_out_frame[21] ({\data_out_frame[21] }), .\Ki[3] (Ki[3]), 
         .\Ki[2] (Ki[2]), .\data_out_frame[20] ({\data_out_frame[20] }), 
         .\data_out_frame[17] ({\data_out_frame[17] }), .pwm_setpoint({pwm_setpoint}), 
         .n59241(n59241), .n59406(n59406), .n58978(n58978), .n29885(n29885), 
         .n29881(n29881), .n29878(n29878), .\data_in_frame[4] ({\data_in_frame[4] }), 
         .n57914(n57914), .n57916(n57916), .n57918(n57918), .\Ki[1] (Ki[1]), 
         .n29861(n29861), .n29858(n29858), .n29855(n29855), .\Kp[15] (Kp[15]), 
         .\Kp[14] (Kp[14]), .n29851(n29851), .\data_in_frame[3][6] (\data_in_frame[3] [6]), 
         .\data_in_frame[3][5] (\data_in_frame[3] [5]), .\Kp[13] (Kp[13]), 
         .\Kp[12] (Kp[12]), .\Kp[11] (Kp[11]), .\Kp[10] (Kp[10]), .encoder0_position_scaled({encoder0_position_scaled}), 
         .\Kp[9] (Kp[9]), .\data_out_frame[15] ({\data_out_frame[15] }), 
         .n59124(n59124), .\Kp[8] (Kp[8]), .n58621(n58621), .\data_out_frame[12] ({\data_out_frame[12] }), 
         .\Kp[7] (Kp[7]), .\data_out_frame[13] ({\data_out_frame[13] }), 
         .n59274(n59274), .n58620(n58620), .\Kp[6] (Kp[6]), .\data_out_frame[14] ({\data_out_frame[14] }), 
         .\Kp[5] (Kp[5]), .\Kp[4] (Kp[4]), .n58671(n58671), .\Kp[3] (Kp[3]), 
         .\Kp[2] (Kp[2]), .n70020(n70020), .reset(reset), .setpoint({setpoint}), 
         .\Kp[1] (Kp[1]), .n2076(n2076), .n25764(n25764), .\data_in_frame[11] ({\data_in_frame[11] }), 
         .IntegralLimit({IntegralLimit}), .n58619(n58619), .n54490(n54490), 
         .\data_out_frame[9] ({\data_out_frame[9] }), .n58495(n58495), .n2217(n2217), 
         .n58618(n58618), .n58617(n58617), .n58616(n58616), .n58615(n58615), 
         .n58614(n58614), .n58613(n58613), .n58612(n58612), .\data_out_frame[10] ({\data_out_frame[10] }), 
         .n58611(n58611), .n58610(n58610), .n58609(n58609), .n58608(n58608), 
         .n58607(n58607), .n58606(n58606), .n58605(n58605), .n58604(n58604), 
         .\data_out_frame[11] ({\data_out_frame[11] }), .n58603(n58603), 
         .n58602(n58602), .n58601(n58601), .n58600(n58600), .n58599(n58599), 
         .n58598(n58598), .n58597(n58597), .n58596(n58596), .n58595(n58595), 
         .n58594(n58594), .n58593(n58593), .n58592(n58592), .n58591(n58591), 
         .n58590(n58590), .n58589(n58589), .n58588(n58588), .\data_in_frame[12] ({\data_in_frame[12] }), 
         .n30494(n30494), .n28975(n28975), .\byte_transmit_counter[2] (byte_transmit_counter[2]), 
         .n58587(n58587), .\data_in_frame[16] ({\data_in_frame[16] }), .deadband({deadband}), 
         .n58586(n58586), .\byte_transmit_counter[1] (byte_transmit_counter[1]), 
         .\byte_transmit_counter[0] (byte_transmit_counter[0]), .n58585(n58585), 
         .n58887(n58887), .\data_out_frame[7] ({\data_out_frame[7] }), .n36(n36), 
         .n26143(n26143), .n26376(n26376), .n58584(n58584), .n58583(n58583), 
         .n58582(n58582), .n58581(n58581), .n58580(n58580), .n58579(n58579), 
         .n58578(n58578), .n58577(n58577), .n58576(n58576), .n58575(n58575), 
         .n58574(n58574), .n58573(n58573), .n30510(n30510), .n28959(n28959), 
         .\data_in_frame[1] ({\data_in_frame[1] }), .n26210(n26210), .n29786(n29786), 
         .\data_in_frame[23] ({\data_in_frame[23] }), .n53515(n53515), .n54620(n54620), 
         .n29771(n29771), .\data_in_frame[0] ({\data_in_frame[0] [7], Open_4, 
         Open_5, Open_6, Open_7, Open_8, \data_in_frame[0] [1], Open_9}), 
         .n29639(n29639), .n29650(n29650), .\data_in_frame[0][3] (\data_in_frame[0] [3]), 
         .n29765(n29765), .n29764(n29764), .n57968(n57968), .n29668(n29668), 
         .n29674(n29674), .n29756(n29756), .\data_in_frame[0][6] (\data_in_frame[0] [6]), 
         .n59055(n59055), .\FRAME_MATCHER.i[0] (\FRAME_MATCHER.i [0]), .n43501(n43501), 
         .n163(n163), .rx_data({rx_data}), .n59027(n59027), .n22(n22_adj_5944), 
         .neopxl_color({neopxl_color}), .n7(n7_adj_5957), .encoder1_position_scaled({encoder1_position_scaled}), 
         .n15(n15_adj_5722), .n15_adj_11(n15), .n19(n19_adj_5843), .\data_out_frame[1][1] (\data_out_frame[1] [1]), 
         .\data_out_frame[3][1] (\data_out_frame[3] [1]), .PWMLimit({PWMLimit}), 
         .n28(n28_adj_5855), .n375(n375), .n376(n376), .n4(n4_adj_5868), 
         .n58572(n58572), .n58571(n58571), .n58570(n58570), .n58569(n58569), 
         .n58568(n58568), .\data_in_frame[6] ({\data_in_frame[6] }), .\data_in_frame[8] ({\data_in_frame[8] }), 
         .n58567(n58567), .n58566(n58566), .n58565(n58565), .n58564(n58564), 
         .n58496(n58496), .n58499(n58499), .\data_out_frame[0][3] (\data_out_frame[0] [3]), 
         .\data_out_frame[1][3] (\data_out_frame[1] [3]), .n28947(n28947), 
         .\data_out_frame[3][3] (\data_out_frame[3] [3]), .n58500(n58500), 
         .n28945(n28945), .n58501(n58501), .n58503(n58503), .\Ki[8] (Ki[8]), 
         .\Ki[9] (Ki[9]), .\Ki[10] (Ki[10]), .\Ki[11] (Ki[11]), .\Ki[12] (Ki[12]), 
         .\Ki[13] (Ki[13]), .n58505(n58505), .\Ki[14] (Ki[14]), .\Ki[15] (Ki[15]), 
         .n58507(n58507), .n58508(n58508), .n58509(n58509), .n58510(n58510), 
         .n58511(n58511), .n58512(n58512), .n58513(n58513), .n71165(n71165), 
         .n71003(n71003), .n58514(n58514), .n58515(n58515), .n58493(n58493), 
         .n58516(n58516), .n58517(n58517), .n28929(n28929), .n28928(n28928), 
         .n58518(n58518), .n58519(n58519), .n58520(n58520), .\data_out_frame[1][6] (\data_out_frame[1] [6]), 
         .\data_out_frame[3][6] (\data_out_frame[3] [6]), .n29643(n29643), 
         .\FRAME_MATCHER.rx_data_ready_prev (\FRAME_MATCHER.rx_data_ready_prev ), 
         .n29642(n29642), .n61932(n61932), .n29638(n29638), .\data_out_frame[1][7] (\data_out_frame[1] [7]), 
         .\data_out_frame[3][7] (\data_out_frame[3] [7]), .n29637(n29637), 
         .current_limit({current_limit}), .n29636(n29636), .control_mode({control_mode}), 
         .n29635(n29635), .n29634(n29634), .n29633(n29633), .n29632(n29632), 
         .n29631(n29631), .n29630(n29630), .n29629(n29629), .n29627(n29627), 
         .n29626(n29626), .n29625(n29625), .n29624(n29624), .n29623(n29623), 
         .n58521(n58521), .\data_out_frame[1][0] (\data_out_frame[1] [0]), 
         .n58522(n58522), .n58523(n58523), .n29621(n29621), .n71225(n71225), 
         .n70991(n70991), .\FRAME_MATCHER.i[3] (\FRAME_MATCHER.i [3]), .\FRAME_MATCHER.i[4] (\FRAME_MATCHER.i [4]), 
         .n8_adj_12(n8_adj_5801), .n29618(n29618), .n29617(n29617), .n29616(n29616), 
         .n29615(n29615), .n29613(n29613), .n29612(n29612), .n29608(n29608), 
         .n29607(n29607), .n29606(n29606), .n29605(n29605), .n29604(n29604), 
         .n29582(n29582), .n29574(n29574), .n29558(n29558), .n29557(n29557), 
         .n29556(n29556), .\Ki[0] (Ki[0]), .\Kp[0] (Kp[0]), .n28921(n28921), 
         .n58524(n58524), .n58525(n58525), .n58526(n58526), .n58527(n58527), 
         .n58528(n58528), .n58529(n58529), .n58530(n58530), .n58531(n58531), 
         .n58532(n58532), .n58533(n58533), .n58534(n58534), .n58535(n58535), 
         .n58536(n58536), .n58492(n58492), .n58537(n58537), .n58538(n58538), 
         .n58539(n58539), .n28903(n28903), .n58540(n58540), .n58541(n58541), 
         .n58494(n58494), .n58542(n58542), .n58543(n58543), .n58544(n58544), 
         .\FRAME_MATCHER.i[5] (\FRAME_MATCHER.i [5]), .tx_active(tx_active), 
         .n58545(n58545), .n28895(n28895), .n28894(n28894), .n58546(n58546), 
         .\data_out_frame[0][4] (\data_out_frame[0] [4]), .n22734(n22734), 
         .\data_out_frame[3][4] (\data_out_frame[3] [4]), .ID({ID}), .\data_out_frame[0][2] (\data_out_frame[0] [2]), 
         .n58670(n58670), .n58669(n58669), .n58668(n58668), .n58667(n58667), 
         .n59299(n59299), .\data_out_frame[26][2] (\data_out_frame[26] [2]), 
         .n30439(n30439), .n30438(n30438), .n30437(n30437), .n30421(n30421), 
         .\data_in_frame[0][0] (\data_in_frame[0] [0]), .n30391(n30391), 
         .n30305(n30305), .n30273(n30273), .n29898(n29898), .n29901(n29901), 
         .n57890(n57890), .n57886(n57886), .n30255(n30255), .n29417(n29417), 
         .n29420(n29420), .n29423(n29423), .n29426(n29426), .n57882(n57882), 
         .n29432(n29432), .n57878(n57878), .\data_in_frame[17] ({\data_in_frame[17] }), 
         .n57876(n57876), .n57874(n57874), .n57872(n57872), .n57868(n57868), 
         .n57864(n57864), .n57860(n57860), .n57856(n57856), .n57852(n57852), 
         .\data_in_frame[18] ({\data_in_frame[18] }), .n57850(n57850), .n29930(n29930), 
         .\data_in_frame[7] ({Open_10, Open_11, \data_in_frame[7] [5:0]}), 
         .n30218(n30218), .n29934(n29934), .n29937(n29937), .n29940(n29940), 
         .n58666(n58666), .n29943(n29943), .n29946(n29946), .n57846(n57846), 
         .n29955(n29955), .n29958(n29958), .n29961(n29961), .n29964(n29964), 
         .n30205(n30205), .n29970(n29970), .n29973(n29973), .n29976(n29976), 
         .n30199(n30199), .n30198(n30198), .n30030(n30030), .n58665(n58665), 
         .n58106(n58106), .n58108(n58108), .n58060(n58060), .n30043(n30043), 
         .n30046(n30046), .n30049(n30049), .n30053(n30053), .n30056(n30056), 
         .n30059(n30059), .n30062(n30062), .n57932(n57932), .n57936(n57936), 
         .n30072(n30072), .n30169(n30169), .n30075(n30075), .n30079(n30079), 
         .n57996(n57996), .n30110(n30110), .n30154(n30154), .n29468(n29468), 
         .\data_out_frame[1][5] (\data_out_frame[1] [5]), .n58664(n58664), 
         .n57842(n57842), .n29474(n29474), .n57838(n57838), .n57834(n57834), 
         .n58663(n58663), .n57986(n57986), .\data_in_frame[20] ({\data_in_frame[20] }), 
         .n57980(n57980), .n29520(n29520), .n29523(n29523), .n57974(n57974), 
         .n29535(n29535), .n29539(n29539), .n29542(n29542), .n29551(n29551), 
         .\data_out_frame[27][2] (\data_out_frame[27] [2]), .n29570(n29570), 
         .n58662(n58662), .n58661(n58661), .n58660(n58660), .n58659(n58659), 
         .n58658(n58658), .n29575(n29575), .n58657(n58657), .n58506(n58506), 
         .n58656(n58656), .n58655(n58655), .n58654(n58654), .n58653(n58653), 
         .n58652(n58652), .n58651(n58651), .n58650(n58650), .n58649(n58649), 
         .n58648(n58648), .n58647(n58647), .n29578(n29578), .n58646(n58646), 
         .n58645(n58645), .n58644(n58644), .n58643(n58643), .n58642(n58642), 
         .n58641(n58641), .n58640(n58640), .n58639(n58639), .n58638(n58638), 
         .n58637(n58637), .n58636(n58636), .n58635(n58635), .n58634(n58634), 
         .n58633(n58633), .n58632(n58632), .n29410(n29410), .n160(n160), 
         .n58547(n58547), .n29405(n29405), .n29403(n29403), .n70997(n70997), 
         .n159(n159), .n58548(n58548), .n58549(n58549), .n58550(n58550), 
         .n58551(n58551), .n58552(n58552), .n58553(n58553), .n58504(n58504), 
         .n58498(n58498), .n58554(n58554), .n58555(n58555), .n58556(n58556), 
         .n58557(n58557), .n58558(n58558), .n58497(n58497), .n58502(n58502), 
         .n58559(n58559), .n58631(n58631), .n58630(n58630), .n58629(n58629), 
         .n58628(n58628), .n58560(n58560), .n58561(n58561), .n58562(n58562), 
         .n58563(n58563), .LED_c(LED_c), .DE_c(DE_c), .n58627(n58627), 
         .n58626(n58626), .n58625(n58625), .n58624(n58624), .\pwm_counter[22] (pwm_counter[22]), 
         .n45(n45), .\pwm_counter[21] (pwm_counter[21]), .n43(n43), .n8_adj_13(n8_adj_5778), 
         .n59638(n59638), .\duty[3] (duty[3]), .\duty[0] (duty[0]), .n260(n260), 
         .n7_adj_14(n7_adj_5826), .n54113(n54113), .n8_adj_15(n8_adj_5798), 
         .n59430(n59430), .n40820(n40820), .n455(n455), .n11597(n11597), 
         .n37330(n37330), .n26282(n26282), .n59007(n59007), .n59215(n59215), 
         .n58805(n58805), .n59153(n59153), .n25700(n25700), .n58928(n58928), 
         .n87(n87), .n75(n75), .n33697(n33697), .n98(n98), .rx_data_ready(rx_data_ready), 
         .Kp_23__N_748(Kp_23__N_748), .n28309(n28309), .n28311(n28311), 
         .n367(n367), .n19_adj_16(n19_adj_5866), .n361(n361), .n31(n31_adj_5871), 
         .n28313(n28313), .n43503(n43503), .n18(n18_adj_5869), .n20(n20_adj_5870), 
         .n230(n230), .n155(n155), .\PID_CONTROLLER.integral_23__N_3715[1] (\PID_CONTROLLER.integral_23__N_3715 [1]), 
         .n161(n161), .n58418(n58418), .n59644(n59644), .n33(n33), .n401(n401), 
         .n4_adj_17(n4_adj_5867), .n26372(n26372), .n28307(n28307), .\current[7] (current[7]), 
         .\current[6] (current[6]), .\current[5] (current[5]), .\current[4] (current[4]), 
         .\current[3] (current[3]), .\current[2] (current[2]), .\current[1] (current[1]), 
         .\current[0] (current[0]), .\current[15] (current[15]), .n456(n456), 
         .n27629(n27629), .\current[11] (current[11]), .\current[10] (current[10]), 
         .\current[9] (current[9]), .\current[8] (current[8]), .n63789(n63789), 
         .n63793(n63793), .n67140(n67140), .n7_adj_18(n7_adj_5956), .n28385(n28385), 
         .n70919(n70919), .r_SM_Main({r_SM_Main_adj_6027}), .tx_o(tx_o), 
         .r_Clock_Count({r_Clock_Count_adj_6028}), .n4938(n4938), .n29(n29_adj_5857), 
         .n23(n23_adj_5860), .\o_Rx_DV_N_3488[12] (o_Rx_DV_N_3488[12]), 
         .\o_Rx_DV_N_3488[24] (o_Rx_DV_N_3488[24]), .n27(n27_adj_5858), 
         .n29581(n29581), .\r_SM_Main_2__N_3536[1] (r_SM_Main_2__N_3536[1]), 
         .n59648(n59648), .n60274(n60274), .n6(n6_adj_5935), .tx_enable(tx_enable), 
         .baudrate({baudrate}), .r_Clock_Count_adj_29({r_Clock_Count}), 
         .\o_Rx_DV_N_3488[2] (o_Rx_DV_N_3488[2]), .\o_Rx_DV_N_3488[1] (o_Rx_DV_N_3488[1]), 
         .\o_Rx_DV_N_3488[3] (o_Rx_DV_N_3488[3]), .\o_Rx_DV_N_3488[4] (o_Rx_DV_N_3488[4]), 
         .\o_Rx_DV_N_3488[5] (o_Rx_DV_N_3488[5]), .\o_Rx_DV_N_3488[6] (o_Rx_DV_N_3488[6]), 
         .\o_Rx_DV_N_3488[8] (o_Rx_DV_N_3488[8]), .\o_Rx_DV_N_3488[7] (o_Rx_DV_N_3488[7]), 
         .\r_Bit_Index[0] (r_Bit_Index[0]), .n61449(n61449), .n62163(n62163), 
         .\r_SM_Main_2__N_3446[1] (r_SM_Main_2__N_3446[1]), .r_Rx_Data(r_Rx_Data), 
         .\r_SM_Main[1]_adj_27 (r_SM_Main[1]), .\r_SM_Main[2]_adj_28 (r_SM_Main[2]), 
         .RX_N_2(RX_N_2), .n25515(n25515), .n62091(n62091), .n60815(n60815), 
         .n62089(n62089), .\o_Rx_DV_N_3488[0] (o_Rx_DV_N_3488[0]), .n4935(n4935), 
         .n27901(n27901), .n59702(n59702), .n62513(n62513), .n62417(n62417), 
         .n62465(n62465), .n62401(n62401), .n30420(n30420), .n54640(n54640), 
         .n30416(n30416), .n62433(n62433), .n30126(n30126), .n30125(n30125), 
         .n30124(n30124), .n30123(n30123), .n30122(n30122), .n30121(n30121), 
         .n30120(n30120), .n62481(n62481), .n58684(n58684), .n62497(n62497), 
         .n62449(n62449), .n27661(n27661)) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(255[22] 280[4])
    SB_LUT4 i15641_3_lut (.I0(b_prev), .I1(b_new[1]), .I2(debounce_cnt_N_3833), 
            .I3(GND_net), .O(n29647));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    defparam i15641_3_lut.LUT_INIT = 16'hacac;
    pwm PWM (.n2873(n2873), .pwm_out(pwm_out), .clk32MHz(clk32MHz), .reset(reset), 
        .\pwm_counter[22] (pwm_counter[22]), .\pwm_counter[21] (pwm_counter[21]), 
        .\pwm_counter[12] (pwm_counter[12]), .pwm_setpoint({pwm_setpoint}), 
        .GND_net(GND_net), .VCC_net(VCC_net), .n25(n25_adj_5864), .n45(n45), 
        .n43(n43)) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(97[6] 102[3])
    SB_LUT4 i1_2_lut_3_lut_adj_2189 (.I0(\data_out_frame[14] [4]), .I1(n59124), 
            .I2(n59452), .I3(GND_net), .O(n6_adj_5924));
    defparam i1_2_lut_3_lut_adj_2189.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_2190 (.I0(\data_out_frame[16] [5]), .I1(\data_out_frame[20] [6]), 
            .I2(\data_out_frame[20] [7]), .I3(GND_net), .O(n59359));
    defparam i1_2_lut_3_lut_adj_2190.LUT_INIT = 16'h9696;
    pll32MHz pll32MHz_inst (.GND_net(GND_net), .clk16MHz(clk16MHz), .VCC_net(VCC_net), 
            .clk32MHz(clk32MHz)) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(34[10] 38[2])
    SB_LUT4 i15642_3_lut (.I0(a_prev), .I1(a_new[1]), .I2(debounce_cnt_N_3833), 
            .I3(GND_net), .O(n29648));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    defparam i15642_3_lut.LUT_INIT = 16'hacac;
    \quadrature_decoder(0)_U0  quad_counter0 (.n1744(n1744), .GND_net(GND_net), 
            .\encoder0_position[30] (encoder0_position[30]), .\encoder0_position[29] (encoder0_position[29]), 
            .ENCODER0_B_N_keep(ENCODER0_B_N), .n1779(clk16MHz), .ENCODER0_A_N_keep(ENCODER0_A_N), 
            .\encoder0_position[28] (encoder0_position[28]), .\encoder0_position[27] (encoder0_position[27]), 
            .\encoder0_position[26] (encoder0_position[26]), .\encoder0_position[25] (encoder0_position[25]), 
            .\encoder0_position[24] (encoder0_position[24]), .b_prev(b_prev), 
            .\a_new[1] (a_new[1]), .\encoder0_position[23] (encoder0_position[23]), 
            .\encoder0_position[22] (encoder0_position[22]), .\encoder0_position[21] (encoder0_position[21]), 
            .\encoder0_position[20] (encoder0_position[20]), .\encoder0_position[19] (encoder0_position[19]), 
            .\encoder0_position[18] (encoder0_position[18]), .\encoder0_position[17] (encoder0_position[17]), 
            .\encoder0_position[16] (encoder0_position[16]), .\encoder0_position[15] (encoder0_position[15]), 
            .\encoder0_position[14] (encoder0_position[14]), .\encoder0_position[13] (encoder0_position[13]), 
            .\encoder0_position[12] (encoder0_position[12]), .\encoder0_position[11] (encoder0_position[11]), 
            .\encoder0_position[10] (encoder0_position[10]), .\encoder0_position[9] (encoder0_position[9]), 
            .\encoder0_position[8] (encoder0_position[8]), .\encoder0_position[7] (encoder0_position[7]), 
            .\encoder0_position[6] (encoder0_position[6]), .\encoder0_position[5] (encoder0_position[5]), 
            .\encoder0_position[4] (encoder0_position[4]), .\encoder0_position[3] (encoder0_position[3]), 
            .\encoder0_position[2] (encoder0_position[2]), .\encoder0_position[1] (encoder0_position[1]), 
            .\encoder0_position[0] (encoder0_position[0]), .VCC_net(VCC_net), 
            .n29648(n29648), .a_prev(a_prev), .n29647(n29647), .n29628(n29628), 
            .n1742(n1742), .position_31__N_3836(position_31__N_3836), .\b_new[1] (b_new[1]), 
            .debounce_cnt_N_3833(debounce_cnt_N_3833)) /* synthesis lattice_noprune=1 */ ;   // verilog/TinyFPGA_B.v(304[27] 310[6])
    SB_LUT4 i15643_3_lut (.I0(a_prev_adj_5770), .I1(a_new_adj_5996[1]), 
            .I2(debounce_cnt_N_3833_adj_5772), .I3(GND_net), .O(n29649));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    defparam i15643_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i2_3_lut_4_lut_adj_2191 (.I0(\data_out_frame[23] [3]), .I1(\data_out_frame[23] [2]), 
            .I2(n53457), .I3(n53546), .O(n54456));
    defparam i2_3_lut_4_lut_adj_2191.LUT_INIT = 16'h6996;
    SB_LUT4 i3_3_lut_4_lut (.I0(\data_out_frame[23] [1]), .I1(\data_out_frame[23] [0]), 
            .I2(\data_out_frame[25] [2]), .I3(n58957), .O(n8_adj_5946));
    defparam i3_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i54470_1_lut (.I0(n43737), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n70164));
    defparam i54470_1_lut.LUT_INIT = 16'h5555;
    TLI4970 tli (.\state[1] (state_adj_6017[1]), .GND_net(GND_net), .clk16MHz(clk16MHz), 
            .VCC_net(VCC_net), .n6(n6), .n5(n5_adj_5733), .n11(n11_adj_5764), 
            .n15(n15_adj_5763), .\state[0] (state_adj_6017[0]), .\data[12] (data_adj_6015[12]), 
            .n29622(n29622), .\data[15] (data_adj_6015[15]), .clk_out(clk_out), 
            .CS_c(CS_c), .CS_CLK_c(CS_CLK_c), .n29602(n29602), .n9(n9_adj_5953), 
            .n29567(n29567), .n29565(n29565), .\current[0] (current[0]), 
            .n29563(n29563), .\data[11] (data_adj_6015[11]), .n29562(n29562), 
            .\data[10] (data_adj_6015[10]), .n29550(n29550), .\data[9] (data_adj_6015[9]), 
            .n29549(n29549), .\data[8] (data_adj_6015[8]), .n29548(n29548), 
            .\data[7] (data_adj_6015[7]), .n29547(n29547), .\data[6] (data_adj_6015[6]), 
            .n29546(n29546), .\data[5] (data_adj_6015[5]), .n29545(n29545), 
            .\data[4] (data_adj_6015[4]), .n29538(n29538), .\data[3] (data_adj_6015[3]), 
            .n29530(n29530), .\data[2] (data_adj_6015[2]), .n29529(n29529), 
            .\data[1] (data_adj_6015[1]), .n25499(n25499), .n4(n4_adj_5934), 
            .n25508(n25508), .n30424(n30424), .\data[0] (data_adj_6015[0]), 
            .n30319(n30319), .\current[1] (current[1]), .n30318(n30318), 
            .\current[2] (current[2]), .n30317(n30317), .\current[3] (current[3]), 
            .n30316(n30316), .\current[4] (current[4]), .n30315(n30315), 
            .\current[5] (current[5]), .n30313(n30313), .\current[6] (current[6]), 
            .n30312(n30312), .\current[7] (current[7]), .n30311(n30311), 
            .\current[8] (current[8]), .n30310(n30310), .\current[9] (current[9]), 
            .n30309(n30309), .\current[10] (current[10]), .n30308(n30308), 
            .\current[11] (current[11]), .n25504(n25504), .n25512(n25512), 
            .n27643(n27643), .\current[15] (current[15]), .n6_adj_7(n6_adj_5762), 
            .n5_adj_8(n5_adj_5734), .n5_adj_9(n5_adj_5824), .n6_adj_10(n6_adj_5759), 
            .state_7__N_4319(state_7__N_4319), .n42981(n42981)) /* synthesis syn_noprune=1, syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(404[11] 410[4])
    SB_LUT4 encoder0_position_30__I_0_i2195_3_lut (.I0(n3224), .I1(n3291), 
            .I2(n3237), .I3(GND_net), .O(n23_adj_5930));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2195_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2191_3_lut (.I0(n3220), .I1(n3287), 
            .I2(n3237), .I3(GND_net), .O(n31_adj_5931));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2191_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2200_3_lut (.I0(n3229), .I1(n3296), 
            .I2(n3237), .I3(GND_net), .O(n13_adj_5926));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2200_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2199_3_lut (.I0(n3228), .I1(n3295), 
            .I2(n3237), .I3(GND_net), .O(n15_adj_5927));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2199_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_2192 (.I0(n3221), .I1(n13_adj_5926), .I2(n3288), 
            .I3(n3237), .O(n62929));
    defparam i1_4_lut_adj_2192.LUT_INIT = 16'heefc;
    SB_LUT4 i16504_2_lut_2_lut_4_lut (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[15] [0]), 
            .O(n30510));   // verilog/coms.v(130[12] 305[6])
    defparam i16504_2_lut_2_lut_4_lut.LUT_INIT = 16'h5555;
    EEPROM eeprom (.n25391(n25391), .\state[0] (state_adj_6008[0]), .\state[1] (state_adj_6008[1]), 
           .enable_slow_N_4213(enable_slow_N_4213), .n5771({n5772}), .ready_prev(ready_prev), 
           .clk16MHz(clk16MHz), .\state[2] (state_adj_6008[2]), .GND_net(GND_net), 
           .n43543(n43543), .\state_7__N_3918[0] (state_7__N_3918[0]), .n42885(n42885), 
           .n29566(n29566), .rw(rw), .n58190(n58190), .data_ready(data_ready), 
           .ID({ID}), .n57800(n57800), .n58002(n58002), .baudrate({baudrate}), 
           .n30330(n30330), .n30329(n30329), .n30328(n30328), .n30327(n30327), 
           .n30326(n30326), .n30325(n30325), .n30324(n30324), .n30323(n30323), 
           .\state[0]_adj_3 (state_adj_6041[0]), .n58751(n58751), .n4(n4_adj_5952), 
           .data({data_adj_6007}), .n61888(n61888), .n25490(n25490), .scl_enable(scl_enable), 
           .\state_7__N_4110[0] (state_7__N_4110[0]), .VCC_net(VCC_net), 
           .scl(scl), .sda_enable(sda_enable), .sda_out(sda_out), .n29573(n29573), 
           .\saved_addr[0] (saved_addr[0]), .n6426(n6426), .n30410(n30410), 
           .n8(n8_adj_5954), .n30134(n30134), .n30133(n30133), .n30132(n30132), 
           .n30131(n30131), .n30130(n30130), .n30129(n30129), .n30128(n30128), 
           .n4_adj_4(n4_adj_5756), .n4_adj_5(n4_adj_5757), .n42994(n42994), 
           .n6(n6_adj_5721), .\state_7__N_4126[3] (state_7__N_4126[3]), 
           .n10(n10_adj_5758), .n25522(n25522), .n25517(n25517), .n10_adj_6(n10_adj_5761)) /* synthesis syn_noprune=1, syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(390[10] 402[6])
    SB_LUT4 encoder0_position_30__I_0_i2190_3_lut (.I0(n3219), .I1(n3286), 
            .I2(n3237), .I3(GND_net), .O(n33_adj_5932));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2190_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2197_3_lut (.I0(n3226), .I1(n3293), 
            .I2(n3237), .I3(GND_net), .O(n19_adj_5929));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2197_3_lut.LUT_INIT = 16'hacac;
    
endmodule
//
// Verilog Description of module \neopixel(CLOCK_SPEED_HZ=16000000) 
//

module \neopixel(CLOCK_SPEED_HZ=16000000)  (VCC_net, timer, clk16MHz, 
            GND_net, state, \neo_pixel_transmitter.t0 , n22979, neopxl_color, 
            bit_ctr, n29595, n27855, \bit_ctr[3] , \bit_ctr[4] , \bit_ctr[1] , 
            n43547, n30238, n30237, n30236, n30235, n30234, n30233, 
            n30232, n30231, n30230, n30224, n30139, n57450, NEOPXL_c, 
            n66810, LED_c, \color_bit_N_502[1] , n53519, n3157) /* synthesis syn_module_defined=1 */ ;
    input VCC_net;
    output [10:0]timer;
    input clk16MHz;
    input GND_net;
    output [1:0]state;
    output [10:0]\neo_pixel_transmitter.t0 ;
    output n22979;
    input [23:0]neopxl_color;
    output [4:0]bit_ctr;
    input n29595;
    output n27855;
    output \bit_ctr[3] ;
    output \bit_ctr[4] ;
    output \bit_ctr[1] ;
    output n43547;
    input n30238;
    input n30237;
    input n30236;
    input n30235;
    input n30234;
    input n30233;
    input n30232;
    input n30231;
    input n30230;
    input n30224;
    input n30139;
    input n57450;
    output NEOPXL_c;
    output n66810;
    input LED_c;
    output \color_bit_N_502[1] ;
    output n53519;
    output n3157;
    
    wire clk16MHz /* synthesis SET_AS_NETWORK=clk16MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    wire [10:0]n13;
    
    wire n51016, \neo_pixel_transmitter.done_N_516 , n58692, \neo_pixel_transmitter.done , 
        start_N_507, n7, start, n51017;
    wire [10:0]one_wire_N_479;
    
    wire n12_adj_5684, n25383, n4, n52740, n59646, n4_adj_5685, 
        n64076, n12_adj_5686, n64216, n39, n61873, n43554, n43633, 
        n64544, n64545, n64536, n64535;
    wire [10:0]n49;
    wire [31:0]n137;
    wire [4:0]bit_ctr_c;   // verilog/neopixel.v(17[11:18])
    
    wire n29097, n70862, n70874, n25471, n43033, n25472, n53544, 
        n66808, n21, n18, n59766, n4_adj_5687, n43537, n61910, 
        n71210, n8, n1, n27845, n28810;
    wire [1:0]state_1__N_440;
    
    wire n27859, n59730, \neo_pixel_transmitter.done_N_524 , n69178, 
        n51025, n51024, n51023, n51022, n51021, n51020, n51019, 
        n51018, n52239, n52238, n52237, n52236, n52235, n52234, 
        n52233, n52232, n52231, n52230;
    wire [5:0]color_bit_N_502;
    
    wire n57_adj_5691, n43665, n6893, n71213, n67135, n59626, n67137, 
        n59754, n69177, n70982, n70985, n2838, n64461, n64460, 
        n4_adj_5692, n64462, n64464, n70877, n70865, n64463, n64465;
    
    SB_CARRY sub_67_add_2_2 (.CI(VCC_net), .I0(timer[0]), .I1(n13[0]), 
            .CO(n51016));
    SB_DFFE \neo_pixel_transmitter.done_96  (.Q(\neo_pixel_transmitter.done ), 
            .C(clk16MHz), .E(n58692), .D(\neo_pixel_transmitter.done_N_516 ));   // verilog/neopixel.v(34[12] 116[6])
    SB_DFFE start_95 (.Q(start), .C(clk16MHz), .E(n7), .D(start_N_507));   // verilog/neopixel.v(34[12] 116[6])
    SB_CARRY sub_67_add_2_3 (.CI(n51016), .I0(timer[1]), .I1(n13[1]), 
            .CO(n51017));
    SB_LUT4 i5_4_lut (.I0(one_wire_N_479[7]), .I1(one_wire_N_479[9]), .I2(one_wire_N_479[4]), 
            .I3(one_wire_N_479[6]), .O(n12_adj_5684));   // verilog/neopixel.v(61[15:42])
    defparam i5_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i6_4_lut (.I0(one_wire_N_479[8]), .I1(n12_adj_5684), .I2(one_wire_N_479[5]), 
            .I3(one_wire_N_479[10]), .O(n25383));   // verilog/neopixel.v(61[15:42])
    defparam i6_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_2_lut (.I0(one_wire_N_479[2]), .I1(n4), .I2(GND_net), .I3(GND_net), 
            .O(n52740));
    defparam i2_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i44008_2_lut (.I0(start), .I1(state[1]), .I2(GND_net), .I3(GND_net), 
            .O(n59646));
    defparam i44008_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut (.I0(one_wire_N_479[2]), .I1(one_wire_N_479[3]), .I2(GND_net), 
            .I3(GND_net), .O(n4_adj_5685));
    defparam i1_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i48391_2_lut (.I0(one_wire_N_479[4]), .I1(n4_adj_5685), .I2(GND_net), 
            .I3(GND_net), .O(n64076));
    defparam i48391_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i3_3_lut (.I0(\neo_pixel_transmitter.done ), .I1(one_wire_N_479[10]), 
            .I2(state[0]), .I3(GND_net), .O(n12_adj_5686));
    defparam i3_3_lut.LUT_INIT = 16'h2121;
    SB_LUT4 i48531_4_lut (.I0(one_wire_N_479[8]), .I1(one_wire_N_479[9]), 
            .I2(one_wire_N_479[6]), .I3(n64076), .O(n64216));
    defparam i48531_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i65_2_lut (.I0(\neo_pixel_transmitter.done ), .I1(state[0]), 
            .I2(GND_net), .I3(GND_net), .O(n39));
    defparam i65_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i8_4_lut (.I0(one_wire_N_479[7]), .I1(n64216), .I2(n12_adj_5686), 
            .I3(one_wire_N_479[5]), .O(n61873));
    defparam i8_4_lut.LUT_INIT = 16'h0010;
    SB_LUT4 i55136_4_lut (.I0(n43554), .I1(n59646), .I2(n61873), .I3(n39), 
            .O(n58692));
    defparam i55136_4_lut.LUT_INIT = 16'hcecf;
    SB_LUT4 sub_67_inv_0_i1_1_lut (.I0(\neo_pixel_transmitter.t0 [0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n13[0]));   // verilog/neopixel.v(101[14:24])
    defparam sub_67_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_2_lut_3_lut (.I0(start), .I1(\neo_pixel_transmitter.done ), 
            .I2(n43633), .I3(GND_net), .O(n22979));   // verilog/neopixel.v(78[18] 98[12])
    defparam i1_2_lut_3_lut.LUT_INIT = 16'hbfbf;
    SB_LUT4 i48850_3_lut (.I0(neopxl_color[16]), .I1(neopxl_color[17]), 
            .I2(bit_ctr[0]), .I3(GND_net), .O(n64544));
    defparam i48850_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48851_3_lut (.I0(neopxl_color[18]), .I1(neopxl_color[19]), 
            .I2(bit_ctr[0]), .I3(GND_net), .O(n64545));
    defparam i48851_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48842_3_lut (.I0(neopxl_color[22]), .I1(neopxl_color[23]), 
            .I2(bit_ctr[0]), .I3(GND_net), .O(n64536));
    defparam i48842_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48841_3_lut (.I0(neopxl_color[20]), .I1(neopxl_color[21]), 
            .I2(bit_ctr[0]), .I3(GND_net), .O(n64535));
    defparam i48841_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF timer_1934__i0 (.Q(timer[0]), .C(clk16MHz), .D(n49[0]));   // verilog/neopixel.v(12[12:21])
    SB_DFF \neo_pixel_transmitter.t0_i0_i0  (.Q(\neo_pixel_transmitter.t0 [0]), 
           .C(clk16MHz), .D(n29595));   // verilog/neopixel.v(34[12] 116[6])
    SB_LUT4 sub_67_inv_0_i2_1_lut (.I0(\neo_pixel_transmitter.t0 [1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n13[1]));   // verilog/neopixel.v(101[14:24])
    defparam sub_67_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_DFFESR bit_ctr_i2 (.Q(bit_ctr_c[2]), .C(clk16MHz), .E(n27855), 
            .D(n137[2]), .R(n29097));   // verilog/neopixel.v(34[12] 116[6])
    SB_DFFESR bit_ctr_i3 (.Q(\bit_ctr[3] ), .C(clk16MHz), .E(n27855), 
            .D(n137[3]), .R(n29097));   // verilog/neopixel.v(34[12] 116[6])
    SB_DFFESR bit_ctr_i4 (.Q(\bit_ctr[4] ), .C(clk16MHz), .E(n27855), 
            .D(n137[4]), .R(n29097));   // verilog/neopixel.v(34[12] 116[6])
    SB_DFF timer_1934__i10 (.Q(timer[10]), .C(clk16MHz), .D(n49[10]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1934__i9 (.Q(timer[9]), .C(clk16MHz), .D(n49[9]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1934__i8 (.Q(timer[8]), .C(clk16MHz), .D(n49[8]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1934__i7 (.Q(timer[7]), .C(clk16MHz), .D(n49[7]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1934__i6 (.Q(timer[6]), .C(clk16MHz), .D(n49[6]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1934__i5 (.Q(timer[5]), .C(clk16MHz), .D(n49[5]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1934__i4 (.Q(timer[4]), .C(clk16MHz), .D(n49[4]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1934__i3 (.Q(timer[3]), .C(clk16MHz), .D(n49[3]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1934__i2 (.Q(timer[2]), .C(clk16MHz), .D(n49[2]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1934__i1 (.Q(timer[1]), .C(clk16MHz), .D(n49[1]));   // verilog/neopixel.v(12[12:21])
    SB_LUT4 bit_ctr_0__bdd_4_lut_55178_4_lut (.I0(bit_ctr[0]), .I1(neopxl_color[6]), 
            .I2(neopxl_color[7]), .I3(\bit_ctr[1] ), .O(n70862));
    defparam bit_ctr_0__bdd_4_lut_55178_4_lut.LUT_INIT = 16'heea0;
    SB_LUT4 bit_ctr_0__bdd_4_lut_55452_4_lut (.I0(bit_ctr[0]), .I1(neopxl_color[2]), 
            .I2(neopxl_color[3]), .I3(\bit_ctr[1] ), .O(n70874));
    defparam bit_ctr_0__bdd_4_lut_55452_4_lut.LUT_INIT = 16'heea0;
    SB_LUT4 i1_2_lut_3_lut_adj_1733 (.I0(n43554), .I1(start), .I2(\neo_pixel_transmitter.done ), 
            .I3(GND_net), .O(n25471));   // verilog/neopixel.v(78[18] 98[12])
    defparam i1_2_lut_3_lut_adj_1733.LUT_INIT = 16'hdfdf;
    SB_LUT4 i1_2_lut_3_lut_adj_1734 (.I0(n43033), .I1(start), .I2(\neo_pixel_transmitter.done ), 
            .I3(GND_net), .O(n25472));   // verilog/neopixel.v(51[18] 71[12])
    defparam i1_2_lut_3_lut_adj_1734.LUT_INIT = 16'hdfdf;
    SB_LUT4 i51114_2_lut_3_lut (.I0(n53544), .I1(\bit_ctr[3] ), .I2(n43547), 
            .I3(GND_net), .O(n66808));   // verilog/neopixel.v(21[26:38])
    defparam i51114_2_lut_3_lut.LUT_INIT = 16'h2828;
    SB_LUT4 i1_4_lut_4_lut (.I0(start), .I1(\neo_pixel_transmitter.done ), 
            .I2(n43033), .I3(n43554), .O(n21));
    defparam i1_4_lut_4_lut.LUT_INIT = 16'h5410;
    SB_LUT4 i1_4_lut_4_lut_adj_1735 (.I0(start), .I1(\neo_pixel_transmitter.done ), 
            .I2(n43554), .I3(n43033), .O(n18));
    defparam i1_4_lut_4_lut_adj_1735.LUT_INIT = 16'h5410;
    SB_LUT4 i2_2_lut_3_lut (.I0(n25383), .I1(one_wire_N_479[2]), .I2(one_wire_N_479[3]), 
            .I3(GND_net), .O(n43033));
    defparam i2_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i50_3_lut_4_lut (.I0(one_wire_N_479[2]), .I1(n4), .I2(one_wire_N_479[3]), 
            .I3(\neo_pixel_transmitter.done ), .O(n59766));
    defparam i50_3_lut_4_lut.LUT_INIT = 16'hfa88;
    SB_LUT4 i1_2_lut_3_lut_adj_1736 (.I0(n25383), .I1(start), .I2(state[1]), 
            .I3(GND_net), .O(n4_adj_5687));
    defparam i1_2_lut_3_lut_adj_1736.LUT_INIT = 16'hfefe;
    SB_DFF \neo_pixel_transmitter.t0_i0_i1  (.Q(\neo_pixel_transmitter.t0 [1]), 
           .C(clk16MHz), .D(n30238));   // verilog/neopixel.v(34[12] 116[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i2  (.Q(\neo_pixel_transmitter.t0 [2]), 
           .C(clk16MHz), .D(n30237));   // verilog/neopixel.v(34[12] 116[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i3  (.Q(\neo_pixel_transmitter.t0 [3]), 
           .C(clk16MHz), .D(n30236));   // verilog/neopixel.v(34[12] 116[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i4  (.Q(\neo_pixel_transmitter.t0 [4]), 
           .C(clk16MHz), .D(n30235));   // verilog/neopixel.v(34[12] 116[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i5  (.Q(\neo_pixel_transmitter.t0 [5]), 
           .C(clk16MHz), .D(n30234));   // verilog/neopixel.v(34[12] 116[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i6  (.Q(\neo_pixel_transmitter.t0 [6]), 
           .C(clk16MHz), .D(n30233));   // verilog/neopixel.v(34[12] 116[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i7  (.Q(\neo_pixel_transmitter.t0 [7]), 
           .C(clk16MHz), .D(n30232));   // verilog/neopixel.v(34[12] 116[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i8  (.Q(\neo_pixel_transmitter.t0 [8]), 
           .C(clk16MHz), .D(n30231));   // verilog/neopixel.v(34[12] 116[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i9  (.Q(\neo_pixel_transmitter.t0 [9]), 
           .C(clk16MHz), .D(n30230));   // verilog/neopixel.v(34[12] 116[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i10  (.Q(\neo_pixel_transmitter.t0 [10]), 
           .C(clk16MHz), .D(n30224));   // verilog/neopixel.v(34[12] 116[6])
    SB_DFF bit_ctr_i1 (.Q(\bit_ctr[1] ), .C(clk16MHz), .D(n30139));   // verilog/neopixel.v(34[12] 116[6])
    SB_DFFE state_i1 (.Q(state[1]), .C(clk16MHz), .E(VCC_net), .D(n57450));   // verilog/neopixel.v(34[12] 116[6])
    SB_LUT4 i3_4_lut_4_lut (.I0(n43537), .I1(state[1]), .I2(state[0]), 
            .I3(\neo_pixel_transmitter.done ), .O(n61910));
    defparam i3_4_lut_4_lut.LUT_INIT = 16'h0004;
    SB_LUT4 bit_ctr_0__bdd_4_lut_4_lut (.I0(bit_ctr[0]), .I1(neopxl_color[10]), 
            .I2(neopxl_color[11]), .I3(\bit_ctr[1] ), .O(n71210));
    defparam bit_ctr_0__bdd_4_lut_4_lut.LUT_INIT = 16'heea0;
    SB_LUT4 i2090_2_lut_3_lut (.I0(bit_ctr_c[2]), .I1(\bit_ctr[1] ), .I2(bit_ctr[0]), 
            .I3(GND_net), .O(n137[2]));   // verilog/neopixel.v(68[23:32])
    defparam i2090_2_lut_3_lut.LUT_INIT = 16'h6a6a;
    SB_LUT4 i3_3_lut_4_lut (.I0(\bit_ctr[3] ), .I1(n43547), .I2(n53544), 
            .I3(bit_ctr[0]), .O(n8));
    defparam i3_3_lut_4_lut.LUT_INIT = 16'hff9f;
    SB_DFFESR bit_ctr_i0 (.Q(bit_ctr[0]), .C(clk16MHz), .E(n27845), .D(n1), 
            .R(n28810));   // verilog/neopixel.v(34[12] 116[6])
    SB_DFFESS state_i0 (.Q(state[0]), .C(clk16MHz), .E(n27859), .D(state_1__N_440[0]), 
            .S(n59730));   // verilog/neopixel.v(34[12] 116[6])
    SB_DFFESR one_wire_99 (.Q(NEOPXL_c), .C(clk16MHz), .E(n69178), .D(\neo_pixel_transmitter.done_N_524 ), 
            .R(n61910));   // verilog/neopixel.v(34[12] 116[6])
    SB_LUT4 sub_67_add_2_12_lut (.I0(GND_net), .I1(timer[10]), .I2(n13[10]), 
            .I3(n51025), .O(one_wire_N_479[10])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_67_add_2_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_67_add_2_11_lut (.I0(GND_net), .I1(timer[9]), .I2(n13[9]), 
            .I3(n51024), .O(one_wire_N_479[9])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_67_add_2_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_67_add_2_11 (.CI(n51024), .I0(timer[9]), .I1(n13[9]), 
            .CO(n51025));
    SB_LUT4 sub_67_add_2_10_lut (.I0(GND_net), .I1(timer[8]), .I2(n13[8]), 
            .I3(n51023), .O(one_wire_N_479[8])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_67_add_2_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_67_add_2_10 (.CI(n51023), .I0(timer[8]), .I1(n13[8]), 
            .CO(n51024));
    SB_LUT4 sub_67_add_2_9_lut (.I0(GND_net), .I1(timer[7]), .I2(n13[7]), 
            .I3(n51022), .O(one_wire_N_479[7])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_67_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_67_add_2_9 (.CI(n51022), .I0(timer[7]), .I1(n13[7]), 
            .CO(n51023));
    SB_LUT4 sub_67_add_2_8_lut (.I0(GND_net), .I1(timer[6]), .I2(n13[6]), 
            .I3(n51021), .O(one_wire_N_479[6])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_67_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_67_add_2_8 (.CI(n51021), .I0(timer[6]), .I1(n13[6]), 
            .CO(n51022));
    SB_LUT4 sub_67_add_2_7_lut (.I0(GND_net), .I1(timer[5]), .I2(n13[5]), 
            .I3(n51020), .O(one_wire_N_479[5])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_67_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_67_add_2_7 (.CI(n51020), .I0(timer[5]), .I1(n13[5]), 
            .CO(n51021));
    SB_LUT4 sub_67_add_2_6_lut (.I0(GND_net), .I1(timer[4]), .I2(n13[4]), 
            .I3(n51019), .O(one_wire_N_479[4])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_67_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_67_add_2_6 (.CI(n51019), .I0(timer[4]), .I1(n13[4]), 
            .CO(n51020));
    SB_LUT4 sub_67_add_2_5_lut (.I0(GND_net), .I1(timer[3]), .I2(n13[3]), 
            .I3(n51018), .O(one_wire_N_479[3])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_67_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_67_add_2_5 (.CI(n51018), .I0(timer[3]), .I1(n13[3]), 
            .CO(n51019));
    SB_LUT4 sub_67_add_2_4_lut (.I0(GND_net), .I1(timer[2]), .I2(n13[2]), 
            .I3(n51017), .O(one_wire_N_479[2])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_67_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_67_add_2_4 (.CI(n51017), .I0(timer[2]), .I1(n13[2]), 
            .CO(n51018));
    SB_LUT4 sub_67_add_2_3_lut (.I0(one_wire_N_479[3]), .I1(timer[1]), .I2(n13[1]), 
            .I3(n51016), .O(n4)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_67_add_2_3_lut.LUT_INIT = 16'h8228;
    SB_LUT4 timer_1934_add_4_12_lut (.I0(GND_net), .I1(GND_net), .I2(timer[10]), 
            .I3(n52239), .O(n49[10])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1934_add_4_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 timer_1934_add_4_11_lut (.I0(GND_net), .I1(GND_net), .I2(timer[9]), 
            .I3(n52238), .O(n49[9])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1934_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1934_add_4_11 (.CI(n52238), .I0(GND_net), .I1(timer[9]), 
            .CO(n52239));
    SB_LUT4 timer_1934_add_4_10_lut (.I0(GND_net), .I1(GND_net), .I2(timer[8]), 
            .I3(n52237), .O(n49[8])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1934_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1934_add_4_10 (.CI(n52237), .I0(GND_net), .I1(timer[8]), 
            .CO(n52238));
    SB_LUT4 timer_1934_add_4_9_lut (.I0(GND_net), .I1(GND_net), .I2(timer[7]), 
            .I3(n52236), .O(n49[7])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1934_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1934_add_4_9 (.CI(n52236), .I0(GND_net), .I1(timer[7]), 
            .CO(n52237));
    SB_LUT4 timer_1934_add_4_8_lut (.I0(GND_net), .I1(GND_net), .I2(timer[6]), 
            .I3(n52235), .O(n49[6])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1934_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1934_add_4_8 (.CI(n52235), .I0(GND_net), .I1(timer[6]), 
            .CO(n52236));
    SB_LUT4 timer_1934_add_4_7_lut (.I0(GND_net), .I1(GND_net), .I2(timer[5]), 
            .I3(n52234), .O(n49[5])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1934_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1934_add_4_7 (.CI(n52234), .I0(GND_net), .I1(timer[5]), 
            .CO(n52235));
    SB_LUT4 timer_1934_add_4_6_lut (.I0(GND_net), .I1(GND_net), .I2(timer[4]), 
            .I3(n52233), .O(n49[4])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1934_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1934_add_4_6 (.CI(n52233), .I0(GND_net), .I1(timer[4]), 
            .CO(n52234));
    SB_LUT4 timer_1934_add_4_5_lut (.I0(GND_net), .I1(GND_net), .I2(timer[3]), 
            .I3(n52232), .O(n49[3])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1934_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1934_add_4_5 (.CI(n52232), .I0(GND_net), .I1(timer[3]), 
            .CO(n52233));
    SB_LUT4 timer_1934_add_4_4_lut (.I0(GND_net), .I1(GND_net), .I2(timer[2]), 
            .I3(n52231), .O(n49[2])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1934_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1934_add_4_4 (.CI(n52231), .I0(GND_net), .I1(timer[2]), 
            .CO(n52232));
    SB_LUT4 timer_1934_add_4_3_lut (.I0(GND_net), .I1(GND_net), .I2(timer[1]), 
            .I3(n52230), .O(n49[1])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1934_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1934_add_4_3 (.CI(n52230), .I0(GND_net), .I1(timer[1]), 
            .CO(n52231));
    SB_LUT4 timer_1934_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(timer[0]), 
            .I3(VCC_net), .O(n49[0])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1934_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_67_inv_0_i3_1_lut (.I0(\neo_pixel_transmitter.t0 [2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n13[2]));   // verilog/neopixel.v(101[14:24])
    defparam sub_67_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i51116_2_lut (.I0(n53544), .I1(color_bit_N_502[2]), .I2(GND_net), 
            .I3(GND_net), .O(n66810));
    defparam i51116_2_lut.LUT_INIT = 16'h2222;
    SB_CARRY timer_1934_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(timer[0]), 
            .CO(n52230));
    SB_LUT4 sub_67_inv_0_i4_1_lut (.I0(\neo_pixel_transmitter.t0 [3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n13[3]));   // verilog/neopixel.v(101[14:24])
    defparam sub_67_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_67_inv_0_i5_1_lut (.I0(\neo_pixel_transmitter.t0 [4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n13[4]));   // verilog/neopixel.v(101[14:24])
    defparam sub_67_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_67_inv_0_i6_1_lut (.I0(\neo_pixel_transmitter.t0 [5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n13[5]));   // verilog/neopixel.v(101[14:24])
    defparam sub_67_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_67_inv_0_i7_1_lut (.I0(\neo_pixel_transmitter.t0 [6]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n13[6]));   // verilog/neopixel.v(101[14:24])
    defparam sub_67_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_67_inv_0_i8_1_lut (.I0(\neo_pixel_transmitter.t0 [7]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n13[7]));   // verilog/neopixel.v(101[14:24])
    defparam sub_67_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_67_inv_0_i9_1_lut (.I0(\neo_pixel_transmitter.t0 [8]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n13[8]));   // verilog/neopixel.v(101[14:24])
    defparam sub_67_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_67_inv_0_i10_1_lut (.I0(\neo_pixel_transmitter.t0 [9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n13[9]));   // verilog/neopixel.v(101[14:24])
    defparam sub_67_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_67_inv_0_i11_1_lut (.I0(\neo_pixel_transmitter.t0 [10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n13[10]));   // verilog/neopixel.v(101[14:24])
    defparam sub_67_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i2097_2_lut_3_lut_4_lut (.I0(bit_ctr_c[2]), .I1(\bit_ctr[1] ), 
            .I2(bit_ctr[0]), .I3(\bit_ctr[3] ), .O(n137[3]));   // verilog/neopixel.v(68[23:32])
    defparam i2097_2_lut_3_lut_4_lut.LUT_INIT = 16'h7f80;
    SB_LUT4 i1_2_lut_4_lut (.I0(state[0]), .I1(n57_adj_5691), .I2(LED_c), 
            .I3(state[1]), .O(n27845));   // verilog/neopixel.v(35[4] 115[11])
    defparam i1_2_lut_4_lut.LUT_INIT = 16'h20ff;
    SB_LUT4 i14804_2_lut_4_lut (.I0(state[0]), .I1(n57_adj_5691), .I2(LED_c), 
            .I3(state[1]), .O(n28810));   // verilog/neopixel.v(35[4] 115[11])
    defparam i14804_2_lut_4_lut.LUT_INIT = 16'h2000;
    SB_LUT4 i1_2_lut_3_lut_adj_1737 (.I0(\bit_ctr[3] ), .I1(n43547), .I2(\bit_ctr[4] ), 
            .I3(GND_net), .O(n53544));
    defparam i1_2_lut_3_lut_adj_1737.LUT_INIT = 16'h7878;
    SB_LUT4 i29765_2_lut_3_lut (.I0(\bit_ctr[3] ), .I1(n43547), .I2(\bit_ctr[4] ), 
            .I3(GND_net), .O(n43665));
    defparam i29765_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i1_2_lut_3_lut_adj_1738 (.I0(\bit_ctr[1] ), .I1(bit_ctr[0]), 
            .I2(bit_ctr_c[2]), .I3(GND_net), .O(color_bit_N_502[2]));
    defparam i1_2_lut_3_lut_adj_1738.LUT_INIT = 16'h1e1e;
    SB_LUT4 i29652_2_lut_3_lut (.I0(\bit_ctr[1] ), .I1(bit_ctr[0]), .I2(bit_ctr_c[2]), 
            .I3(GND_net), .O(n43547));
    defparam i29652_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i2104_3_lut_4_lut (.I0(bit_ctr_c[2]), .I1(n6893), .I2(\bit_ctr[3] ), 
            .I3(\bit_ctr[4] ), .O(n137[4]));   // verilog/neopixel.v(68[23:32])
    defparam i2104_3_lut_4_lut.LUT_INIT = 16'h7f80;
    SB_LUT4 i1_2_lut_adj_1739 (.I0(\bit_ctr[1] ), .I1(bit_ctr[0]), .I2(GND_net), 
            .I3(GND_net), .O(\color_bit_N_502[1] ));
    defparam i1_2_lut_adj_1739.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1740 (.I0(\bit_ctr[3] ), .I1(n43547), .I2(GND_net), 
            .I3(GND_net), .O(n53519));
    defparam i1_2_lut_adj_1740.LUT_INIT = 16'h6666;
    SB_LUT4 i1077_4_lut (.I0(\color_bit_N_502[1] ), .I1(n43665), .I2(n8), 
            .I3(color_bit_N_502[2]), .O(n57_adj_5691));   // verilog/neopixel.v(21[26:38])
    defparam i1077_4_lut.LUT_INIT = 16'h3332;
    SB_LUT4 i2085_2_lut (.I0(\bit_ctr[1] ), .I1(bit_ctr[0]), .I2(GND_net), 
            .I3(GND_net), .O(n6893));   // verilog/neopixel.v(68[23:32])
    defparam i2085_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i15091_2_lut (.I0(n27855), .I1(state[1]), .I2(GND_net), .I3(GND_net), 
            .O(n29097));   // verilog/neopixel.v(34[12] 116[6])
    defparam i15091_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_3_lut (.I0(n27845), .I1(n22979), .I2(state[1]), .I3(GND_net), 
            .O(n27855));
    defparam i1_3_lut.LUT_INIT = 16'ha2a2;
    SB_LUT4 i29643_3_lut (.I0(one_wire_N_479[8]), .I1(one_wire_N_479[10]), 
            .I2(one_wire_N_479[9]), .I3(GND_net), .O(n43537));
    defparam i29643_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i43917_4_lut (.I0(n25383), .I1(n52740), .I2(n4_adj_5685), 
            .I3(state[0]), .O(n43633));   // verilog/neopixel.v(35[4] 115[11])
    defparam i43917_4_lut.LUT_INIT = 16'hfaee;
    SB_LUT4 n71210_bdd_4_lut (.I0(n71210), .I1(neopxl_color[9]), .I2(neopxl_color[8]), 
            .I3(\color_bit_N_502[1] ), .O(n71213));
    defparam n71210_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i51656_2_lut (.I0(\neo_pixel_transmitter.done ), .I1(state[0]), 
            .I2(GND_net), .I3(GND_net), .O(n67135));
    defparam i51656_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i43988_3_lut (.I0(\neo_pixel_transmitter.done ), .I1(start), 
            .I2(n43633), .I3(GND_net), .O(n59626));
    defparam i43988_3_lut.LUT_INIT = 16'hecec;
    SB_LUT4 i15_4_lut (.I0(n59626), .I1(n67135), .I2(state[1]), .I3(n43537), 
            .O(n7));
    defparam i15_4_lut.LUT_INIT = 16'h3a0a;
    SB_LUT4 i54374_2_lut (.I0(start), .I1(state[1]), .I2(GND_net), .I3(GND_net), 
            .O(start_N_507));   // verilog/neopixel.v(35[4] 115[11])
    defparam i54374_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 i51516_2_lut (.I0(n25383), .I1(start), .I2(GND_net), .I3(GND_net), 
            .O(n67137));
    defparam i51516_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i51_4_lut (.I0(n67137), .I1(n43537), .I2(state[1]), .I3(n4_adj_5685), 
            .O(n59754));
    defparam i51_4_lut.LUT_INIT = 16'hcfca;
    SB_LUT4 i53483_4_lut (.I0(n59754), .I1(n59646), .I2(\neo_pixel_transmitter.done ), 
            .I3(n43554), .O(n69177));
    defparam i53483_4_lut.LUT_INIT = 16'hfaca;
    SB_LUT4 i53484_4_lut (.I0(n69177), .I1(n59766), .I2(state[0]), .I3(n4_adj_5687), 
            .O(n69178));
    defparam i53484_4_lut.LUT_INIT = 16'h0535;
    SB_LUT4 color_bit_N_502_1__bdd_4_lut (.I0(\color_bit_N_502[1] ), .I1(n64535), 
            .I2(n64536), .I3(color_bit_N_502[2]), .O(n70982));
    defparam color_bit_N_502_1__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n70982_bdd_4_lut (.I0(n70982), .I1(n64545), .I2(n64544), .I3(color_bit_N_502[2]), 
            .O(n70985));
    defparam n70982_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i2_1_lut (.I0(\neo_pixel_transmitter.done ), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(\neo_pixel_transmitter.done_N_524 ));
    defparam i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 state_1__I_0_i3_3_lut_3_lut (.I0(start), .I1(\neo_pixel_transmitter.done ), 
            .I2(state[1]), .I3(GND_net), .O(\neo_pixel_transmitter.done_N_516 ));   // verilog/neopixel.v(35[4] 115[11])
    defparam state_1__I_0_i3_3_lut_3_lut.LUT_INIT = 16'hc1c1;
    SB_LUT4 i602_2_lut (.I0(n43537), .I1(\neo_pixel_transmitter.done ), 
            .I2(GND_net), .I3(GND_net), .O(n2838));   // verilog/neopixel.v(102[9] 110[12])
    defparam i602_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 i15_4_lut_adj_1741 (.I0(n22979), .I1(n2838), .I2(state[1]), 
            .I3(state[0]), .O(n59730));   // verilog/neopixel.v(34[12] 116[6])
    defparam i15_4_lut_adj_1741.LUT_INIT = 16'h0535;
    SB_LUT4 i20_4_lut (.I0(n22979), .I1(n2838), .I2(state[1]), .I3(state[0]), 
            .O(n27859));
    defparam i20_4_lut.LUT_INIT = 16'hf535;
    SB_LUT4 i48767_3_lut (.I0(neopxl_color[14]), .I1(neopxl_color[15]), 
            .I2(bit_ctr[0]), .I3(GND_net), .O(n64461));
    defparam i48767_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48766_3_lut (.I0(neopxl_color[12]), .I1(neopxl_color[13]), 
            .I2(bit_ctr[0]), .I3(GND_net), .O(n64460));
    defparam i48766_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i54307_4_lut (.I0(state[1]), .I1(state[0]), .I2(n21), .I3(n18), 
            .O(n4_adj_5692));
    defparam i54307_4_lut.LUT_INIT = 16'h5410;
    SB_LUT4 i2_3_lut (.I0(start), .I1(n4_adj_5692), .I2(state[1]), .I3(GND_net), 
            .O(n3157));
    defparam i2_3_lut.LUT_INIT = 16'hcece;
    SB_LUT4 i48768_4_lut (.I0(n64461), .I1(n70985), .I2(n53544), .I3(n53519), 
            .O(n64462));
    defparam i48768_4_lut.LUT_INIT = 16'haca0;
    SB_LUT4 i48770_4_lut (.I0(n64462), .I1(n64460), .I2(n53544), .I3(\color_bit_N_502[1] ), 
            .O(n64464));
    defparam i48770_4_lut.LUT_INIT = 16'haaca;
    SB_LUT4 i48769_3_lut (.I0(n70877), .I1(n70865), .I2(color_bit_N_502[2]), 
            .I3(GND_net), .O(n64463));
    defparam i48769_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48771_3_lut (.I0(n64464), .I1(n71213), .I2(n66810), .I3(GND_net), 
            .O(n64465));
    defparam i48771_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i28922_4_lut (.I0(n64465), .I1(n57_adj_5691), .I2(n64463), 
            .I3(n66808), .O(state_1__N_440[0]));   // verilog/neopixel.v(39[18] 44[12])
    defparam i28922_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i29659_2_lut_3_lut (.I0(one_wire_N_479[2]), .I1(n4), .I2(n25383), 
            .I3(GND_net), .O(n43554));
    defparam i29659_2_lut_3_lut.LUT_INIT = 16'hf8f8;
    SB_LUT4 state_1__I_0_102_Mux_0_i1_4_lut (.I0(n25471), .I1(n25472), .I2(state[0]), 
            .I3(bit_ctr[0]), .O(n1));   // verilog/neopixel.v(35[4] 115[11])
    defparam state_1__I_0_102_Mux_0_i1_4_lut.LUT_INIT = 16'hca35;
    SB_LUT4 n70874_bdd_4_lut (.I0(n70874), .I1(neopxl_color[1]), .I2(neopxl_color[0]), 
            .I3(\color_bit_N_502[1] ), .O(n70877));
    defparam n70874_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n70862_bdd_4_lut (.I0(n70862), .I1(neopxl_color[5]), .I2(neopxl_color[4]), 
            .I3(\color_bit_N_502[1] ), .O(n70865));
    defparam n70862_bdd_4_lut.LUT_INIT = 16'haad8;
    
endmodule
//
// Verilog Description of module motorControl
//

module motorControl (GND_net, control_update, duty, clk16MHz, reset, 
            \Ki[11] , \PID_CONTROLLER.integral_23__N_3715[0] , \Kp[7] , 
            \Kp[1] , \Kp[0] , \Kp[8] , \Kp[9] , n43055, \Kp[10] , 
            \Kp[13] , \Kp[2] , IntegralLimit, \Kp[11] , n155, \PID_CONTROLLER.integral_23__N_3715[15] , 
            \Ki[1] , \PID_CONTROLLER.integral_23__N_3715[14] , \Ki[0] , 
            n367, VCC_net, n375, n376, \Kp[12] , \PID_CONTROLLER.integral , 
            \Ki[2] , \Kp[3] , \Kp[14] , n53, \Kp[4] , \Kp[15] , 
            \Kp[5] , \Kp[6] , \Ki[12] , \Ki[13] , PWMLimit, \Ki[14] , 
            \Ki[15] , \Ki[4] , n4, setpoint, n16, n3, n18, \motor_state[21] , 
            \motor_state[20] , \motor_state[19] , \Ki[5] , \motor_state[18] , 
            n28, \PID_CONTROLLER.integral_23__N_3715[13] , \PID_CONTROLLER.integral_23__N_3715[12] , 
            \Ki[3] , n214, \PID_CONTROLLER.integral_23__N_3715[16] , n29560, 
            \Ki[6] , \Ki[7] , \Ki[8] , \Ki[9] , \Ki[10] , \PID_CONTROLLER.integral_23__N_3715[11] , 
            \motor_state[17] , \PID_CONTROLLER.integral_23__N_3715[10] , 
            n30387, n30386, n30385, n30384, n30383, n30382, n30381, 
            n30380, n30379, n30378, n30377, n30376, n30374, n30372, 
            n30371, n30370, n30369, n30368, n30367, n30366, n30365, 
            n30364, n30363, \PID_CONTROLLER.integral_23__N_3715[9] , \PID_CONTROLLER.integral_23__N_3715[20] , 
            n36816, n20183, \PID_CONTROLLER.integral_23__N_3715[8] , \PID_CONTROLLER.integral_23__N_3715[23] , 
            n20, \motor_state[15] , \motor_state[14] , n490, n417, 
            n20136, n344, \motor_state[13] , n20137, n271, n20138, 
            n198, \PID_CONTROLLER.integral_23__N_3715[7] , \motor_state[12] , 
            n56, n125, \motor_state[11] , n455, n456, \motor_state[10] , 
            \motor_state[9] , \motor_state[8] , \motor_state[7] , n41635, 
            \motor_state[5] , \motor_state[4] , \motor_state[3] , \motor_state[2] , 
            \motor_state[1] , \motor_state[0] , n401, n33, n361, \PID_CONTROLLER.integral_23__N_3715[6] , 
            \PID_CONTROLLER.integral_23__N_3715[5] , deadband, n38, n110, 
            \PID_CONTROLLER.integral_23__N_3715[4] , \PID_CONTROLLER.integral_23__N_3715[3] , 
            \PID_CONTROLLER.integral_23__N_3715[21] , n37330, n11597, 
            n131, n204, n4_adj_30, n20182, n31, \PID_CONTROLLER.integral_23__N_3715[22] , 
            n20_adj_31, n212, n213, \PID_CONTROLLER.integral_23__N_3715[2] , 
            n219, n230, n19, \PID_CONTROLLER.integral_23__N_3715[1] , 
            n4_adj_32, n20181, n6, n36845, n20209, n6_adj_33, n27629) /* synthesis syn_module_defined=1 */ ;
    input GND_net;
    output control_update;
    output [23:0]duty;
    input clk16MHz;
    input reset;
    input \Ki[11] ;
    output \PID_CONTROLLER.integral_23__N_3715[0] ;
    input \Kp[7] ;
    input \Kp[1] ;
    input \Kp[0] ;
    input \Kp[8] ;
    input \Kp[9] ;
    output n43055;
    input \Kp[10] ;
    input \Kp[13] ;
    input \Kp[2] ;
    input [23:0]IntegralLimit;
    input \Kp[11] ;
    output n155;
    output \PID_CONTROLLER.integral_23__N_3715[15] ;
    input \Ki[1] ;
    output \PID_CONTROLLER.integral_23__N_3715[14] ;
    input \Ki[0] ;
    output n367;
    input VCC_net;
    output n375;
    output n376;
    input \Kp[12] ;
    output [23:0]\PID_CONTROLLER.integral ;
    input \Ki[2] ;
    input \Kp[3] ;
    input \Kp[14] ;
    input n53;
    input \Kp[4] ;
    input \Kp[15] ;
    input \Kp[5] ;
    input \Kp[6] ;
    input \Ki[12] ;
    input \Ki[13] ;
    input [23:0]PWMLimit;
    input \Ki[14] ;
    input \Ki[15] ;
    input \Ki[4] ;
    input n4;
    input [23:0]setpoint;
    input n16;
    input n3;
    output n18;
    input \motor_state[21] ;
    input \motor_state[20] ;
    input \motor_state[19] ;
    input \Ki[5] ;
    input \motor_state[18] ;
    output n28;
    output \PID_CONTROLLER.integral_23__N_3715[13] ;
    input \PID_CONTROLLER.integral_23__N_3715[12] ;
    input \Ki[3] ;
    output n214;
    output \PID_CONTROLLER.integral_23__N_3715[16] ;
    input n29560;
    input \Ki[6] ;
    input \Ki[7] ;
    input \Ki[8] ;
    input \Ki[9] ;
    input \Ki[10] ;
    output \PID_CONTROLLER.integral_23__N_3715[11] ;
    input \motor_state[17] ;
    output \PID_CONTROLLER.integral_23__N_3715[10] ;
    input n30387;
    input n30386;
    input n30385;
    input n30384;
    input n30383;
    input n30382;
    input n30381;
    input n30380;
    input n30379;
    input n30378;
    input n30377;
    input n30376;
    input n30374;
    input n30372;
    input n30371;
    input n30370;
    input n30369;
    input n30368;
    input n30367;
    input n30366;
    input n30365;
    input n30364;
    input n30363;
    output \PID_CONTROLLER.integral_23__N_3715[9] ;
    output \PID_CONTROLLER.integral_23__N_3715[20] ;
    input n36816;
    output n20183;
    output \PID_CONTROLLER.integral_23__N_3715[8] ;
    output \PID_CONTROLLER.integral_23__N_3715[23] ;
    input n20;
    input \motor_state[15] ;
    input \motor_state[14] ;
    input n490;
    input n417;
    input n20136;
    input n344;
    input \motor_state[13] ;
    input n20137;
    input n271;
    input n20138;
    input n198;
    output \PID_CONTROLLER.integral_23__N_3715[7] ;
    input \motor_state[12] ;
    input n56;
    input n125;
    input \motor_state[11] ;
    output n455;
    output n456;
    input \motor_state[10] ;
    input \motor_state[9] ;
    input \motor_state[8] ;
    input \motor_state[7] ;
    input n41635;
    input \motor_state[5] ;
    input \motor_state[4] ;
    input \motor_state[3] ;
    input \motor_state[2] ;
    input \motor_state[1] ;
    input \motor_state[0] ;
    output n401;
    output n33;
    output n361;
    output \PID_CONTROLLER.integral_23__N_3715[6] ;
    output \PID_CONTROLLER.integral_23__N_3715[5] ;
    input [23:0]deadband;
    input n38;
    input n110;
    output \PID_CONTROLLER.integral_23__N_3715[4] ;
    output \PID_CONTROLLER.integral_23__N_3715[3] ;
    output \PID_CONTROLLER.integral_23__N_3715[21] ;
    input n37330;
    output n11597;
    input n131;
    input n204;
    output n4_adj_30;
    output n20182;
    input n31;
    output \PID_CONTROLLER.integral_23__N_3715[22] ;
    input n20_adj_31;
    output n212;
    output n213;
    output \PID_CONTROLLER.integral_23__N_3715[2] ;
    output n219;
    output n230;
    input n19;
    input \PID_CONTROLLER.integral_23__N_3715[1] ;
    input n4_adj_32;
    input n20181;
    input n6;
    input n36845;
    output n20209;
    input n6_adj_33;
    input n27629;
    
    wire clk16MHz /* synthesis SET_AS_NETWORK=clk16MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    
    wire n13, n11, n9, n67196, n68872, n51427;
    wire [14:0]n17517;
    
    wire n314, n51428, n19_c, n17, n15, n68864;
    wire [23:0]n182;
    wire [23:0]n1;
    
    wire n51157, n51083;
    wire [43:0]n257;
    wire [47:0]n49;
    
    wire n51084;
    wire [15:0]n16974;
    
    wire n241, n51426, n51546;
    wire [7:0]n19847;
    
    wire n189, n51547, n25, n23, n21, n69778;
    wire [23:0]n51;
    wire [21:0]n12096;
    wire [20:0]n13158;
    
    wire n51645, n804;
    wire [23:0]n55;
    
    wire n539, n31_c, n29, n27, n69213, n95, n51158, n37, n35, 
        n33_c, n69853, n43, n16_c, n6_c, n69394, n26, n69395, 
        n612, n8, n45, n24, n68096, n68048, n68024, n68942, 
        n68259;
    wire [23:0]n130;
    
    wire n4_c, n69357, n69358, n685, n758, n68070, n68066, n51646;
    wire [8:0]n19689;
    
    wire n47, n116_adj_5143, n51644;
    wire [31:0]counter;   // verilog/motorControl.v(21[11:18])
    
    wire n18_c, n12, n61767, n30, n28_c, n51156;
    wire [18:0]n14921;
    wire [17:0]n15680;
    
    wire n51545, n168, n51425, n51544;
    wire [23:0]n352;
    
    wire n51082, counter_31__N_3714, n29_adj_5144, n27_adj_5145, n30_adj_5146, 
        n10_adj_5147, n68063, n69728, n10_adj_5148, n68261, n51543, 
        n9_adj_5149, n950, n51542, n51155, n69920, n61348, n69921, 
        n1099, n51643, n1108, n51541, n1026, n51642, n1035, n51540, 
        n51154, n39, n69890, n962, n51539, n41, n68051, n51153, 
        n51152, n889, n51538, n69583, n953, n51641, n831, n51151, 
        n816, n51537, n880, n51640, n51081, n181;
    wire [23:0]n207;
    
    wire n743, n51536, n807, n51639, n68267, n69788, n670, n51535, 
        n51080, n51150, n597, n51534, n524, n51533, n51149, n734, 
        n51638, n451, n51532, n51148, n378, n51531, n661, n51637, 
        n305, n51530, n51079, n51078, n51077, n51147, n51076, 
        n51146, n232, n51529, n588, n51636, n51145, n159, n51528, 
        n17_adj_5159, n86, n51144, n51075, n515, n51635, n442, 
        n51634, n51143, n51074, n369_adj_5161, n51633, n51142;
    wire [6:0]n19971;
    wire [5:0]n20065;
    
    wire n560, n51410, n51073, n487, n51409, n296_adj_5164, n51632, 
        n414, n51408, n51072, n223, n51631, n341_adj_5165, n51407, 
        n268, n51406, n150, n51630, n904, n8_adj_5166, n77, n51071, 
        n195_adj_5167, n51405;
    wire [19:0]n14082;
    
    wire n51629, n51070, n977, n80, n11_adj_5168, n1050, n1023, 
        n51628, n122_adj_5169, n51627, n51626;
    wire [5:0]n20004;
    
    wire n61804, n490_c, n51985;
    wire [4:0]n20087;
    
    wire n417_c, n51984, n51625;
    wire [13:0]n17996;
    
    wire n1120, n51404, n51624;
    wire [11:0]n18778;
    wire [10:0]n19089;
    
    wire n910, n51279, n51069, n1047, n51403, n344_adj_5170, n51983, 
        n837, n51278, n51068, n764, n51277, n1102, n51623, n974, 
        n51402, n691, n51276, n51067, n271_c, n51982, n618, n51275;
    wire [16:0]n16363;
    
    wire n51510, n901, n51401, n51509, n198_adj_5171, n51981, n51508, 
        n545, n51274, n51066, n1029, n51622, n828, n51400, n472, 
        n51273, n1111, n51507, n51065, n153_adj_5172, n956, n51621, 
        n755, n51399, n1038, n51506, n399, n51272, n51064, n51063, 
        n326, n51271, n965, n51505, n51062, n682, n51398, n883, 
        n51620, n253, n51270, n892, n51504, n609, n51397, n819, 
        n51503, n180, n51269, n536, n51396, n51061, n746, n51502, 
        n38_c, n107_adj_5173, n51060, n463, n51395, n56_c, n125_c, 
        n51059, n390, n51394, n673, n51501, n51058, n810, n51619, 
        n600, n51500, n317, n51393, n737, n51618, n527, n51499, 
        n244, n51392;
    wire [0:0]n11637;
    
    wire n51701, n664, n51617, n171, n51391, n51700, n454, n51498, 
        n51699, n29_adj_5174, n98, n591, n51616, n381, n51497, 
        n51057, n51698, n51056, n308, n51496, n518, n51615, n1096, 
        n51055, n226, n235, n51495, n51054, n51053, n51697, n51052, 
        n299_adj_5176, n445, n51614, n162, n51494, n20_adj_5177, 
        n89, n372_adj_5178, n51613, n51696, n51051, n51695, n51694, 
        n51612, n51050, n51049, n293_adj_5179, n877, n950_adj_5180;
    wire [23:0]n1_adj_5682;
    
    wire n1023_adj_5181, n1096_adj_5182, n51611, n51693, n27_adj_5183, 
        n29_adj_5184, n338_adj_5185, n15_adj_5186, n9_adj_5187, n13_adj_5188, 
        n51610, n110_adj_5189, n51692, n11_adj_5190, n41_adj_5191, 
        n183_adj_5192;
    wire [12:0]n18415;
    
    wire n51377, n51376, n69325, n51375, n51048, n256, n69326, 
        n51374, n67907, n68768, n6_adj_5195, n8_adj_5196, n51691, 
        n51047, n68289, n69259, n329, n402, n25_adj_5199, n33_adj_5200, 
        n475, n51373, n51046, n51372, n548;
    wire [31:0]n57;
    
    wire n52331, n52330, n51371, n52329, n51045, n52328, n621, 
        n51370, n51044, n694, n52327, n767, n840, n52326, n466, 
        n51369, n393, n51368, n52325, n52324, n320, n51367, n50735, 
        n63605, n877_adj_5211, n51690, n52323, n411, n52322;
    wire [2:0]n20185;
    
    wire n4_adj_5214, n366_adj_5215, n347_adj_5216, n6_adj_5217, n59071, 
        n51043, n247, n51366, n63601, n62, n50749, n61580, n63591, 
        n71499, n63595, n8_adj_5219, n6_adj_5220, n41_adj_5221, n183_adj_5222, 
        n256_adj_5223, n329_adj_5225, n402_adj_5226, n475_adj_5227, 
        n548_adj_5228, n387, n621_adj_5229, n694_adj_5230, n767_adj_5231, 
        n52321, n840_adj_5233, n107_adj_5234, n180_adj_5235, n253_adj_5236, 
        n326_adj_5237, n399_adj_5238, n472_adj_5239, n545_adj_5240, 
        n618_adj_5241, n691_adj_5242, n764_adj_5243, n837_adj_5258, 
        n910_adj_5259, n122_adj_5260, n52320, n52319, n53_adj_5261, 
        n195_adj_5262, n51042, n52318, n268_adj_5263, n52317, n341_adj_5264, 
        n414_adj_5265, n487_adj_5266, n560_adj_5267, n104, n67202, 
        n52316, n35_adj_5270, n177, n67423, n250, n323, n396, 
        n460, n804_adj_5273, n51689, n174, n51365, n731, n51688, 
        n658, n51687, n469, n52315, n32_adj_5275, n101, n542, 
        n52314, n262, n615, n688, n585, n51686, n52313, n533, 
        n761, n512, n51685, n335, n834, n630, n51477, n557, 
        n51476, n907, n980, n52312;
    wire [23:0]n432;
    
    wire n67830, n101_adj_5277, n32_adj_5278, n606, n174_adj_5279, 
        n484, n51475, n439, n51684, n247_adj_5280, n320_adj_5281, 
        n52311, n52310, n393_adj_5282, n466_adj_5283, n539_adj_5284, 
        n51683, n612_adj_5285, n67844, n685_adj_5286, n52309, n51474, 
        n758_adj_5287, n52308, n831_adj_5288, n904_adj_5289, n977_adj_5290, 
        n1050_adj_5291, n52307, n52306, n119_adj_5292, n50_adj_5293, 
        n52305, n52304, n52303, n192_adj_5294, n265, n338_adj_5295, 
        n411_adj_5297, n484_adj_5298, n557_adj_5299, n51210, n408, 
        n630_adj_5300, n51209, n51208, n52302;
    wire [9:0]n19352;
    
    wire n52705, n52704, n98_adj_5301, n52703, n51207, n52702, n29_adj_5302, 
        n679, n171_adj_5303, n244_adj_5304, n317_adj_5305, n390_adj_5306, 
        n52701, n463_adj_5307, n52700, n752, n52699, n536_adj_5308, 
        n52698, n609_adj_5309, n51206, n52697, n52696, n825;
    wire [0:0]n12213;
    wire [21:0]n12720;
    
    wire n52695, n52694, n682_adj_5310, n51041, n51473, n52693, 
        n52692, n755_adj_5313, n52691, n481, n52690, n52689, n52688, 
        n52687, n52301, n52686, n828_adj_5315, n51040, n51205, n52685, 
        n52684, n51682, n901_adj_5316, n898, n52683, n974_adj_5317, 
        n971, n731_adj_5318, n52682, n658_adj_5319, n52681, n554, 
        n51204, n585_adj_5322, n52680, n512_adj_5323, n52679, n439_adj_5324, 
        n52678, n366_adj_5325, n52677, n293_adj_5326, n52676, n220, 
        n52675, n147_adj_5327, n52674, n220_adj_5328, n51681, n5_adj_5329, 
        n74, n1047_adj_5330;
    wire [20:0]n13685;
    
    wire n52673, n52672, n265_adj_5331, n51472, n52671, n51203, 
        n51039, n147_adj_5333, n51680, n52670, n52669, n52668, n51202, 
        n192_adj_5335, n51471, n52667, n61429, n51352;
    wire [4:0]n20133;
    
    wire n51351, n1099_adj_5338, n52666, n51201, n1026_adj_5341, n52665, 
        n5_adj_5342, n74_adj_5343, n51200, n953_adj_5345, n52664, 
        n880_adj_5346, n52663, n50_adj_5347, n119_adj_5348, n807_adj_5349, 
        n52662, n51350;
    wire [9:0]n19493;
    
    wire n770, n51679, n734_adj_5351, n52661, n697, n51678, n51199, 
        n661_adj_5353, n52660, n51038, n51198, n588_adj_5356, n52659, 
        n51470, n515_adj_5357, n52658, n1120_adj_5358, n51349, n624, 
        n51677, n51348, n442_adj_5361, n52657, n51197, n369_adj_5363, 
        n52656, n95_adj_5364, n551, n51676, n51196, n51037, n51195, 
        n478, n51675, n405, n51674, n51469, n296_adj_5369, n52655, 
        n980_adj_5370, n51347, n51194, n223_adj_5372, n52654, n26_adj_5373, 
        n150_adj_5374, n52653, n51193, n1114, n51468, n907_adj_5376, 
        n51346, n168_adj_5377, n627, n8_adj_5378, n77_adj_5379, n332_adj_5380, 
        n51673, n51192;
    wire [19:0]n14563;
    
    wire n52652, n51590, n51589, n52651, n1041, n51467, n52650, 
        n52649, n52648, n834_adj_5383, n51345, n52647, n761_adj_5384, 
        n51344, n51191, n1102_adj_5386, n52646, n51190, n1029_adj_5388, 
        n52645, n968, n51466, n956_adj_5389, n52644, n883_adj_5390, 
        n52643, n688_adj_5391, n51343, n895, n51465, n51189, n810_adj_5394, 
        n52642, n737_adj_5395, n52641, n664_adj_5396, n52640, n615_adj_5397, 
        n51342, n591_adj_5398, n52639, n518_adj_5399, n52638, n51588, 
        n259, n51672, n445_adj_5400, n52637, n51036, n372_adj_5401, 
        n52636, n299_adj_5402, n52635, n186_adj_5403, n51671, n226_adj_5404, 
        n52634, n153_adj_5405, n52633, n51587, n11_adj_5406, n80_adj_5407, 
        n822, n51464, n542_adj_5408, n51341, n51188;
    wire [18:0]n15359;
    
    wire n52632, n52631, n469_adj_5410, n51340, n241_adj_5411, n52630, 
        n52629, n52628, n1105, n52627, n44_adj_5413, n113_adj_5414, 
        n749, n51463, n1032, n52626, n396_adj_5415, n51339, n51586, 
        n47_adj_5416;
    wire [23:0]n1_adj_5683;
    
    wire n51187;
    wire [23:0]n59;
    
    wire n51186, n51035, n1105_adj_5419, n51585, n676, n51462, n51034, 
        n323_adj_5420, n51338, n250_adj_5421, n51337, n314_adj_5422, 
        n51185, n603, n51461, n51184, n177_adj_5426, n51336, n35_adj_5427, 
        n104_adj_5428, n51033, n387_adj_5429, n959, n52625, n51183, 
        n886, n52624, n51182, n813, n52623, n51181, n740, n52622, 
        n530, n51460, n1032_adj_5433, n51584, n51032, n667, n52621, 
        n457, n51459, n594, n52620, n521, n52619, n959_adj_5434, 
        n51583, n51180, n51179, n384_adj_5438, n51458, n448_adj_5439, 
        n52618, n51031, n375_adj_5440, n52617, n302, n52616, n51178, 
        n229, n52615, n51030, n311, n51457, n156_adj_5442, n52614, 
        n886_adj_5443, n51582, n14_adj_5444, n83, n813_adj_5445, n51581;
    wire [17:0]n16077;
    
    wire n52613, n52612, n740_adj_5446, n51580, n52611, n238, n51456, 
        n667_adj_5447, n51579, n51177, n52610, n51029, n165_adj_5449, 
        n51455, n1108_adj_5450, n52609, n594_adj_5451, n51578, n1035_adj_5452, 
        n52608, n521_adj_5453, n51577, n23_adj_5454, n92, n962_adj_5455, 
        n52607, n448_adj_5456, n51576, n51176, n51028, n889_adj_5459, 
        n52606, n1044, n51175, n375_adj_5461, n51575, n816_adj_5462, 
        n52605, n743_adj_5463, n52604, n51027, n51174, n302_adj_5465, 
        n51574, n670_adj_5466, n52603, n51026, n229_adj_5467, n51573, 
        n156_adj_5468, n51572, n597_adj_5469, n52602, n51173, n524_adj_5472, 
        n52601, n51172, n51094, n451_adj_5474, n52600, n51093, n14_adj_5475, 
        n83_adj_5476, n51171, n51170, n51092, n460_adj_5480, n51169, 
        n51091, n51168, n51090, n378_adj_5483, n52599, n51167, n305_adj_5486, 
        n52598, n232_adj_5487, n52597, n51089, n159_adj_5488, n52596, 
        n17_adj_5489, n86_adj_5490;
    wire [8:0]n19571;
    
    wire n770_adj_5491, n52595, n697_adj_5492, n52594, n624_adj_5493, 
        n52593, n551_adj_5494, n52592, n478_adj_5495, n52591, n51166, 
        n405_adj_5497, n52590, n332_adj_5498, n52589, n533_adj_5499, 
        n259_adj_5500, n52588, n186_adj_5501, n52587, n44_adj_5502, 
        n113_adj_5503;
    wire [16:0]n16721;
    
    wire n52586, n52585, n606_adj_5504, n52584, n51165, n1111_adj_5506, 
        n52583, n1038_adj_5507, n52582, n965_adj_5508, n52581, n679_adj_5509, 
        n892_adj_5510, n52580, n819_adj_5511, n52579, n746_adj_5512, 
        n52578, n37313, n673_adj_5515, n52577, n600_adj_5516, n52576, 
        n51088, n527_adj_5517, n52575, n454_adj_5518, n52574, n381_adj_5519, 
        n52573, n308_adj_5520, n52572, n51087, n235_adj_5521, n52571, 
        n162_adj_5522, n52570, n51164, n20_adj_5524, n89_adj_5525;
    wire [15:0]n17295;
    
    wire n52569, n52568, n51163, n1114_adj_5527, n52567, n1041_adj_5528, 
        n52566, n968_adj_5529, n52565, n895_adj_5530, n52564, n822_adj_5531, 
        n52563, n51162, n749_adj_5533, n52562, n676_adj_5534, n52561, 
        n752_adj_5535, n51161, n603_adj_5537, n52560, n51086, n530_adj_5538, 
        n52559, n457_adj_5539, n52558, n51160, n384_adj_5541, n52557, 
        n51085, n311_adj_5542, n52556, n825_adj_5543, n898_adj_5544, 
        n971_adj_5545, n1044_adj_5546, n238_adj_5547, n52555, n165_adj_5548, 
        n52554, n23_adj_5549, n92_adj_5550;
    wire [7:0]n19750;
    
    wire n700, n52553, n627_adj_5551, n52552, n1117, n51439, n554_adj_5552, 
        n52551, n700_adj_5553, n51553, n481_adj_5554, n52550, n408_adj_5555, 
        n52549, n116_adj_5556, n47_adj_5557, n335_adj_5558, n52548, 
        n189_adj_5559, n1117_adj_5560, n262_adj_5561, n52547, n51438, 
        n52546;
    wire [14:0]n17803;
    
    wire n52545, n52544, n52543, n52542, n52541, n52540, n52539, 
        n52538, n52537, n52536, n52535, n51437, n52534, n52533, 
        n52532, n51552, n52531;
    wire [13:0]n18249;
    
    wire n52530, n52529, n51551, n51436, n52528, n51435, n52527, 
        n52526, n51550, n52525, n52524, n51434, n52523, n52522, 
        n51433, n52521, n52520, n51650, n52519, n52518, n52517, 
        n51432;
    wire [6:0]n19893;
    
    wire n52516, n51549, n52515, n52514, n52513, n51159, n52512, 
        n52511, n52510;
    wire [12:0]n18637;
    
    wire n52509, n52508, n52507, n52506, n52505, n52504, n52503, 
        n52502, n52501, n52500, n52499, n52498, n52497, n51649, 
        n51431;
    wire [11:0]n18971;
    
    wire n52496, n52495, n51648, n52494, n51548, n52493, n51430, 
        n52492, n52491, n52490, n52489, n51429, n52488, n52487, 
        n52486, n52485, n52484, n52483, n52482, n52481, n52480, 
        n52479;
    wire [10:0]n19255;
    
    wire n52478, n52477, n52476, n52475, n52474, n52473, n52472, 
        n52471, n52470, n52469, n52468, n52467, n52466, n52465, 
        n52464, n52463, n52462, n52461, n52460, n51647, n52459, 
        n52458, n67952, n67962, n67494, n6_adj_5564;
    wire [2:0]n20207;
    
    wire n50890, n69824, n11595, n67885, n67891, n61943, n6_adj_5565, 
        n67871, n27827, n27822, n4_adj_5566, n27817, n62_adj_5567, 
        n27812, n27807, n27802, n41_adj_5571, n39_adj_5572, n68012, 
        n45_adj_5573, n43_adj_5574, n37_adj_5575, n6_adj_5576, n29_adj_5577, 
        n31_adj_5578, n21_adj_5579, n23_adj_5580, n25_adj_5581, n17_adj_5582, 
        n9_adj_5583, n35_adj_5584, n33_adj_5585, n11_adj_5586, n13_adj_5587, 
        n15_adj_5588, n27_adj_5589, n41_adj_5590, n37_adj_5591, n39_adj_5592, 
        n35_adj_5593, n23_adj_5594, n21_adj_5595, n67893, n67887, 
        n26_adj_5597, n28_adj_5598, n24_adj_5599, n22_adj_5600, n32_adj_5601, 
        n69736, n69737, n69628, n69472, n69827, n68293, n69906, 
        n69907, n405_adj_5603, n67946, n68798, n71315, n68786, n71309, 
        n67942, n68794, n71330, n68792, n71325, n16_adj_5605, n67909, 
        n8_adj_5607, n24_adj_5608, n67950, n71323, n67948, n71351, 
        n69175, n71348, n68796, n27797, n69478, n67933, n27792, 
        n71313, n69169, n27787, n71341, n69724, n71304, n69939, 
        n71301, n67978, n12_adj_5611, n10_adj_5612, n30_adj_5613, 
        n68832, n68828, n69770, n69191, n69851, n69343, n16_adj_5615, 
        n8_adj_5616, n24_adj_5617, n67984, n69344, n67954, n69255, 
        n68269, n12_adj_5618, n69329, n69330, n27782, n27777, n67921, 
        n71336, n10_adj_5620, n30_adj_5621, n67923, n69734, n68281, 
        n69926, n69927, n6_adj_5622, n69333, n69334, n27772, n67913, 
        n71298, n69257, n68279, n27767, n69884, n67915, n27762, 
        n69587, n27757, n27752, n68287, n4_adj_5623, n69339, n69340, 
        n27747, n67969, n69732, n68271, n69924, n69925, n69886, 
        n67956, n69585, n27742, n68277, n69790, n69792, n27737, 
        n63567, n27732, n27727, n27722, n39_adj_5625, n41_adj_5626;
    wire [1:0]n20216;
    
    wire n45_adj_5627, n43_adj_5628, n37_adj_5629, n23_adj_5630, n25_adj_5631, 
        n29_adj_5632, n31_adj_5633, n35_adj_5634, n11_adj_5635, n13_adj_5636, 
        n27_adj_5637, n15_adj_5638, n33_adj_5639, n9_adj_5640, n17_adj_5641, 
        n140_adj_5642, n63559, n19_adj_5643, n63581, n21_adj_5644, 
        n67858, n4_adj_5645, n50839, n67850, n12_adj_5646, n63561, 
        n10_adj_5647, n61017, n30_adj_5648, n68736, n68732, n69700, 
        n69141, n69819, n8_adj_5649, n69319, n16_adj_5651, n8_adj_5652, 
        n24_adj_5653, n69320, n67834, n69263, n68295, n69317, n69318, 
        n67846, n69738, n68297, n69928, n69929, n69880, n67836, 
        n69591, n68303, n69796, n69797, n41_adj_5654, n39_adj_5655, 
        n45_adj_5656, n43_adj_5657, n29_adj_5658, n31_adj_5659, n23_adj_5660, 
        n25_adj_5661, n37_adj_5662, n35_adj_5663, n33_adj_5664, n9_adj_5665, 
        n17_adj_5666, n19_adj_5667, n21_adj_5668, n11_adj_5669, n13_adj_5670, 
        n15_adj_5671, n27_adj_5672, n67458, n67445, n12_adj_5673, 
        n10_adj_5674, n30_adj_5675, n68388, n68376, n69613, n68964, 
        n69798, n16_adj_5676, n69251, n69252, n8_adj_5677, n24_adj_5678, 
        n67234, n68940, n68255, n4_adj_5679, n69037, n69038, n67431, 
        n69825, n68257, n69966, n69967, n69933, n67281, n69579, 
        n40_adj_5680, n69581, n12_adj_5681;
    
    SB_LUT4 i53178_4_lut (.I0(n13), .I1(n11), .I2(n9), .I3(n67196), 
            .O(n68872));
    defparam i53178_4_lut.LUT_INIT = 16'heeef;
    SB_CARRY add_6292_5 (.CI(n51427), .I0(n17517[2]), .I1(n314), .CO(n51428));
    SB_LUT4 i53170_4_lut (.I0(n19_c), .I1(n17), .I2(n15), .I3(n68872), 
            .O(n68864));
    defparam i53170_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 unary_minus_13_add_3_18_lut (.I0(GND_net), .I1(GND_net), .I2(n1[16]), 
            .I3(n51157), .O(n182[16])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_18_14 (.CI(n51083), .I0(n257[12]), .I1(n49[12]), .CO(n51084));
    SB_LUT4 add_6292_4_lut (.I0(GND_net), .I1(n17517[1]), .I2(n241), .I3(n51426), 
            .O(n16974[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6292_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6478_3 (.CI(n51546), .I0(n19847[0]), .I1(n189), .CO(n51547));
    SB_LUT4 i54084_4_lut (.I0(n25), .I1(n23), .I2(n21), .I3(n68864), 
            .O(n69778));
    defparam i54084_4_lut.LUT_INIT = 16'hfffe;
    SB_DFFER result__i0 (.Q(duty[0]), .C(clk16MHz), .E(control_update), 
            .D(n51[0]), .R(reset));   // verilog/motorControl.v(41[14] 62[8])
    SB_LUT4 add_6037_18_lut (.I0(GND_net), .I1(n13158[15]), .I2(GND_net), 
            .I3(n51645), .O(n12096[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6037_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6292_4 (.CI(n51426), .I0(n17517[1]), .I1(n241), .CO(n51427));
    SB_LUT4 mult_17_i541_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3715[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n804));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i541_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i363_2_lut (.I0(\Kp[7] ), .I1(n55[13]), .I2(GND_net), 
            .I3(GND_net), .O(n539));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i363_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i53519_4_lut (.I0(n31_c), .I1(n29), .I2(n27), .I3(n69778), 
            .O(n69213));
    defparam i53519_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 mult_16_i65_2_lut (.I0(\Kp[1] ), .I1(n55[11]), .I2(GND_net), 
            .I3(GND_net), .O(n95));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i65_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY unary_minus_13_add_3_18 (.CI(n51157), .I0(GND_net), .I1(n1[16]), 
            .CO(n51158));
    SB_LUT4 i54159_4_lut (.I0(n37), .I1(n35), .I2(n33_c), .I3(n69213), 
            .O(n69853));
    defparam i54159_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 LessThan_12_i16_3_lut (.I0(n182[9]), .I1(n182[21]), .I2(n43), 
            .I3(GND_net), .O(n16_c));   // verilog/motorControl.v(48[21:44])
    defparam LessThan_12_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53700_3_lut (.I0(n6_c), .I1(n182[10]), .I2(n21), .I3(GND_net), 
            .O(n69394));   // verilog/motorControl.v(48[21:44])
    defparam i53700_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_16_i18_2_lut (.I0(\Kp[0] ), .I1(n55[12]), .I2(GND_net), 
            .I3(GND_net), .O(n26));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i18_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i53701_3_lut (.I0(n69394), .I1(n182[11]), .I2(n23), .I3(GND_net), 
            .O(n69395));   // verilog/motorControl.v(48[21:44])
    defparam i53701_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_16_i412_2_lut (.I0(\Kp[8] ), .I1(n55[13]), .I2(GND_net), 
            .I3(GND_net), .O(n612));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i412_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_12_i8_3_lut (.I0(n182[4]), .I1(n182[8]), .I2(n17), 
            .I3(GND_net), .O(n8));   // verilog/motorControl.v(48[21:44])
    defparam LessThan_12_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_12_i24_3_lut (.I0(n16_c), .I1(n182[22]), .I2(n45), 
            .I3(GND_net), .O(n24));   // verilog/motorControl.v(48[21:44])
    defparam LessThan_12_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52354_4_lut (.I0(n43), .I1(n25), .I2(n23), .I3(n68096), 
            .O(n68048));
    defparam i52354_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i53248_4_lut (.I0(n24), .I1(n8), .I2(n45), .I3(n68024), 
            .O(n68942));   // verilog/motorControl.v(48[21:44])
    defparam i53248_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i52565_3_lut (.I0(n69395), .I1(n182[12]), .I2(n25), .I3(GND_net), 
            .O(n68259));   // verilog/motorControl.v(48[21:44])
    defparam i52565_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_12_i4_4_lut (.I0(n130[0]), .I1(n182[1]), .I2(n130[1]), 
            .I3(n182[0]), .O(n4_c));   // verilog/motorControl.v(48[21:44])
    defparam LessThan_12_i4_4_lut.LUT_INIT = 16'h4d0c;
    SB_LUT4 i53663_3_lut (.I0(n4_c), .I1(n182[13]), .I2(n27), .I3(GND_net), 
            .O(n69357));   // verilog/motorControl.v(48[21:44])
    defparam i53663_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53664_3_lut (.I0(n69357), .I1(n182[14]), .I2(n29), .I3(GND_net), 
            .O(n69358));   // verilog/motorControl.v(48[21:44])
    defparam i53664_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_16_i461_2_lut (.I0(\Kp[9] ), .I1(n55[13]), .I2(GND_net), 
            .I3(GND_net), .O(n685));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i461_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i29162_1_lut (.I0(duty[0]), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n43055));   // verilog/motorControl.v(41[14] 62[8])
    defparam i29162_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_16_i510_2_lut (.I0(\Kp[10] ), .I1(n55[13]), .I2(GND_net), 
            .I3(GND_net), .O(n758));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i510_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i52372_4_lut (.I0(n33_c), .I1(n31_c), .I2(n29), .I3(n68070), 
            .O(n68066));
    defparam i52372_4_lut.LUT_INIT = 16'haaab;
    SB_CARRY add_6037_18 (.CI(n51645), .I0(n13158[15]), .I1(GND_net), 
            .CO(n51646));
    SB_LUT4 add_6478_2_lut (.I0(GND_net), .I1(n47), .I2(n116_adj_5143), 
            .I3(GND_net), .O(n19689[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6478_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6037_17_lut (.I0(GND_net), .I1(n13158[14]), .I2(GND_net), 
            .I3(n51644), .O(n12096[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6037_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6478_2 (.CI(GND_net), .I0(n47), .I1(n116_adj_5143), .CO(n51546));
    SB_LUT4 i1_2_lut (.I0(counter[23]), .I1(counter[24]), .I2(GND_net), 
            .I3(GND_net), .O(n18_c));
    defparam i1_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i5_4_lut (.I0(counter[1]), .I1(counter[4]), .I2(counter[5]), 
            .I3(counter[6]), .O(n12));
    defparam i5_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i6_4_lut (.I0(counter[3]), .I1(n12), .I2(counter[2]), .I3(counter[0]), 
            .O(n61767));
    defparam i6_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_4_lut (.I0(counter[15]), .I1(counter[19]), .I2(counter[25]), 
            .I3(n18_c), .O(n30));
    defparam i13_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i11_4_lut (.I0(counter[21]), .I1(counter[27]), .I2(counter[26]), 
            .I3(counter[30]), .O(n28_c));
    defparam i11_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 unary_minus_13_add_3_17_lut (.I0(GND_net), .I1(GND_net), .I2(n1[15]), 
            .I3(n51156), .O(n182[15])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6187_20_lut (.I0(GND_net), .I1(n15680[17]), .I2(GND_net), 
            .I3(n51545), .O(n14921[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6187_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6292_3_lut (.I0(GND_net), .I1(n17517[0]), .I2(n168), .I3(n51425), 
            .O(n16974[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6292_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6187_19_lut (.I0(GND_net), .I1(n15680[16]), .I2(GND_net), 
            .I3(n51544), .O(n14921[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6187_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6187_19 (.CI(n51544), .I0(n15680[16]), .I1(GND_net), 
            .CO(n51545));
    SB_LUT4 add_18_13_lut (.I0(GND_net), .I1(n257[11]), .I2(n49[11]), 
            .I3(n51082), .O(n352[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_13_lut.LUT_INIT = 16'hC33C;
    SB_DFF control_update_37 (.Q(control_update), .C(clk16MHz), .D(counter_31__N_3714));   // verilog/motorControl.v(23[10] 30[6])
    SB_CARRY add_6292_3 (.CI(n51425), .I0(n17517[0]), .I1(n168), .CO(n51426));
    SB_LUT4 i12_4_lut (.I0(counter[20]), .I1(counter[22]), .I2(counter[14]), 
            .I3(counter[18]), .O(n29_adj_5144));
    defparam i12_4_lut.LUT_INIT = 16'hfffe;
    SB_CARRY unary_minus_13_add_3_17 (.CI(n51156), .I0(GND_net), .I1(n1[15]), 
            .CO(n51157));
    SB_LUT4 i10_4_lut (.I0(counter[29]), .I1(counter[28]), .I2(counter[17]), 
            .I3(counter[16]), .O(n27_adj_5145));
    defparam i10_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i54034_4_lut (.I0(n30_adj_5146), .I1(n10_adj_5147), .I2(n35), 
            .I3(n68063), .O(n69728));   // verilog/motorControl.v(48[21:44])
    defparam i54034_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i4_4_lut (.I0(counter[13]), .I1(counter[9]), .I2(counter[10]), 
            .I3(counter[11]), .O(n10_adj_5148));
    defparam i4_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 add_6292_2_lut (.I0(GND_net), .I1(n26), .I2(n95), .I3(GND_net), 
            .O(n16974[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6292_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6037_17 (.CI(n51644), .I0(n13158[14]), .I1(GND_net), 
            .CO(n51645));
    SB_LUT4 i52567_3_lut (.I0(n69358), .I1(n182[15]), .I2(n31_c), .I3(GND_net), 
            .O(n68261));   // verilog/motorControl.v(48[21:44])
    defparam i52567_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_6187_18_lut (.I0(GND_net), .I1(n15680[15]), .I2(GND_net), 
            .I3(n51543), .O(n14921[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6187_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i3_4_lut (.I0(counter[12]), .I1(n61767), .I2(counter[8]), 
            .I3(counter[7]), .O(n9_adj_5149));
    defparam i3_4_lut.LUT_INIT = 16'ha8a0;
    SB_CARRY add_6187_18 (.CI(n51543), .I0(n15680[15]), .I1(GND_net), 
            .CO(n51544));
    SB_LUT4 mult_16_i639_2_lut (.I0(\Kp[13] ), .I1(n55[4]), .I2(GND_net), 
            .I3(GND_net), .O(n950));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i639_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6187_17_lut (.I0(GND_net), .I1(n15680[14]), .I2(GND_net), 
            .I3(n51542), .O(n14921[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6187_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_13_add_3_16_lut (.I0(GND_net), .I1(GND_net), .I2(n1[14]), 
            .I3(n51155), .O(n182[14])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i54226_4_lut (.I0(n68261), .I1(n69728), .I2(n35), .I3(n68066), 
            .O(n69920));   // verilog/motorControl.v(48[21:44])
    defparam i54226_4_lut.LUT_INIT = 16'hccca;
    SB_CARRY add_6292_2 (.CI(GND_net), .I0(n26), .I1(n95), .CO(n51425));
    SB_LUT4 i16_4_lut (.I0(n27_adj_5145), .I1(n29_adj_5144), .I2(n28_c), 
            .I3(n30), .O(n61348));
    defparam i16_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i29155_4_lut (.I0(n61348), .I1(counter[31]), .I2(n9_adj_5149), 
            .I3(n10_adj_5148), .O(counter_31__N_3714));   // verilog/motorControl.v(26[8:41])
    defparam i29155_4_lut.LUT_INIT = 16'h3222;
    SB_LUT4 i54227_3_lut (.I0(n69920), .I1(n182[18]), .I2(n37), .I3(GND_net), 
            .O(n69921));   // verilog/motorControl.v(48[21:44])
    defparam i54227_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_18_13 (.CI(n51082), .I0(n257[11]), .I1(n49[11]), .CO(n51083));
    SB_LUT4 add_6037_16_lut (.I0(GND_net), .I1(n13158[13]), .I2(n1099), 
            .I3(n51643), .O(n12096[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6037_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i114_2_lut (.I0(\Kp[2] ), .I1(n55[11]), .I2(GND_net), 
            .I3(GND_net), .O(n168));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i114_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6187_17 (.CI(n51542), .I0(n15680[14]), .I1(GND_net), 
            .CO(n51543));
    SB_LUT4 add_6187_16_lut (.I0(GND_net), .I1(n15680[13]), .I2(n1108), 
            .I3(n51541), .O(n14921[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6187_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6187_16 (.CI(n51541), .I0(n15680[13]), .I1(n1108), .CO(n51542));
    SB_CARRY add_6037_16 (.CI(n51643), .I0(n13158[13]), .I1(n1099), .CO(n51644));
    SB_LUT4 add_6037_15_lut (.I0(GND_net), .I1(n13158[12]), .I2(n1026), 
            .I3(n51642), .O(n12096[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6037_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6187_15_lut (.I0(GND_net), .I1(n15680[12]), .I2(n1035), 
            .I3(n51540), .O(n14921[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6187_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_13_inv_0_i16_1_lut (.I0(IntegralLimit[15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[15]));   // verilog/motorControl.v(49[22:36])
    defparam unary_minus_13_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY unary_minus_13_add_3_16 (.CI(n51155), .I0(GND_net), .I1(n1[14]), 
            .CO(n51156));
    SB_CARRY add_6187_15 (.CI(n51540), .I0(n15680[12]), .I1(n1035), .CO(n51541));
    SB_LUT4 unary_minus_13_add_3_15_lut (.I0(GND_net), .I1(GND_net), .I2(n1[13]), 
            .I3(n51154), .O(n182[13])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i54196_3_lut (.I0(n69921), .I1(n182[19]), .I2(n39), .I3(GND_net), 
            .O(n69890));   // verilog/motorControl.v(48[21:44])
    defparam i54196_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_6187_14_lut (.I0(GND_net), .I1(n15680[11]), .I2(n962), 
            .I3(n51539), .O(n14921[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6187_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i52357_4_lut (.I0(n43), .I1(n41), .I2(n39), .I3(n69853), 
            .O(n68051));
    defparam i52357_4_lut.LUT_INIT = 16'haaab;
    SB_CARRY unary_minus_13_add_3_15 (.CI(n51154), .I0(GND_net), .I1(n1[13]), 
            .CO(n51155));
    SB_CARRY add_6037_15 (.CI(n51642), .I0(n13158[12]), .I1(n1026), .CO(n51643));
    SB_CARRY add_6187_14 (.CI(n51539), .I0(n15680[11]), .I1(n962), .CO(n51540));
    SB_LUT4 unary_minus_13_add_3_14_lut (.I0(GND_net), .I1(GND_net), .I2(n1[12]), 
            .I3(n51153), .O(n182[12])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_13_add_3_14 (.CI(n51153), .I0(GND_net), .I1(n1[12]), 
            .CO(n51154));
    SB_LUT4 unary_minus_13_add_3_13_lut (.I0(GND_net), .I1(GND_net), .I2(n1[11]), 
            .I3(n51152), .O(n182[11])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6187_13_lut (.I0(GND_net), .I1(n15680[10]), .I2(n889), 
            .I3(n51538), .O(n14921[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6187_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i53889_4_lut (.I0(n68259), .I1(n68942), .I2(n45), .I3(n68048), 
            .O(n69583));   // verilog/motorControl.v(48[21:44])
    defparam i53889_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 add_6037_14_lut (.I0(GND_net), .I1(n13158[11]), .I2(n953), 
            .I3(n51641), .O(n12096[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6037_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_13_add_3_13 (.CI(n51152), .I0(GND_net), .I1(n1[11]), 
            .CO(n51153));
    SB_LUT4 mult_16_i559_2_lut (.I0(\Kp[11] ), .I1(n55[13]), .I2(GND_net), 
            .I3(GND_net), .O(n831));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i559_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_13_add_3_12_lut (.I0(GND_net), .I1(GND_net), .I2(n1[10]), 
            .I3(n51151), .O(n182[10])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6187_13 (.CI(n51538), .I0(n15680[10]), .I1(n889), .CO(n51539));
    SB_CARRY add_6037_14 (.CI(n51641), .I0(n13158[11]), .I1(n953), .CO(n51642));
    SB_LUT4 add_6187_12_lut (.I0(GND_net), .I1(n15680[9]), .I2(n816), 
            .I3(n51537), .O(n14921[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6187_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_13_add_3_12 (.CI(n51151), .I0(GND_net), .I1(n1[10]), 
            .CO(n51152));
    SB_LUT4 add_6037_13_lut (.I0(GND_net), .I1(n13158[10]), .I2(n880), 
            .I3(n51640), .O(n12096[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6037_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_18_12_lut (.I0(GND_net), .I1(n257[10]), .I2(n49[10]), 
            .I3(n51081), .O(n352[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6187_12 (.CI(n51537), .I0(n15680[9]), .I1(n816), .CO(n51538));
    SB_LUT4 mux_14_i16_3_lut (.I0(n130[15]), .I1(n182[15]), .I2(n181), 
            .I3(GND_net), .O(n207[15]));   // verilog/motorControl.v(48[18] 50[12])
    defparam mux_14_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_15_i16_3_lut (.I0(n207[15]), .I1(IntegralLimit[15]), .I2(n155), 
            .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3715[15] ));   // verilog/motorControl.v(48[18] 50[12])
    defparam mux_15_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_6037_13 (.CI(n51640), .I0(n13158[10]), .I1(n880), .CO(n51641));
    SB_LUT4 mult_17_i79_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3715[14] ), 
            .I2(GND_net), .I3(GND_net), .O(n116_adj_5143));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i79_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_18_12 (.CI(n51081), .I0(n257[10]), .I1(n49[10]), .CO(n51082));
    SB_LUT4 add_6187_11_lut (.I0(GND_net), .I1(n15680[8]), .I2(n743), 
            .I3(n51536), .O(n14921[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6187_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6187_11 (.CI(n51536), .I0(n15680[8]), .I1(n743), .CO(n51537));
    SB_LUT4 add_6037_12_lut (.I0(GND_net), .I1(n13158[9]), .I2(n807), 
            .I3(n51639), .O(n12096[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6037_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i52573_3_lut (.I0(n69890), .I1(n182[20]), .I2(n41), .I3(GND_net), 
            .O(n68267));   // verilog/motorControl.v(48[21:44])
    defparam i52573_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_17_i32_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3715[15] ), 
            .I2(GND_net), .I3(GND_net), .O(n47));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i32_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i54094_4_lut (.I0(n68267), .I1(n69583), .I2(n45), .I3(n68051), 
            .O(n69788));   // verilog/motorControl.v(48[21:44])
    defparam i54094_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 add_6187_10_lut (.I0(GND_net), .I1(n15680[7]), .I2(n670), 
            .I3(n51535), .O(n14921[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6187_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_18_11_lut (.I0(GND_net), .I1(n257[9]), .I2(n49[9]), .I3(n51080), 
            .O(n367)) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6187_10 (.CI(n51535), .I0(n15680[7]), .I1(n670), .CO(n51536));
    SB_LUT4 unary_minus_13_add_3_11_lut (.I0(GND_net), .I1(GND_net), .I2(n1[9]), 
            .I3(n51150), .O(n182[9])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_18_11 (.CI(n51080), .I0(n257[9]), .I1(n49[9]), .CO(n51081));
    SB_LUT4 add_6187_9_lut (.I0(GND_net), .I1(n15680[6]), .I2(n597), .I3(n51534), 
            .O(n14921[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6187_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_13_add_3_11 (.CI(n51150), .I0(GND_net), .I1(n1[9]), 
            .CO(n51151));
    SB_CARRY add_6037_12 (.CI(n51639), .I0(n13158[9]), .I1(n807), .CO(n51640));
    SB_CARRY add_6187_9 (.CI(n51534), .I0(n15680[6]), .I1(n597), .CO(n51535));
    SB_LUT4 add_6187_8_lut (.I0(GND_net), .I1(n15680[5]), .I2(n524), .I3(n51533), 
            .O(n14921[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6187_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6187_8 (.CI(n51533), .I0(n15680[5]), .I1(n524), .CO(n51534));
    SB_LUT4 unary_minus_13_add_3_10_lut (.I0(GND_net), .I1(GND_net), .I2(n1[8]), 
            .I3(n51149), .O(n182[8])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6037_11_lut (.I0(GND_net), .I1(n13158[8]), .I2(n734), 
            .I3(n51638), .O(n12096[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6037_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6187_7_lut (.I0(GND_net), .I1(n15680[4]), .I2(n451), .I3(n51532), 
            .O(n14921[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6187_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6187_7 (.CI(n51532), .I0(n15680[4]), .I1(n451), .CO(n51533));
    SB_CARRY unary_minus_13_add_3_10 (.CI(n51149), .I0(GND_net), .I1(n1[8]), 
            .CO(n51150));
    SB_LUT4 unary_minus_13_add_3_9_lut (.I0(GND_net), .I1(GND_net), .I2(n1[7]), 
            .I3(n51148), .O(n182[7])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6187_6_lut (.I0(GND_net), .I1(n15680[3]), .I2(n378), .I3(n51531), 
            .O(n14921[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6187_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6037_11 (.CI(n51638), .I0(n13158[8]), .I1(n734), .CO(n51639));
    SB_LUT4 add_6037_10_lut (.I0(GND_net), .I1(n13158[7]), .I2(n661), 
            .I3(n51637), .O(n12096[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6037_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6187_6 (.CI(n51531), .I0(n15680[3]), .I1(n378), .CO(n51532));
    SB_LUT4 add_6187_5_lut (.I0(GND_net), .I1(n15680[2]), .I2(n305), .I3(n51530), 
            .O(n14921[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6187_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_18_10_lut (.I0(GND_net), .I1(n257[8]), .I2(n49[8]), .I3(n51079), 
            .O(n352[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6187_5 (.CI(n51530), .I0(n15680[2]), .I1(n305), .CO(n51531));
    SB_CARRY add_18_10 (.CI(n51079), .I0(n257[8]), .I1(n49[8]), .CO(n51080));
    SB_LUT4 add_18_9_lut (.I0(GND_net), .I1(n257[7]), .I2(n49[7]), .I3(n51078), 
            .O(n352[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_18_9 (.CI(n51078), .I0(n257[7]), .I1(n49[7]), .CO(n51079));
    SB_LUT4 add_18_8_lut (.I0(GND_net), .I1(n257[6]), .I2(n49[6]), .I3(n51077), 
            .O(n352[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_13_add_3_9 (.CI(n51148), .I0(GND_net), .I1(n1[7]), 
            .CO(n51149));
    SB_CARRY add_18_8 (.CI(n51077), .I0(n257[6]), .I1(n49[6]), .CO(n51078));
    SB_LUT4 unary_minus_13_add_3_8_lut (.I0(GND_net), .I1(GND_net), .I2(n1[6]), 
            .I3(n51147), .O(n182[6])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_18_7_lut (.I0(GND_net), .I1(n257[5]), .I2(n49[5]), .I3(n51076), 
            .O(n352[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_13_add_3_8 (.CI(n51147), .I0(GND_net), .I1(n1[6]), 
            .CO(n51148));
    SB_LUT4 i54095_3_lut (.I0(n69788), .I1(n130[23]), .I2(n182[23]), .I3(GND_net), 
            .O(n181));   // verilog/motorControl.v(48[21:44])
    defparam i54095_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 unary_minus_13_add_3_7_lut (.I0(GND_net), .I1(GND_net), .I2(n1[5]), 
            .I3(n51146), .O(n182[5])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_18_7 (.CI(n51076), .I0(n257[5]), .I1(n49[5]), .CO(n51077));
    SB_LUT4 add_6187_4_lut (.I0(GND_net), .I1(n15680[1]), .I2(n232), .I3(n51529), 
            .O(n14921[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6187_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6037_10 (.CI(n51637), .I0(n13158[7]), .I1(n661), .CO(n51638));
    SB_LUT4 add_6037_9_lut (.I0(GND_net), .I1(n13158[6]), .I2(n588), .I3(n51636), 
            .O(n12096[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6037_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_13_add_3_7 (.CI(n51146), .I0(GND_net), .I1(n1[5]), 
            .CO(n51147));
    SB_CARRY add_6187_4 (.CI(n51529), .I0(n15680[1]), .I1(n232), .CO(n51530));
    SB_LUT4 unary_minus_13_add_3_6_lut (.I0(GND_net), .I1(GND_net), .I2(n1[4]), 
            .I3(n51145), .O(n182[4])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6187_3_lut (.I0(GND_net), .I1(n15680[0]), .I2(n159), .I3(n51528), 
            .O(n14921[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6187_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6037_9 (.CI(n51636), .I0(n13158[6]), .I1(n588), .CO(n51637));
    SB_CARRY unary_minus_13_add_3_6 (.CI(n51145), .I0(GND_net), .I1(n1[4]), 
            .CO(n51146));
    SB_CARRY add_6187_3 (.CI(n51528), .I0(n15680[0]), .I1(n159), .CO(n51529));
    SB_LUT4 add_6187_2_lut (.I0(GND_net), .I1(n17_adj_5159), .I2(n86), 
            .I3(GND_net), .O(n14921[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6187_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_13_add_3_5_lut (.I0(GND_net), .I1(GND_net), .I2(n1[3]), 
            .I3(n51144), .O(n182[3])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_18_6_lut (.I0(GND_net), .I1(n257[4]), .I2(n49[4]), .I3(n51075), 
            .O(n352[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6187_2 (.CI(GND_net), .I0(n17_adj_5159), .I1(n86), .CO(n51528));
    SB_LUT4 add_6037_8_lut (.I0(GND_net), .I1(n13158[5]), .I2(n515), .I3(n51635), 
            .O(n12096[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6037_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6037_8 (.CI(n51635), .I0(n13158[5]), .I1(n515), .CO(n51636));
    SB_LUT4 add_6037_7_lut (.I0(GND_net), .I1(n13158[4]), .I2(n442), .I3(n51634), 
            .O(n12096[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6037_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_18_6 (.CI(n51075), .I0(n257[4]), .I1(n49[4]), .CO(n51076));
    SB_CARRY unary_minus_13_add_3_5 (.CI(n51144), .I0(GND_net), .I1(n1[3]), 
            .CO(n51145));
    SB_CARRY add_6037_7 (.CI(n51634), .I0(n13158[4]), .I1(n442), .CO(n51635));
    SB_LUT4 unary_minus_13_add_3_4_lut (.I0(GND_net), .I1(GND_net), .I2(n1[2]), 
            .I3(n51143), .O(n182[2])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_18_5_lut (.I0(GND_net), .I1(n257[3]), .I2(n49[3]), .I3(n51074), 
            .O(n352[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6037_6_lut (.I0(GND_net), .I1(n13158[3]), .I2(n369_adj_5161), 
            .I3(n51633), .O(n12096[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6037_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_13_add_3_4 (.CI(n51143), .I0(GND_net), .I1(n1[2]), 
            .CO(n51144));
    SB_LUT4 unary_minus_13_add_3_3_lut (.I0(GND_net), .I1(GND_net), .I2(n1[1]), 
            .I3(n51142), .O(n182[1])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6508_8_lut (.I0(GND_net), .I1(n20065[5]), .I2(n560), .I3(n51410), 
            .O(n19971[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6508_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_18_5 (.CI(n51074), .I0(n257[3]), .I1(n49[3]), .CO(n51075));
    SB_CARRY unary_minus_13_add_3_3 (.CI(n51142), .I0(GND_net), .I1(n1[1]), 
            .CO(n51143));
    SB_LUT4 mux_14_i15_3_lut (.I0(n130[14]), .I1(n182[14]), .I2(n181), 
            .I3(GND_net), .O(n207[14]));   // verilog/motorControl.v(48[18] 50[12])
    defparam mux_14_i15_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_13_add_3_2_lut (.I0(GND_net), .I1(GND_net), .I2(n1[0]), 
            .I3(VCC_net), .O(n182[0])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_13_add_3_2 (.CI(VCC_net), .I0(GND_net), .I1(n1[0]), 
            .CO(n51142));
    SB_LUT4 add_18_4_lut (.I0(GND_net), .I1(n257[2]), .I2(n49[2]), .I3(n51073), 
            .O(n352[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6037_6 (.CI(n51633), .I0(n13158[3]), .I1(n369_adj_5161), 
            .CO(n51634));
    SB_LUT4 add_6508_7_lut (.I0(GND_net), .I1(n20065[4]), .I2(n487), .I3(n51409), 
            .O(n19971[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6508_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6037_5_lut (.I0(GND_net), .I1(n13158[2]), .I2(n296_adj_5164), 
            .I3(n51632), .O(n12096[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6037_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6508_7 (.CI(n51409), .I0(n20065[4]), .I1(n487), .CO(n51410));
    SB_CARRY add_6037_5 (.CI(n51632), .I0(n13158[2]), .I1(n296_adj_5164), 
            .CO(n51633));
    SB_LUT4 add_6508_6_lut (.I0(GND_net), .I1(n20065[3]), .I2(n414), .I3(n51408), 
            .O(n19971[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6508_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_18_4 (.CI(n51073), .I0(n257[2]), .I1(n49[2]), .CO(n51074));
    SB_LUT4 add_18_3_lut (.I0(GND_net), .I1(n257[1]), .I2(n49[1]), .I3(n51072), 
            .O(n375)) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6508_6 (.CI(n51408), .I0(n20065[3]), .I1(n414), .CO(n51409));
    SB_LUT4 add_6037_4_lut (.I0(GND_net), .I1(n13158[1]), .I2(n223), .I3(n51631), 
            .O(n12096[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6037_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6508_5_lut (.I0(GND_net), .I1(n20065[2]), .I2(n341_adj_5165), 
            .I3(n51407), .O(n19971[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6508_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6508_5 (.CI(n51407), .I0(n20065[2]), .I1(n341_adj_5165), 
            .CO(n51408));
    SB_CARRY add_6037_4 (.CI(n51631), .I0(n13158[1]), .I1(n223), .CO(n51632));
    SB_CARRY add_18_3 (.CI(n51072), .I0(n257[1]), .I1(n49[1]), .CO(n51073));
    SB_LUT4 add_6508_4_lut (.I0(GND_net), .I1(n20065[1]), .I2(n268), .I3(n51406), 
            .O(n19971[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6508_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_18_2_lut (.I0(GND_net), .I1(n257[0]), .I2(n49[0]), .I3(GND_net), 
            .O(n376)) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6037_3_lut (.I0(GND_net), .I1(n13158[0]), .I2(n150), .I3(n51630), 
            .O(n12096[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6037_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_18_2 (.CI(GND_net), .I0(n257[0]), .I1(n49[0]), .CO(n51072));
    SB_CARRY add_6508_4 (.CI(n51406), .I0(n20065[1]), .I1(n268), .CO(n51407));
    SB_LUT4 mult_16_i608_2_lut (.I0(\Kp[12] ), .I1(n55[13]), .I2(GND_net), 
            .I3(GND_net), .O(n904));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i608_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6037_3 (.CI(n51630), .I0(n13158[0]), .I1(n150), .CO(n51631));
    SB_LUT4 add_6037_2_lut (.I0(GND_net), .I1(n8_adj_5166), .I2(n77), 
            .I3(GND_net), .O(n12096[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6037_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_9_25_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [23]), 
            .I2(n55[23]), .I3(n51071), .O(n130[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_15_i15_3_lut (.I0(n207[14]), .I1(IntegralLimit[14]), .I2(n155), 
            .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3715[14] ));   // verilog/motorControl.v(48[18] 50[12])
    defparam mux_15_i15_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_6037_2 (.CI(GND_net), .I0(n8_adj_5166), .I1(n77), .CO(n51630));
    SB_LUT4 add_6508_3_lut (.I0(GND_net), .I1(n20065[0]), .I2(n195_adj_5167), 
            .I3(n51405), .O(n19971[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6508_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6106_22_lut (.I0(GND_net), .I1(n14082[19]), .I2(GND_net), 
            .I3(n51629), .O(n13158[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6106_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_9_24_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [22]), 
            .I2(n55[23]), .I3(n51070), .O(n130[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_i128_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3715[14] ), 
            .I2(GND_net), .I3(GND_net), .O(n189));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i128_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i657_2_lut (.I0(\Kp[13] ), .I1(n55[13]), .I2(GND_net), 
            .I3(GND_net), .O(n977));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i657_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i55_2_lut (.I0(\Kp[1] ), .I1(n55[6]), .I2(GND_net), 
            .I3(GND_net), .O(n80));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i55_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i8_2_lut (.I0(\Kp[0] ), .I1(n55[7]), .I2(GND_net), 
            .I3(GND_net), .O(n11_adj_5168));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i8_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i163_2_lut (.I0(\Kp[3] ), .I1(n55[11]), .I2(GND_net), 
            .I3(GND_net), .O(n241));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i163_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_13_inv_0_i17_1_lut (.I0(IntegralLimit[16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[16]));   // verilog/motorControl.v(49[22:36])
    defparam unary_minus_13_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_16_i706_2_lut (.I0(\Kp[14] ), .I1(n55[13]), .I2(GND_net), 
            .I3(GND_net), .O(n1050));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i706_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i688_2_lut (.I0(\Kp[14] ), .I1(n55[4]), .I2(GND_net), 
            .I3(GND_net), .O(n1023));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i688_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6106_21_lut (.I0(GND_net), .I1(n14082[18]), .I2(GND_net), 
            .I3(n51628), .O(n13158[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6106_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6106_21 (.CI(n51628), .I0(n14082[18]), .I1(GND_net), 
            .CO(n51629));
    SB_CARRY add_6508_3 (.CI(n51405), .I0(n20065[0]), .I1(n195_adj_5167), 
            .CO(n51406));
    SB_LUT4 add_6508_2_lut (.I0(GND_net), .I1(n53), .I2(n122_adj_5169), 
            .I3(GND_net), .O(n19971[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6508_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6106_20_lut (.I0(GND_net), .I1(n14082[17]), .I2(GND_net), 
            .I3(n51627), .O(n13158[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6106_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6508_2 (.CI(GND_net), .I0(n53), .I1(n122_adj_5169), .CO(n51405));
    SB_CARRY add_6106_20 (.CI(n51627), .I0(n14082[17]), .I1(GND_net), 
            .CO(n51628));
    SB_LUT4 add_6106_19_lut (.I0(GND_net), .I1(n14082[16]), .I2(GND_net), 
            .I3(n51626), .O(n13158[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6106_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6106_19 (.CI(n51626), .I0(n14082[16]), .I1(GND_net), 
            .CO(n51627));
    SB_LUT4 add_6512_7_lut (.I0(GND_net), .I1(n61804), .I2(n490_c), .I3(n51985), 
            .O(n20004[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6512_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6512_6_lut (.I0(GND_net), .I1(n20087[3]), .I2(n417_c), 
            .I3(n51984), .O(n20004[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6512_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6106_18_lut (.I0(GND_net), .I1(n14082[15]), .I2(GND_net), 
            .I3(n51625), .O(n13158[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6106_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6106_18 (.CI(n51625), .I0(n14082[15]), .I1(GND_net), 
            .CO(n51626));
    SB_CARRY add_9_24 (.CI(n51070), .I0(\PID_CONTROLLER.integral [22]), 
            .I1(n55[23]), .CO(n51071));
    SB_LUT4 add_6323_16_lut (.I0(GND_net), .I1(n17996[13]), .I2(n1120), 
            .I3(n51404), .O(n17517[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6323_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6106_17_lut (.I0(GND_net), .I1(n14082[14]), .I2(GND_net), 
            .I3(n51624), .O(n13158[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6106_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6404_13_lut (.I0(GND_net), .I1(n19089[10]), .I2(n910), 
            .I3(n51279), .O(n18778[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6404_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_9_23_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [21]), 
            .I2(n55[23]), .I3(n51069), .O(n130[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_9_23 (.CI(n51069), .I0(\PID_CONTROLLER.integral [21]), 
            .I1(n55[23]), .CO(n51070));
    SB_LUT4 add_6323_15_lut (.I0(GND_net), .I1(n17996[12]), .I2(n1047), 
            .I3(n51403), .O(n17517[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6323_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6106_17 (.CI(n51624), .I0(n14082[14]), .I1(GND_net), 
            .CO(n51625));
    SB_CARRY add_6512_6 (.CI(n51984), .I0(n20087[3]), .I1(n417_c), .CO(n51985));
    SB_CARRY add_6323_15 (.CI(n51403), .I0(n17996[12]), .I1(n1047), .CO(n51404));
    SB_LUT4 add_6512_5_lut (.I0(GND_net), .I1(n20087[2]), .I2(n344_adj_5170), 
            .I3(n51983), .O(n20004[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6512_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6512_5 (.CI(n51983), .I0(n20087[2]), .I1(n344_adj_5170), 
            .CO(n51984));
    SB_LUT4 add_6404_12_lut (.I0(GND_net), .I1(n19089[9]), .I2(n837), 
            .I3(n51278), .O(n18778[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6404_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6404_12 (.CI(n51278), .I0(n19089[9]), .I1(n837), .CO(n51279));
    SB_LUT4 add_9_22_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [20]), 
            .I2(n55[23]), .I3(n51068), .O(n130[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6404_11_lut (.I0(GND_net), .I1(n19089[8]), .I2(n764), 
            .I3(n51277), .O(n18778[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6404_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6404_11 (.CI(n51277), .I0(n19089[8]), .I1(n764), .CO(n51278));
    SB_LUT4 add_6106_16_lut (.I0(GND_net), .I1(n14082[13]), .I2(n1102), 
            .I3(n51623), .O(n13158[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6106_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6323_14_lut (.I0(GND_net), .I1(n17996[11]), .I2(n974), 
            .I3(n51402), .O(n17517[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6323_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_9_22 (.CI(n51068), .I0(\PID_CONTROLLER.integral [20]), 
            .I1(n55[23]), .CO(n51069));
    SB_LUT4 add_6404_10_lut (.I0(GND_net), .I1(n19089[7]), .I2(n691), 
            .I3(n51276), .O(n18778[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6404_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_9_21_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [19]), 
            .I2(n55[23]), .I3(n51067), .O(n130[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6404_10 (.CI(n51276), .I0(n19089[7]), .I1(n691), .CO(n51277));
    SB_LUT4 add_6512_4_lut (.I0(GND_net), .I1(n20087[1]), .I2(n271_c), 
            .I3(n51982), .O(n20004[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6512_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6512_4 (.CI(n51982), .I0(n20087[1]), .I1(n271_c), .CO(n51983));
    SB_LUT4 add_6404_9_lut (.I0(GND_net), .I1(n19089[6]), .I2(n618), .I3(n51275), 
            .O(n18778[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6404_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6106_16 (.CI(n51623), .I0(n14082[13]), .I1(n1102), .CO(n51624));
    SB_LUT4 add_6224_19_lut (.I0(GND_net), .I1(n16363[16]), .I2(GND_net), 
            .I3(n51510), .O(n15680[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6224_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6323_14 (.CI(n51402), .I0(n17996[11]), .I1(n974), .CO(n51403));
    SB_LUT4 add_6323_13_lut (.I0(GND_net), .I1(n17996[10]), .I2(n901), 
            .I3(n51401), .O(n17517[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6323_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6224_18_lut (.I0(GND_net), .I1(n16363[15]), .I2(GND_net), 
            .I3(n51509), .O(n15680[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6224_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6512_3_lut (.I0(GND_net), .I1(n20087[0]), .I2(n198_adj_5171), 
            .I3(n51981), .O(n20004[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6512_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6224_18 (.CI(n51509), .I0(n16363[15]), .I1(GND_net), 
            .CO(n51510));
    SB_CARRY add_6404_9 (.CI(n51275), .I0(n19089[6]), .I1(n618), .CO(n51276));
    SB_CARRY add_6323_13 (.CI(n51401), .I0(n17996[10]), .I1(n901), .CO(n51402));
    SB_LUT4 add_6224_17_lut (.I0(GND_net), .I1(n16363[14]), .I2(GND_net), 
            .I3(n51508), .O(n15680[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6224_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6404_8_lut (.I0(GND_net), .I1(n19089[5]), .I2(n545), .I3(n51274), 
            .O(n18778[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6404_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_9_21 (.CI(n51067), .I0(\PID_CONTROLLER.integral [19]), 
            .I1(n55[23]), .CO(n51068));
    SB_LUT4 add_9_20_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [18]), 
            .I2(n55[22]), .I3(n51066), .O(n130[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6106_15_lut (.I0(GND_net), .I1(n14082[12]), .I2(n1029), 
            .I3(n51622), .O(n13158[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6106_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6323_12_lut (.I0(GND_net), .I1(n17996[9]), .I2(n828), 
            .I3(n51400), .O(n17517[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6323_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6404_8 (.CI(n51274), .I0(n19089[5]), .I1(n545), .CO(n51275));
    SB_LUT4 add_6404_7_lut (.I0(GND_net), .I1(n19089[4]), .I2(n472), .I3(n51273), 
            .O(n18778[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6404_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6224_17 (.CI(n51508), .I0(n16363[14]), .I1(GND_net), 
            .CO(n51509));
    SB_LUT4 add_6224_16_lut (.I0(GND_net), .I1(n16363[13]), .I2(n1111), 
            .I3(n51507), .O(n15680[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6224_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_9_20 (.CI(n51066), .I0(\PID_CONTROLLER.integral [18]), 
            .I1(n55[22]), .CO(n51067));
    SB_LUT4 add_9_19_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [17]), 
            .I2(n55[21]), .I3(n51065), .O(n130[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i104_2_lut (.I0(\Kp[2] ), .I1(n55[6]), .I2(GND_net), 
            .I3(GND_net), .O(n153_adj_5172));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i104_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6106_15 (.CI(n51622), .I0(n14082[12]), .I1(n1029), .CO(n51623));
    SB_CARRY add_6404_7 (.CI(n51273), .I0(n19089[4]), .I1(n472), .CO(n51274));
    SB_CARRY add_6224_16 (.CI(n51507), .I0(n16363[13]), .I1(n1111), .CO(n51508));
    SB_CARRY add_6323_12 (.CI(n51400), .I0(n17996[9]), .I1(n828), .CO(n51401));
    SB_LUT4 add_6106_14_lut (.I0(GND_net), .I1(n14082[11]), .I2(n956), 
            .I3(n51621), .O(n13158[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6106_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i212_2_lut (.I0(\Kp[4] ), .I1(n55[11]), .I2(GND_net), 
            .I3(GND_net), .O(n314));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i212_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6106_14 (.CI(n51621), .I0(n14082[11]), .I1(n956), .CO(n51622));
    SB_CARRY add_9_19 (.CI(n51065), .I0(\PID_CONTROLLER.integral [17]), 
            .I1(n55[21]), .CO(n51066));
    SB_LUT4 add_6323_11_lut (.I0(GND_net), .I1(n17996[8]), .I2(n755), 
            .I3(n51399), .O(n17517[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6323_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6224_15_lut (.I0(GND_net), .I1(n16363[12]), .I2(n1038), 
            .I3(n51506), .O(n15680[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6224_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6404_6_lut (.I0(GND_net), .I1(n19089[3]), .I2(n399), .I3(n51272), 
            .O(n18778[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6404_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_9_18_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [16]), 
            .I2(n55[20]), .I3(n51064), .O(n130[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_9_18 (.CI(n51064), .I0(\PID_CONTROLLER.integral [16]), 
            .I1(n55[20]), .CO(n51065));
    SB_LUT4 add_9_17_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [15]), 
            .I2(n55[19]), .I3(n51063), .O(n130[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6404_6 (.CI(n51272), .I0(n19089[3]), .I1(n399), .CO(n51273));
    SB_CARRY add_6323_11 (.CI(n51399), .I0(n17996[8]), .I1(n755), .CO(n51400));
    SB_LUT4 add_6404_5_lut (.I0(GND_net), .I1(n19089[2]), .I2(n326), .I3(n51271), 
            .O(n18778[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6404_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6224_15 (.CI(n51506), .I0(n16363[12]), .I1(n1038), .CO(n51507));
    SB_LUT4 add_6224_14_lut (.I0(GND_net), .I1(n16363[11]), .I2(n965), 
            .I3(n51505), .O(n15680[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6224_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_9_17 (.CI(n51063), .I0(\PID_CONTROLLER.integral [15]), 
            .I1(n55[19]), .CO(n51064));
    SB_LUT4 add_9_16_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [14]), 
            .I2(n55[18]), .I3(n51062), .O(n130[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6224_14 (.CI(n51505), .I0(n16363[11]), .I1(n965), .CO(n51506));
    SB_CARRY add_6404_5 (.CI(n51271), .I0(n19089[2]), .I1(n326), .CO(n51272));
    SB_LUT4 add_6323_10_lut (.I0(GND_net), .I1(n17996[7]), .I2(n682), 
            .I3(n51398), .O(n17517[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6323_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6106_13_lut (.I0(GND_net), .I1(n14082[10]), .I2(n883), 
            .I3(n51620), .O(n13158[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6106_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6404_4_lut (.I0(GND_net), .I1(n19089[1]), .I2(n253), .I3(n51270), 
            .O(n18778[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6404_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6224_13_lut (.I0(GND_net), .I1(n16363[10]), .I2(n892), 
            .I3(n51504), .O(n15680[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6224_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6323_10 (.CI(n51398), .I0(n17996[7]), .I1(n682), .CO(n51399));
    SB_LUT4 add_6323_9_lut (.I0(GND_net), .I1(n17996[6]), .I2(n609), .I3(n51397), 
            .O(n17517[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6323_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6404_4 (.CI(n51270), .I0(n19089[1]), .I1(n253), .CO(n51271));
    SB_CARRY add_6224_13 (.CI(n51504), .I0(n16363[10]), .I1(n892), .CO(n51505));
    SB_CARRY add_6512_3 (.CI(n51981), .I0(n20087[0]), .I1(n198_adj_5171), 
            .CO(n51982));
    SB_CARRY add_9_16 (.CI(n51062), .I0(\PID_CONTROLLER.integral [14]), 
            .I1(n55[18]), .CO(n51063));
    SB_LUT4 add_6224_12_lut (.I0(GND_net), .I1(n16363[9]), .I2(n819), 
            .I3(n51503), .O(n15680[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6224_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6404_3_lut (.I0(GND_net), .I1(n19089[0]), .I2(n180), .I3(n51269), 
            .O(n18778[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6404_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6323_9 (.CI(n51397), .I0(n17996[6]), .I1(n609), .CO(n51398));
    SB_CARRY add_6224_12 (.CI(n51503), .I0(n16363[9]), .I1(n819), .CO(n51504));
    SB_LUT4 add_6323_8_lut (.I0(GND_net), .I1(n17996[5]), .I2(n536), .I3(n51396), 
            .O(n17517[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6323_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6404_3 (.CI(n51269), .I0(n19089[0]), .I1(n180), .CO(n51270));
    SB_LUT4 add_9_15_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [13]), 
            .I2(n55[17]), .I3(n51061), .O(n130[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6224_11_lut (.I0(GND_net), .I1(n16363[8]), .I2(n746), 
            .I3(n51502), .O(n15680[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6224_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_9_15 (.CI(n51061), .I0(\PID_CONTROLLER.integral [13]), 
            .I1(n55[17]), .CO(n51062));
    SB_CARRY add_6323_8 (.CI(n51396), .I0(n17996[5]), .I1(n536), .CO(n51397));
    SB_LUT4 add_6404_2_lut (.I0(GND_net), .I1(n38_c), .I2(n107_adj_5173), 
            .I3(GND_net), .O(n18778[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6404_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6404_2 (.CI(GND_net), .I0(n38_c), .I1(n107_adj_5173), 
            .CO(n51269));
    SB_LUT4 add_9_14_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [12]), 
            .I2(n55[16]), .I3(n51060), .O(n130[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6323_7_lut (.I0(GND_net), .I1(n17996[4]), .I2(n463), .I3(n51395), 
            .O(n17517[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6323_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6512_2_lut (.I0(GND_net), .I1(n56_c), .I2(n125_c), .I3(GND_net), 
            .O(n20004[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6512_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_9_14 (.CI(n51060), .I0(\PID_CONTROLLER.integral [12]), 
            .I1(n55[16]), .CO(n51061));
    SB_CARRY add_6323_7 (.CI(n51395), .I0(n17996[4]), .I1(n463), .CO(n51396));
    SB_LUT4 add_9_13_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [11]), 
            .I2(n55[15]), .I3(n51059), .O(n130[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_9_13 (.CI(n51059), .I0(\PID_CONTROLLER.integral [11]), 
            .I1(n55[15]), .CO(n51060));
    SB_LUT4 add_6323_6_lut (.I0(GND_net), .I1(n17996[3]), .I2(n390), .I3(n51394), 
            .O(n17517[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6323_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6224_11 (.CI(n51502), .I0(n16363[8]), .I1(n746), .CO(n51503));
    SB_LUT4 add_6224_10_lut (.I0(GND_net), .I1(n16363[7]), .I2(n673), 
            .I3(n51501), .O(n15680[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6224_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_9_12_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [10]), 
            .I2(n55[14]), .I3(n51058), .O(n130[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6106_13 (.CI(n51620), .I0(n14082[10]), .I1(n883), .CO(n51621));
    SB_LUT4 add_6106_12_lut (.I0(GND_net), .I1(n14082[9]), .I2(n810), 
            .I3(n51619), .O(n13158[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6106_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6224_10 (.CI(n51501), .I0(n16363[7]), .I1(n673), .CO(n51502));
    SB_LUT4 add_6224_9_lut (.I0(GND_net), .I1(n16363[6]), .I2(n600), .I3(n51500), 
            .O(n15680[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6224_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6323_6 (.CI(n51394), .I0(n17996[3]), .I1(n390), .CO(n51395));
    SB_CARRY add_6106_12 (.CI(n51619), .I0(n14082[9]), .I1(n810), .CO(n51620));
    SB_LUT4 add_6323_5_lut (.I0(GND_net), .I1(n17996[2]), .I2(n317), .I3(n51393), 
            .O(n17517[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6323_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6106_11_lut (.I0(GND_net), .I1(n14082[8]), .I2(n737), 
            .I3(n51618), .O(n13158[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6106_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6512_2 (.CI(GND_net), .I0(n56_c), .I1(n125_c), .CO(n51981));
    SB_CARRY add_6323_5 (.CI(n51393), .I0(n17996[2]), .I1(n317), .CO(n51394));
    SB_CARRY add_6224_9 (.CI(n51500), .I0(n16363[6]), .I1(n600), .CO(n51501));
    SB_LUT4 add_6224_8_lut (.I0(GND_net), .I1(n16363[5]), .I2(n527), .I3(n51499), 
            .O(n15680[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6224_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6323_4_lut (.I0(GND_net), .I1(n17996[1]), .I2(n244), .I3(n51392), 
            .O(n17517[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6323_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6323_4 (.CI(n51392), .I0(n17996[1]), .I1(n244), .CO(n51393));
    SB_CARRY add_6106_11 (.CI(n51618), .I0(n14082[8]), .I1(n737), .CO(n51619));
    SB_LUT4 mult_16_add_1221_24_lut (.I0(n55[23]), .I1(n12096[21]), .I2(GND_net), 
            .I3(n51701), .O(n11637[0])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_16_add_1221_24_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_6106_10_lut (.I0(GND_net), .I1(n14082[7]), .I2(n664), 
            .I3(n51617), .O(n13158[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6106_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6323_3_lut (.I0(GND_net), .I1(n17996[0]), .I2(n171), .I3(n51391), 
            .O(n17517[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6323_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6323_3 (.CI(n51391), .I0(n17996[0]), .I1(n171), .CO(n51392));
    SB_CARRY add_6106_10 (.CI(n51617), .I0(n14082[7]), .I1(n664), .CO(n51618));
    SB_LUT4 mult_16_add_1221_23_lut (.I0(GND_net), .I1(n12096[20]), .I2(GND_net), 
            .I3(n51700), .O(n257[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_16_add_1221_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6224_8 (.CI(n51499), .I0(n16363[5]), .I1(n527), .CO(n51500));
    SB_CARRY mult_16_add_1221_23 (.CI(n51700), .I0(n12096[20]), .I1(GND_net), 
            .CO(n51701));
    SB_LUT4 add_6224_7_lut (.I0(GND_net), .I1(n16363[4]), .I2(n454), .I3(n51498), 
            .O(n15680[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6224_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_add_1221_22_lut (.I0(GND_net), .I1(n12096[19]), .I2(GND_net), 
            .I3(n51699), .O(n257[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_16_add_1221_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6323_2_lut (.I0(GND_net), .I1(n29_adj_5174), .I2(n98), 
            .I3(GND_net), .O(n17517[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6323_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6106_9_lut (.I0(GND_net), .I1(n14082[6]), .I2(n591), .I3(n51616), 
            .O(n13158[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6106_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6224_7 (.CI(n51498), .I0(n16363[4]), .I1(n454), .CO(n51499));
    SB_CARRY add_9_12 (.CI(n51058), .I0(\PID_CONTROLLER.integral [10]), 
            .I1(n55[14]), .CO(n51059));
    SB_LUT4 add_6224_6_lut (.I0(GND_net), .I1(n16363[3]), .I2(n381), .I3(n51497), 
            .O(n15680[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6224_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_9_11_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(n55[13]), .I3(n51057), .O(n130[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_16_add_1221_22 (.CI(n51699), .I0(n12096[19]), .I1(GND_net), 
            .CO(n51700));
    SB_CARRY add_6323_2 (.CI(GND_net), .I0(n29_adj_5174), .I1(n98), .CO(n51391));
    SB_CARRY add_9_11 (.CI(n51057), .I0(\PID_CONTROLLER.integral [9]), .I1(n55[13]), 
            .CO(n51058));
    SB_CARRY add_6106_9 (.CI(n51616), .I0(n14082[6]), .I1(n591), .CO(n51617));
    SB_LUT4 mult_16_add_1221_21_lut (.I0(GND_net), .I1(n12096[18]), .I2(GND_net), 
            .I3(n51698), .O(n257[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_16_add_1221_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6224_6 (.CI(n51497), .I0(n16363[3]), .I1(n381), .CO(n51498));
    SB_LUT4 add_9_10_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(n55[12]), .I3(n51056), .O(n130[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6224_5_lut (.I0(GND_net), .I1(n16363[2]), .I2(n308), .I3(n51496), 
            .O(n15680[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6224_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6106_8_lut (.I0(GND_net), .I1(n14082[5]), .I2(n518), .I3(n51615), 
            .O(n13158[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6106_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_9_10 (.CI(n51056), .I0(\PID_CONTROLLER.integral [8]), .I1(n55[12]), 
            .CO(n51057));
    SB_CARRY mult_16_add_1221_21 (.CI(n51698), .I0(n12096[18]), .I1(GND_net), 
            .CO(n51699));
    SB_LUT4 mult_16_i737_2_lut (.I0(\Kp[15] ), .I1(n55[4]), .I2(GND_net), 
            .I3(GND_net), .O(n1096));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i737_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_9_9_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(n55[11]), .I3(n51055), .O(n130[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_9_9 (.CI(n51055), .I0(\PID_CONTROLLER.integral [7]), .I1(n55[11]), 
            .CO(n51056));
    SB_LUT4 mult_16_i153_2_lut (.I0(\Kp[3] ), .I1(n55[6]), .I2(GND_net), 
            .I3(GND_net), .O(n226));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i153_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6106_8 (.CI(n51615), .I0(n14082[5]), .I1(n518), .CO(n51616));
    SB_CARRY add_6224_5 (.CI(n51496), .I0(n16363[2]), .I1(n308), .CO(n51497));
    SB_LUT4 add_6224_4_lut (.I0(GND_net), .I1(n16363[1]), .I2(n235), .I3(n51495), 
            .O(n15680[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6224_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_9_8_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(n55[10]), .I3(n51054), .O(n130[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6224_4 (.CI(n51495), .I0(n16363[1]), .I1(n235), .CO(n51496));
    SB_CARRY add_9_8 (.CI(n51054), .I0(\PID_CONTROLLER.integral [6]), .I1(n55[10]), 
            .CO(n51055));
    SB_LUT4 add_9_7_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(n55[9]), .I3(n51053), .O(n130[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_9_7 (.CI(n51053), .I0(\PID_CONTROLLER.integral [5]), .I1(n55[9]), 
            .CO(n51054));
    SB_LUT4 mult_16_add_1221_20_lut (.I0(GND_net), .I1(n12096[17]), .I2(GND_net), 
            .I3(n51697), .O(n257[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_16_add_1221_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_9_6_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(n55[8]), .I3(n51052), .O(n130[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i202_2_lut (.I0(\Kp[4] ), .I1(n55[6]), .I2(GND_net), 
            .I3(GND_net), .O(n299_adj_5176));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i202_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6106_7_lut (.I0(GND_net), .I1(n14082[4]), .I2(n445), .I3(n51614), 
            .O(n13158[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6106_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6224_3_lut (.I0(GND_net), .I1(n16363[0]), .I2(n162), .I3(n51494), 
            .O(n15680[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6224_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6224_3 (.CI(n51494), .I0(n16363[0]), .I1(n162), .CO(n51495));
    SB_CARRY mult_16_add_1221_20 (.CI(n51697), .I0(n12096[17]), .I1(GND_net), 
            .CO(n51698));
    SB_LUT4 add_6224_2_lut (.I0(GND_net), .I1(n20_adj_5177), .I2(n89), 
            .I3(GND_net), .O(n15680[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6224_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_9_6 (.CI(n51052), .I0(\PID_CONTROLLER.integral [4]), .I1(n55[8]), 
            .CO(n51053));
    SB_CARRY add_6106_7 (.CI(n51614), .I0(n14082[4]), .I1(n445), .CO(n51615));
    SB_LUT4 add_6106_6_lut (.I0(GND_net), .I1(n14082[3]), .I2(n372_adj_5178), 
            .I3(n51613), .O(n13158[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6106_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6224_2 (.CI(GND_net), .I0(n20_adj_5177), .I1(n89), .CO(n51494));
    SB_LUT4 mult_16_add_1221_19_lut (.I0(GND_net), .I1(n12096[16]), .I2(GND_net), 
            .I3(n51696), .O(n257[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_16_add_1221_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_16_add_1221_19 (.CI(n51696), .I0(n12096[16]), .I1(GND_net), 
            .CO(n51697));
    SB_LUT4 add_9_5_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(n55[7]), .I3(n51051), .O(n130[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6106_6 (.CI(n51613), .I0(n14082[3]), .I1(n372_adj_5178), 
            .CO(n51614));
    SB_CARRY add_9_5 (.CI(n51051), .I0(\PID_CONTROLLER.integral [3]), .I1(n55[7]), 
            .CO(n51052));
    SB_LUT4 mult_16_i251_2_lut (.I0(\Kp[5] ), .I1(n55[6]), .I2(GND_net), 
            .I3(GND_net), .O(n372_adj_5178));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i251_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i61_2_lut (.I0(\Kp[1] ), .I1(n55[9]), .I2(GND_net), 
            .I3(GND_net), .O(n89));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i61_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i14_2_lut (.I0(\Kp[0] ), .I1(n55[10]), .I2(GND_net), 
            .I3(GND_net), .O(n20_adj_5177));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i14_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_add_1221_18_lut (.I0(GND_net), .I1(n12096[15]), .I2(GND_net), 
            .I3(n51695), .O(n257[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_16_add_1221_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i110_2_lut (.I0(\Kp[2] ), .I1(n55[9]), .I2(GND_net), 
            .I3(GND_net), .O(n162));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i110_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i300_2_lut (.I0(\Kp[6] ), .I1(n55[6]), .I2(GND_net), 
            .I3(GND_net), .O(n445));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i300_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mult_16_add_1221_18 (.CI(n51695), .I0(n12096[15]), .I1(GND_net), 
            .CO(n51696));
    SB_LUT4 mult_16_add_1221_17_lut (.I0(GND_net), .I1(n12096[14]), .I2(GND_net), 
            .I3(n51694), .O(n257[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_16_add_1221_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6106_5_lut (.I0(GND_net), .I1(n14082[2]), .I2(n299_adj_5176), 
            .I3(n51612), .O(n13158[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6106_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_9_4_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(n55[6]), .I3(n51050), .O(n130[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6106_5 (.CI(n51612), .I0(n14082[2]), .I1(n299_adj_5176), 
            .CO(n51613));
    SB_CARRY add_9_4 (.CI(n51050), .I0(\PID_CONTROLLER.integral [2]), .I1(n55[6]), 
            .CO(n51051));
    SB_LUT4 add_9_3_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(n55[5]), .I3(n51049), .O(n130[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_16_add_1221_17 (.CI(n51694), .I0(n12096[14]), .I1(GND_net), 
            .CO(n51695));
    SB_CARRY add_9_3 (.CI(n51049), .I0(\PID_CONTROLLER.integral [1]), .I1(n55[5]), 
            .CO(n51050));
    SB_LUT4 mult_16_i198_2_lut (.I0(\Kp[4] ), .I1(n55[4]), .I2(GND_net), 
            .I3(GND_net), .O(n293_adj_5179));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i198_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i590_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3715[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n877));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i590_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i639_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3715[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n950_adj_5180));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i639_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i159_2_lut (.I0(\Kp[3] ), .I1(n55[9]), .I2(GND_net), 
            .I3(GND_net), .O(n235));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i159_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_26_inv_0_i19_1_lut (.I0(PWMLimit[18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5682[18]));   // verilog/motorControl.v(56[22:31])
    defparam unary_minus_26_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_17_i688_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3715[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n1023_adj_5181));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i688_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i349_2_lut (.I0(\Kp[7] ), .I1(n55[6]), .I2(GND_net), 
            .I3(GND_net), .O(n518));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i349_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i737_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3715[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n1096_adj_5182));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i737_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i208_2_lut (.I0(\Kp[4] ), .I1(n55[9]), .I2(GND_net), 
            .I3(GND_net), .O(n308));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i208_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6106_4_lut (.I0(GND_net), .I1(n14082[1]), .I2(n226), .I3(n51611), 
            .O(n13158[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6106_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_add_1221_16_lut (.I0(GND_net), .I1(n12096[13]), .I2(n1096), 
            .I3(n51693), .O(n257[15])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_16_add_1221_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6106_4 (.CI(n51611), .I0(n14082[1]), .I1(n226), .CO(n51612));
    SB_LUT4 mult_16_i257_2_lut (.I0(\Kp[5] ), .I1(n55[9]), .I2(GND_net), 
            .I3(GND_net), .O(n381));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i257_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_23_i27_2_lut (.I0(PWMLimit[13]), .I1(n352[13]), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_5183));   // verilog/motorControl.v(53[14:29])
    defparam LessThan_23_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_23_i29_2_lut (.I0(PWMLimit[14]), .I1(n352[14]), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_5184));   // verilog/motorControl.v(53[14:29])
    defparam LessThan_23_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_17_i228_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3715[15] ), 
            .I2(GND_net), .I3(GND_net), .O(n338_adj_5185));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i228_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_23_i15_2_lut (.I0(PWMLimit[7]), .I1(n352[7]), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_5186));   // verilog/motorControl.v(53[14:29])
    defparam LessThan_23_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_23_i9_2_lut (.I0(PWMLimit[4]), .I1(n352[4]), .I2(GND_net), 
            .I3(GND_net), .O(n9_adj_5187));   // verilog/motorControl.v(53[14:29])
    defparam LessThan_23_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_23_i13_2_lut (.I0(PWMLimit[6]), .I1(n352[6]), .I2(GND_net), 
            .I3(GND_net), .O(n13_adj_5188));   // verilog/motorControl.v(53[14:29])
    defparam LessThan_23_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_6106_3_lut (.I0(GND_net), .I1(n14082[0]), .I2(n153_adj_5172), 
            .I3(n51610), .O(n13158[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6106_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i75_2_lut (.I0(\Kp[1] ), .I1(n55[16]), .I2(GND_net), 
            .I3(GND_net), .O(n110_adj_5189));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i75_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mult_16_add_1221_16 (.CI(n51693), .I0(n12096[13]), .I1(n1096), 
            .CO(n51694));
    SB_LUT4 add_9_2_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [0]), 
            .I2(n55[4]), .I3(GND_net), .O(n130[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_add_1221_15_lut (.I0(GND_net), .I1(n12096[12]), .I2(n1023), 
            .I3(n51692), .O(n257[14])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_16_add_1221_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_23_i11_2_lut (.I0(PWMLimit[5]), .I1(n352[5]), .I2(GND_net), 
            .I3(GND_net), .O(n11_adj_5190));   // verilog/motorControl.v(53[14:29])
    defparam LessThan_23_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_16_i28_2_lut (.I0(\Kp[0] ), .I1(n55[17]), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_5191));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i28_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i398_2_lut (.I0(\Kp[8] ), .I1(n55[6]), .I2(GND_net), 
            .I3(GND_net), .O(n591));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i398_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i124_2_lut (.I0(\Kp[2] ), .I1(n55[16]), .I2(GND_net), 
            .I3(GND_net), .O(n183_adj_5192));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i124_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_9_2 (.CI(GND_net), .I0(\PID_CONTROLLER.integral [0]), .I1(n55[4]), 
            .CO(n51049));
    SB_LUT4 add_6352_15_lut (.I0(GND_net), .I1(n18415[12]), .I2(n1050), 
            .I3(n51377), .O(n17996[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6352_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6106_3 (.CI(n51610), .I0(n14082[0]), .I1(n153_adj_5172), 
            .CO(n51611));
    SB_LUT4 add_6106_2_lut (.I0(GND_net), .I1(n11_adj_5168), .I2(n80), 
            .I3(GND_net), .O(n13158[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6106_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6352_14_lut (.I0(GND_net), .I1(n18415[11]), .I2(n977), 
            .I3(n51376), .O(n17996[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6352_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i53631_3_lut (.I0(n4), .I1(n352[5]), .I2(n11_adj_5190), .I3(GND_net), 
            .O(n69325));   // verilog/motorControl.v(53[14:29])
    defparam i53631_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_16_i67_2_lut (.I0(\Kp[1] ), .I1(n55[12]), .I2(GND_net), 
            .I3(GND_net), .O(n98));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i67_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i20_2_lut (.I0(\Kp[0] ), .I1(n55[13]), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_5174));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i20_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6352_14 (.CI(n51376), .I0(n18415[11]), .I1(n977), .CO(n51377));
    SB_LUT4 add_6352_13_lut (.I0(GND_net), .I1(n18415[10]), .I2(n904), 
            .I3(n51375), .O(n17996[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6352_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_8_add_2_25_lut (.I0(GND_net), .I1(setpoint[23]), .I2(n16), 
            .I3(n51048), .O(n55[23])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_8_add_2_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6352_13 (.CI(n51375), .I0(n18415[10]), .I1(n904), .CO(n51376));
    SB_LUT4 mult_16_i173_2_lut (.I0(\Kp[3] ), .I1(n55[16]), .I2(GND_net), 
            .I3(GND_net), .O(n256));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i173_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i53632_3_lut (.I0(n69325), .I1(n352[6]), .I2(n13_adj_5188), 
            .I3(GND_net), .O(n69326));   // verilog/motorControl.v(53[14:29])
    defparam i53632_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_6352_12_lut (.I0(GND_net), .I1(n18415[9]), .I2(n831), 
            .I3(n51374), .O(n17996[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6352_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i53074_4_lut (.I0(n13_adj_5188), .I1(n11_adj_5190), .I2(n9_adj_5187), 
            .I3(n67907), .O(n68768));
    defparam i53074_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 LessThan_23_i8_3_lut (.I0(n6_adj_5195), .I1(n352[4]), .I2(n9_adj_5187), 
            .I3(GND_net), .O(n8_adj_5196));   // verilog/motorControl.v(53[14:29])
    defparam LessThan_23_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_26_inv_0_i20_1_lut (.I0(PWMLimit[19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5682[19]));   // verilog/motorControl.v(56[22:31])
    defparam unary_minus_26_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_16_i306_2_lut (.I0(\Kp[6] ), .I1(n55[9]), .I2(GND_net), 
            .I3(GND_net), .O(n454));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i306_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mult_16_add_1221_15 (.CI(n51692), .I0(n12096[12]), .I1(n1023), 
            .CO(n51693));
    SB_LUT4 mult_16_add_1221_14_lut (.I0(GND_net), .I1(n12096[11]), .I2(n950), 
            .I3(n51691), .O(n257[13])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_16_add_1221_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_8_add_2_24_lut (.I0(GND_net), .I1(setpoint[22]), .I2(n3), 
            .I3(n51047), .O(n55[22])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_8_add_2_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6106_2 (.CI(GND_net), .I0(n11_adj_5168), .I1(n80), .CO(n51610));
    SB_LUT4 i52595_3_lut (.I0(n69326), .I1(n352[7]), .I2(n15_adj_5186), 
            .I3(GND_net), .O(n68289));   // verilog/motorControl.v(53[14:29])
    defparam i52595_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53565_4_lut (.I0(n68289), .I1(n8_adj_5196), .I2(n15_adj_5186), 
            .I3(n68768), .O(n69259));   // verilog/motorControl.v(53[14:29])
    defparam i53565_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 mult_16_i222_2_lut (.I0(\Kp[4] ), .I1(n55[16]), .I2(GND_net), 
            .I3(GND_net), .O(n329));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i222_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i116_2_lut (.I0(\Kp[2] ), .I1(n55[12]), .I2(GND_net), 
            .I3(GND_net), .O(n171));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i116_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i53566_3_lut (.I0(n69259), .I1(n352[8]), .I2(PWMLimit[8]), 
            .I3(GND_net), .O(n18));   // verilog/motorControl.v(53[14:29])
    defparam i53566_3_lut.LUT_INIT = 16'h8e8e;
    SB_CARRY add_6352_12 (.CI(n51374), .I0(n18415[9]), .I1(n831), .CO(n51375));
    SB_LUT4 mult_16_i271_2_lut (.I0(\Kp[5] ), .I1(n55[16]), .I2(GND_net), 
            .I3(GND_net), .O(n402));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i271_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_23_i25_2_lut (.I0(PWMLimit[12]), .I1(n352[12]), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_5199));   // verilog/motorControl.v(53[14:29])
    defparam LessThan_23_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_23_i33_2_lut (.I0(PWMLimit[16]), .I1(n352[16]), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_5200));   // verilog/motorControl.v(53[14:29])
    defparam LessThan_23_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_16_i320_2_lut (.I0(\Kp[6] ), .I1(n55[16]), .I2(GND_net), 
            .I3(GND_net), .O(n475));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i320_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i447_2_lut (.I0(\Kp[9] ), .I1(n55[6]), .I2(GND_net), 
            .I3(GND_net), .O(n664));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i447_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mult_16_add_1221_14 (.CI(n51691), .I0(n12096[11]), .I1(n950), 
            .CO(n51692));
    SB_CARRY sub_8_add_2_24 (.CI(n51047), .I0(setpoint[22]), .I1(n3), 
            .CO(n51048));
    SB_LUT4 add_6352_11_lut (.I0(GND_net), .I1(n18415[8]), .I2(n758), 
            .I3(n51373), .O(n17996[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6352_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6352_11 (.CI(n51373), .I0(n18415[8]), .I1(n758), .CO(n51374));
    SB_LUT4 sub_8_add_2_23_lut (.I0(GND_net), .I1(setpoint[21]), .I2(\motor_state[21] ), 
            .I3(n51046), .O(n55[21])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_8_add_2_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6352_10_lut (.I0(GND_net), .I1(n18415[7]), .I2(n685), 
            .I3(n51372), .O(n17996[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6352_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i165_2_lut (.I0(\Kp[3] ), .I1(n55[12]), .I2(GND_net), 
            .I3(GND_net), .O(n244));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i165_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i355_2_lut (.I0(\Kp[7] ), .I1(n55[9]), .I2(GND_net), 
            .I3(GND_net), .O(n527));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i355_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i496_2_lut (.I0(\Kp[10] ), .I1(n55[6]), .I2(GND_net), 
            .I3(GND_net), .O(n737));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i496_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i369_2_lut (.I0(\Kp[7] ), .I1(n55[16]), .I2(GND_net), 
            .I3(GND_net), .O(n548));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i369_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6352_10 (.CI(n51372), .I0(n18415[7]), .I1(n685), .CO(n51373));
    SB_LUT4 mult_16_i214_2_lut (.I0(\Kp[4] ), .I1(n55[12]), .I2(GND_net), 
            .I3(GND_net), .O(n317));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i214_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 counter_1939_add_4_33_lut (.I0(GND_net), .I1(GND_net), .I2(counter[31]), 
            .I3(n52331), .O(n57[31])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1939_add_4_33_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 counter_1939_add_4_32_lut (.I0(GND_net), .I1(GND_net), .I2(counter[30]), 
            .I3(n52330), .O(n57[30])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1939_add_4_32_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i404_2_lut (.I0(\Kp[8] ), .I1(n55[9]), .I2(GND_net), 
            .I3(GND_net), .O(n600));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i404_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i545_2_lut (.I0(\Kp[11] ), .I1(n55[6]), .I2(GND_net), 
            .I3(GND_net), .O(n810));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i545_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY counter_1939_add_4_32 (.CI(n52330), .I0(GND_net), .I1(counter[30]), 
            .CO(n52331));
    SB_LUT4 add_6352_9_lut (.I0(GND_net), .I1(n18415[6]), .I2(n612), .I3(n51371), 
            .O(n17996[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6352_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6352_9 (.CI(n51371), .I0(n18415[6]), .I1(n612), .CO(n51372));
    SB_CARRY sub_8_add_2_23 (.CI(n51046), .I0(setpoint[21]), .I1(\motor_state[21] ), 
            .CO(n51047));
    SB_LUT4 mult_16_i453_2_lut (.I0(\Kp[9] ), .I1(n55[9]), .I2(GND_net), 
            .I3(GND_net), .O(n673));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i453_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i263_2_lut (.I0(\Kp[5] ), .I1(n55[12]), .I2(GND_net), 
            .I3(GND_net), .O(n390));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i263_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 counter_1939_add_4_31_lut (.I0(GND_net), .I1(GND_net), .I2(counter[29]), 
            .I3(n52329), .O(n57[29])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1939_add_4_31_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_8_add_2_22_lut (.I0(GND_net), .I1(setpoint[20]), .I2(\motor_state[20] ), 
            .I3(n51045), .O(n55[20])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_8_add_2_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_8_add_2_22 (.CI(n51045), .I0(setpoint[20]), .I1(\motor_state[20] ), 
            .CO(n51046));
    SB_CARRY counter_1939_add_4_31 (.CI(n52329), .I0(GND_net), .I1(counter[29]), 
            .CO(n52330));
    SB_LUT4 counter_1939_add_4_30_lut (.I0(GND_net), .I1(GND_net), .I2(counter[28]), 
            .I3(n52328), .O(n57[28])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1939_add_4_30_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i418_2_lut (.I0(\Kp[8] ), .I1(n55[16]), .I2(GND_net), 
            .I3(GND_net), .O(n621));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i418_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_26_inv_0_i21_1_lut (.I0(PWMLimit[20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5682[20]));   // verilog/motorControl.v(56[22:31])
    defparam unary_minus_26_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_6352_8_lut (.I0(GND_net), .I1(n18415[5]), .I2(n539), .I3(n51370), 
            .O(n17996[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6352_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_8_add_2_21_lut (.I0(GND_net), .I1(setpoint[19]), .I2(\motor_state[19] ), 
            .I3(n51044), .O(n55[19])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_8_add_2_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i467_2_lut (.I0(\Kp[9] ), .I1(n55[16]), .I2(GND_net), 
            .I3(GND_net), .O(n694));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i467_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY counter_1939_add_4_30 (.CI(n52328), .I0(GND_net), .I1(counter[28]), 
            .CO(n52329));
    SB_CARRY add_6352_8 (.CI(n51370), .I0(n18415[5]), .I1(n539), .CO(n51371));
    SB_LUT4 counter_1939_add_4_29_lut (.I0(GND_net), .I1(GND_net), .I2(counter[27]), 
            .I3(n52327), .O(n57[27])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1939_add_4_29_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i516_2_lut (.I0(\Kp[10] ), .I1(n55[16]), .I2(GND_net), 
            .I3(GND_net), .O(n767));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i516_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i565_2_lut (.I0(\Kp[11] ), .I1(n55[16]), .I2(GND_net), 
            .I3(GND_net), .O(n840));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i565_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY counter_1939_add_4_29 (.CI(n52327), .I0(GND_net), .I1(counter[27]), 
            .CO(n52328));
    SB_LUT4 mult_16_i85_2_lut (.I0(\Kp[1] ), .I1(n55[21]), .I2(GND_net), 
            .I3(GND_net), .O(n125_c));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i85_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i38_2_lut (.I0(\Kp[0] ), .I1(n55[22]), .I2(GND_net), 
            .I3(GND_net), .O(n56_c));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i38_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i312_2_lut (.I0(\Kp[6] ), .I1(n55[12]), .I2(GND_net), 
            .I3(GND_net), .O(n463));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i312_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i73_2_lut (.I0(\Kp[1] ), .I1(n55[15]), .I2(GND_net), 
            .I3(GND_net), .O(n107_adj_5173));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i73_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i26_2_lut (.I0(\Kp[0] ), .I1(n55[16]), .I2(GND_net), 
            .I3(GND_net), .O(n38_c));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i26_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i502_2_lut (.I0(\Kp[10] ), .I1(n55[9]), .I2(GND_net), 
            .I3(GND_net), .O(n746));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i502_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_26_inv_0_i22_1_lut (.I0(PWMLimit[21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5682[21]));   // verilog/motorControl.v(56[22:31])
    defparam unary_minus_26_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_26_inv_0_i23_1_lut (.I0(PWMLimit[22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5682[22]));   // verilog/motorControl.v(56[22:31])
    defparam unary_minus_26_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 counter_1939_add_4_28_lut (.I0(GND_net), .I1(GND_net), .I2(counter[26]), 
            .I3(n52326), .O(n57[26])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1939_add_4_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_1939_add_4_28 (.CI(n52326), .I0(GND_net), .I1(counter[26]), 
            .CO(n52327));
    SB_LUT4 mult_16_i361_2_lut (.I0(\Kp[7] ), .I1(n55[12]), .I2(GND_net), 
            .I3(GND_net), .O(n536));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i361_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i122_2_lut (.I0(\Kp[2] ), .I1(n55[15]), .I2(GND_net), 
            .I3(GND_net), .O(n180));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i122_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i551_2_lut (.I0(\Kp[11] ), .I1(n55[9]), .I2(GND_net), 
            .I3(GND_net), .O(n819));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i551_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_26_inv_0_i24_1_lut (.I0(PWMLimit[23]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5682[23]));   // verilog/motorControl.v(56[22:31])
    defparam unary_minus_26_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_16_i410_2_lut (.I0(\Kp[8] ), .I1(n55[12]), .I2(GND_net), 
            .I3(GND_net), .O(n609));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i410_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i600_2_lut (.I0(\Kp[12] ), .I1(n55[9]), .I2(GND_net), 
            .I3(GND_net), .O(n892));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i600_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i171_2_lut (.I0(\Kp[3] ), .I1(n55[15]), .I2(GND_net), 
            .I3(GND_net), .O(n253));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i171_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6352_7_lut (.I0(GND_net), .I1(n18415[4]), .I2(n466), .I3(n51369), 
            .O(n17996[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6352_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i594_2_lut (.I0(\Kp[12] ), .I1(n55[6]), .I2(GND_net), 
            .I3(GND_net), .O(n883));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i594_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6352_7 (.CI(n51369), .I0(n18415[4]), .I1(n466), .CO(n51370));
    SB_LUT4 mult_16_i459_2_lut (.I0(\Kp[9] ), .I1(n55[12]), .I2(GND_net), 
            .I3(GND_net), .O(n682));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i459_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i649_2_lut (.I0(\Kp[13] ), .I1(n55[9]), .I2(GND_net), 
            .I3(GND_net), .O(n965));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i649_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6352_6_lut (.I0(GND_net), .I1(n18415[3]), .I2(n393), .I3(n51368), 
            .O(n17996[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6352_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 counter_1939_add_4_27_lut (.I0(GND_net), .I1(GND_net), .I2(counter[25]), 
            .I3(n52325), .O(n57[25])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1939_add_4_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6352_6 (.CI(n51368), .I0(n18415[3]), .I1(n393), .CO(n51369));
    SB_CARRY counter_1939_add_4_27 (.CI(n52325), .I0(GND_net), .I1(counter[25]), 
            .CO(n52326));
    SB_LUT4 mult_16_i220_2_lut (.I0(\Kp[4] ), .I1(n55[15]), .I2(GND_net), 
            .I3(GND_net), .O(n326));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i220_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 counter_1939_add_4_26_lut (.I0(GND_net), .I1(GND_net), .I2(counter[24]), 
            .I3(n52324), .O(n57[24])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1939_add_4_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i269_2_lut (.I0(\Kp[5] ), .I1(n55[15]), .I2(GND_net), 
            .I3(GND_net), .O(n399));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i269_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i698_2_lut (.I0(\Kp[14] ), .I1(n55[9]), .I2(GND_net), 
            .I3(GND_net), .O(n1038));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i698_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i508_2_lut (.I0(\Kp[10] ), .I1(n55[12]), .I2(GND_net), 
            .I3(GND_net), .O(n755));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i508_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i643_2_lut (.I0(\Kp[13] ), .I1(n55[6]), .I2(GND_net), 
            .I3(GND_net), .O(n956));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i643_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i747_2_lut (.I0(\Kp[15] ), .I1(n55[9]), .I2(GND_net), 
            .I3(GND_net), .O(n1111));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i747_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i318_2_lut (.I0(\Kp[6] ), .I1(n55[15]), .I2(GND_net), 
            .I3(GND_net), .O(n472));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i318_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i557_2_lut (.I0(\Kp[11] ), .I1(n55[12]), .I2(GND_net), 
            .I3(GND_net), .O(n828));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i557_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i692_2_lut (.I0(\Kp[14] ), .I1(n55[6]), .I2(GND_net), 
            .I3(GND_net), .O(n1029));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i692_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i367_2_lut (.I0(\Kp[7] ), .I1(n55[15]), .I2(GND_net), 
            .I3(GND_net), .O(n545));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i367_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i134_2_lut (.I0(\Kp[2] ), .I1(n55[21]), .I2(GND_net), 
            .I3(GND_net), .O(n198_adj_5171));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i134_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i606_2_lut (.I0(\Kp[12] ), .I1(n55[12]), .I2(GND_net), 
            .I3(GND_net), .O(n901));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i606_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i416_2_lut (.I0(\Kp[8] ), .I1(n55[15]), .I2(GND_net), 
            .I3(GND_net), .O(n618));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i416_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i183_2_lut (.I0(\Kp[3] ), .I1(n55[21]), .I2(GND_net), 
            .I3(GND_net), .O(n271_c));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i183_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6352_5_lut (.I0(GND_net), .I1(n18415[2]), .I2(n320), .I3(n51367), 
            .O(n17996[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6352_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut (.I0(n55[23]), .I1(\Kp[2] ), .I2(n50735), .I3(n55[22]), 
            .O(n63605));   // verilog/motorControl.v(51[18:24])
    defparam i1_4_lut.LUT_INIT = 16'h6ca0;
    SB_LUT4 mult_16_add_1221_13_lut (.I0(GND_net), .I1(n12096[10]), .I2(n877_adj_5211), 
            .I3(n51690), .O(n257[12])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_16_add_1221_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_1939_add_4_26 (.CI(n52324), .I0(GND_net), .I1(counter[24]), 
            .CO(n52325));
    SB_LUT4 counter_1939_add_4_25_lut (.I0(GND_net), .I1(GND_net), .I2(counter[23]), 
            .I3(n52323), .O(n57[23])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1939_add_4_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i465_2_lut (.I0(\Kp[9] ), .I1(n55[15]), .I2(GND_net), 
            .I3(GND_net), .O(n691));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i465_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i277_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3715[15] ), 
            .I2(GND_net), .I3(GND_net), .O(n411));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i277_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i655_2_lut (.I0(\Kp[13] ), .I1(n55[12]), .I2(GND_net), 
            .I3(GND_net), .O(n974));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i655_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i741_2_lut (.I0(\Kp[15] ), .I1(n55[6]), .I2(GND_net), 
            .I3(GND_net), .O(n1102));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i741_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY counter_1939_add_4_25 (.CI(n52323), .I0(GND_net), .I1(counter[23]), 
            .CO(n52324));
    SB_LUT4 mult_16_i514_2_lut (.I0(\Kp[10] ), .I1(n55[15]), .I2(GND_net), 
            .I3(GND_net), .O(n764));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i514_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i563_2_lut (.I0(\Kp[11] ), .I1(n55[15]), .I2(GND_net), 
            .I3(GND_net), .O(n837));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i563_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i232_2_lut (.I0(\Kp[4] ), .I1(n55[21]), .I2(GND_net), 
            .I3(GND_net), .O(n344_adj_5170));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i232_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 counter_1939_add_4_24_lut (.I0(GND_net), .I1(GND_net), .I2(counter[22]), 
            .I3(n52322), .O(n57[22])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1939_add_4_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1717 (.I0(n55[22]), .I1(n20185[1]), .I2(n4_adj_5214), 
            .I3(\Kp[3] ), .O(n20087[2]));   // verilog/motorControl.v(51[18:24])
    defparam i1_4_lut_adj_1717.LUT_INIT = 16'hc66c;
    SB_LUT4 mult_16_i704_2_lut (.I0(\Kp[14] ), .I1(n55[12]), .I2(GND_net), 
            .I3(GND_net), .O(n1047));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i704_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i612_2_lut (.I0(\Kp[12] ), .I1(n55[15]), .I2(GND_net), 
            .I3(GND_net), .O(n910));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i612_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i247_2_lut (.I0(\Kp[5] ), .I1(n55[4]), .I2(GND_net), 
            .I3(GND_net), .O(n366_adj_5215));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i247_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i753_2_lut (.I0(\Kp[15] ), .I1(n55[12]), .I2(GND_net), 
            .I3(GND_net), .O(n1120));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i753_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY sub_8_add_2_21 (.CI(n51044), .I0(setpoint[19]), .I1(\motor_state[19] ), 
            .CO(n51045));
    SB_LUT4 mult_16_i281_2_lut (.I0(\Kp[5] ), .I1(n55[21]), .I2(GND_net), 
            .I3(GND_net), .O(n417_c));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i281_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i234_2_lut (.I0(\Kp[4] ), .I1(n55[22]), .I2(GND_net), 
            .I3(GND_net), .O(n347_adj_5216));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i234_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut_adj_1718 (.I0(n20185[1]), .I1(n6_adj_5217), .I2(n347_adj_5216), 
            .I3(n59071), .O(n20087[3]));   // verilog/motorControl.v(51[18:24])
    defparam i1_4_lut_adj_1718.LUT_INIT = 16'h6996;
    SB_LUT4 sub_8_add_2_20_lut (.I0(GND_net), .I1(setpoint[18]), .I2(\motor_state[18] ), 
            .I3(n51043), .O(n55[18])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_8_add_2_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6352_5 (.CI(n51367), .I0(n18415[2]), .I1(n320), .CO(n51368));
    SB_LUT4 add_6352_4_lut (.I0(GND_net), .I1(n18415[1]), .I2(n247), .I3(n51366), 
            .O(n17996[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6352_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_3_lut (.I0(\Kp[0] ), .I1(\Kp[2] ), .I2(\Kp[1] ), .I3(GND_net), 
            .O(n63601));   // verilog/motorControl.v(51[18:24])
    defparam i1_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i1_2_lut_adj_1719 (.I0(n63601), .I1(n55[23]), .I2(GND_net), 
            .I3(GND_net), .O(n4_adj_5214));   // verilog/motorControl.v(51[18:24])
    defparam i1_2_lut_adj_1719.LUT_INIT = 16'h8888;
    SB_LUT4 i36937_4_lut (.I0(n20185[1]), .I1(\Kp[3] ), .I2(n4_adj_5214), 
            .I3(n55[22]), .O(n6_adj_5217));   // verilog/motorControl.v(51[18:24])
    defparam i36937_4_lut.LUT_INIT = 16'he800;
    SB_LUT4 mult_16_i40_2_lut (.I0(\Kp[0] ), .I1(n55[23]), .I2(GND_net), 
            .I3(GND_net), .O(n62));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i40_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i36876_2_lut (.I0(\Kp[0] ), .I1(\Kp[1] ), .I2(GND_net), .I3(GND_net), 
            .O(n50735));   // verilog/motorControl.v(51[18:24])
    defparam i36876_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_3_lut_3_lut (.I0(n376), .I1(PWMLimit[0]), .I2(PWMLimit[1]), 
            .I3(GND_net), .O(n28));   // verilog/motorControl.v(51[18:38])
    defparam i1_3_lut_3_lut.LUT_INIT = 16'hd0d0;
    SB_LUT4 i48297_3_lut (.I0(n55[23]), .I1(n63601), .I2(\Kp[3] ), .I3(GND_net), 
            .O(n59071));   // verilog/motorControl.v(51[18:24])
    defparam i48297_3_lut.LUT_INIT = 16'h2828;
    SB_LUT4 i37068_3_lut (.I0(n55[23]), .I1(n50749), .I2(n61580), .I3(GND_net), 
            .O(n20185[1]));   // verilog/motorControl.v(51[18:24])
    defparam i37068_3_lut.LUT_INIT = 16'h6c6c;
    SB_LUT4 mult_16_i330_2_lut (.I0(\Kp[6] ), .I1(n55[21]), .I2(GND_net), 
            .I3(GND_net), .O(n490_c));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i330_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut_adj_1720 (.I0(n55[23]), .I1(\Kp[5] ), .I2(n61580), 
            .I3(n55[22]), .O(n63591));   // verilog/motorControl.v(51[18:24])
    defparam i1_4_lut_adj_1720.LUT_INIT = 16'hc60a;
    SB_LUT4 i1_rep_257_2_lut (.I0(n20185[1]), .I1(n59071), .I2(GND_net), 
            .I3(GND_net), .O(n71499));   // verilog/motorControl.v(51[18:24])
    defparam i1_rep_257_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1721 (.I0(n50749), .I1(n63591), .I2(\Kp[4] ), 
            .I3(n55[23]), .O(n63595));   // verilog/motorControl.v(51[18:24])
    defparam i1_4_lut_adj_1721.LUT_INIT = 16'h9666;
    SB_LUT4 i36945_4_lut (.I0(n71499), .I1(\Kp[4] ), .I2(n6_adj_5217), 
            .I3(n55[22]), .O(n8_adj_5219));   // verilog/motorControl.v(51[18:24])
    defparam i36945_4_lut.LUT_INIT = 16'he8a0;
    SB_LUT4 i36898_4_lut (.I0(n20185[1]), .I1(\Kp[3] ), .I2(n63601), .I3(n55[23]), 
            .O(n6_adj_5220));   // verilog/motorControl.v(51[18:24])
    defparam i36898_4_lut.LUT_INIT = 16'he800;
    SB_LUT4 i1_4_lut_adj_1722 (.I0(n6_adj_5220), .I1(n8_adj_5219), .I2(n63595), 
            .I3(n59071), .O(n61804));   // verilog/motorControl.v(51[18:24])
    defparam i1_4_lut_adj_1722.LUT_INIT = 16'h6996;
    SB_LUT4 mult_17_i28_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3715[13] ), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_5221));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i28_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i124_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3715[12] ), 
            .I2(GND_net), .I3(GND_net), .O(n183_adj_5222));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i124_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i173_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3715[12] ), 
            .I2(GND_net), .I3(GND_net), .O(n256_adj_5223));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i173_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_14_i18_3_lut (.I0(n130[17]), .I1(n182[17]), .I2(n181), 
            .I3(GND_net), .O(n214));   // verilog/motorControl.v(48[18] 50[12])
    defparam mux_14_i18_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_17_i83_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3715[16] ), 
            .I2(GND_net), .I3(GND_net), .O(n122_adj_5169));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i83_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i222_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3715[12] ), 
            .I2(GND_net), .I3(GND_net), .O(n329_adj_5225));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i222_2_lut.LUT_INIT = 16'h8888;
    SB_DFFR \PID_CONTROLLER.integral_i0_i0  (.Q(\PID_CONTROLLER.integral [0]), 
            .C(clk16MHz), .D(n29560), .R(reset));   // verilog/motorControl.v(41[14] 62[8])
    SB_LUT4 mult_17_i271_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3715[12] ), 
            .I2(GND_net), .I3(GND_net), .O(n402_adj_5226));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i271_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i320_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3715[12] ), 
            .I2(GND_net), .I3(GND_net), .O(n475_adj_5227));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i320_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i369_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3715[12] ), 
            .I2(GND_net), .I3(GND_net), .O(n548_adj_5228));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i369_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i261_2_lut (.I0(\Kp[5] ), .I1(n55[11]), .I2(GND_net), 
            .I3(GND_net), .O(n387));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i261_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i418_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3715[12] ), 
            .I2(GND_net), .I3(GND_net), .O(n621_adj_5229));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i418_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i467_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3715[12] ), 
            .I2(GND_net), .I3(GND_net), .O(n694_adj_5230));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i467_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY sub_8_add_2_20 (.CI(n51043), .I0(setpoint[18]), .I1(\motor_state[18] ), 
            .CO(n51044));
    SB_CARRY counter_1939_add_4_24 (.CI(n52322), .I0(GND_net), .I1(counter[22]), 
            .CO(n52323));
    SB_LUT4 mult_17_i516_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3715[12] ), 
            .I2(GND_net), .I3(GND_net), .O(n767_adj_5231));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i516_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 counter_1939_add_4_23_lut (.I0(GND_net), .I1(GND_net), .I2(counter[21]), 
            .I3(n52321), .O(n57[21])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1939_add_4_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_i565_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3715[12] ), 
            .I2(GND_net), .I3(GND_net), .O(n840_adj_5233));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i565_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY counter_1939_add_4_23 (.CI(n52321), .I0(GND_net), .I1(counter[21]), 
            .CO(n52322));
    SB_LUT4 mult_17_i73_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3715[11] ), 
            .I2(GND_net), .I3(GND_net), .O(n107_adj_5234));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i73_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i122_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3715[11] ), 
            .I2(GND_net), .I3(GND_net), .O(n180_adj_5235));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i122_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i171_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3715[11] ), 
            .I2(GND_net), .I3(GND_net), .O(n253_adj_5236));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i171_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i220_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3715[11] ), 
            .I2(GND_net), .I3(GND_net), .O(n326_adj_5237));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i220_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i269_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3715[11] ), 
            .I2(GND_net), .I3(GND_net), .O(n399_adj_5238));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i269_2_lut.LUT_INIT = 16'h8888;
    SB_DFFSR counter_1939__i0 (.Q(counter[0]), .C(clk16MHz), .D(n57[0]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(24[16:25])
    SB_LUT4 mult_17_i318_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3715[11] ), 
            .I2(GND_net), .I3(GND_net), .O(n472_adj_5239));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i318_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i367_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3715[11] ), 
            .I2(GND_net), .I3(GND_net), .O(n545_adj_5240));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i367_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i416_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3715[11] ), 
            .I2(GND_net), .I3(GND_net), .O(n618_adj_5241));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i416_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i465_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3715[11] ), 
            .I2(GND_net), .I3(GND_net), .O(n691_adj_5242));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i465_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i514_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3715[11] ), 
            .I2(GND_net), .I3(GND_net), .O(n764_adj_5243));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i514_2_lut.LUT_INIT = 16'h8888;
    SB_DFFSR counter_1939__i31 (.Q(counter[31]), .C(clk16MHz), .D(n57[31]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_1939__i30 (.Q(counter[30]), .C(clk16MHz), .D(n57[30]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_1939__i29 (.Q(counter[29]), .C(clk16MHz), .D(n57[29]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_1939__i28 (.Q(counter[28]), .C(clk16MHz), .D(n57[28]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_1939__i27 (.Q(counter[27]), .C(clk16MHz), .D(n57[27]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_1939__i26 (.Q(counter[26]), .C(clk16MHz), .D(n57[26]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_1939__i25 (.Q(counter[25]), .C(clk16MHz), .D(n57[25]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_1939__i24 (.Q(counter[24]), .C(clk16MHz), .D(n57[24]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_1939__i23 (.Q(counter[23]), .C(clk16MHz), .D(n57[23]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_1939__i22 (.Q(counter[22]), .C(clk16MHz), .D(n57[22]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_1939__i21 (.Q(counter[21]), .C(clk16MHz), .D(n57[21]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_1939__i20 (.Q(counter[20]), .C(clk16MHz), .D(n57[20]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_1939__i19 (.Q(counter[19]), .C(clk16MHz), .D(n57[19]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_1939__i18 (.Q(counter[18]), .C(clk16MHz), .D(n57[18]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_1939__i17 (.Q(counter[17]), .C(clk16MHz), .D(n57[17]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_1939__i16 (.Q(counter[16]), .C(clk16MHz), .D(n57[16]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_1939__i15 (.Q(counter[15]), .C(clk16MHz), .D(n57[15]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_1939__i14 (.Q(counter[14]), .C(clk16MHz), .D(n57[14]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_1939__i13 (.Q(counter[13]), .C(clk16MHz), .D(n57[13]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_1939__i12 (.Q(counter[12]), .C(clk16MHz), .D(n57[12]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_1939__i11 (.Q(counter[11]), .C(clk16MHz), .D(n57[11]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_1939__i10 (.Q(counter[10]), .C(clk16MHz), .D(n57[10]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_1939__i9 (.Q(counter[9]), .C(clk16MHz), .D(n57[9]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_1939__i8 (.Q(counter[8]), .C(clk16MHz), .D(n57[8]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_1939__i7 (.Q(counter[7]), .C(clk16MHz), .D(n57[7]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_1939__i6 (.Q(counter[6]), .C(clk16MHz), .D(n57[6]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_1939__i5 (.Q(counter[5]), .C(clk16MHz), .D(n57[5]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_1939__i4 (.Q(counter[4]), .C(clk16MHz), .D(n57[4]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_1939__i3 (.Q(counter[3]), .C(clk16MHz), .D(n57[3]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_1939__i2 (.Q(counter[2]), .C(clk16MHz), .D(n57[2]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_1939__i1 (.Q(counter[1]), .C(clk16MHz), .D(n57[1]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(24[16:25])
    SB_DFFER result__i23 (.Q(duty[23]), .C(clk16MHz), .E(control_update), 
            .D(n51[23]), .R(reset));   // verilog/motorControl.v(41[14] 62[8])
    SB_LUT4 mult_17_i563_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3715[11] ), 
            .I2(GND_net), .I3(GND_net), .O(n837_adj_5258));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i563_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i132_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3715[16] ), 
            .I2(GND_net), .I3(GND_net), .O(n195_adj_5167));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i132_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i52369_2_lut_4_lut (.I0(n130[16]), .I1(n182[16]), .I2(n130[7]), 
            .I3(n182[7]), .O(n68063));
    defparam i52369_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 mult_17_i612_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3715[11] ), 
            .I2(GND_net), .I3(GND_net), .O(n910_adj_5259));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i612_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i53_2_lut (.I0(\Kp[1] ), .I1(n55[5]), .I2(GND_net), 
            .I3(GND_net), .O(n77));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i53_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i6_2_lut (.I0(\Kp[0] ), .I1(n55[6]), .I2(GND_net), 
            .I3(GND_net), .O(n8_adj_5166));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i6_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i83_2_lut (.I0(\Kp[1] ), .I1(n55[20]), .I2(GND_net), 
            .I3(GND_net), .O(n122_adj_5260));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i83_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 counter_1939_add_4_22_lut (.I0(GND_net), .I1(GND_net), .I2(counter[20]), 
            .I3(n52320), .O(n57[20])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1939_add_4_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_1939_add_4_22 (.CI(n52320), .I0(GND_net), .I1(counter[20]), 
            .CO(n52321));
    SB_LUT4 counter_1939_add_4_21_lut (.I0(GND_net), .I1(GND_net), .I2(counter[19]), 
            .I3(n52319), .O(n57[19])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1939_add_4_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i36_2_lut (.I0(\Kp[0] ), .I1(n55[21]), .I2(GND_net), 
            .I3(GND_net), .O(n53_adj_5261));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i36_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i132_2_lut (.I0(\Kp[2] ), .I1(n55[20]), .I2(GND_net), 
            .I3(GND_net), .O(n195_adj_5262));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i132_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 sub_8_add_2_19_lut (.I0(GND_net), .I1(setpoint[17]), .I2(\motor_state[17] ), 
            .I3(n51042), .O(n55[17])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_8_add_2_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_1939_add_4_21 (.CI(n52319), .I0(GND_net), .I1(counter[19]), 
            .CO(n52320));
    SB_LUT4 counter_1939_add_4_20_lut (.I0(GND_net), .I1(GND_net), .I2(counter[18]), 
            .I3(n52318), .O(n57[18])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1939_add_4_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i181_2_lut (.I0(\Kp[3] ), .I1(n55[20]), .I2(GND_net), 
            .I3(GND_net), .O(n268_adj_5263));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i181_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i102_2_lut (.I0(\Kp[2] ), .I1(n55[5]), .I2(GND_net), 
            .I3(GND_net), .O(n150));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i102_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY counter_1939_add_4_20 (.CI(n52318), .I0(GND_net), .I1(counter[18]), 
            .CO(n52319));
    SB_LUT4 counter_1939_add_4_19_lut (.I0(GND_net), .I1(GND_net), .I2(counter[17]), 
            .I3(n52317), .O(n57[17])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1939_add_4_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_1939_add_4_19 (.CI(n52317), .I0(GND_net), .I1(counter[17]), 
            .CO(n52318));
    SB_LUT4 mux_14_i1_3_lut (.I0(n130[0]), .I1(n182[0]), .I2(n181), .I3(GND_net), 
            .O(n207[0]));   // verilog/motorControl.v(48[18] 50[12])
    defparam mux_14_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_15_i1_3_lut (.I0(n207[0]), .I1(IntegralLimit[0]), .I2(n155), 
            .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3715[0] ));   // verilog/motorControl.v(48[18] 50[12])
    defparam mux_15_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_16_i230_2_lut (.I0(\Kp[4] ), .I1(n55[20]), .I2(GND_net), 
            .I3(GND_net), .O(n341_adj_5264));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i230_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i2_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3715[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n49[0]));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i2_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i2_2_lut (.I0(\Kp[0] ), .I1(n55[4]), .I2(GND_net), 
            .I3(GND_net), .O(n257[0]));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i2_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i279_2_lut (.I0(\Kp[5] ), .I1(n55[20]), .I2(GND_net), 
            .I3(GND_net), .O(n414_adj_5265));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i279_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i328_2_lut (.I0(\Kp[6] ), .I1(n55[20]), .I2(GND_net), 
            .I3(GND_net), .O(n487_adj_5266));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i328_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i377_2_lut (.I0(\Kp[7] ), .I1(n55[20]), .I2(GND_net), 
            .I3(GND_net), .O(n560_adj_5267));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i377_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i181_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3715[16] ), 
            .I2(GND_net), .I3(GND_net), .O(n268));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i181_2_lut.LUT_INIT = 16'h8888;
    SB_DFFER result__i22 (.Q(duty[22]), .C(clk16MHz), .E(control_update), 
            .D(n51[22]), .R(reset));   // verilog/motorControl.v(41[14] 62[8])
    SB_LUT4 mult_17_i71_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3715[10] ), 
            .I2(GND_net), .I3(GND_net), .O(n104));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i71_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i51508_2_lut_4_lut (.I0(IntegralLimit[21]), .I1(n130[21]), .I2(IntegralLimit[9]), 
            .I3(n130[9]), .O(n67202));
    defparam i51508_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 mult_17_i230_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3715[16] ), 
            .I2(GND_net), .I3(GND_net), .O(n341_adj_5165));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i230_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i151_2_lut (.I0(\Kp[3] ), .I1(n55[5]), .I2(GND_net), 
            .I3(GND_net), .O(n223));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i151_2_lut.LUT_INIT = 16'h8888;
    SB_DFFER result__i21 (.Q(duty[21]), .C(clk16MHz), .E(control_update), 
            .D(n51[21]), .R(reset));   // verilog/motorControl.v(41[14] 62[8])
    SB_DFFER result__i20 (.Q(duty[20]), .C(clk16MHz), .E(control_update), 
            .D(n51[20]), .R(reset));   // verilog/motorControl.v(41[14] 62[8])
    SB_DFFER result__i19 (.Q(duty[19]), .C(clk16MHz), .E(control_update), 
            .D(n51[19]), .R(reset));   // verilog/motorControl.v(41[14] 62[8])
    SB_CARRY add_6352_4 (.CI(n51366), .I0(n18415[1]), .I1(n247), .CO(n51367));
    SB_LUT4 mult_17_i279_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3715[16] ), 
            .I2(GND_net), .I3(GND_net), .O(n414));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i279_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 counter_1939_add_4_18_lut (.I0(GND_net), .I1(GND_net), .I2(counter[16]), 
            .I3(n52316), .O(n57[16])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1939_add_4_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_16_add_1221_13 (.CI(n51690), .I0(n12096[10]), .I1(n877_adj_5211), 
            .CO(n51691));
    SB_LUT4 mult_17_i24_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3715[11] ), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_5270));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i24_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY counter_1939_add_4_18 (.CI(n52316), .I0(GND_net), .I1(counter[16]), 
            .CO(n52317));
    SB_LUT4 mult_17_i120_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3715[10] ), 
            .I2(GND_net), .I3(GND_net), .O(n177));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i120_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i51729_2_lut_4_lut (.I0(IntegralLimit[16]), .I1(n130[16]), .I2(IntegralLimit[7]), 
            .I3(n130[7]), .O(n67423));
    defparam i51729_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_DFFER result__i18 (.Q(duty[18]), .C(clk16MHz), .E(control_update), 
            .D(n51[18]), .R(reset));   // verilog/motorControl.v(41[14] 62[8])
    SB_DFFER result__i17 (.Q(duty[17]), .C(clk16MHz), .E(control_update), 
            .D(n51[17]), .R(reset));   // verilog/motorControl.v(41[14] 62[8])
    SB_DFFER result__i16 (.Q(duty[16]), .C(clk16MHz), .E(control_update), 
            .D(n51[16]), .R(reset));   // verilog/motorControl.v(41[14] 62[8])
    SB_LUT4 mult_17_i169_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3715[10] ), 
            .I2(GND_net), .I3(GND_net), .O(n250));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i169_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i218_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3715[10] ), 
            .I2(GND_net), .I3(GND_net), .O(n323));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i218_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i267_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3715[10] ), 
            .I2(GND_net), .I3(GND_net), .O(n396));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i267_2_lut.LUT_INIT = 16'h8888;
    SB_DFFER result__i15 (.Q(duty[15]), .C(clk16MHz), .E(control_update), 
            .D(n51[15]), .R(reset));   // verilog/motorControl.v(41[14] 62[8])
    SB_DFFER result__i14 (.Q(duty[14]), .C(clk16MHz), .E(control_update), 
            .D(n51[14]), .R(reset));   // verilog/motorControl.v(41[14] 62[8])
    SB_LUT4 mult_16_i310_2_lut (.I0(\Kp[6] ), .I1(n55[11]), .I2(GND_net), 
            .I3(GND_net), .O(n460));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i310_2_lut.LUT_INIT = 16'h8888;
    SB_DFFER result__i13 (.Q(duty[13]), .C(clk16MHz), .E(control_update), 
            .D(n51[13]), .R(reset));   // verilog/motorControl.v(41[14] 62[8])
    SB_DFFER result__i12 (.Q(duty[12]), .C(clk16MHz), .E(control_update), 
            .D(n51[12]), .R(reset));   // verilog/motorControl.v(41[14] 62[8])
    SB_DFFER result__i11 (.Q(duty[11]), .C(clk16MHz), .E(control_update), 
            .D(n51[11]), .R(reset));   // verilog/motorControl.v(41[14] 62[8])
    SB_DFFER result__i10 (.Q(duty[10]), .C(clk16MHz), .E(control_update), 
            .D(n51[10]), .R(reset));   // verilog/motorControl.v(41[14] 62[8])
    SB_DFFER result__i9 (.Q(duty[9]), .C(clk16MHz), .E(control_update), 
            .D(n51[9]), .R(reset));   // verilog/motorControl.v(41[14] 62[8])
    SB_DFFER result__i8 (.Q(duty[8]), .C(clk16MHz), .E(control_update), 
            .D(n51[8]), .R(reset));   // verilog/motorControl.v(41[14] 62[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i1  (.Q(\PID_CONTROLLER.integral [1]), 
            .C(clk16MHz), .D(n30387), .R(reset));   // verilog/motorControl.v(41[14] 62[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i2  (.Q(\PID_CONTROLLER.integral [2]), 
            .C(clk16MHz), .D(n30386), .R(reset));   // verilog/motorControl.v(41[14] 62[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i3  (.Q(\PID_CONTROLLER.integral [3]), 
            .C(clk16MHz), .D(n30385), .R(reset));   // verilog/motorControl.v(41[14] 62[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i4  (.Q(\PID_CONTROLLER.integral [4]), 
            .C(clk16MHz), .D(n30384), .R(reset));   // verilog/motorControl.v(41[14] 62[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i5  (.Q(\PID_CONTROLLER.integral [5]), 
            .C(clk16MHz), .D(n30383), .R(reset));   // verilog/motorControl.v(41[14] 62[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i6  (.Q(\PID_CONTROLLER.integral [6]), 
            .C(clk16MHz), .D(n30382), .R(reset));   // verilog/motorControl.v(41[14] 62[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i7  (.Q(\PID_CONTROLLER.integral [7]), 
            .C(clk16MHz), .D(n30381), .R(reset));   // verilog/motorControl.v(41[14] 62[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i8  (.Q(\PID_CONTROLLER.integral [8]), 
            .C(clk16MHz), .D(n30380), .R(reset));   // verilog/motorControl.v(41[14] 62[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i9  (.Q(\PID_CONTROLLER.integral [9]), 
            .C(clk16MHz), .D(n30379), .R(reset));   // verilog/motorControl.v(41[14] 62[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i10  (.Q(\PID_CONTROLLER.integral [10]), 
            .C(clk16MHz), .D(n30378), .R(reset));   // verilog/motorControl.v(41[14] 62[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i11  (.Q(\PID_CONTROLLER.integral [11]), 
            .C(clk16MHz), .D(n30377), .R(reset));   // verilog/motorControl.v(41[14] 62[8])
    SB_LUT4 mult_16_add_1221_12_lut (.I0(GND_net), .I1(n12096[9]), .I2(n804_adj_5273), 
            .I3(n51689), .O(n257[11])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_16_add_1221_12_lut.LUT_INIT = 16'hC33C;
    SB_DFFR \PID_CONTROLLER.integral_i0_i12  (.Q(\PID_CONTROLLER.integral [12]), 
            .C(clk16MHz), .D(n30376), .R(reset));   // verilog/motorControl.v(41[14] 62[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i13  (.Q(\PID_CONTROLLER.integral [13]), 
            .C(clk16MHz), .D(n30374), .R(reset));   // verilog/motorControl.v(41[14] 62[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i14  (.Q(\PID_CONTROLLER.integral [14]), 
            .C(clk16MHz), .D(n30372), .R(reset));   // verilog/motorControl.v(41[14] 62[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i15  (.Q(\PID_CONTROLLER.integral [15]), 
            .C(clk16MHz), .D(n30371), .R(reset));   // verilog/motorControl.v(41[14] 62[8])
    SB_CARRY mult_16_add_1221_12 (.CI(n51689), .I0(n12096[9]), .I1(n804_adj_5273), 
            .CO(n51690));
    SB_DFFR \PID_CONTROLLER.integral_i0_i16  (.Q(\PID_CONTROLLER.integral [16]), 
            .C(clk16MHz), .D(n30370), .R(reset));   // verilog/motorControl.v(41[14] 62[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i17  (.Q(\PID_CONTROLLER.integral [17]), 
            .C(clk16MHz), .D(n30369), .R(reset));   // verilog/motorControl.v(41[14] 62[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i18  (.Q(\PID_CONTROLLER.integral [18]), 
            .C(clk16MHz), .D(n30368), .R(reset));   // verilog/motorControl.v(41[14] 62[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i19  (.Q(\PID_CONTROLLER.integral [19]), 
            .C(clk16MHz), .D(n30367), .R(reset));   // verilog/motorControl.v(41[14] 62[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i20  (.Q(\PID_CONTROLLER.integral [20]), 
            .C(clk16MHz), .D(n30366), .R(reset));   // verilog/motorControl.v(41[14] 62[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i21  (.Q(\PID_CONTROLLER.integral [21]), 
            .C(clk16MHz), .D(n30365), .R(reset));   // verilog/motorControl.v(41[14] 62[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i22  (.Q(\PID_CONTROLLER.integral [22]), 
            .C(clk16MHz), .D(n30364), .R(reset));   // verilog/motorControl.v(41[14] 62[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i23  (.Q(\PID_CONTROLLER.integral [23]), 
            .C(clk16MHz), .D(n30363), .R(reset));   // verilog/motorControl.v(41[14] 62[8])
    SB_DFFER result__i7 (.Q(duty[7]), .C(clk16MHz), .E(control_update), 
            .D(n51[7]), .R(reset));   // verilog/motorControl.v(41[14] 62[8])
    SB_DFFER result__i6 (.Q(duty[6]), .C(clk16MHz), .E(control_update), 
            .D(n51[6]), .R(reset));   // verilog/motorControl.v(41[14] 62[8])
    SB_DFFER result__i5 (.Q(duty[5]), .C(clk16MHz), .E(control_update), 
            .D(n51[5]), .R(reset));   // verilog/motorControl.v(41[14] 62[8])
    SB_DFFER result__i4 (.Q(duty[4]), .C(clk16MHz), .E(control_update), 
            .D(n51[4]), .R(reset));   // verilog/motorControl.v(41[14] 62[8])
    SB_DFFER result__i3 (.Q(duty[3]), .C(clk16MHz), .E(control_update), 
            .D(n51[3]), .R(reset));   // verilog/motorControl.v(41[14] 62[8])
    SB_DFFER result__i2 (.Q(duty[2]), .C(clk16MHz), .E(control_update), 
            .D(n51[2]), .R(reset));   // verilog/motorControl.v(41[14] 62[8])
    SB_LUT4 add_6352_3_lut (.I0(GND_net), .I1(n18415[0]), .I2(n174), .I3(n51365), 
            .O(n17996[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6352_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_add_1221_11_lut (.I0(GND_net), .I1(n12096[8]), .I2(n731), 
            .I3(n51688), .O(n257[10])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_16_add_1221_11_lut.LUT_INIT = 16'hC33C;
    SB_DFFER result__i1 (.Q(duty[1]), .C(clk16MHz), .E(control_update), 
            .D(n51[1]), .R(reset));   // verilog/motorControl.v(41[14] 62[8])
    SB_CARRY mult_16_add_1221_11 (.CI(n51688), .I0(n12096[8]), .I1(n731), 
            .CO(n51689));
    SB_LUT4 mult_16_add_1221_10_lut (.I0(GND_net), .I1(n12096[7]), .I2(n658), 
            .I3(n51687), .O(n257[9])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_16_add_1221_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6352_3 (.CI(n51365), .I0(n18415[0]), .I1(n174), .CO(n51366));
    SB_LUT4 mult_16_i200_2_lut (.I0(\Kp[4] ), .I1(n55[5]), .I2(GND_net), 
            .I3(GND_net), .O(n296_adj_5164));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i200_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i316_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3715[10] ), 
            .I2(GND_net), .I3(GND_net), .O(n469));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i316_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i328_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3715[16] ), 
            .I2(GND_net), .I3(GND_net), .O(n487));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i328_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 counter_1939_add_4_17_lut (.I0(GND_net), .I1(GND_net), .I2(counter[15]), 
            .I3(n52315), .O(n57[15])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1939_add_4_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6352_2_lut (.I0(GND_net), .I1(n32_adj_5275), .I2(n101), 
            .I3(GND_net), .O(n17996[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6352_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6352_2 (.CI(GND_net), .I0(n32_adj_5275), .I1(n101), .CO(n51365));
    SB_LUT4 mult_17_i365_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3715[10] ), 
            .I2(GND_net), .I3(GND_net), .O(n542));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i365_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_13_inv_0_i1_1_lut (.I0(IntegralLimit[0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[0]));   // verilog/motorControl.v(49[22:36])
    defparam unary_minus_13_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY counter_1939_add_4_17 (.CI(n52315), .I0(GND_net), .I1(counter[15]), 
            .CO(n52316));
    SB_CARRY mult_16_add_1221_10 (.CI(n51687), .I0(n12096[7]), .I1(n658), 
            .CO(n51688));
    SB_LUT4 counter_1939_add_4_16_lut (.I0(GND_net), .I1(GND_net), .I2(counter[14]), 
            .I3(n52314), .O(n57[14])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1939_add_4_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_14_i17_3_lut (.I0(n130[16]), .I1(n182[16]), .I2(n181), 
            .I3(GND_net), .O(n207[16]));   // verilog/motorControl.v(48[18] 50[12])
    defparam mux_14_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_17_i177_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3715[14] ), 
            .I2(GND_net), .I3(GND_net), .O(n262));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i177_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_15_i17_3_lut (.I0(n207[16]), .I1(IntegralLimit[16]), .I2(n155), 
            .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3715[16] ));   // verilog/motorControl.v(48[18] 50[12])
    defparam mux_15_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_17_i377_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3715[16] ), 
            .I2(GND_net), .I3(GND_net), .O(n560));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i377_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i414_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3715[10] ), 
            .I2(GND_net), .I3(GND_net), .O(n615));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i414_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_13_inv_0_i18_1_lut (.I0(IntegralLimit[17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[17]));   // verilog/motorControl.v(49[22:36])
    defparam unary_minus_13_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY counter_1939_add_4_16 (.CI(n52314), .I0(GND_net), .I1(counter[14]), 
            .CO(n52315));
    SB_LUT4 mult_17_i463_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3715[10] ), 
            .I2(GND_net), .I3(GND_net), .O(n688));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i463_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_add_1221_9_lut (.I0(GND_net), .I1(n12096[6]), .I2(n585), 
            .I3(n51686), .O(n257[8])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_16_add_1221_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 counter_1939_add_4_15_lut (.I0(GND_net), .I1(GND_net), .I2(counter[13]), 
            .I3(n52313), .O(n57[13])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1939_add_4_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_13_inv_0_i2_1_lut (.I0(IntegralLimit[1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[1]));   // verilog/motorControl.v(49[22:36])
    defparam unary_minus_13_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_16_i359_2_lut (.I0(\Kp[7] ), .I1(n55[11]), .I2(GND_net), 
            .I3(GND_net), .O(n533));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i359_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i249_2_lut (.I0(\Kp[5] ), .I1(n55[5]), .I2(GND_net), 
            .I3(GND_net), .O(n369_adj_5161));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i249_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_13_inv_0_i3_1_lut (.I0(IntegralLimit[2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[2]));   // verilog/motorControl.v(49[22:36])
    defparam unary_minus_13_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY mult_16_add_1221_9 (.CI(n51686), .I0(n12096[6]), .I1(n585), 
            .CO(n51687));
    SB_LUT4 mult_17_i512_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3715[10] ), 
            .I2(GND_net), .I3(GND_net), .O(n761));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i512_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_add_1221_8_lut (.I0(GND_net), .I1(n12096[5]), .I2(n512), 
            .I3(n51685), .O(n257[7])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_16_add_1221_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i298_2_lut (.I0(\Kp[6] ), .I1(n55[5]), .I2(GND_net), 
            .I3(GND_net), .O(n442));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i298_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mult_16_add_1221_8 (.CI(n51685), .I0(n12096[5]), .I1(n512), 
            .CO(n51686));
    SB_LUT4 mult_16_i347_2_lut (.I0(\Kp[7] ), .I1(n55[5]), .I2(GND_net), 
            .I3(GND_net), .O(n515));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i347_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i226_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3715[14] ), 
            .I2(GND_net), .I3(GND_net), .O(n335));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i226_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i561_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3715[10] ), 
            .I2(GND_net), .I3(GND_net), .O(n834));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i561_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_13_inv_0_i4_1_lut (.I0(IntegralLimit[3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[3]));   // verilog/motorControl.v(49[22:36])
    defparam unary_minus_13_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY counter_1939_add_4_15 (.CI(n52313), .I0(GND_net), .I1(counter[13]), 
            .CO(n52314));
    SB_LUT4 add_6494_9_lut (.I0(GND_net), .I1(n19971[6]), .I2(n630), .I3(n51477), 
            .O(n19847[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6494_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_8_add_2_19 (.CI(n51042), .I0(setpoint[17]), .I1(\motor_state[17] ), 
            .CO(n51043));
    SB_LUT4 add_6494_8_lut (.I0(GND_net), .I1(n19971[5]), .I2(n557), .I3(n51476), 
            .O(n19847[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6494_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_i610_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3715[10] ), 
            .I2(GND_net), .I3(GND_net), .O(n907));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i610_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i59_2_lut (.I0(\Kp[1] ), .I1(n55[8]), .I2(GND_net), 
            .I3(GND_net), .O(n86));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i59_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i12_2_lut (.I0(\Kp[0] ), .I1(n55[9]), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_5159));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i12_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i659_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3715[10] ), 
            .I2(GND_net), .I3(GND_net), .O(n980));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i659_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 counter_1939_add_4_14_lut (.I0(GND_net), .I1(GND_net), .I2(counter[12]), 
            .I3(n52312), .O(n57[12])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1939_add_4_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i52136_2_lut_4_lut (.I0(n352[21]), .I1(n432[21]), .I2(n367), 
            .I3(n432[9]), .O(n67830));
    defparam i52136_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 mult_16_i108_2_lut (.I0(\Kp[2] ), .I1(n55[8]), .I2(GND_net), 
            .I3(GND_net), .O(n159));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i108_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i69_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3715[9] ), 
            .I2(GND_net), .I3(GND_net), .O(n101_adj_5277));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i69_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i22_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3715[10] ), 
            .I2(GND_net), .I3(GND_net), .O(n32_adj_5278));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i22_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_13_inv_0_i5_1_lut (.I0(IntegralLimit[4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[4]));   // verilog/motorControl.v(49[22:36])
    defparam unary_minus_13_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_16_i396_2_lut (.I0(\Kp[8] ), .I1(n55[5]), .I2(GND_net), 
            .I3(GND_net), .O(n588));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i396_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i157_2_lut (.I0(\Kp[3] ), .I1(n55[8]), .I2(GND_net), 
            .I3(GND_net), .O(n232));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i157_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i408_2_lut (.I0(\Kp[8] ), .I1(n55[11]), .I2(GND_net), 
            .I3(GND_net), .O(n606));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i408_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i118_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3715[9] ), 
            .I2(GND_net), .I3(GND_net), .O(n174_adj_5279));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i118_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6494_8 (.CI(n51476), .I0(n19971[5]), .I1(n557), .CO(n51477));
    SB_LUT4 add_6494_7_lut (.I0(GND_net), .I1(n19971[4]), .I2(n484), .I3(n51475), 
            .O(n19847[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6494_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_1939_add_4_14 (.CI(n52312), .I0(GND_net), .I1(counter[12]), 
            .CO(n52313));
    SB_LUT4 mult_16_add_1221_7_lut (.I0(GND_net), .I1(n12096[4]), .I2(n439), 
            .I3(n51684), .O(n257[6])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_16_add_1221_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_i167_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3715[9] ), 
            .I2(GND_net), .I3(GND_net), .O(n247_adj_5280));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i167_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i216_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3715[9] ), 
            .I2(GND_net), .I3(GND_net), .O(n320_adj_5281));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i216_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 counter_1939_add_4_13_lut (.I0(GND_net), .I1(GND_net), .I2(counter[11]), 
            .I3(n52311), .O(n57[11])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1939_add_4_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_16_add_1221_7 (.CI(n51684), .I0(n12096[4]), .I1(n439), 
            .CO(n51685));
    SB_CARRY counter_1939_add_4_13 (.CI(n52311), .I0(GND_net), .I1(counter[11]), 
            .CO(n52312));
    SB_LUT4 counter_1939_add_4_12_lut (.I0(GND_net), .I1(GND_net), .I2(counter[10]), 
            .I3(n52310), .O(n57[10])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1939_add_4_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_1939_add_4_12 (.CI(n52310), .I0(GND_net), .I1(counter[10]), 
            .CO(n52311));
    SB_LUT4 mult_17_i265_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3715[9] ), 
            .I2(GND_net), .I3(GND_net), .O(n393_adj_5282));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i265_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i314_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3715[9] ), 
            .I2(GND_net), .I3(GND_net), .O(n466_adj_5283));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i314_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i363_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3715[9] ), 
            .I2(GND_net), .I3(GND_net), .O(n539_adj_5284));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i363_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i296_2_lut (.I0(\Kp[6] ), .I1(n55[4]), .I2(GND_net), 
            .I3(GND_net), .O(n439));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i296_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i326_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3715[15] ), 
            .I2(GND_net), .I3(GND_net), .O(n484));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i326_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_add_1221_6_lut (.I0(GND_net), .I1(n12096[3]), .I2(n366_adj_5215), 
            .I3(n51683), .O(n257[5])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_16_add_1221_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_i412_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3715[9] ), 
            .I2(GND_net), .I3(GND_net), .O(n612_adj_5285));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i412_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6494_7 (.CI(n51475), .I0(n19971[4]), .I1(n484), .CO(n51476));
    SB_LUT4 i52150_2_lut_4_lut (.I0(n352[16]), .I1(n432[16]), .I2(n352[7]), 
            .I3(n432[7]), .O(n67844));
    defparam i52150_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 mult_17_i461_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3715[9] ), 
            .I2(GND_net), .I3(GND_net), .O(n685_adj_5286));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i461_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 counter_1939_add_4_11_lut (.I0(GND_net), .I1(GND_net), .I2(counter[9]), 
            .I3(n52309), .O(n57[9])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1939_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6494_6_lut (.I0(GND_net), .I1(n19971[3]), .I2(n411), .I3(n51474), 
            .O(n19847[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6494_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_i510_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3715[9] ), 
            .I2(GND_net), .I3(GND_net), .O(n758_adj_5287));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i510_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY counter_1939_add_4_11 (.CI(n52309), .I0(GND_net), .I1(counter[9]), 
            .CO(n52310));
    SB_LUT4 counter_1939_add_4_10_lut (.I0(GND_net), .I1(GND_net), .I2(counter[8]), 
            .I3(n52308), .O(n57[8])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1939_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_i559_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3715[9] ), 
            .I2(GND_net), .I3(GND_net), .O(n831_adj_5288));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i559_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_13_inv_0_i6_1_lut (.I0(IntegralLimit[5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[5]));   // verilog/motorControl.v(49[22:36])
    defparam unary_minus_13_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_17_i608_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3715[9] ), 
            .I2(GND_net), .I3(GND_net), .O(n904_adj_5289));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i608_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY counter_1939_add_4_10 (.CI(n52308), .I0(GND_net), .I1(counter[8]), 
            .CO(n52309));
    SB_LUT4 mult_17_i657_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3715[9] ), 
            .I2(GND_net), .I3(GND_net), .O(n977_adj_5290));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i657_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i706_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3715[9] ), 
            .I2(GND_net), .I3(GND_net), .O(n1050_adj_5291));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i706_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 counter_1939_add_4_9_lut (.I0(GND_net), .I1(GND_net), .I2(counter[7]), 
            .I3(n52307), .O(n57[7])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1939_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_1939_add_4_9 (.CI(n52307), .I0(GND_net), .I1(counter[7]), 
            .CO(n52308));
    SB_LUT4 counter_1939_add_4_8_lut (.I0(GND_net), .I1(GND_net), .I2(counter[6]), 
            .I3(n52306), .O(n57[6])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1939_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i81_2_lut (.I0(\Kp[1] ), .I1(n55[19]), .I2(GND_net), 
            .I3(GND_net), .O(n119_adj_5292));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i81_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i34_2_lut (.I0(\Kp[0] ), .I1(n55[20]), .I2(GND_net), 
            .I3(GND_net), .O(n50_adj_5293));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i34_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i375_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3715[15] ), 
            .I2(GND_net), .I3(GND_net), .O(n557));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i375_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY counter_1939_add_4_8 (.CI(n52306), .I0(GND_net), .I1(counter[6]), 
            .CO(n52307));
    SB_LUT4 counter_1939_add_4_7_lut (.I0(GND_net), .I1(GND_net), .I2(counter[5]), 
            .I3(n52305), .O(n57[5])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1939_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_i424_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3715[15] ), 
            .I2(GND_net), .I3(GND_net), .O(n630));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i424_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY counter_1939_add_4_7 (.CI(n52305), .I0(GND_net), .I1(counter[5]), 
            .CO(n52306));
    SB_LUT4 counter_1939_add_4_6_lut (.I0(GND_net), .I1(GND_net), .I2(counter[4]), 
            .I3(n52304), .O(n57[4])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1939_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_1939_add_4_6 (.CI(n52304), .I0(GND_net), .I1(counter[4]), 
            .CO(n52305));
    SB_LUT4 counter_1939_add_4_5_lut (.I0(GND_net), .I1(GND_net), .I2(counter[3]), 
            .I3(n52303), .O(n57[3])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1939_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_1939_add_4_5 (.CI(n52303), .I0(GND_net), .I1(counter[3]), 
            .CO(n52304));
    SB_LUT4 mult_16_i130_2_lut (.I0(\Kp[2] ), .I1(n55[19]), .I2(GND_net), 
            .I3(GND_net), .O(n192_adj_5294));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i130_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i179_2_lut (.I0(\Kp[3] ), .I1(n55[19]), .I2(GND_net), 
            .I3(GND_net), .O(n265));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i179_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i228_2_lut (.I0(\Kp[4] ), .I1(n55[19]), .I2(GND_net), 
            .I3(GND_net), .O(n338_adj_5295));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i228_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_13_inv_0_i19_1_lut (.I0(IntegralLimit[18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[18]));   // verilog/motorControl.v(49[22:36])
    defparam unary_minus_13_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_16_i277_2_lut (.I0(\Kp[5] ), .I1(n55[19]), .I2(GND_net), 
            .I3(GND_net), .O(n411_adj_5297));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i277_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i345_2_lut (.I0(\Kp[7] ), .I1(n55[4]), .I2(GND_net), 
            .I3(GND_net), .O(n512));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i345_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_13_inv_0_i7_1_lut (.I0(IntegralLimit[6]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[6]));   // verilog/motorControl.v(49[22:36])
    defparam unary_minus_13_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_16_i326_2_lut (.I0(\Kp[6] ), .I1(n55[19]), .I2(GND_net), 
            .I3(GND_net), .O(n484_adj_5298));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i326_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i375_2_lut (.I0(\Kp[7] ), .I1(n55[19]), .I2(GND_net), 
            .I3(GND_net), .O(n557_adj_5299));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i375_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i206_2_lut (.I0(\Kp[4] ), .I1(n55[8]), .I2(GND_net), 
            .I3(GND_net), .O(n305));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i206_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i37028_2_lut_4_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3715[20] ), 
            .I2(n36816), .I3(\Ki[1] ), .O(n20183));   // verilog/motorControl.v(51[27:38])
    defparam i37028_2_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 unary_minus_26_add_3_25_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5682[23]), 
            .I3(n51210), .O(n432[23])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6494_6 (.CI(n51474), .I0(n19971[3]), .I1(n411), .CO(n51475));
    SB_LUT4 mult_16_i445_2_lut (.I0(\Kp[9] ), .I1(n55[5]), .I2(GND_net), 
            .I3(GND_net), .O(n661));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i445_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i255_2_lut (.I0(\Kp[5] ), .I1(n55[8]), .I2(GND_net), 
            .I3(GND_net), .O(n378));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i255_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i394_2_lut (.I0(\Kp[8] ), .I1(n55[4]), .I2(GND_net), 
            .I3(GND_net), .O(n585));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i394_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_13_inv_0_i8_1_lut (.I0(IntegralLimit[7]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[7]));   // verilog/motorControl.v(49[22:36])
    defparam unary_minus_13_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_16_i304_2_lut (.I0(\Kp[6] ), .I1(n55[8]), .I2(GND_net), 
            .I3(GND_net), .O(n451));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i304_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i494_2_lut (.I0(\Kp[10] ), .I1(n55[5]), .I2(GND_net), 
            .I3(GND_net), .O(n734));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i494_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_13_inv_0_i9_1_lut (.I0(IntegralLimit[8]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[8]));   // verilog/motorControl.v(49[22:36])
    defparam unary_minus_13_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_16_i353_2_lut (.I0(\Kp[7] ), .I1(n55[8]), .I2(GND_net), 
            .I3(GND_net), .O(n524));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i353_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i275_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3715[14] ), 
            .I2(GND_net), .I3(GND_net), .O(n408));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i275_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i424_2_lut (.I0(\Kp[8] ), .I1(n55[19]), .I2(GND_net), 
            .I3(GND_net), .O(n630_adj_5300));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i424_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_26_add_3_24_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5682[22]), 
            .I3(n51209), .O(n432[22])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_26_add_3_24 (.CI(n51209), .I0(GND_net), .I1(n1_adj_5682[22]), 
            .CO(n51210));
    SB_LUT4 unary_minus_26_add_3_23_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5682[21]), 
            .I3(n51208), .O(n432[21])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_26_add_3_23 (.CI(n51208), .I0(GND_net), .I1(n1_adj_5682[21]), 
            .CO(n51209));
    SB_LUT4 counter_1939_add_4_4_lut (.I0(GND_net), .I1(GND_net), .I2(counter[2]), 
            .I3(n52302), .O(n57[2])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1939_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6427_12_lut (.I0(GND_net), .I1(n19352[9]), .I2(n840), 
            .I3(n52705), .O(n19089[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6427_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6427_11_lut (.I0(GND_net), .I1(n19352[8]), .I2(n767), 
            .I3(n52704), .O(n19089[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6427_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_i67_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3715[8] ), 
            .I2(GND_net), .I3(GND_net), .O(n98_adj_5301));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i67_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6427_11 (.CI(n52704), .I0(n19352[8]), .I1(n767), .CO(n52705));
    SB_LUT4 mult_16_i402_2_lut (.I0(\Kp[8] ), .I1(n55[8]), .I2(GND_net), 
            .I3(GND_net), .O(n597));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i402_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_13_inv_0_i10_1_lut (.I0(IntegralLimit[9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[9]));   // verilog/motorControl.v(49[22:36])
    defparam unary_minus_13_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_16_i451_2_lut (.I0(\Kp[9] ), .I1(n55[8]), .I2(GND_net), 
            .I3(GND_net), .O(n670));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i451_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6427_10_lut (.I0(GND_net), .I1(n19352[7]), .I2(n694), 
            .I3(n52703), .O(n19089[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6427_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_26_add_3_22_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5682[20]), 
            .I3(n51207), .O(n432[20])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6427_10 (.CI(n52703), .I0(n19352[7]), .I1(n694), .CO(n52704));
    SB_LUT4 add_6427_9_lut (.I0(GND_net), .I1(n19352[6]), .I2(n621), .I3(n52702), 
            .O(n19089[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6427_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_26_add_3_22 (.CI(n51207), .I0(GND_net), .I1(n1_adj_5682[20]), 
            .CO(n51208));
    SB_LUT4 mult_17_i20_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3715[9] ), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_5302));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i20_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i457_2_lut (.I0(\Kp[9] ), .I1(n55[11]), .I2(GND_net), 
            .I3(GND_net), .O(n679));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i457_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i116_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3715[8] ), 
            .I2(GND_net), .I3(GND_net), .O(n171_adj_5303));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i116_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i165_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3715[8] ), 
            .I2(GND_net), .I3(GND_net), .O(n244_adj_5304));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i165_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i214_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3715[8] ), 
            .I2(GND_net), .I3(GND_net), .O(n317_adj_5305));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i214_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6427_9 (.CI(n52702), .I0(n19352[6]), .I1(n621), .CO(n52703));
    SB_LUT4 mult_17_i263_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3715[8] ), 
            .I2(GND_net), .I3(GND_net), .O(n390_adj_5306));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i263_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6427_8_lut (.I0(GND_net), .I1(n19352[5]), .I2(n548), .I3(n52701), 
            .O(n19089[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6427_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6427_8 (.CI(n52701), .I0(n19352[5]), .I1(n548), .CO(n52702));
    SB_LUT4 mult_17_i312_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3715[8] ), 
            .I2(GND_net), .I3(GND_net), .O(n463_adj_5307));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i312_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6427_7_lut (.I0(GND_net), .I1(n19352[4]), .I2(n475), .I3(n52700), 
            .O(n19089[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6427_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6427_7 (.CI(n52700), .I0(n19352[4]), .I1(n475), .CO(n52701));
    SB_LUT4 mult_16_i506_2_lut (.I0(\Kp[10] ), .I1(n55[11]), .I2(GND_net), 
            .I3(GND_net), .O(n752));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i506_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6427_6_lut (.I0(GND_net), .I1(n19352[3]), .I2(n402), .I3(n52699), 
            .O(n19089[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6427_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6427_6 (.CI(n52699), .I0(n19352[3]), .I1(n402), .CO(n52700));
    SB_LUT4 mult_17_i361_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3715[8] ), 
            .I2(GND_net), .I3(GND_net), .O(n536_adj_5308));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i361_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6427_5_lut (.I0(GND_net), .I1(n19352[2]), .I2(n329), .I3(n52698), 
            .O(n19089[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6427_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_i410_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3715[8] ), 
            .I2(GND_net), .I3(GND_net), .O(n609_adj_5309));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i410_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6427_5 (.CI(n52698), .I0(n19352[2]), .I1(n329), .CO(n52699));
    SB_LUT4 unary_minus_26_add_3_21_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5682[19]), 
            .I3(n51206), .O(n432[19])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6427_4_lut (.I0(GND_net), .I1(n19352[1]), .I2(n256), .I3(n52697), 
            .O(n19089[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6427_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6427_4 (.CI(n52697), .I0(n19352[1]), .I1(n256), .CO(n52698));
    SB_LUT4 mult_16_i543_2_lut (.I0(\Kp[11] ), .I1(n55[5]), .I2(GND_net), 
            .I3(GND_net), .O(n807));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i543_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6427_3_lut (.I0(GND_net), .I1(n19352[0]), .I2(n183_adj_5192), 
            .I3(n52696), .O(n19089[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6427_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i555_2_lut (.I0(\Kp[11] ), .I1(n55[11]), .I2(GND_net), 
            .I3(GND_net), .O(n825));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i555_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6427_3 (.CI(n52696), .I0(n19352[0]), .I1(n183_adj_5192), 
            .CO(n52697));
    SB_LUT4 add_6427_2_lut (.I0(GND_net), .I1(n41_adj_5191), .I2(n110_adj_5189), 
            .I3(GND_net), .O(n19089[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6427_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6427_2 (.CI(GND_net), .I0(n41_adj_5191), .I1(n110_adj_5189), 
            .CO(n52696));
    SB_LUT4 mult_17_add_1225_24_lut (.I0(\PID_CONTROLLER.integral_23__N_3715[23] ), 
            .I1(n12720[21]), .I2(GND_net), .I3(n52695), .O(n12213[0])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1225_24_lut.LUT_INIT = 16'h6996;
    SB_LUT4 mult_17_add_1225_23_lut (.I0(GND_net), .I1(n12720[20]), .I2(GND_net), 
            .I3(n52694), .O(n49[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1225_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_i459_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3715[8] ), 
            .I2(GND_net), .I3(GND_net), .O(n682_adj_5310));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i459_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 sub_8_add_2_18_lut (.I0(GND_net), .I1(setpoint[16]), .I2(n20), 
            .I3(n51041), .O(n55[16])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_8_add_2_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_17_add_1225_23 (.CI(n52694), .I0(n12720[20]), .I1(GND_net), 
            .CO(n52695));
    SB_LUT4 add_6494_5_lut (.I0(GND_net), .I1(n19971[2]), .I2(n338_adj_5185), 
            .I3(n51473), .O(n19847[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6494_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_add_1225_22_lut (.I0(GND_net), .I1(n12720[19]), .I2(GND_net), 
            .I3(n52693), .O(n49[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1225_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_17_add_1225_22 (.CI(n52693), .I0(n12720[19]), .I1(GND_net), 
            .CO(n52694));
    SB_LUT4 mult_17_add_1225_21_lut (.I0(GND_net), .I1(n12720[18]), .I2(GND_net), 
            .I3(n52692), .O(n49[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1225_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_i508_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3715[8] ), 
            .I2(GND_net), .I3(GND_net), .O(n755_adj_5313));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i508_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mult_17_add_1225_21 (.CI(n52692), .I0(n12720[18]), .I1(GND_net), 
            .CO(n52693));
    SB_CARRY mult_16_add_1221_6 (.CI(n51683), .I0(n12096[3]), .I1(n366_adj_5215), 
            .CO(n51684));
    SB_LUT4 mult_17_add_1225_20_lut (.I0(GND_net), .I1(n12720[17]), .I2(GND_net), 
            .I3(n52691), .O(n49[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1225_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_26_add_3_21 (.CI(n51206), .I0(GND_net), .I1(n1_adj_5682[19]), 
            .CO(n51207));
    SB_CARRY mult_17_add_1225_20 (.CI(n52691), .I0(n12720[17]), .I1(GND_net), 
            .CO(n52692));
    SB_LUT4 mult_17_i324_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3715[14] ), 
            .I2(GND_net), .I3(GND_net), .O(n481));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i324_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_add_1225_19_lut (.I0(GND_net), .I1(n12720[16]), .I2(GND_net), 
            .I3(n52690), .O(n49[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1225_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_17_add_1225_19 (.CI(n52690), .I0(n12720[16]), .I1(GND_net), 
            .CO(n52691));
    SB_LUT4 mult_17_add_1225_18_lut (.I0(GND_net), .I1(n12720[15]), .I2(GND_net), 
            .I3(n52689), .O(n49[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1225_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_17_add_1225_18 (.CI(n52689), .I0(n12720[15]), .I1(GND_net), 
            .CO(n52690));
    SB_LUT4 mult_17_add_1225_17_lut (.I0(GND_net), .I1(n12720[14]), .I2(GND_net), 
            .I3(n52688), .O(n49[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1225_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_17_add_1225_17 (.CI(n52688), .I0(n12720[14]), .I1(GND_net), 
            .CO(n52689));
    SB_LUT4 mult_17_add_1225_16_lut (.I0(GND_net), .I1(n12720[13]), .I2(n1096_adj_5182), 
            .I3(n52687), .O(n49[15])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1225_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_17_add_1225_16 (.CI(n52687), .I0(n12720[13]), .I1(n1096_adj_5182), 
            .CO(n52688));
    SB_CARRY sub_8_add_2_18 (.CI(n51041), .I0(setpoint[16]), .I1(n20), 
            .CO(n51042));
    SB_CARRY counter_1939_add_4_4 (.CI(n52302), .I0(GND_net), .I1(counter[2]), 
            .CO(n52303));
    SB_LUT4 counter_1939_add_4_3_lut (.I0(GND_net), .I1(GND_net), .I2(counter[1]), 
            .I3(n52301), .O(n57[1])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1939_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_add_1225_15_lut (.I0(GND_net), .I1(n12720[12]), .I2(n1023_adj_5181), 
            .I3(n52686), .O(n49[14])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1225_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_17_add_1225_15 (.CI(n52686), .I0(n12720[12]), .I1(n1023_adj_5181), 
            .CO(n52687));
    SB_CARRY counter_1939_add_4_3 (.CI(n52301), .I0(GND_net), .I1(counter[1]), 
            .CO(n52302));
    SB_LUT4 mult_17_i557_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3715[8] ), 
            .I2(GND_net), .I3(GND_net), .O(n828_adj_5315));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i557_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 sub_8_add_2_17_lut (.I0(GND_net), .I1(setpoint[15]), .I2(\motor_state[15] ), 
            .I3(n51040), .O(n55[15])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_8_add_2_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_26_add_3_20_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5682[18]), 
            .I3(n51205), .O(n432[18])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6494_5 (.CI(n51473), .I0(n19971[2]), .I1(n338_adj_5185), 
            .CO(n51474));
    SB_LUT4 mult_17_add_1225_14_lut (.I0(GND_net), .I1(n12720[11]), .I2(n950_adj_5180), 
            .I3(n52685), .O(n49[13])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1225_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_17_add_1225_14 (.CI(n52685), .I0(n12720[11]), .I1(n950_adj_5180), 
            .CO(n52686));
    SB_LUT4 mult_17_add_1225_13_lut (.I0(GND_net), .I1(n12720[10]), .I2(n877), 
            .I3(n52684), .O(n49[12])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1225_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_add_1221_5_lut (.I0(GND_net), .I1(n12096[2]), .I2(n293_adj_5179), 
            .I3(n51682), .O(n257[4])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_16_add_1221_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_17_add_1225_13 (.CI(n52684), .I0(n12720[10]), .I1(n877), 
            .CO(n52685));
    SB_LUT4 mult_17_i606_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3715[8] ), 
            .I2(GND_net), .I3(GND_net), .O(n901_adj_5316));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i606_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i604_2_lut (.I0(\Kp[12] ), .I1(n55[11]), .I2(GND_net), 
            .I3(GND_net), .O(n898));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i604_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_add_1225_12_lut (.I0(GND_net), .I1(n12720[9]), .I2(n804), 
            .I3(n52683), .O(n49[11])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1225_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_i655_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3715[8] ), 
            .I2(GND_net), .I3(GND_net), .O(n974_adj_5317));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i655_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i653_2_lut (.I0(\Kp[13] ), .I1(n55[11]), .I2(GND_net), 
            .I3(GND_net), .O(n971));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i653_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mult_17_add_1225_12 (.CI(n52683), .I0(n12720[9]), .I1(n804), 
            .CO(n52684));
    SB_LUT4 mult_16_i500_2_lut (.I0(\Kp[10] ), .I1(n55[8]), .I2(GND_net), 
            .I3(GND_net), .O(n743));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i500_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_add_1225_11_lut (.I0(GND_net), .I1(n12720[8]), .I2(n731_adj_5318), 
            .I3(n52682), .O(n49[10])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1225_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_26_add_3_20 (.CI(n51205), .I0(GND_net), .I1(n1_adj_5682[18]), 
            .CO(n51206));
    SB_CARRY mult_17_add_1225_11 (.CI(n52682), .I0(n12720[8]), .I1(n731_adj_5318), 
            .CO(n52683));
    SB_LUT4 mult_17_add_1225_10_lut (.I0(GND_net), .I1(n12720[7]), .I2(n658_adj_5319), 
            .I3(n52681), .O(n49[9])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1225_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_i373_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3715[14] ), 
            .I2(GND_net), .I3(GND_net), .O(n554));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i373_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_26_add_3_19_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5682[17]), 
            .I3(n51204), .O(n432[17])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_17_add_1225_10 (.CI(n52681), .I0(n12720[7]), .I1(n658_adj_5319), 
            .CO(n52682));
    SB_LUT4 mult_17_add_1225_9_lut (.I0(GND_net), .I1(n12720[6]), .I2(n585_adj_5322), 
            .I3(n52680), .O(n49[8])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1225_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_17_add_1225_9 (.CI(n52680), .I0(n12720[6]), .I1(n585_adj_5322), 
            .CO(n52681));
    SB_LUT4 mult_17_add_1225_8_lut (.I0(GND_net), .I1(n12720[5]), .I2(n512_adj_5323), 
            .I3(n52679), .O(n49[7])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1225_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_17_add_1225_8 (.CI(n52679), .I0(n12720[5]), .I1(n512_adj_5323), 
            .CO(n52680));
    SB_LUT4 mult_17_add_1225_7_lut (.I0(GND_net), .I1(n12720[4]), .I2(n439_adj_5324), 
            .I3(n52678), .O(n49[6])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1225_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_17_add_1225_7 (.CI(n52678), .I0(n12720[4]), .I1(n439_adj_5324), 
            .CO(n52679));
    SB_LUT4 mult_17_add_1225_6_lut (.I0(GND_net), .I1(n12720[3]), .I2(n366_adj_5325), 
            .I3(n52677), .O(n49[5])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1225_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_17_add_1225_6 (.CI(n52677), .I0(n12720[3]), .I1(n366_adj_5325), 
            .CO(n52678));
    SB_LUT4 mult_17_add_1225_5_lut (.I0(GND_net), .I1(n12720[2]), .I2(n293_adj_5326), 
            .I3(n52676), .O(n49[4])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1225_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_17_add_1225_5 (.CI(n52676), .I0(n12720[2]), .I1(n293_adj_5326), 
            .CO(n52677));
    SB_LUT4 mult_17_add_1225_4_lut (.I0(GND_net), .I1(n12720[1]), .I2(n220), 
            .I3(n52675), .O(n49[3])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1225_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_17_add_1225_4 (.CI(n52675), .I0(n12720[1]), .I1(n220), 
            .CO(n52676));
    SB_CARRY mult_16_add_1221_5 (.CI(n51682), .I0(n12096[2]), .I1(n293_adj_5179), 
            .CO(n51683));
    SB_LUT4 mult_17_add_1225_3_lut (.I0(GND_net), .I1(n12720[0]), .I2(n147_adj_5327), 
            .I3(n52674), .O(n49[2])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1225_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_add_1221_4_lut (.I0(GND_net), .I1(n12096[1]), .I2(n220_adj_5328), 
            .I3(n51681), .O(n257[3])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_16_add_1221_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_17_add_1225_3 (.CI(n52674), .I0(n12720[0]), .I1(n147_adj_5327), 
            .CO(n52675));
    SB_LUT4 mult_17_add_1225_2_lut (.I0(GND_net), .I1(n5_adj_5329), .I2(n74), 
            .I3(GND_net), .O(n49[1])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1225_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_i704_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3715[8] ), 
            .I2(GND_net), .I3(GND_net), .O(n1047_adj_5330));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i704_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mult_17_add_1225_2 (.CI(GND_net), .I0(n5_adj_5329), .I1(n74), 
            .CO(n52674));
    SB_CARRY mult_16_add_1221_4 (.CI(n51681), .I0(n12096[1]), .I1(n220_adj_5328), 
            .CO(n51682));
    SB_LUT4 add_6087_23_lut (.I0(GND_net), .I1(n13685[20]), .I2(GND_net), 
            .I3(n52673), .O(n12720[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6087_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6087_22_lut (.I0(GND_net), .I1(n13685[19]), .I2(GND_net), 
            .I3(n52672), .O(n12720[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6087_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_8_add_2_17 (.CI(n51040), .I0(setpoint[15]), .I1(\motor_state[15] ), 
            .CO(n51041));
    SB_LUT4 counter_1939_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(counter[0]), 
            .I3(VCC_net), .O(n57[0])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1939_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_1939_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(counter[0]), 
            .CO(n52301));
    SB_LUT4 add_6494_4_lut (.I0(GND_net), .I1(n19971[1]), .I2(n265_adj_5331), 
            .I3(n51472), .O(n19847[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6494_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6087_22 (.CI(n52672), .I0(n13685[19]), .I1(GND_net), 
            .CO(n52673));
    SB_CARRY unary_minus_26_add_3_19 (.CI(n51204), .I0(GND_net), .I1(n1_adj_5682[17]), 
            .CO(n51205));
    SB_LUT4 add_6087_21_lut (.I0(GND_net), .I1(n13685[18]), .I2(GND_net), 
            .I3(n52671), .O(n12720[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6087_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_26_add_3_18_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5682[16]), 
            .I3(n51203), .O(n432[16])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_8_add_2_16_lut (.I0(GND_net), .I1(setpoint[14]), .I2(\motor_state[14] ), 
            .I3(n51039), .O(n55[14])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_8_add_2_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_26_add_3_18 (.CI(n51203), .I0(GND_net), .I1(n1_adj_5682[16]), 
            .CO(n51204));
    SB_CARRY add_6087_21 (.CI(n52671), .I0(n13685[18]), .I1(GND_net), 
            .CO(n52672));
    SB_LUT4 mult_16_add_1221_3_lut (.I0(GND_net), .I1(n12096[0]), .I2(n147_adj_5333), 
            .I3(n51680), .O(n257[2])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_16_add_1221_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6087_20_lut (.I0(GND_net), .I1(n13685[17]), .I2(GND_net), 
            .I3(n52670), .O(n12720[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6087_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6087_20 (.CI(n52670), .I0(n13685[17]), .I1(GND_net), 
            .CO(n52671));
    SB_LUT4 add_6087_19_lut (.I0(GND_net), .I1(n13685[16]), .I2(GND_net), 
            .I3(n52669), .O(n12720[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6087_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i592_2_lut (.I0(\Kp[12] ), .I1(n55[5]), .I2(GND_net), 
            .I3(GND_net), .O(n880));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i592_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6087_19 (.CI(n52669), .I0(n13685[16]), .I1(GND_net), 
            .CO(n52670));
    SB_LUT4 add_6087_18_lut (.I0(GND_net), .I1(n13685[15]), .I2(GND_net), 
            .I3(n52668), .O(n12720[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6087_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_26_add_3_17_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5682[15]), 
            .I3(n51202), .O(n432[15])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6087_18 (.CI(n52668), .I0(n13685[15]), .I1(GND_net), 
            .CO(n52669));
    SB_CARRY add_6494_4 (.CI(n51472), .I0(n19971[1]), .I1(n265_adj_5331), 
            .CO(n51473));
    SB_LUT4 add_6494_3_lut (.I0(GND_net), .I1(n19971[0]), .I2(n192_adj_5335), 
            .I3(n51471), .O(n19847[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6494_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6087_17_lut (.I0(GND_net), .I1(n13685[14]), .I2(GND_net), 
            .I3(n52667), .O(n12720[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6087_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6087_17 (.CI(n52667), .I0(n13685[14]), .I1(GND_net), 
            .CO(n52668));
    SB_LUT4 add_6520_7_lut (.I0(GND_net), .I1(n61429), .I2(n490), .I3(n51352), 
            .O(n20065[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6520_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_26_add_3_17 (.CI(n51202), .I0(GND_net), .I1(n1_adj_5682[15]), 
            .CO(n51203));
    SB_LUT4 add_6520_6_lut (.I0(GND_net), .I1(n20133[3]), .I2(n417), .I3(n51351), 
            .O(n20065[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6520_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_16_add_1221_3 (.CI(n51680), .I0(n12096[0]), .I1(n147_adj_5333), 
            .CO(n51681));
    SB_LUT4 add_6087_16_lut (.I0(GND_net), .I1(n13685[13]), .I2(n1099_adj_5338), 
            .I3(n52666), .O(n12720[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6087_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6520_6 (.CI(n51351), .I0(n20133[3]), .I1(n417), .CO(n51352));
    SB_LUT4 unary_minus_26_add_3_16_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5682[14]), 
            .I3(n51201), .O(n432[14])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6087_16 (.CI(n52666), .I0(n13685[13]), .I1(n1099_adj_5338), 
            .CO(n52667));
    SB_LUT4 add_6087_15_lut (.I0(GND_net), .I1(n13685[12]), .I2(n1026_adj_5341), 
            .I3(n52665), .O(n12720[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6087_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_add_1221_2_lut (.I0(GND_net), .I1(n5_adj_5342), .I2(n74_adj_5343), 
            .I3(GND_net), .O(n257[1])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_16_add_1221_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6087_15 (.CI(n52665), .I0(n13685[12]), .I1(n1026_adj_5341), 
            .CO(n52666));
    SB_CARRY unary_minus_26_add_3_16 (.CI(n51201), .I0(GND_net), .I1(n1_adj_5682[14]), 
            .CO(n51202));
    SB_LUT4 unary_minus_26_add_3_15_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5682[13]), 
            .I3(n51200), .O(n432[13])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6087_14_lut (.I0(GND_net), .I1(n13685[11]), .I2(n953_adj_5345), 
            .I3(n52664), .O(n12720[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6087_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6087_14 (.CI(n52664), .I0(n13685[11]), .I1(n953_adj_5345), 
            .CO(n52665));
    SB_CARRY sub_8_add_2_16 (.CI(n51039), .I0(setpoint[14]), .I1(\motor_state[14] ), 
            .CO(n51040));
    SB_CARRY unary_minus_26_add_3_15 (.CI(n51200), .I0(GND_net), .I1(n1_adj_5682[13]), 
            .CO(n51201));
    SB_CARRY mult_16_add_1221_2 (.CI(GND_net), .I0(n5_adj_5342), .I1(n74_adj_5343), 
            .CO(n51680));
    SB_LUT4 add_6087_13_lut (.I0(GND_net), .I1(n13685[10]), .I2(n880_adj_5346), 
            .I3(n52663), .O(n12720[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6087_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6087_13 (.CI(n52663), .I0(n13685[10]), .I1(n880_adj_5346), 
            .CO(n52664));
    SB_CARRY add_6494_3 (.CI(n51471), .I0(n19971[0]), .I1(n192_adj_5335), 
            .CO(n51472));
    SB_LUT4 add_6494_2_lut (.I0(GND_net), .I1(n50_adj_5347), .I2(n119_adj_5348), 
            .I3(GND_net), .O(n19847[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6494_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6087_12_lut (.I0(GND_net), .I1(n13685[9]), .I2(n807_adj_5349), 
            .I3(n52662), .O(n12720[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6087_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6087_12 (.CI(n52662), .I0(n13685[9]), .I1(n807_adj_5349), 
            .CO(n52663));
    SB_LUT4 add_6520_5_lut (.I0(GND_net), .I1(n20136), .I2(n344), .I3(n51350), 
            .O(n20065[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6520_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6460_11_lut (.I0(GND_net), .I1(n19689[8]), .I2(n770), 
            .I3(n51679), .O(n19493[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6460_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6087_11_lut (.I0(GND_net), .I1(n13685[8]), .I2(n734_adj_5351), 
            .I3(n52661), .O(n12720[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6087_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6087_11 (.CI(n52661), .I0(n13685[8]), .I1(n734_adj_5351), 
            .CO(n52662));
    SB_LUT4 add_6460_10_lut (.I0(GND_net), .I1(n19689[7]), .I2(n697), 
            .I3(n51678), .O(n19493[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6460_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_26_add_3_14_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5682[12]), 
            .I3(n51199), .O(n432[12])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6087_10_lut (.I0(GND_net), .I1(n13685[7]), .I2(n661_adj_5353), 
            .I3(n52660), .O(n12720[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6087_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_26_add_3_14 (.CI(n51199), .I0(GND_net), .I1(n1_adj_5682[12]), 
            .CO(n51200));
    SB_LUT4 sub_8_add_2_15_lut (.I0(GND_net), .I1(setpoint[13]), .I2(\motor_state[13] ), 
            .I3(n51038), .O(n55[13])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_8_add_2_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_26_add_3_13_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5682[11]), 
            .I3(n51198), .O(n432[11])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6087_10 (.CI(n52660), .I0(n13685[7]), .I1(n661_adj_5353), 
            .CO(n52661));
    SB_CARRY add_6520_5 (.CI(n51350), .I0(n20136), .I1(n344), .CO(n51351));
    SB_LUT4 add_6087_9_lut (.I0(GND_net), .I1(n13685[6]), .I2(n588_adj_5356), 
            .I3(n52659), .O(n12720[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6087_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i549_2_lut (.I0(\Kp[11] ), .I1(n55[8]), .I2(GND_net), 
            .I3(GND_net), .O(n816));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i549_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY sub_8_add_2_15 (.CI(n51038), .I0(setpoint[13]), .I1(\motor_state[13] ), 
            .CO(n51039));
    SB_CARRY add_6494_2 (.CI(GND_net), .I0(n50_adj_5347), .I1(n119_adj_5348), 
            .CO(n51471));
    SB_LUT4 add_6259_18_lut (.I0(GND_net), .I1(n16974[15]), .I2(GND_net), 
            .I3(n51470), .O(n16363[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6259_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6087_9 (.CI(n52659), .I0(n13685[6]), .I1(n588_adj_5356), 
            .CO(n52660));
    SB_LUT4 add_6087_8_lut (.I0(GND_net), .I1(n13685[5]), .I2(n515_adj_5357), 
            .I3(n52658), .O(n12720[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6087_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_i753_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3715[8] ), 
            .I2(GND_net), .I3(GND_net), .O(n1120_adj_5358));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i753_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6520_4_lut (.I0(GND_net), .I1(n20137), .I2(n271), .I3(n51349), 
            .O(n20065[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6520_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6460_10 (.CI(n51678), .I0(n19689[7]), .I1(n697), .CO(n51679));
    SB_LUT4 add_6460_9_lut (.I0(GND_net), .I1(n19689[6]), .I2(n624), .I3(n51677), 
            .O(n19493[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6460_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6520_4 (.CI(n51349), .I0(n20137), .I1(n271), .CO(n51350));
    SB_LUT4 add_6520_3_lut (.I0(GND_net), .I1(n20138), .I2(n198), .I3(n51348), 
            .O(n20065[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6520_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_26_add_3_13 (.CI(n51198), .I0(GND_net), .I1(n1_adj_5682[11]), 
            .CO(n51199));
    SB_CARRY add_6087_8 (.CI(n52658), .I0(n13685[5]), .I1(n515_adj_5357), 
            .CO(n52659));
    SB_LUT4 add_6087_7_lut (.I0(GND_net), .I1(n13685[4]), .I2(n442_adj_5361), 
            .I3(n52657), .O(n12720[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6087_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_26_add_3_12_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5682[10]), 
            .I3(n51197), .O(n432[10])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_26_add_3_12 (.CI(n51197), .I0(GND_net), .I1(n1_adj_5682[10]), 
            .CO(n51198));
    SB_CARRY add_6087_7 (.CI(n52657), .I0(n13685[4]), .I1(n442_adj_5361), 
            .CO(n52658));
    SB_CARRY add_6460_9 (.CI(n51677), .I0(n19689[6]), .I1(n624), .CO(n51678));
    SB_LUT4 add_6087_6_lut (.I0(GND_net), .I1(n13685[3]), .I2(n369_adj_5363), 
            .I3(n52656), .O(n12720[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6087_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_i65_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3715[7] ), 
            .I2(GND_net), .I3(GND_net), .O(n95_adj_5364));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i65_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6460_8_lut (.I0(GND_net), .I1(n19689[5]), .I2(n551), .I3(n51676), 
            .O(n19493[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6460_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_26_add_3_11_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5682[9]), 
            .I3(n51196), .O(n432[9])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6460_8 (.CI(n51676), .I0(n19689[5]), .I1(n551), .CO(n51677));
    SB_CARRY unary_minus_26_add_3_11 (.CI(n51196), .I0(GND_net), .I1(n1_adj_5682[9]), 
            .CO(n51197));
    SB_LUT4 sub_8_add_2_14_lut (.I0(GND_net), .I1(setpoint[12]), .I2(\motor_state[12] ), 
            .I3(n51037), .O(n55[12])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_8_add_2_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_26_add_3_10_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5682[8]), 
            .I3(n51195), .O(n432[8])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_8_add_2_14 (.CI(n51037), .I0(setpoint[12]), .I1(\motor_state[12] ), 
            .CO(n51038));
    SB_LUT4 add_6460_7_lut (.I0(GND_net), .I1(n19689[4]), .I2(n478), .I3(n51675), 
            .O(n19493[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6460_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6520_3 (.CI(n51348), .I0(n20138), .I1(n198), .CO(n51349));
    SB_CARRY add_6460_7 (.CI(n51675), .I0(n19689[4]), .I1(n478), .CO(n51676));
    SB_LUT4 add_6520_2_lut (.I0(GND_net), .I1(n56), .I2(n125), .I3(GND_net), 
            .O(n20065[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6520_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6460_6_lut (.I0(GND_net), .I1(n19689[3]), .I2(n405), .I3(n51674), 
            .O(n19493[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6460_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6259_17_lut (.I0(GND_net), .I1(n16974[14]), .I2(GND_net), 
            .I3(n51469), .O(n16363[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6259_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6520_2 (.CI(GND_net), .I0(n56), .I1(n125), .CO(n51348));
    SB_CARRY add_6460_6 (.CI(n51674), .I0(n19689[3]), .I1(n405), .CO(n51675));
    SB_CARRY add_6259_17 (.CI(n51469), .I0(n16974[14]), .I1(GND_net), 
            .CO(n51470));
    SB_CARRY add_6087_6 (.CI(n52656), .I0(n13685[3]), .I1(n369_adj_5363), 
            .CO(n52657));
    SB_LUT4 add_6087_5_lut (.I0(GND_net), .I1(n13685[2]), .I2(n296_adj_5369), 
            .I3(n52655), .O(n12720[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6087_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_26_add_3_10 (.CI(n51195), .I0(GND_net), .I1(n1_adj_5682[8]), 
            .CO(n51196));
    SB_LUT4 add_6379_14_lut (.I0(GND_net), .I1(n18778[11]), .I2(n980_adj_5370), 
            .I3(n51347), .O(n18415[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6379_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_26_add_3_9_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5682[7]), 
            .I3(n51194), .O(n432[7])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6087_5 (.CI(n52655), .I0(n13685[2]), .I1(n296_adj_5369), 
            .CO(n52656));
    SB_LUT4 add_6087_4_lut (.I0(GND_net), .I1(n13685[1]), .I2(n223_adj_5372), 
            .I3(n52654), .O(n12720[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6087_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6087_4 (.CI(n52654), .I0(n13685[1]), .I1(n223_adj_5372), 
            .CO(n52655));
    SB_LUT4 mult_17_i18_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3715[8] ), 
            .I2(GND_net), .I3(GND_net), .O(n26_adj_5373));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i18_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY unary_minus_26_add_3_9 (.CI(n51194), .I0(GND_net), .I1(n1_adj_5682[7]), 
            .CO(n51195));
    SB_LUT4 add_6087_3_lut (.I0(GND_net), .I1(n13685[0]), .I2(n150_adj_5374), 
            .I3(n52653), .O(n12720[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6087_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_26_add_3_8_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5682[6]), 
            .I3(n51193), .O(n432[6])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6259_16_lut (.I0(GND_net), .I1(n16974[13]), .I2(n1114), 
            .I3(n51468), .O(n16363[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6259_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6379_13_lut (.I0(GND_net), .I1(n18778[10]), .I2(n907_adj_5376), 
            .I3(n51346), .O(n18415[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6379_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6087_3 (.CI(n52653), .I0(n13685[0]), .I1(n150_adj_5374), 
            .CO(n52654));
    SB_LUT4 mult_17_i114_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3715[7] ), 
            .I2(GND_net), .I3(GND_net), .O(n168_adj_5377));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i114_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i422_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3715[14] ), 
            .I2(GND_net), .I3(GND_net), .O(n627));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i422_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6087_2_lut (.I0(GND_net), .I1(n8_adj_5378), .I2(n77_adj_5379), 
            .I3(GND_net), .O(n12720[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6087_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6259_16 (.CI(n51468), .I0(n16974[13]), .I1(n1114), .CO(n51469));
    SB_CARRY unary_minus_26_add_3_8 (.CI(n51193), .I0(GND_net), .I1(n1_adj_5682[6]), 
            .CO(n51194));
    SB_CARRY add_6087_2 (.CI(GND_net), .I0(n8_adj_5378), .I1(n77_adj_5379), 
            .CO(n52653));
    SB_LUT4 add_6460_5_lut (.I0(GND_net), .I1(n19689[2]), .I2(n332_adj_5380), 
            .I3(n51673), .O(n19493[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6460_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_26_add_3_7_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5682[5]), 
            .I3(n51192), .O(n432[5])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6130_22_lut (.I0(GND_net), .I1(n14563[19]), .I2(GND_net), 
            .I3(n52652), .O(n13685[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6130_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6148_21_lut (.I0(GND_net), .I1(n14921[18]), .I2(GND_net), 
            .I3(n51590), .O(n14082[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6148_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6148_20_lut (.I0(GND_net), .I1(n14921[17]), .I2(GND_net), 
            .I3(n51589), .O(n14082[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6148_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6130_21_lut (.I0(GND_net), .I1(n14563[18]), .I2(GND_net), 
            .I3(n52651), .O(n13685[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6130_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6130_21 (.CI(n52651), .I0(n14563[18]), .I1(GND_net), 
            .CO(n52652));
    SB_LUT4 add_6259_15_lut (.I0(GND_net), .I1(n16974[12]), .I2(n1041), 
            .I3(n51467), .O(n16363[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6259_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6130_20_lut (.I0(GND_net), .I1(n14563[17]), .I2(GND_net), 
            .I3(n52650), .O(n13685[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6130_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6148_20 (.CI(n51589), .I0(n14921[17]), .I1(GND_net), 
            .CO(n51590));
    SB_CARRY add_6130_20 (.CI(n52650), .I0(n14563[17]), .I1(GND_net), 
            .CO(n52651));
    SB_CARRY add_6460_5 (.CI(n51673), .I0(n19689[2]), .I1(n332_adj_5380), 
            .CO(n51674));
    SB_CARRY add_6379_13 (.CI(n51346), .I0(n18778[10]), .I1(n907_adj_5376), 
            .CO(n51347));
    SB_CARRY add_6259_15 (.CI(n51467), .I0(n16974[12]), .I1(n1041), .CO(n51468));
    SB_LUT4 add_6130_19_lut (.I0(GND_net), .I1(n14563[16]), .I2(GND_net), 
            .I3(n52649), .O(n13685[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6130_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6130_19 (.CI(n52649), .I0(n14563[16]), .I1(GND_net), 
            .CO(n52650));
    SB_LUT4 add_6130_18_lut (.I0(GND_net), .I1(n14563[15]), .I2(GND_net), 
            .I3(n52648), .O(n13685[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6130_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6379_12_lut (.I0(GND_net), .I1(n18778[9]), .I2(n834_adj_5383), 
            .I3(n51345), .O(n18415[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6379_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_26_add_3_7 (.CI(n51192), .I0(GND_net), .I1(n1_adj_5682[5]), 
            .CO(n51193));
    SB_CARRY add_6379_12 (.CI(n51345), .I0(n18778[9]), .I1(n834_adj_5383), 
            .CO(n51346));
    SB_CARRY add_6130_18 (.CI(n52648), .I0(n14563[15]), .I1(GND_net), 
            .CO(n52649));
    SB_LUT4 add_6130_17_lut (.I0(GND_net), .I1(n14563[14]), .I2(GND_net), 
            .I3(n52647), .O(n13685[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6130_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6130_17 (.CI(n52647), .I0(n14563[14]), .I1(GND_net), 
            .CO(n52648));
    SB_LUT4 add_6379_11_lut (.I0(GND_net), .I1(n18778[8]), .I2(n761_adj_5384), 
            .I3(n51344), .O(n18415[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6379_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_26_add_3_6_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5682[4]), 
            .I3(n51191), .O(n432[4])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6379_11 (.CI(n51344), .I0(n18778[8]), .I1(n761_adj_5384), 
            .CO(n51345));
    SB_CARRY unary_minus_26_add_3_6 (.CI(n51191), .I0(GND_net), .I1(n1_adj_5682[4]), 
            .CO(n51192));
    SB_LUT4 add_6130_16_lut (.I0(GND_net), .I1(n14563[13]), .I2(n1102_adj_5386), 
            .I3(n52646), .O(n13685[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6130_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_26_add_3_5_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5682[3]), 
            .I3(n51190), .O(n432[3])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6130_16 (.CI(n52646), .I0(n14563[13]), .I1(n1102_adj_5386), 
            .CO(n52647));
    SB_LUT4 add_6130_15_lut (.I0(GND_net), .I1(n14563[12]), .I2(n1029_adj_5388), 
            .I3(n52645), .O(n13685[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6130_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6130_15 (.CI(n52645), .I0(n14563[12]), .I1(n1029_adj_5388), 
            .CO(n52646));
    SB_LUT4 add_6259_14_lut (.I0(GND_net), .I1(n16974[11]), .I2(n968), 
            .I3(n51466), .O(n16363[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6259_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6259_14 (.CI(n51466), .I0(n16974[11]), .I1(n968), .CO(n51467));
    SB_LUT4 add_6130_14_lut (.I0(GND_net), .I1(n14563[11]), .I2(n956_adj_5389), 
            .I3(n52644), .O(n13685[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6130_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6130_14 (.CI(n52644), .I0(n14563[11]), .I1(n956_adj_5389), 
            .CO(n52645));
    SB_LUT4 add_6130_13_lut (.I0(GND_net), .I1(n14563[10]), .I2(n883_adj_5390), 
            .I3(n52643), .O(n13685[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6130_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6379_10_lut (.I0(GND_net), .I1(n18778[7]), .I2(n688_adj_5391), 
            .I3(n51343), .O(n18415[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6379_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6259_13_lut (.I0(GND_net), .I1(n16974[10]), .I2(n895), 
            .I3(n51465), .O(n16363[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6259_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_26_add_3_5 (.CI(n51190), .I0(GND_net), .I1(n1_adj_5682[3]), 
            .CO(n51191));
    SB_CARRY add_6379_10 (.CI(n51343), .I0(n18778[7]), .I1(n688_adj_5391), 
            .CO(n51344));
    SB_CARRY add_6130_13 (.CI(n52643), .I0(n14563[10]), .I1(n883_adj_5390), 
            .CO(n52644));
    SB_LUT4 unary_minus_26_add_3_4_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5682[2]), 
            .I3(n51189), .O(n432[2])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6130_12_lut (.I0(GND_net), .I1(n14563[9]), .I2(n810_adj_5394), 
            .I3(n52642), .O(n13685[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6130_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6130_12 (.CI(n52642), .I0(n14563[9]), .I1(n810_adj_5394), 
            .CO(n52643));
    SB_LUT4 add_6130_11_lut (.I0(GND_net), .I1(n14563[8]), .I2(n737_adj_5395), 
            .I3(n52641), .O(n13685[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6130_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6130_11 (.CI(n52641), .I0(n14563[8]), .I1(n737_adj_5395), 
            .CO(n52642));
    SB_LUT4 add_6130_10_lut (.I0(GND_net), .I1(n14563[7]), .I2(n664_adj_5396), 
            .I3(n52640), .O(n13685[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6130_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6379_9_lut (.I0(GND_net), .I1(n18778[6]), .I2(n615_adj_5397), 
            .I3(n51342), .O(n18415[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6379_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6130_10 (.CI(n52640), .I0(n14563[7]), .I1(n664_adj_5396), 
            .CO(n52641));
    SB_CARRY unary_minus_26_add_3_4 (.CI(n51189), .I0(GND_net), .I1(n1_adj_5682[2]), 
            .CO(n51190));
    SB_LUT4 add_6130_9_lut (.I0(GND_net), .I1(n14563[6]), .I2(n591_adj_5398), 
            .I3(n52639), .O(n13685[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6130_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6130_9 (.CI(n52639), .I0(n14563[6]), .I1(n591_adj_5398), 
            .CO(n52640));
    SB_LUT4 add_6130_8_lut (.I0(GND_net), .I1(n14563[5]), .I2(n518_adj_5399), 
            .I3(n52638), .O(n13685[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6130_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6130_8 (.CI(n52638), .I0(n14563[5]), .I1(n518_adj_5399), 
            .CO(n52639));
    SB_LUT4 add_6148_19_lut (.I0(GND_net), .I1(n14921[16]), .I2(GND_net), 
            .I3(n51588), .O(n14082[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6148_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6460_4_lut (.I0(GND_net), .I1(n19689[1]), .I2(n259), .I3(n51672), 
            .O(n19493[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6460_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6130_7_lut (.I0(GND_net), .I1(n14563[4]), .I2(n445_adj_5400), 
            .I3(n52637), .O(n13685[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6130_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6130_7 (.CI(n52637), .I0(n14563[4]), .I1(n445_adj_5400), 
            .CO(n52638));
    SB_CARRY add_6460_4 (.CI(n51672), .I0(n19689[1]), .I1(n259), .CO(n51673));
    SB_LUT4 sub_8_add_2_13_lut (.I0(GND_net), .I1(setpoint[11]), .I2(\motor_state[11] ), 
            .I3(n51036), .O(n55[11])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_8_add_2_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6379_9 (.CI(n51342), .I0(n18778[6]), .I1(n615_adj_5397), 
            .CO(n51343));
    SB_CARRY add_6148_19 (.CI(n51588), .I0(n14921[16]), .I1(GND_net), 
            .CO(n51589));
    SB_LUT4 add_6130_6_lut (.I0(GND_net), .I1(n14563[3]), .I2(n372_adj_5401), 
            .I3(n52636), .O(n13685[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6130_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6130_6 (.CI(n52636), .I0(n14563[3]), .I1(n372_adj_5401), 
            .CO(n52637));
    SB_LUT4 add_6130_5_lut (.I0(GND_net), .I1(n14563[2]), .I2(n299_adj_5402), 
            .I3(n52635), .O(n13685[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6130_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6130_5 (.CI(n52635), .I0(n14563[2]), .I1(n299_adj_5402), 
            .CO(n52636));
    SB_LUT4 add_6460_3_lut (.I0(GND_net), .I1(n19689[0]), .I2(n186_adj_5403), 
            .I3(n51671), .O(n19493[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6460_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6259_13 (.CI(n51465), .I0(n16974[10]), .I1(n895), .CO(n51466));
    SB_LUT4 add_6130_4_lut (.I0(GND_net), .I1(n14563[1]), .I2(n226_adj_5404), 
            .I3(n52634), .O(n13685[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6130_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6130_4 (.CI(n52634), .I0(n14563[1]), .I1(n226_adj_5404), 
            .CO(n52635));
    SB_LUT4 add_6130_3_lut (.I0(GND_net), .I1(n14563[0]), .I2(n153_adj_5405), 
            .I3(n52633), .O(n13685[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6130_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6148_18_lut (.I0(GND_net), .I1(n14921[15]), .I2(GND_net), 
            .I3(n51587), .O(n14082[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6148_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6130_3 (.CI(n52633), .I0(n14563[0]), .I1(n153_adj_5405), 
            .CO(n52634));
    SB_LUT4 add_6130_2_lut (.I0(GND_net), .I1(n11_adj_5406), .I2(n80_adj_5407), 
            .I3(GND_net), .O(n13685[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6130_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6259_12_lut (.I0(GND_net), .I1(n16974[9]), .I2(n822), 
            .I3(n51464), .O(n16363[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6259_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6379_8_lut (.I0(GND_net), .I1(n18778[5]), .I2(n542_adj_5408), 
            .I3(n51341), .O(n18415[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6379_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_26_add_3_3_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5682[1]), 
            .I3(n51188), .O(n455)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6379_8 (.CI(n51341), .I0(n18778[5]), .I1(n542_adj_5408), 
            .CO(n51342));
    SB_CARRY add_6130_2 (.CI(GND_net), .I0(n11_adj_5406), .I1(n80_adj_5407), 
            .CO(n52633));
    SB_LUT4 add_6170_21_lut (.I0(GND_net), .I1(n15359[18]), .I2(GND_net), 
            .I3(n52632), .O(n14563[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6170_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6170_20_lut (.I0(GND_net), .I1(n15359[17]), .I2(GND_net), 
            .I3(n52631), .O(n14563[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6170_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6170_20 (.CI(n52631), .I0(n15359[17]), .I1(GND_net), 
            .CO(n52632));
    SB_LUT4 add_6379_7_lut (.I0(GND_net), .I1(n18778[4]), .I2(n469_adj_5410), 
            .I3(n51340), .O(n18415[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6379_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_i163_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3715[7] ), 
            .I2(GND_net), .I3(GND_net), .O(n241_adj_5411));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i163_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY unary_minus_26_add_3_3 (.CI(n51188), .I0(GND_net), .I1(n1_adj_5682[1]), 
            .CO(n51189));
    SB_LUT4 add_6170_19_lut (.I0(GND_net), .I1(n15359[16]), .I2(GND_net), 
            .I3(n52630), .O(n14563[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6170_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6170_19 (.CI(n52630), .I0(n15359[16]), .I1(GND_net), 
            .CO(n52631));
    SB_LUT4 add_6170_18_lut (.I0(GND_net), .I1(n15359[15]), .I2(GND_net), 
            .I3(n52629), .O(n14563[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6170_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6379_7 (.CI(n51340), .I0(n18778[4]), .I1(n469_adj_5410), 
            .CO(n51341));
    SB_LUT4 unary_minus_13_inv_0_i11_1_lut (.I0(IntegralLimit[10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[10]));   // verilog/motorControl.v(49[22:36])
    defparam unary_minus_13_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_6170_18 (.CI(n52629), .I0(n15359[15]), .I1(GND_net), 
            .CO(n52630));
    SB_LUT4 add_6170_17_lut (.I0(GND_net), .I1(n15359[14]), .I2(GND_net), 
            .I3(n52628), .O(n14563[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6170_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6170_17 (.CI(n52628), .I0(n15359[14]), .I1(GND_net), 
            .CO(n52629));
    SB_LUT4 add_6170_16_lut (.I0(GND_net), .I1(n15359[13]), .I2(n1105), 
            .I3(n52627), .O(n14563[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6170_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_26_add_3_2_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5682[0]), 
            .I3(VCC_net), .O(n456)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_26_add_3_2 (.CI(VCC_net), .I0(GND_net), .I1(n1_adj_5682[0]), 
            .CO(n51188));
    SB_CARRY add_6460_3 (.CI(n51671), .I0(n19689[0]), .I1(n186_adj_5403), 
            .CO(n51672));
    SB_LUT4 add_6460_2_lut (.I0(GND_net), .I1(n44_adj_5413), .I2(n113_adj_5414), 
            .I3(GND_net), .O(n19493[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6460_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6259_12 (.CI(n51464), .I0(n16974[9]), .I1(n822), .CO(n51465));
    SB_CARRY add_6170_16 (.CI(n52627), .I0(n15359[13]), .I1(n1105), .CO(n52628));
    SB_LUT4 add_6259_11_lut (.I0(GND_net), .I1(n16974[8]), .I2(n749), 
            .I3(n51463), .O(n16363[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6259_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6170_15_lut (.I0(GND_net), .I1(n15359[12]), .I2(n1032), 
            .I3(n52626), .O(n14563[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6170_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6379_6_lut (.I0(GND_net), .I1(n18778[3]), .I2(n396_adj_5415), 
            .I3(n51339), .O(n18415[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6379_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6379_6 (.CI(n51339), .I0(n18778[3]), .I1(n396_adj_5415), 
            .CO(n51340));
    SB_CARRY add_6148_18 (.CI(n51587), .I0(n14921[15]), .I1(GND_net), 
            .CO(n51588));
    SB_LUT4 add_6148_17_lut (.I0(GND_net), .I1(n14921[14]), .I2(GND_net), 
            .I3(n51586), .O(n14082[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6148_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_20_add_3_25_lut (.I0(n352[23]), .I1(GND_net), .I2(n1_adj_5683[23]), 
            .I3(n51187), .O(n47_adj_5416)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_25_lut.LUT_INIT = 16'h6996;
    SB_CARRY sub_8_add_2_13 (.CI(n51036), .I0(setpoint[11]), .I1(\motor_state[11] ), 
            .CO(n51037));
    SB_LUT4 unary_minus_20_add_3_24_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5683[22]), 
            .I3(n51186), .O(n59[22])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_8_add_2_12_lut (.I0(GND_net), .I1(setpoint[10]), .I2(\motor_state[10] ), 
            .I3(n51035), .O(n55[10])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_8_add_2_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6148_17 (.CI(n51586), .I0(n14921[14]), .I1(GND_net), 
            .CO(n51587));
    SB_LUT4 add_6148_16_lut (.I0(GND_net), .I1(n14921[13]), .I2(n1105_adj_5419), 
            .I3(n51585), .O(n14082[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6148_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_8_add_2_12 (.CI(n51035), .I0(setpoint[10]), .I1(\motor_state[10] ), 
            .CO(n51036));
    SB_CARRY add_6259_11 (.CI(n51463), .I0(n16974[8]), .I1(n749), .CO(n51464));
    SB_LUT4 add_6259_10_lut (.I0(GND_net), .I1(n16974[7]), .I2(n676), 
            .I3(n51462), .O(n16363[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6259_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6259_10 (.CI(n51462), .I0(n16974[7]), .I1(n676), .CO(n51463));
    SB_CARRY unary_minus_20_add_3_24 (.CI(n51186), .I0(GND_net), .I1(n1_adj_5683[22]), 
            .CO(n51187));
    SB_LUT4 sub_8_add_2_11_lut (.I0(GND_net), .I1(setpoint[9]), .I2(\motor_state[9] ), 
            .I3(n51034), .O(n55[9])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_8_add_2_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6379_5_lut (.I0(GND_net), .I1(n18778[2]), .I2(n323_adj_5420), 
            .I3(n51338), .O(n18415[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6379_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6379_5 (.CI(n51338), .I0(n18778[2]), .I1(n323_adj_5420), 
            .CO(n51339));
    SB_LUT4 add_6379_4_lut (.I0(GND_net), .I1(n18778[1]), .I2(n250_adj_5421), 
            .I3(n51337), .O(n18415[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6379_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_i212_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3715[7] ), 
            .I2(GND_net), .I3(GND_net), .O(n314_adj_5422));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i212_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY sub_8_add_2_11 (.CI(n51034), .I0(setpoint[9]), .I1(\motor_state[9] ), 
            .CO(n51035));
    SB_LUT4 unary_minus_20_add_3_23_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5683[21]), 
            .I3(n51185), .O(n59[21])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_23 (.CI(n51185), .I0(GND_net), .I1(n1_adj_5683[21]), 
            .CO(n51186));
    SB_LUT4 add_6259_9_lut (.I0(GND_net), .I1(n16974[6]), .I2(n603), .I3(n51461), 
            .O(n16363[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6259_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_20_add_3_22_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5683[20]), 
            .I3(n51184), .O(n59[20])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_22 (.CI(n51184), .I0(GND_net), .I1(n1_adj_5683[20]), 
            .CO(n51185));
    SB_CARRY add_6379_4 (.CI(n51337), .I0(n18778[1]), .I1(n250_adj_5421), 
            .CO(n51338));
    SB_CARRY add_6259_9 (.CI(n51461), .I0(n16974[6]), .I1(n603), .CO(n51462));
    SB_LUT4 add_6379_3_lut (.I0(GND_net), .I1(n18778[0]), .I2(n177_adj_5426), 
            .I3(n51336), .O(n18415[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6379_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6379_3 (.CI(n51336), .I0(n18778[0]), .I1(n177_adj_5426), 
            .CO(n51337));
    SB_LUT4 add_6379_2_lut (.I0(GND_net), .I1(n35_adj_5427), .I2(n104_adj_5428), 
            .I3(GND_net), .O(n18415[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6379_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6170_15 (.CI(n52626), .I0(n15359[12]), .I1(n1032), .CO(n52627));
    SB_CARRY add_6148_16 (.CI(n51585), .I0(n14921[13]), .I1(n1105_adj_5419), 
            .CO(n51586));
    SB_LUT4 sub_8_add_2_10_lut (.I0(GND_net), .I1(setpoint[8]), .I2(\motor_state[8] ), 
            .I3(n51033), .O(n55[8])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_8_add_2_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_i261_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3715[7] ), 
            .I2(GND_net), .I3(GND_net), .O(n387_adj_5429));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i261_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6170_14_lut (.I0(GND_net), .I1(n15359[11]), .I2(n959), 
            .I3(n52625), .O(n14563[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6170_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6170_14 (.CI(n52625), .I0(n15359[11]), .I1(n959), .CO(n52626));
    SB_LUT4 unary_minus_20_add_3_21_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5683[19]), 
            .I3(n51183), .O(n59[19])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6170_13_lut (.I0(GND_net), .I1(n15359[10]), .I2(n886), 
            .I3(n52624), .O(n14563[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6170_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6170_13 (.CI(n52624), .I0(n15359[10]), .I1(n886), .CO(n52625));
    SB_CARRY unary_minus_20_add_3_21 (.CI(n51183), .I0(GND_net), .I1(n1_adj_5683[19]), 
            .CO(n51184));
    SB_LUT4 unary_minus_20_add_3_20_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5683[18]), 
            .I3(n51182), .O(n59[18])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_20 (.CI(n51182), .I0(GND_net), .I1(n1_adj_5683[18]), 
            .CO(n51183));
    SB_LUT4 add_6170_12_lut (.I0(GND_net), .I1(n15359[9]), .I2(n813), 
            .I3(n52623), .O(n14563[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6170_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6379_2 (.CI(GND_net), .I0(n35_adj_5427), .I1(n104_adj_5428), 
            .CO(n51336));
    SB_LUT4 unary_minus_20_add_3_19_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5683[17]), 
            .I3(n51181), .O(n59[17])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_19 (.CI(n51181), .I0(GND_net), .I1(n1_adj_5683[17]), 
            .CO(n51182));
    SB_CARRY add_6170_12 (.CI(n52623), .I0(n15359[9]), .I1(n813), .CO(n52624));
    SB_CARRY add_6460_2 (.CI(GND_net), .I0(n44_adj_5413), .I1(n113_adj_5414), 
            .CO(n51671));
    SB_CARRY sub_8_add_2_10 (.CI(n51033), .I0(setpoint[8]), .I1(\motor_state[8] ), 
            .CO(n51034));
    SB_LUT4 add_6170_11_lut (.I0(GND_net), .I1(n15359[8]), .I2(n740), 
            .I3(n52622), .O(n14563[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6170_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6259_8_lut (.I0(GND_net), .I1(n16974[5]), .I2(n530), .I3(n51460), 
            .O(n16363[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6259_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6148_15_lut (.I0(GND_net), .I1(n14921[12]), .I2(n1032_adj_5433), 
            .I3(n51584), .O(n14082[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6148_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6259_8 (.CI(n51460), .I0(n16974[5]), .I1(n530), .CO(n51461));
    SB_CARRY add_6170_11 (.CI(n52622), .I0(n15359[8]), .I1(n740), .CO(n52623));
    SB_LUT4 sub_8_add_2_9_lut (.I0(GND_net), .I1(setpoint[7]), .I2(\motor_state[7] ), 
            .I3(n51032), .O(n55[7])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_8_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6148_15 (.CI(n51584), .I0(n14921[12]), .I1(n1032_adj_5433), 
            .CO(n51585));
    SB_LUT4 add_6170_10_lut (.I0(GND_net), .I1(n15359[7]), .I2(n667), 
            .I3(n52621), .O(n14563[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6170_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6259_7_lut (.I0(GND_net), .I1(n16974[4]), .I2(n457), .I3(n51459), 
            .O(n16363[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6259_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6170_10 (.CI(n52621), .I0(n15359[7]), .I1(n667), .CO(n52622));
    SB_CARRY sub_8_add_2_9 (.CI(n51032), .I0(setpoint[7]), .I1(\motor_state[7] ), 
            .CO(n51033));
    SB_LUT4 add_6170_9_lut (.I0(GND_net), .I1(n15359[6]), .I2(n594), .I3(n52620), 
            .O(n14563[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6170_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6259_7 (.CI(n51459), .I0(n16974[4]), .I1(n457), .CO(n51460));
    SB_CARRY add_6170_9 (.CI(n52620), .I0(n15359[6]), .I1(n594), .CO(n52621));
    SB_LUT4 add_6170_8_lut (.I0(GND_net), .I1(n15359[5]), .I2(n521), .I3(n52619), 
            .O(n14563[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6170_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6148_14_lut (.I0(GND_net), .I1(n14921[11]), .I2(n959_adj_5434), 
            .I3(n51583), .O(n14082[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6148_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_20_add_3_18_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5683[16]), 
            .I3(n51180), .O(n59[16])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6148_14 (.CI(n51583), .I0(n14921[11]), .I1(n959_adj_5434), 
            .CO(n51584));
    SB_CARRY add_6170_8 (.CI(n52619), .I0(n15359[5]), .I1(n521), .CO(n52620));
    SB_CARRY unary_minus_20_add_3_18 (.CI(n51180), .I0(GND_net), .I1(n1_adj_5683[16]), 
            .CO(n51181));
    SB_LUT4 unary_minus_20_add_3_17_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5683[15]), 
            .I3(n51179), .O(n59[15])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6259_6_lut (.I0(GND_net), .I1(n16974[3]), .I2(n384_adj_5438), 
            .I3(n51458), .O(n16363[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6259_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6170_7_lut (.I0(GND_net), .I1(n15359[4]), .I2(n448_adj_5439), 
            .I3(n52618), .O(n14563[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6170_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_8_add_2_8_lut (.I0(GND_net), .I1(setpoint[6]), .I2(n41635), 
            .I3(n51031), .O(n55[6])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_8_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6170_7 (.CI(n52618), .I0(n15359[4]), .I1(n448_adj_5439), 
            .CO(n52619));
    SB_LUT4 add_6170_6_lut (.I0(GND_net), .I1(n15359[3]), .I2(n375_adj_5440), 
            .I3(n52617), .O(n14563[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6170_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_17 (.CI(n51179), .I0(GND_net), .I1(n1_adj_5683[15]), 
            .CO(n51180));
    SB_CARRY add_6170_6 (.CI(n52617), .I0(n15359[3]), .I1(n375_adj_5440), 
            .CO(n52618));
    SB_LUT4 add_6170_5_lut (.I0(GND_net), .I1(n15359[2]), .I2(n302), .I3(n52616), 
            .O(n14563[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6170_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6259_6 (.CI(n51458), .I0(n16974[3]), .I1(n384_adj_5438), 
            .CO(n51459));
    SB_LUT4 unary_minus_20_add_3_16_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5683[14]), 
            .I3(n51178), .O(n59[14])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6170_5 (.CI(n52616), .I0(n15359[2]), .I1(n302), .CO(n52617));
    SB_LUT4 add_6170_4_lut (.I0(GND_net), .I1(n15359[1]), .I2(n229), .I3(n52615), 
            .O(n14563[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6170_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_8_add_2_8 (.CI(n51031), .I0(setpoint[6]), .I1(n41635), 
            .CO(n51032));
    SB_LUT4 sub_8_add_2_7_lut (.I0(GND_net), .I1(setpoint[5]), .I2(\motor_state[5] ), 
            .I3(n51030), .O(n55[5])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_8_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6170_4 (.CI(n52615), .I0(n15359[1]), .I1(n229), .CO(n52616));
    SB_LUT4 add_6259_5_lut (.I0(GND_net), .I1(n16974[2]), .I2(n311), .I3(n51457), 
            .O(n16363[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6259_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6170_3_lut (.I0(GND_net), .I1(n15359[0]), .I2(n156_adj_5442), 
            .I3(n52614), .O(n14563[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6170_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6170_3 (.CI(n52614), .I0(n15359[0]), .I1(n156_adj_5442), 
            .CO(n52615));
    SB_LUT4 add_6148_13_lut (.I0(GND_net), .I1(n14921[10]), .I2(n886_adj_5443), 
            .I3(n51582), .O(n14082[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6148_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6170_2_lut (.I0(GND_net), .I1(n14_adj_5444), .I2(n83), 
            .I3(GND_net), .O(n14563[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6170_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6148_13 (.CI(n51582), .I0(n14921[10]), .I1(n886_adj_5443), 
            .CO(n51583));
    SB_CARRY unary_minus_20_add_3_16 (.CI(n51178), .I0(GND_net), .I1(n1_adj_5683[14]), 
            .CO(n51179));
    SB_LUT4 add_6148_12_lut (.I0(GND_net), .I1(n14921[9]), .I2(n813_adj_5445), 
            .I3(n51581), .O(n14082[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6148_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6170_2 (.CI(GND_net), .I0(n14_adj_5444), .I1(n83), .CO(n52614));
    SB_LUT4 add_6208_20_lut (.I0(GND_net), .I1(n16077[17]), .I2(GND_net), 
            .I3(n52613), .O(n15359[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6208_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6208_19_lut (.I0(GND_net), .I1(n16077[16]), .I2(GND_net), 
            .I3(n52612), .O(n15359[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6208_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_8_add_2_7 (.CI(n51030), .I0(setpoint[5]), .I1(\motor_state[5] ), 
            .CO(n51031));
    SB_CARRY add_6148_12 (.CI(n51581), .I0(n14921[9]), .I1(n813_adj_5445), 
            .CO(n51582));
    SB_CARRY add_6259_5 (.CI(n51457), .I0(n16974[2]), .I1(n311), .CO(n51458));
    SB_CARRY add_6208_19 (.CI(n52612), .I0(n16077[16]), .I1(GND_net), 
            .CO(n52613));
    SB_LUT4 add_6148_11_lut (.I0(GND_net), .I1(n14921[8]), .I2(n740_adj_5446), 
            .I3(n51580), .O(n14082[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6148_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6208_18_lut (.I0(GND_net), .I1(n16077[15]), .I2(GND_net), 
            .I3(n52611), .O(n15359[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6208_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6259_4_lut (.I0(GND_net), .I1(n16974[1]), .I2(n238), .I3(n51456), 
            .O(n16363[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6259_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6148_11 (.CI(n51580), .I0(n14921[8]), .I1(n740_adj_5446), 
            .CO(n51581));
    SB_CARRY add_6208_18 (.CI(n52611), .I0(n16077[15]), .I1(GND_net), 
            .CO(n52612));
    SB_CARRY add_6259_4 (.CI(n51456), .I0(n16974[1]), .I1(n238), .CO(n51457));
    SB_LUT4 add_6148_10_lut (.I0(GND_net), .I1(n14921[7]), .I2(n667_adj_5447), 
            .I3(n51579), .O(n14082[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6148_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_20_add_3_15_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5683[13]), 
            .I3(n51177), .O(n59[13])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6208_17_lut (.I0(GND_net), .I1(n16077[14]), .I2(GND_net), 
            .I3(n52610), .O(n15359[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6208_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6208_17 (.CI(n52610), .I0(n16077[14]), .I1(GND_net), 
            .CO(n52611));
    SB_LUT4 sub_8_add_2_6_lut (.I0(GND_net), .I1(setpoint[4]), .I2(\motor_state[4] ), 
            .I3(n51029), .O(n55[4])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_8_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6259_3_lut (.I0(GND_net), .I1(n16974[0]), .I2(n165_adj_5449), 
            .I3(n51455), .O(n16363[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6259_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6208_16_lut (.I0(GND_net), .I1(n16077[13]), .I2(n1108_adj_5450), 
            .I3(n52609), .O(n15359[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6208_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6148_10 (.CI(n51579), .I0(n14921[7]), .I1(n667_adj_5447), 
            .CO(n51580));
    SB_CARRY add_6208_16 (.CI(n52609), .I0(n16077[13]), .I1(n1108_adj_5450), 
            .CO(n52610));
    SB_LUT4 add_6148_9_lut (.I0(GND_net), .I1(n14921[6]), .I2(n594_adj_5451), 
            .I3(n51578), .O(n14082[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6148_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6208_15_lut (.I0(GND_net), .I1(n16077[12]), .I2(n1035_adj_5452), 
            .I3(n52608), .O(n15359[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6208_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6148_9 (.CI(n51578), .I0(n14921[6]), .I1(n594_adj_5451), 
            .CO(n51579));
    SB_CARRY unary_minus_20_add_3_15 (.CI(n51177), .I0(GND_net), .I1(n1_adj_5683[13]), 
            .CO(n51178));
    SB_LUT4 add_6148_8_lut (.I0(GND_net), .I1(n14921[5]), .I2(n521_adj_5453), 
            .I3(n51577), .O(n14082[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6148_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6148_8 (.CI(n51577), .I0(n14921[5]), .I1(n521_adj_5453), 
            .CO(n51578));
    SB_CARRY add_6208_15 (.CI(n52608), .I0(n16077[12]), .I1(n1035_adj_5452), 
            .CO(n52609));
    SB_CARRY add_6259_3 (.CI(n51455), .I0(n16974[0]), .I1(n165_adj_5449), 
            .CO(n51456));
    SB_LUT4 add_6259_2_lut (.I0(GND_net), .I1(n23_adj_5454), .I2(n92), 
            .I3(GND_net), .O(n16363[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6259_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6208_14_lut (.I0(GND_net), .I1(n16077[11]), .I2(n962_adj_5455), 
            .I3(n52607), .O(n15359[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6208_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6208_14 (.CI(n52607), .I0(n16077[11]), .I1(n962_adj_5455), 
            .CO(n52608));
    SB_LUT4 add_6148_7_lut (.I0(GND_net), .I1(n14921[4]), .I2(n448_adj_5456), 
            .I3(n51576), .O(n14082[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6148_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_20_add_3_14_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5683[12]), 
            .I3(n51176), .O(n59[12])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_8_add_2_6 (.CI(n51029), .I0(setpoint[4]), .I1(\motor_state[4] ), 
            .CO(n51030));
    SB_CARRY sub_8_add_2_5 (.CI(n51028), .I0(setpoint[3]), .I1(\motor_state[3] ), 
            .CO(n51029));
    SB_CARRY unary_minus_20_add_3_14 (.CI(n51176), .I0(GND_net), .I1(n1_adj_5683[12]), 
            .CO(n51177));
    SB_CARRY add_6148_7 (.CI(n51576), .I0(n14921[4]), .I1(n448_adj_5456), 
            .CO(n51577));
    SB_CARRY add_6259_2 (.CI(GND_net), .I0(n23_adj_5454), .I1(n92), .CO(n51455));
    SB_LUT4 add_6208_13_lut (.I0(GND_net), .I1(n16077[10]), .I2(n889_adj_5459), 
            .I3(n52606), .O(n15359[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6208_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6208_13 (.CI(n52606), .I0(n16077[10]), .I1(n889_adj_5459), 
            .CO(n52607));
    SB_LUT4 mult_16_i702_2_lut (.I0(\Kp[14] ), .I1(n55[11]), .I2(GND_net), 
            .I3(GND_net), .O(n1044));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i702_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_20_add_3_13_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5683[11]), 
            .I3(n51175), .O(n59[11])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6148_6_lut (.I0(GND_net), .I1(n14921[3]), .I2(n375_adj_5461), 
            .I3(n51575), .O(n14082[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6148_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6148_6 (.CI(n51575), .I0(n14921[3]), .I1(n375_adj_5461), 
            .CO(n51576));
    SB_LUT4 add_6208_12_lut (.I0(GND_net), .I1(n16077[9]), .I2(n816_adj_5462), 
            .I3(n52605), .O(n15359[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6208_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_13 (.CI(n51175), .I0(GND_net), .I1(n1_adj_5683[11]), 
            .CO(n51176));
    SB_CARRY add_6208_12 (.CI(n52605), .I0(n16077[9]), .I1(n816_adj_5462), 
            .CO(n52606));
    SB_LUT4 add_6208_11_lut (.I0(GND_net), .I1(n16077[8]), .I2(n743_adj_5463), 
            .I3(n52604), .O(n15359[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6208_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_8_add_2_4 (.CI(n51027), .I0(setpoint[2]), .I1(\motor_state[2] ), 
            .CO(n51028));
    SB_LUT4 unary_minus_20_add_3_12_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5683[10]), 
            .I3(n51174), .O(n59[10])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_12 (.CI(n51174), .I0(GND_net), .I1(n1_adj_5683[10]), 
            .CO(n51175));
    SB_LUT4 add_6148_5_lut (.I0(GND_net), .I1(n14921[2]), .I2(n302_adj_5465), 
            .I3(n51574), .O(n14082[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6148_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6208_11 (.CI(n52604), .I0(n16077[8]), .I1(n743_adj_5463), 
            .CO(n52605));
    SB_LUT4 add_6208_10_lut (.I0(GND_net), .I1(n16077[7]), .I2(n670_adj_5466), 
            .I3(n52603), .O(n15359[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6208_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6208_10 (.CI(n52603), .I0(n16077[7]), .I1(n670_adj_5466), 
            .CO(n52604));
    SB_CARRY sub_8_add_2_3 (.CI(n51026), .I0(setpoint[1]), .I1(\motor_state[1] ), 
            .CO(n51027));
    SB_CARRY add_6148_5 (.CI(n51574), .I0(n14921[2]), .I1(n302_adj_5465), 
            .CO(n51575));
    SB_LUT4 add_6148_4_lut (.I0(GND_net), .I1(n14921[1]), .I2(n229_adj_5467), 
            .I3(n51573), .O(n14082[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6148_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6148_4 (.CI(n51573), .I0(n14921[1]), .I1(n229_adj_5467), 
            .CO(n51574));
    SB_LUT4 add_6148_3_lut (.I0(GND_net), .I1(n14921[0]), .I2(n156_adj_5468), 
            .I3(n51572), .O(n14082[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6148_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6208_9_lut (.I0(GND_net), .I1(n16077[6]), .I2(n597_adj_5469), 
            .I3(n52602), .O(n15359[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6208_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_8_add_2_2 (.CI(VCC_net), .I0(setpoint[0]), .I1(\motor_state[0] ), 
            .CO(n51026));
    SB_LUT4 unary_minus_20_add_3_11_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5683[9]), 
            .I3(n51173), .O(n59[9])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_11 (.CI(n51173), .I0(GND_net), .I1(n1_adj_5683[9]), 
            .CO(n51174));
    SB_CARRY add_6208_9 (.CI(n52602), .I0(n16077[6]), .I1(n597_adj_5469), 
            .CO(n52603));
    SB_LUT4 add_6208_8_lut (.I0(GND_net), .I1(n16077[5]), .I2(n524_adj_5472), 
            .I3(n52601), .O(n15359[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6208_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_20_add_3_10_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5683[8]), 
            .I3(n51172), .O(n59[8])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_18_25_lut (.I0(GND_net), .I1(n11637[0]), .I2(n12213[0]), 
            .I3(n51094), .O(n352[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6208_8 (.CI(n52601), .I0(n16077[5]), .I1(n524_adj_5472), 
            .CO(n52602));
    SB_LUT4 add_6208_7_lut (.I0(GND_net), .I1(n16077[4]), .I2(n451_adj_5474), 
            .I3(n52600), .O(n15359[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6208_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_10 (.CI(n51172), .I0(GND_net), .I1(n1_adj_5683[8]), 
            .CO(n51173));
    SB_LUT4 add_18_24_lut (.I0(GND_net), .I1(n257[22]), .I2(n49[22]), 
            .I3(n51093), .O(n352[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6148_3 (.CI(n51572), .I0(n14921[0]), .I1(n156_adj_5468), 
            .CO(n51573));
    SB_CARRY add_6208_7 (.CI(n52600), .I0(n16077[4]), .I1(n451_adj_5474), 
            .CO(n52601));
    SB_CARRY add_18_24 (.CI(n51093), .I0(n257[22]), .I1(n49[22]), .CO(n51094));
    SB_LUT4 add_6148_2_lut (.I0(GND_net), .I1(n14_adj_5475), .I2(n83_adj_5476), 
            .I3(GND_net), .O(n14082[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6148_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6148_2 (.CI(GND_net), .I0(n14_adj_5475), .I1(n83_adj_5476), 
            .CO(n51572));
    SB_LUT4 unary_minus_20_add_3_9_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5683[7]), 
            .I3(n51171), .O(n59[7])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_9 (.CI(n51171), .I0(GND_net), .I1(n1_adj_5683[7]), 
            .CO(n51172));
    SB_LUT4 unary_minus_20_add_3_8_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5683[6]), 
            .I3(n51170), .O(n59[6])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_8 (.CI(n51170), .I0(GND_net), .I1(n1_adj_5683[6]), 
            .CO(n51171));
    SB_LUT4 add_18_23_lut (.I0(GND_net), .I1(n257[21]), .I2(n49[21]), 
            .I3(n51092), .O(n352[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_18_23 (.CI(n51092), .I0(n257[21]), .I1(n49[21]), .CO(n51093));
    SB_LUT4 mult_17_i310_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3715[7] ), 
            .I2(GND_net), .I3(GND_net), .O(n460_adj_5480));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i310_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_20_add_3_7_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5683[5]), 
            .I3(n51169), .O(n59[5])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_18_22_lut (.I0(GND_net), .I1(n257[20]), .I2(n49[20]), 
            .I3(n51091), .O(n352[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_7 (.CI(n51169), .I0(GND_net), .I1(n1_adj_5683[5]), 
            .CO(n51170));
    SB_LUT4 unary_minus_20_add_3_6_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5683[4]), 
            .I3(n51168), .O(n59[4])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_18_22 (.CI(n51091), .I0(n257[20]), .I1(n49[20]), .CO(n51092));
    SB_LUT4 add_18_21_lut (.I0(GND_net), .I1(n257[19]), .I2(n49[19]), 
            .I3(n51090), .O(n352[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_18_21 (.CI(n51090), .I0(n257[19]), .I1(n49[19]), .CO(n51091));
    SB_CARRY unary_minus_20_add_3_6 (.CI(n51168), .I0(GND_net), .I1(n1_adj_5683[4]), 
            .CO(n51169));
    SB_LUT4 add_6208_6_lut (.I0(GND_net), .I1(n16077[3]), .I2(n378_adj_5483), 
            .I3(n52599), .O(n15359[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6208_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_20_add_3_5_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5683[3]), 
            .I3(n51167), .O(n59[3])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6208_6 (.CI(n52599), .I0(n16077[3]), .I1(n378_adj_5483), 
            .CO(n52600));
    SB_LUT4 add_6208_5_lut (.I0(GND_net), .I1(n16077[2]), .I2(n305_adj_5486), 
            .I3(n52598), .O(n15359[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6208_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6208_5 (.CI(n52598), .I0(n16077[2]), .I1(n305_adj_5486), 
            .CO(n52599));
    SB_CARRY unary_minus_20_add_3_5 (.CI(n51167), .I0(GND_net), .I1(n1_adj_5683[3]), 
            .CO(n51168));
    SB_LUT4 add_6208_4_lut (.I0(GND_net), .I1(n16077[1]), .I2(n232_adj_5487), 
            .I3(n52597), .O(n15359[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6208_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_18_20_lut (.I0(GND_net), .I1(n257[18]), .I2(n49[18]), 
            .I3(n51089), .O(n352[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6208_4 (.CI(n52597), .I0(n16077[1]), .I1(n232_adj_5487), 
            .CO(n52598));
    SB_LUT4 add_6208_3_lut (.I0(GND_net), .I1(n16077[0]), .I2(n159_adj_5488), 
            .I3(n52596), .O(n15359[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6208_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6208_3 (.CI(n52596), .I0(n16077[0]), .I1(n159_adj_5488), 
            .CO(n52597));
    SB_LUT4 add_6208_2_lut (.I0(GND_net), .I1(n17_adj_5489), .I2(n86_adj_5490), 
            .I3(GND_net), .O(n15359[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6208_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6208_2 (.CI(GND_net), .I0(n17_adj_5489), .I1(n86_adj_5490), 
            .CO(n52596));
    SB_LUT4 add_6448_11_lut (.I0(GND_net), .I1(n19571[8]), .I2(n770_adj_5491), 
            .I3(n52595), .O(n19352[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6448_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6448_10_lut (.I0(GND_net), .I1(n19571[7]), .I2(n697_adj_5492), 
            .I3(n52594), .O(n19352[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6448_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6448_10 (.CI(n52594), .I0(n19571[7]), .I1(n697_adj_5492), 
            .CO(n52595));
    SB_LUT4 add_6448_9_lut (.I0(GND_net), .I1(n19571[6]), .I2(n624_adj_5493), 
            .I3(n52593), .O(n19352[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6448_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6448_9 (.CI(n52593), .I0(n19571[6]), .I1(n624_adj_5493), 
            .CO(n52594));
    SB_LUT4 add_6448_8_lut (.I0(GND_net), .I1(n19571[5]), .I2(n551_adj_5494), 
            .I3(n52592), .O(n19352[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6448_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6448_8 (.CI(n52592), .I0(n19571[5]), .I1(n551_adj_5494), 
            .CO(n52593));
    SB_LUT4 add_6448_7_lut (.I0(GND_net), .I1(n19571[4]), .I2(n478_adj_5495), 
            .I3(n52591), .O(n19352[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6448_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6448_7 (.CI(n52591), .I0(n19571[4]), .I1(n478_adj_5495), 
            .CO(n52592));
    SB_CARRY add_18_20 (.CI(n51089), .I0(n257[18]), .I1(n49[18]), .CO(n51090));
    SB_LUT4 unary_minus_20_add_3_4_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5683[2]), 
            .I3(n51166), .O(n59[2])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6448_6_lut (.I0(GND_net), .I1(n19571[3]), .I2(n405_adj_5497), 
            .I3(n52590), .O(n19352[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6448_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6448_6 (.CI(n52590), .I0(n19571[3]), .I1(n405_adj_5497), 
            .CO(n52591));
    SB_LUT4 add_6448_5_lut (.I0(GND_net), .I1(n19571[2]), .I2(n332_adj_5498), 
            .I3(n52589), .O(n19352[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6448_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6448_5 (.CI(n52589), .I0(n19571[2]), .I1(n332_adj_5498), 
            .CO(n52590));
    SB_LUT4 mult_17_i359_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3715[7] ), 
            .I2(GND_net), .I3(GND_net), .O(n533_adj_5499));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i359_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6448_4_lut (.I0(GND_net), .I1(n19571[1]), .I2(n259_adj_5500), 
            .I3(n52588), .O(n19352[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6448_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_4 (.CI(n51166), .I0(GND_net), .I1(n1_adj_5683[2]), 
            .CO(n51167));
    SB_CARRY add_6448_4 (.CI(n52588), .I0(n19571[1]), .I1(n259_adj_5500), 
            .CO(n52589));
    SB_LUT4 add_6448_3_lut (.I0(GND_net), .I1(n19571[0]), .I2(n186_adj_5501), 
            .I3(n52587), .O(n19352[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6448_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6448_3 (.CI(n52587), .I0(n19571[0]), .I1(n186_adj_5501), 
            .CO(n52588));
    SB_LUT4 add_6448_2_lut (.I0(GND_net), .I1(n44_adj_5502), .I2(n113_adj_5503), 
            .I3(GND_net), .O(n19352[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6448_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6448_2 (.CI(GND_net), .I0(n44_adj_5502), .I1(n113_adj_5503), 
            .CO(n52587));
    SB_LUT4 add_6244_19_lut (.I0(GND_net), .I1(n16721[16]), .I2(GND_net), 
            .I3(n52586), .O(n16077[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6244_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6244_18_lut (.I0(GND_net), .I1(n16721[15]), .I2(GND_net), 
            .I3(n52585), .O(n16077[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6244_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6244_18 (.CI(n52585), .I0(n16721[15]), .I1(GND_net), 
            .CO(n52586));
    SB_LUT4 mult_17_i408_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3715[7] ), 
            .I2(GND_net), .I3(GND_net), .O(n606_adj_5504));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i408_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6244_17_lut (.I0(GND_net), .I1(n16721[14]), .I2(GND_net), 
            .I3(n52584), .O(n16077[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6244_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6244_17 (.CI(n52584), .I0(n16721[14]), .I1(GND_net), 
            .CO(n52585));
    SB_LUT4 unary_minus_20_add_3_3_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5683[1]), 
            .I3(n51165), .O(n401)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6244_16_lut (.I0(GND_net), .I1(n16721[13]), .I2(n1111_adj_5506), 
            .I3(n52583), .O(n16077[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6244_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6244_16 (.CI(n52583), .I0(n16721[13]), .I1(n1111_adj_5506), 
            .CO(n52584));
    SB_LUT4 add_6244_15_lut (.I0(GND_net), .I1(n16721[12]), .I2(n1038_adj_5507), 
            .I3(n52582), .O(n16077[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6244_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6244_15 (.CI(n52582), .I0(n16721[12]), .I1(n1038_adj_5507), 
            .CO(n52583));
    SB_LUT4 add_6244_14_lut (.I0(GND_net), .I1(n16721[11]), .I2(n965_adj_5508), 
            .I3(n52581), .O(n16077[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6244_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_i457_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3715[7] ), 
            .I2(GND_net), .I3(GND_net), .O(n679_adj_5509));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i457_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY unary_minus_20_add_3_3 (.CI(n51165), .I0(GND_net), .I1(n1_adj_5683[1]), 
            .CO(n51166));
    SB_CARRY add_6244_14 (.CI(n52581), .I0(n16721[11]), .I1(n965_adj_5508), 
            .CO(n52582));
    SB_LUT4 add_6244_13_lut (.I0(GND_net), .I1(n16721[10]), .I2(n892_adj_5510), 
            .I3(n52580), .O(n16077[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6244_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6244_13 (.CI(n52580), .I0(n16721[10]), .I1(n892_adj_5510), 
            .CO(n52581));
    SB_LUT4 add_6244_12_lut (.I0(GND_net), .I1(n16721[9]), .I2(n819_adj_5511), 
            .I3(n52579), .O(n16077[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6244_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6244_12 (.CI(n52579), .I0(n16721[9]), .I1(n819_adj_5511), 
            .CO(n52580));
    SB_LUT4 add_6244_11_lut (.I0(GND_net), .I1(n16721[8]), .I2(n746_adj_5512), 
            .I3(n52578), .O(n16077[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6244_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6244_11 (.CI(n52578), .I0(n16721[8]), .I1(n746_adj_5512), 
            .CO(n52579));
    SB_LUT4 unary_minus_20_add_3_2_lut (.I0(n37313), .I1(GND_net), .I2(n1_adj_5683[0]), 
            .I3(VCC_net), .O(n33)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_2_lut.LUT_INIT = 16'h8228;
    SB_LUT4 add_6244_10_lut (.I0(GND_net), .I1(n16721[7]), .I2(n673_adj_5515), 
            .I3(n52577), .O(n16077[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6244_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6244_10 (.CI(n52577), .I0(n16721[7]), .I1(n673_adj_5515), 
            .CO(n52578));
    SB_LUT4 add_6244_9_lut (.I0(GND_net), .I1(n16721[6]), .I2(n600_adj_5516), 
            .I3(n52576), .O(n16077[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6244_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_18_19_lut (.I0(GND_net), .I1(n257[17]), .I2(n49[17]), 
            .I3(n51088), .O(n352[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6244_9 (.CI(n52576), .I0(n16721[6]), .I1(n600_adj_5516), 
            .CO(n52577));
    SB_LUT4 add_6244_8_lut (.I0(GND_net), .I1(n16721[5]), .I2(n527_adj_5517), 
            .I3(n52575), .O(n16077[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6244_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6244_8 (.CI(n52575), .I0(n16721[5]), .I1(n527_adj_5517), 
            .CO(n52576));
    SB_LUT4 add_6244_7_lut (.I0(GND_net), .I1(n16721[4]), .I2(n454_adj_5518), 
            .I3(n52574), .O(n16077[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6244_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_18_19 (.CI(n51088), .I0(n257[17]), .I1(n49[17]), .CO(n51089));
    SB_CARRY add_6244_7 (.CI(n52574), .I0(n16721[4]), .I1(n454_adj_5518), 
            .CO(n52575));
    SB_LUT4 add_6244_6_lut (.I0(GND_net), .I1(n16721[3]), .I2(n381_adj_5519), 
            .I3(n52573), .O(n16077[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6244_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6244_6 (.CI(n52573), .I0(n16721[3]), .I1(n381_adj_5519), 
            .CO(n52574));
    SB_CARRY unary_minus_20_add_3_2 (.CI(VCC_net), .I0(GND_net), .I1(n1_adj_5683[0]), 
            .CO(n51165));
    SB_LUT4 add_6244_5_lut (.I0(GND_net), .I1(n16721[2]), .I2(n308_adj_5520), 
            .I3(n52572), .O(n16077[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6244_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6244_5 (.CI(n52572), .I0(n16721[2]), .I1(n308_adj_5520), 
            .CO(n52573));
    SB_LUT4 add_18_18_lut (.I0(GND_net), .I1(n257[16]), .I2(n49[16]), 
            .I3(n51087), .O(n352[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6244_4_lut (.I0(GND_net), .I1(n16721[1]), .I2(n235_adj_5521), 
            .I3(n52571), .O(n16077[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6244_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6244_4 (.CI(n52571), .I0(n16721[1]), .I1(n235_adj_5521), 
            .CO(n52572));
    SB_LUT4 add_6244_3_lut (.I0(GND_net), .I1(n16721[0]), .I2(n162_adj_5522), 
            .I3(n52570), .O(n16077[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6244_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_13_add_3_25_lut (.I0(GND_net), .I1(GND_net), .I2(n1[23]), 
            .I3(n51164), .O(n182[23])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_18_18 (.CI(n51087), .I0(n257[16]), .I1(n49[16]), .CO(n51088));
    SB_CARRY add_6244_3 (.CI(n52570), .I0(n16721[0]), .I1(n162_adj_5522), 
            .CO(n52571));
    SB_LUT4 add_6244_2_lut (.I0(GND_net), .I1(n20_adj_5524), .I2(n89_adj_5525), 
            .I3(GND_net), .O(n16077[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6244_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6244_2 (.CI(GND_net), .I0(n20_adj_5524), .I1(n89_adj_5525), 
            .CO(n52570));
    SB_LUT4 add_6278_18_lut (.I0(GND_net), .I1(n17295[15]), .I2(GND_net), 
            .I3(n52569), .O(n16721[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6278_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6278_17_lut (.I0(GND_net), .I1(n17295[14]), .I2(GND_net), 
            .I3(n52568), .O(n16721[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6278_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6278_17 (.CI(n52568), .I0(n17295[14]), .I1(GND_net), 
            .CO(n52569));
    SB_LUT4 unary_minus_13_add_3_24_lut (.I0(GND_net), .I1(GND_net), .I2(n1[22]), 
            .I3(n51163), .O(n182[22])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6278_16_lut (.I0(GND_net), .I1(n17295[13]), .I2(n1114_adj_5527), 
            .I3(n52567), .O(n16721[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6278_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6278_16 (.CI(n52567), .I0(n17295[13]), .I1(n1114_adj_5527), 
            .CO(n52568));
    SB_CARRY unary_minus_13_add_3_24 (.CI(n51163), .I0(GND_net), .I1(n1[22]), 
            .CO(n51164));
    SB_LUT4 add_6278_15_lut (.I0(GND_net), .I1(n17295[12]), .I2(n1041_adj_5528), 
            .I3(n52566), .O(n16721[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6278_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6278_15 (.CI(n52566), .I0(n17295[12]), .I1(n1041_adj_5528), 
            .CO(n52567));
    SB_LUT4 add_6278_14_lut (.I0(GND_net), .I1(n17295[11]), .I2(n968_adj_5529), 
            .I3(n52565), .O(n16721[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6278_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6278_14 (.CI(n52565), .I0(n17295[11]), .I1(n968_adj_5529), 
            .CO(n52566));
    SB_LUT4 add_6278_13_lut (.I0(GND_net), .I1(n17295[10]), .I2(n895_adj_5530), 
            .I3(n52564), .O(n16721[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6278_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6278_13 (.CI(n52564), .I0(n17295[10]), .I1(n895_adj_5530), 
            .CO(n52565));
    SB_LUT4 add_6278_12_lut (.I0(GND_net), .I1(n17295[9]), .I2(n822_adj_5531), 
            .I3(n52563), .O(n16721[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6278_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_13_add_3_23_lut (.I0(GND_net), .I1(GND_net), .I2(n1[21]), 
            .I3(n51162), .O(n182[21])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_13_add_3_23 (.CI(n51162), .I0(GND_net), .I1(n1[21]), 
            .CO(n51163));
    SB_CARRY add_6278_12 (.CI(n52563), .I0(n17295[9]), .I1(n822_adj_5531), 
            .CO(n52564));
    SB_LUT4 add_6278_11_lut (.I0(GND_net), .I1(n17295[8]), .I2(n749_adj_5533), 
            .I3(n52562), .O(n16721[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6278_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6278_11 (.CI(n52562), .I0(n17295[8]), .I1(n749_adj_5533), 
            .CO(n52563));
    SB_LUT4 add_6278_10_lut (.I0(GND_net), .I1(n17295[7]), .I2(n676_adj_5534), 
            .I3(n52561), .O(n16721[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6278_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_i506_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3715[7] ), 
            .I2(GND_net), .I3(GND_net), .O(n752_adj_5535));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i506_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_13_add_3_22_lut (.I0(GND_net), .I1(GND_net), .I2(n1[20]), 
            .I3(n51161), .O(n182[20])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6278_10 (.CI(n52561), .I0(n17295[7]), .I1(n676_adj_5534), 
            .CO(n52562));
    SB_LUT4 add_6278_9_lut (.I0(GND_net), .I1(n17295[6]), .I2(n603_adj_5537), 
            .I3(n52560), .O(n16721[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6278_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_18_17_lut (.I0(GND_net), .I1(n257[15]), .I2(n49[15]), 
            .I3(n51086), .O(n361)) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6278_9 (.CI(n52560), .I0(n17295[6]), .I1(n603_adj_5537), 
            .CO(n52561));
    SB_LUT4 add_6278_8_lut (.I0(GND_net), .I1(n17295[5]), .I2(n530_adj_5538), 
            .I3(n52559), .O(n16721[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6278_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6278_8 (.CI(n52559), .I0(n17295[5]), .I1(n530_adj_5538), 
            .CO(n52560));
    SB_CARRY unary_minus_13_add_3_22 (.CI(n51161), .I0(GND_net), .I1(n1[20]), 
            .CO(n51162));
    SB_CARRY add_18_17 (.CI(n51086), .I0(n257[15]), .I1(n49[15]), .CO(n51087));
    SB_LUT4 add_6278_7_lut (.I0(GND_net), .I1(n17295[4]), .I2(n457_adj_5539), 
            .I3(n52558), .O(n16721[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6278_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_13_add_3_21_lut (.I0(GND_net), .I1(GND_net), .I2(n1[19]), 
            .I3(n51160), .O(n182[19])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6278_7 (.CI(n52558), .I0(n17295[4]), .I1(n457_adj_5539), 
            .CO(n52559));
    SB_LUT4 add_6278_6_lut (.I0(GND_net), .I1(n17295[3]), .I2(n384_adj_5541), 
            .I3(n52557), .O(n16721[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6278_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_18_16_lut (.I0(GND_net), .I1(n257[14]), .I2(n49[14]), 
            .I3(n51085), .O(n352[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6278_6 (.CI(n52557), .I0(n17295[3]), .I1(n384_adj_5541), 
            .CO(n52558));
    SB_LUT4 add_6278_5_lut (.I0(GND_net), .I1(n17295[2]), .I2(n311_adj_5542), 
            .I3(n52556), .O(n16721[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6278_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_18_16 (.CI(n51085), .I0(n257[14]), .I1(n49[14]), .CO(n51086));
    SB_CARRY add_6278_5 (.CI(n52556), .I0(n17295[2]), .I1(n311_adj_5542), 
            .CO(n52557));
    SB_LUT4 mult_17_i555_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3715[7] ), 
            .I2(GND_net), .I3(GND_net), .O(n825_adj_5543));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i555_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i604_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3715[7] ), 
            .I2(GND_net), .I3(GND_net), .O(n898_adj_5544));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i604_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i653_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3715[7] ), 
            .I2(GND_net), .I3(GND_net), .O(n971_adj_5545));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i653_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i702_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3715[7] ), 
            .I2(GND_net), .I3(GND_net), .O(n1044_adj_5546));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i702_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6278_4_lut (.I0(GND_net), .I1(n17295[1]), .I2(n238_adj_5547), 
            .I3(n52555), .O(n16721[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6278_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6278_4 (.CI(n52555), .I0(n17295[1]), .I1(n238_adj_5547), 
            .CO(n52556));
    SB_LUT4 add_6278_3_lut (.I0(GND_net), .I1(n17295[0]), .I2(n165_adj_5548), 
            .I3(n52554), .O(n16721[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6278_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6278_3 (.CI(n52554), .I0(n17295[0]), .I1(n165_adj_5548), 
            .CO(n52555));
    SB_LUT4 add_6278_2_lut (.I0(GND_net), .I1(n23_adj_5549), .I2(n92_adj_5550), 
            .I3(GND_net), .O(n16721[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6278_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6278_2 (.CI(GND_net), .I0(n23_adj_5549), .I1(n92_adj_5550), 
            .CO(n52554));
    SB_LUT4 add_6467_10_lut (.I0(GND_net), .I1(n19750[7]), .I2(n700), 
            .I3(n52553), .O(n19571[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6467_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6467_9_lut (.I0(GND_net), .I1(n19750[6]), .I2(n627_adj_5551), 
            .I3(n52552), .O(n19571[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6467_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6467_9 (.CI(n52552), .I0(n19750[6]), .I1(n627_adj_5551), 
            .CO(n52553));
    SB_LUT4 mult_17_i751_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3715[7] ), 
            .I2(GND_net), .I3(GND_net), .O(n1117));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i751_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6292_17_lut (.I0(GND_net), .I1(n17517[14]), .I2(GND_net), 
            .I3(n51439), .O(n16974[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6292_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6467_8_lut (.I0(GND_net), .I1(n19750[5]), .I2(n554_adj_5552), 
            .I3(n52551), .O(n19571[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6467_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6478_10_lut (.I0(GND_net), .I1(n19847[7]), .I2(n700_adj_5553), 
            .I3(n51553), .O(n19689[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6478_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6467_8 (.CI(n52551), .I0(n19750[5]), .I1(n554_adj_5552), 
            .CO(n52552));
    SB_LUT4 add_6467_7_lut (.I0(GND_net), .I1(n19750[4]), .I2(n481_adj_5554), 
            .I3(n52550), .O(n19571[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6467_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6467_7 (.CI(n52550), .I0(n19750[4]), .I1(n481_adj_5554), 
            .CO(n52551));
    SB_LUT4 add_6467_6_lut (.I0(GND_net), .I1(n19750[3]), .I2(n408_adj_5555), 
            .I3(n52549), .O(n19571[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6467_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i79_2_lut (.I0(\Kp[1] ), .I1(n55[18]), .I2(GND_net), 
            .I3(GND_net), .O(n116_adj_5556));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i79_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i32_2_lut (.I0(\Kp[0] ), .I1(n55[19]), .I2(GND_net), 
            .I3(GND_net), .O(n47_adj_5557));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i32_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6467_6 (.CI(n52549), .I0(n19750[3]), .I1(n408_adj_5555), 
            .CO(n52550));
    SB_LUT4 add_6467_5_lut (.I0(GND_net), .I1(n19750[2]), .I2(n335_adj_5558), 
            .I3(n52548), .O(n19571[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6467_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i128_2_lut (.I0(\Kp[2] ), .I1(n55[18]), .I2(GND_net), 
            .I3(GND_net), .O(n189_adj_5559));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i128_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i751_2_lut (.I0(\Kp[15] ), .I1(n55[11]), .I2(GND_net), 
            .I3(GND_net), .O(n1117_adj_5560));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i751_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i177_2_lut (.I0(\Kp[3] ), .I1(n55[18]), .I2(GND_net), 
            .I3(GND_net), .O(n262_adj_5561));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i177_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i226_2_lut (.I0(\Kp[4] ), .I1(n55[18]), .I2(GND_net), 
            .I3(GND_net), .O(n335_adj_5558));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i226_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i275_2_lut (.I0(\Kp[5] ), .I1(n55[18]), .I2(GND_net), 
            .I3(GND_net), .O(n408_adj_5555));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i275_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i324_2_lut (.I0(\Kp[6] ), .I1(n55[18]), .I2(GND_net), 
            .I3(GND_net), .O(n481_adj_5554));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i324_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6467_5 (.CI(n52548), .I0(n19750[2]), .I1(n335_adj_5558), 
            .CO(n52549));
    SB_LUT4 add_6467_4_lut (.I0(GND_net), .I1(n19750[1]), .I2(n262_adj_5561), 
            .I3(n52547), .O(n19571[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6467_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_i471_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3715[14] ), 
            .I2(GND_net), .I3(GND_net), .O(n700_adj_5553));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i471_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i373_2_lut (.I0(\Kp[7] ), .I1(n55[18]), .I2(GND_net), 
            .I3(GND_net), .O(n554_adj_5552));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i373_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i422_2_lut (.I0(\Kp[8] ), .I1(n55[18]), .I2(GND_net), 
            .I3(GND_net), .O(n627_adj_5551));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i422_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6467_4 (.CI(n52547), .I0(n19750[1]), .I1(n262_adj_5561), 
            .CO(n52548));
    SB_LUT4 mult_16_i471_2_lut (.I0(\Kp[9] ), .I1(n55[18]), .I2(GND_net), 
            .I3(GND_net), .O(n700));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i471_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6292_16_lut (.I0(GND_net), .I1(n17517[13]), .I2(n1117_adj_5560), 
            .I3(n51438), .O(n16974[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6292_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6467_3_lut (.I0(GND_net), .I1(n19750[0]), .I2(n189_adj_5559), 
            .I3(n52546), .O(n19571[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6467_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6467_3 (.CI(n52546), .I0(n19750[0]), .I1(n189_adj_5559), 
            .CO(n52547));
    SB_LUT4 add_6467_2_lut (.I0(GND_net), .I1(n47_adj_5557), .I2(n116_adj_5556), 
            .I3(GND_net), .O(n19571[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6467_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6467_2 (.CI(GND_net), .I0(n47_adj_5557), .I1(n116_adj_5556), 
            .CO(n52546));
    SB_LUT4 add_6310_17_lut (.I0(GND_net), .I1(n17803[14]), .I2(GND_net), 
            .I3(n52545), .O(n17295[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6310_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6310_16_lut (.I0(GND_net), .I1(n17803[13]), .I2(n1117), 
            .I3(n52544), .O(n17295[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6310_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6310_16 (.CI(n52544), .I0(n17803[13]), .I1(n1117), .CO(n52545));
    SB_LUT4 add_6310_15_lut (.I0(GND_net), .I1(n17803[12]), .I2(n1044_adj_5546), 
            .I3(n52543), .O(n17295[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6310_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6310_15 (.CI(n52543), .I0(n17803[12]), .I1(n1044_adj_5546), 
            .CO(n52544));
    SB_LUT4 add_6310_14_lut (.I0(GND_net), .I1(n17803[11]), .I2(n971_adj_5545), 
            .I3(n52542), .O(n17295[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6310_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6310_14 (.CI(n52542), .I0(n17803[11]), .I1(n971_adj_5545), 
            .CO(n52543));
    SB_LUT4 add_6310_13_lut (.I0(GND_net), .I1(n17803[10]), .I2(n898_adj_5544), 
            .I3(n52541), .O(n17295[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6310_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6310_13 (.CI(n52541), .I0(n17803[10]), .I1(n898_adj_5544), 
            .CO(n52542));
    SB_LUT4 add_6310_12_lut (.I0(GND_net), .I1(n17803[9]), .I2(n825_adj_5543), 
            .I3(n52540), .O(n17295[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6310_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6310_12 (.CI(n52540), .I0(n17803[9]), .I1(n825_adj_5543), 
            .CO(n52541));
    SB_LUT4 add_6310_11_lut (.I0(GND_net), .I1(n17803[8]), .I2(n752_adj_5535), 
            .I3(n52539), .O(n17295[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6310_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6310_11 (.CI(n52539), .I0(n17803[8]), .I1(n752_adj_5535), 
            .CO(n52540));
    SB_LUT4 add_6310_10_lut (.I0(GND_net), .I1(n17803[7]), .I2(n679_adj_5509), 
            .I3(n52538), .O(n17295[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6310_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6310_10 (.CI(n52538), .I0(n17803[7]), .I1(n679_adj_5509), 
            .CO(n52539));
    SB_LUT4 mult_17_i63_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3715[6] ), 
            .I2(GND_net), .I3(GND_net), .O(n92_adj_5550));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i63_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i16_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3715[7] ), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_5549));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i16_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i112_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3715[6] ), 
            .I2(GND_net), .I3(GND_net), .O(n165_adj_5548));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i112_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6310_9_lut (.I0(GND_net), .I1(n17803[6]), .I2(n606_adj_5504), 
            .I3(n52537), .O(n17295[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6310_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_i161_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3715[6] ), 
            .I2(GND_net), .I3(GND_net), .O(n238_adj_5547));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i161_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i210_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3715[6] ), 
            .I2(GND_net), .I3(GND_net), .O(n311_adj_5542));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i210_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i259_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3715[6] ), 
            .I2(GND_net), .I3(GND_net), .O(n384_adj_5541));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i259_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6310_9 (.CI(n52537), .I0(n17803[6]), .I1(n606_adj_5504), 
            .CO(n52538));
    SB_LUT4 unary_minus_13_inv_0_i20_1_lut (.I0(IntegralLimit[19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[19]));   // verilog/motorControl.v(49[22:36])
    defparam unary_minus_13_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_6310_8_lut (.I0(GND_net), .I1(n17803[5]), .I2(n533_adj_5499), 
            .I3(n52536), .O(n17295[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6310_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6310_8 (.CI(n52536), .I0(n17803[5]), .I1(n533_adj_5499), 
            .CO(n52537));
    SB_LUT4 add_6310_7_lut (.I0(GND_net), .I1(n17803[4]), .I2(n460_adj_5480), 
            .I3(n52535), .O(n17295[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6310_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_i308_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3715[6] ), 
            .I2(GND_net), .I3(GND_net), .O(n457_adj_5539));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i308_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6292_16 (.CI(n51438), .I0(n17517[13]), .I1(n1117_adj_5560), 
            .CO(n51439));
    SB_CARRY add_6310_7 (.CI(n52535), .I0(n17803[4]), .I1(n460_adj_5480), 
            .CO(n52536));
    SB_LUT4 add_6292_15_lut (.I0(GND_net), .I1(n17517[12]), .I2(n1044), 
            .I3(n51437), .O(n16974[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6292_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6310_6_lut (.I0(GND_net), .I1(n17803[3]), .I2(n387_adj_5429), 
            .I3(n52534), .O(n17295[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6310_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6310_6 (.CI(n52534), .I0(n17803[3]), .I1(n387_adj_5429), 
            .CO(n52535));
    SB_LUT4 add_6310_5_lut (.I0(GND_net), .I1(n17803[2]), .I2(n314_adj_5422), 
            .I3(n52533), .O(n17295[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6310_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6310_5 (.CI(n52533), .I0(n17803[2]), .I1(n314_adj_5422), 
            .CO(n52534));
    SB_LUT4 add_6310_4_lut (.I0(GND_net), .I1(n17803[1]), .I2(n241_adj_5411), 
            .I3(n52532), .O(n17295[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6310_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6478_9_lut (.I0(GND_net), .I1(n19847[6]), .I2(n627), .I3(n51552), 
            .O(n19689[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6478_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6292_15 (.CI(n51437), .I0(n17517[12]), .I1(n1044), .CO(n51438));
    SB_LUT4 mult_17_i357_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3715[6] ), 
            .I2(GND_net), .I3(GND_net), .O(n530_adj_5538));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i357_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i406_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3715[6] ), 
            .I2(GND_net), .I3(GND_net), .O(n603_adj_5537));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i406_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_13_inv_0_i21_1_lut (.I0(IntegralLimit[20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[20]));   // verilog/motorControl.v(49[22:36])
    defparam unary_minus_13_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_6310_4 (.CI(n52532), .I0(n17803[1]), .I1(n241_adj_5411), 
            .CO(n52533));
    SB_LUT4 add_6310_3_lut (.I0(GND_net), .I1(n17803[0]), .I2(n168_adj_5377), 
            .I3(n52531), .O(n17295[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6310_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6478_9 (.CI(n51552), .I0(n19847[6]), .I1(n627), .CO(n51553));
    SB_CARRY add_6310_3 (.CI(n52531), .I0(n17803[0]), .I1(n168_adj_5377), 
            .CO(n52532));
    SB_LUT4 add_6310_2_lut (.I0(GND_net), .I1(n26_adj_5373), .I2(n95_adj_5364), 
            .I3(GND_net), .O(n17295[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6310_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6310_2 (.CI(GND_net), .I0(n26_adj_5373), .I1(n95_adj_5364), 
            .CO(n52531));
    SB_LUT4 add_6340_16_lut (.I0(GND_net), .I1(n18249[13]), .I2(n1120_adj_5358), 
            .I3(n52530), .O(n17803[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6340_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6340_15_lut (.I0(GND_net), .I1(n18249[12]), .I2(n1047_adj_5330), 
            .I3(n52529), .O(n17803[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6340_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6478_8_lut (.I0(GND_net), .I1(n19847[5]), .I2(n554), .I3(n51551), 
            .O(n19689[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6478_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6292_14_lut (.I0(GND_net), .I1(n17517[11]), .I2(n971), 
            .I3(n51436), .O(n16974[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6292_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6292_14 (.CI(n51436), .I0(n17517[11]), .I1(n971), .CO(n51437));
    SB_CARRY add_6340_15 (.CI(n52529), .I0(n18249[12]), .I1(n1047_adj_5330), 
            .CO(n52530));
    SB_LUT4 add_6340_14_lut (.I0(GND_net), .I1(n18249[11]), .I2(n974_adj_5317), 
            .I3(n52528), .O(n17803[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6340_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6292_13_lut (.I0(GND_net), .I1(n17517[10]), .I2(n898), 
            .I3(n51435), .O(n16974[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6292_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6340_14 (.CI(n52528), .I0(n18249[11]), .I1(n974_adj_5317), 
            .CO(n52529));
    SB_LUT4 add_6340_13_lut (.I0(GND_net), .I1(n18249[10]), .I2(n901_adj_5316), 
            .I3(n52527), .O(n17803[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6340_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6478_8 (.CI(n51551), .I0(n19847[5]), .I1(n554), .CO(n51552));
    SB_CARRY add_6340_13 (.CI(n52527), .I0(n18249[10]), .I1(n901_adj_5316), 
            .CO(n52528));
    SB_LUT4 add_6340_12_lut (.I0(GND_net), .I1(n18249[9]), .I2(n828_adj_5315), 
            .I3(n52526), .O(n17803[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6340_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6340_12 (.CI(n52526), .I0(n18249[9]), .I1(n828_adj_5315), 
            .CO(n52527));
    SB_LUT4 add_6478_7_lut (.I0(GND_net), .I1(n19847[4]), .I2(n481), .I3(n51550), 
            .O(n19689[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6478_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6340_11_lut (.I0(GND_net), .I1(n18249[8]), .I2(n755_adj_5313), 
            .I3(n52525), .O(n17803[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6340_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6292_13 (.CI(n51435), .I0(n17517[10]), .I1(n898), .CO(n51436));
    SB_CARRY add_6340_11 (.CI(n52525), .I0(n18249[8]), .I1(n755_adj_5313), 
            .CO(n52526));
    SB_LUT4 add_6340_10_lut (.I0(GND_net), .I1(n18249[7]), .I2(n682_adj_5310), 
            .I3(n52524), .O(n17803[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6340_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6340_10 (.CI(n52524), .I0(n18249[7]), .I1(n682_adj_5310), 
            .CO(n52525));
    SB_CARRY unary_minus_13_add_3_21 (.CI(n51160), .I0(GND_net), .I1(n1[19]), 
            .CO(n51161));
    SB_LUT4 add_6292_12_lut (.I0(GND_net), .I1(n17517[9]), .I2(n825), 
            .I3(n51434), .O(n16974[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6292_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6340_9_lut (.I0(GND_net), .I1(n18249[6]), .I2(n609_adj_5309), 
            .I3(n52523), .O(n17803[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6340_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6340_9 (.CI(n52523), .I0(n18249[6]), .I1(n609_adj_5309), 
            .CO(n52524));
    SB_CARRY add_6292_12 (.CI(n51434), .I0(n17517[9]), .I1(n825), .CO(n51435));
    SB_LUT4 add_6340_8_lut (.I0(GND_net), .I1(n18249[5]), .I2(n536_adj_5308), 
            .I3(n52522), .O(n17803[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6340_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6292_11_lut (.I0(GND_net), .I1(n17517[8]), .I2(n752), 
            .I3(n51433), .O(n16974[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6292_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6340_8 (.CI(n52522), .I0(n18249[5]), .I1(n536_adj_5308), 
            .CO(n52523));
    SB_LUT4 add_6340_7_lut (.I0(GND_net), .I1(n18249[4]), .I2(n463_adj_5307), 
            .I3(n52521), .O(n17803[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6340_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6340_7 (.CI(n52521), .I0(n18249[4]), .I1(n463_adj_5307), 
            .CO(n52522));
    SB_LUT4 add_6340_6_lut (.I0(GND_net), .I1(n18249[3]), .I2(n390_adj_5306), 
            .I3(n52520), .O(n17803[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6340_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6037_23_lut (.I0(GND_net), .I1(n13158[20]), .I2(GND_net), 
            .I3(n51650), .O(n12096[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6037_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6340_6 (.CI(n52520), .I0(n18249[3]), .I1(n390_adj_5306), 
            .CO(n52521));
    SB_LUT4 add_6340_5_lut (.I0(GND_net), .I1(n18249[2]), .I2(n317_adj_5305), 
            .I3(n52519), .O(n17803[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6340_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6478_7 (.CI(n51550), .I0(n19847[4]), .I1(n481), .CO(n51551));
    SB_CARRY add_6340_5 (.CI(n52519), .I0(n18249[2]), .I1(n317_adj_5305), 
            .CO(n52520));
    SB_LUT4 add_6340_4_lut (.I0(GND_net), .I1(n18249[1]), .I2(n244_adj_5304), 
            .I3(n52518), .O(n17803[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6340_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6340_4 (.CI(n52518), .I0(n18249[1]), .I1(n244_adj_5304), 
            .CO(n52519));
    SB_CARRY add_6292_11 (.CI(n51433), .I0(n17517[8]), .I1(n752), .CO(n51434));
    SB_LUT4 add_6340_3_lut (.I0(GND_net), .I1(n18249[0]), .I2(n171_adj_5303), 
            .I3(n52517), .O(n17803[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6340_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6340_3 (.CI(n52517), .I0(n18249[0]), .I1(n171_adj_5303), 
            .CO(n52518));
    SB_LUT4 add_6292_10_lut (.I0(GND_net), .I1(n17517[7]), .I2(n679), 
            .I3(n51432), .O(n16974[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6292_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6340_2_lut (.I0(GND_net), .I1(n29_adj_5302), .I2(n98_adj_5301), 
            .I3(GND_net), .O(n17803[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6340_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6340_2 (.CI(GND_net), .I0(n29_adj_5302), .I1(n98_adj_5301), 
            .CO(n52517));
    SB_LUT4 add_6484_9_lut (.I0(GND_net), .I1(n19893[6]), .I2(n630_adj_5300), 
            .I3(n52516), .O(n19750[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6484_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6478_6_lut (.I0(GND_net), .I1(n19847[3]), .I2(n408), .I3(n51549), 
            .O(n19689[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6478_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6484_8_lut (.I0(GND_net), .I1(n19893[5]), .I2(n557_adj_5299), 
            .I3(n52515), .O(n19750[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6484_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6484_8 (.CI(n52515), .I0(n19893[5]), .I1(n557_adj_5299), 
            .CO(n52516));
    SB_LUT4 add_6484_7_lut (.I0(GND_net), .I1(n19893[4]), .I2(n484_adj_5298), 
            .I3(n52514), .O(n19750[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6484_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6484_7 (.CI(n52514), .I0(n19893[4]), .I1(n484_adj_5298), 
            .CO(n52515));
    SB_LUT4 add_6484_6_lut (.I0(GND_net), .I1(n19893[3]), .I2(n411_adj_5297), 
            .I3(n52513), .O(n19750[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6484_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6484_6 (.CI(n52513), .I0(n19893[3]), .I1(n411_adj_5297), 
            .CO(n52514));
    SB_LUT4 unary_minus_13_add_3_20_lut (.I0(GND_net), .I1(GND_net), .I2(n1[18]), 
            .I3(n51159), .O(n182[18])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6484_5_lut (.I0(GND_net), .I1(n19893[2]), .I2(n338_adj_5295), 
            .I3(n52512), .O(n19750[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6484_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6484_5 (.CI(n52512), .I0(n19893[2]), .I1(n338_adj_5295), 
            .CO(n52513));
    SB_LUT4 add_6484_4_lut (.I0(GND_net), .I1(n19893[1]), .I2(n265), .I3(n52511), 
            .O(n19750[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6484_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6292_10 (.CI(n51432), .I0(n17517[7]), .I1(n679), .CO(n51433));
    SB_LUT4 mult_17_i455_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3715[6] ), 
            .I2(GND_net), .I3(GND_net), .O(n676_adj_5534));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i455_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i504_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3715[6] ), 
            .I2(GND_net), .I3(GND_net), .O(n749_adj_5533));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i504_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6484_4 (.CI(n52511), .I0(n19893[1]), .I1(n265), .CO(n52512));
    SB_LUT4 add_6484_3_lut (.I0(GND_net), .I1(n19893[0]), .I2(n192_adj_5294), 
            .I3(n52510), .O(n19750[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6484_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6484_3 (.CI(n52510), .I0(n19893[0]), .I1(n192_adj_5294), 
            .CO(n52511));
    SB_LUT4 unary_minus_13_inv_0_i22_1_lut (.I0(IntegralLimit[21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[21]));   // verilog/motorControl.v(49[22:36])
    defparam unary_minus_13_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_16_i641_2_lut (.I0(\Kp[13] ), .I1(n55[5]), .I2(GND_net), 
            .I3(GND_net), .O(n953));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i641_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6484_2_lut (.I0(GND_net), .I1(n50_adj_5293), .I2(n119_adj_5292), 
            .I3(GND_net), .O(n19750[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6484_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6484_2 (.CI(GND_net), .I0(n50_adj_5293), .I1(n119_adj_5292), 
            .CO(n52510));
    SB_LUT4 mult_17_i553_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3715[6] ), 
            .I2(GND_net), .I3(GND_net), .O(n822_adj_5531));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i553_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i602_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3715[6] ), 
            .I2(GND_net), .I3(GND_net), .O(n895_adj_5530));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i602_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i598_2_lut (.I0(\Kp[12] ), .I1(n55[8]), .I2(GND_net), 
            .I3(GND_net), .O(n889));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i598_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6368_15_lut (.I0(GND_net), .I1(n18637[12]), .I2(n1050_adj_5291), 
            .I3(n52509), .O(n18249[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6368_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6368_14_lut (.I0(GND_net), .I1(n18637[11]), .I2(n977_adj_5290), 
            .I3(n52508), .O(n18249[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6368_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_13_inv_0_i12_1_lut (.I0(IntegralLimit[11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[11]));   // verilog/motorControl.v(49[22:36])
    defparam unary_minus_13_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_13_inv_0_i13_1_lut (.I0(IntegralLimit[12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[12]));   // verilog/motorControl.v(49[22:36])
    defparam unary_minus_13_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_17_i651_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3715[6] ), 
            .I2(GND_net), .I3(GND_net), .O(n968_adj_5529));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i651_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i647_2_lut (.I0(\Kp[13] ), .I1(n55[8]), .I2(GND_net), 
            .I3(GND_net), .O(n962));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i647_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i700_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3715[6] ), 
            .I2(GND_net), .I3(GND_net), .O(n1041_adj_5528));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i700_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i749_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3715[6] ), 
            .I2(GND_net), .I3(GND_net), .O(n1114_adj_5527));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i749_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_13_inv_0_i23_1_lut (.I0(IntegralLimit[22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[22]));   // verilog/motorControl.v(49[22:36])
    defparam unary_minus_13_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_13_inv_0_i14_1_lut (.I0(IntegralLimit[13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[13]));   // verilog/motorControl.v(49[22:36])
    defparam unary_minus_13_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_6368_14 (.CI(n52508), .I0(n18637[11]), .I1(n977_adj_5290), 
            .CO(n52509));
    SB_LUT4 mult_16_i696_2_lut (.I0(\Kp[14] ), .I1(n55[8]), .I2(GND_net), 
            .I3(GND_net), .O(n1035));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i696_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i690_2_lut (.I0(\Kp[14] ), .I1(n55[5]), .I2(GND_net), 
            .I3(GND_net), .O(n1026));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i690_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6368_13_lut (.I0(GND_net), .I1(n18637[10]), .I2(n904_adj_5289), 
            .I3(n52507), .O(n18249[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6368_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6368_13 (.CI(n52507), .I0(n18637[10]), .I1(n904_adj_5289), 
            .CO(n52508));
    SB_LUT4 add_6368_12_lut (.I0(GND_net), .I1(n18637[9]), .I2(n831_adj_5288), 
            .I3(n52506), .O(n18249[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6368_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6368_12 (.CI(n52506), .I0(n18637[9]), .I1(n831_adj_5288), 
            .CO(n52507));
    SB_LUT4 add_6368_11_lut (.I0(GND_net), .I1(n18637[8]), .I2(n758_adj_5287), 
            .I3(n52505), .O(n18249[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6368_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6368_11 (.CI(n52505), .I0(n18637[8]), .I1(n758_adj_5287), 
            .CO(n52506));
    SB_LUT4 add_6368_10_lut (.I0(GND_net), .I1(n18637[7]), .I2(n685_adj_5286), 
            .I3(n52504), .O(n18249[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6368_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_i61_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3715[5] ), 
            .I2(GND_net), .I3(GND_net), .O(n89_adj_5525));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i61_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i14_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3715[6] ), 
            .I2(GND_net), .I3(GND_net), .O(n20_adj_5524));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i14_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6368_10 (.CI(n52504), .I0(n18637[7]), .I1(n685_adj_5286), 
            .CO(n52505));
    SB_LUT4 add_6368_9_lut (.I0(GND_net), .I1(n18637[6]), .I2(n612_adj_5285), 
            .I3(n52503), .O(n18249[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6368_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6368_9 (.CI(n52503), .I0(n18637[6]), .I1(n612_adj_5285), 
            .CO(n52504));
    SB_LUT4 add_6368_8_lut (.I0(GND_net), .I1(n18637[5]), .I2(n539_adj_5284), 
            .I3(n52502), .O(n18249[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6368_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6368_8 (.CI(n52502), .I0(n18637[5]), .I1(n539_adj_5284), 
            .CO(n52503));
    SB_LUT4 add_6368_7_lut (.I0(GND_net), .I1(n18637[4]), .I2(n466_adj_5283), 
            .I3(n52501), .O(n18249[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6368_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6368_7 (.CI(n52501), .I0(n18637[4]), .I1(n466_adj_5283), 
            .CO(n52502));
    SB_LUT4 unary_minus_13_inv_0_i24_1_lut (.I0(IntegralLimit[23]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[23]));   // verilog/motorControl.v(49[22:36])
    defparam unary_minus_13_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_6368_6_lut (.I0(GND_net), .I1(n18637[3]), .I2(n393_adj_5282), 
            .I3(n52500), .O(n18249[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6368_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6368_6 (.CI(n52500), .I0(n18637[3]), .I1(n393_adj_5282), 
            .CO(n52501));
    SB_LUT4 add_6368_5_lut (.I0(GND_net), .I1(n18637[2]), .I2(n320_adj_5281), 
            .I3(n52499), .O(n18249[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6368_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6368_5 (.CI(n52499), .I0(n18637[2]), .I1(n320_adj_5281), 
            .CO(n52500));
    SB_LUT4 add_6368_4_lut (.I0(GND_net), .I1(n18637[1]), .I2(n247_adj_5280), 
            .I3(n52498), .O(n18249[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6368_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_i110_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3715[5] ), 
            .I2(GND_net), .I3(GND_net), .O(n162_adj_5522));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i110_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i159_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3715[5] ), 
            .I2(GND_net), .I3(GND_net), .O(n235_adj_5521));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i159_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6368_4 (.CI(n52498), .I0(n18637[1]), .I1(n247_adj_5280), 
            .CO(n52499));
    SB_LUT4 add_6368_3_lut (.I0(GND_net), .I1(n18637[0]), .I2(n174_adj_5279), 
            .I3(n52497), .O(n18249[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6368_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6368_3 (.CI(n52497), .I0(n18637[0]), .I1(n174_adj_5279), 
            .CO(n52498));
    SB_LUT4 mult_17_i208_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3715[5] ), 
            .I2(GND_net), .I3(GND_net), .O(n308_adj_5520));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i208_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6037_22_lut (.I0(GND_net), .I1(n13158[19]), .I2(GND_net), 
            .I3(n51649), .O(n12096[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6037_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_i257_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3715[5] ), 
            .I2(GND_net), .I3(GND_net), .O(n381_adj_5519));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i257_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i306_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3715[5] ), 
            .I2(GND_net), .I3(GND_net), .O(n454_adj_5518));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i306_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i355_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3715[5] ), 
            .I2(GND_net), .I3(GND_net), .O(n527_adj_5517));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i355_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6478_6 (.CI(n51549), .I0(n19847[3]), .I1(n408), .CO(n51550));
    SB_LUT4 add_6292_9_lut (.I0(GND_net), .I1(n17517[6]), .I2(n606), .I3(n51431), 
            .O(n16974[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6292_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6037_22 (.CI(n51649), .I0(n13158[19]), .I1(GND_net), 
            .CO(n51650));
    SB_LUT4 add_6368_2_lut (.I0(GND_net), .I1(n32_adj_5278), .I2(n101_adj_5277), 
            .I3(GND_net), .O(n18249[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6368_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6368_2 (.CI(GND_net), .I0(n32_adj_5278), .I1(n101_adj_5277), 
            .CO(n52497));
    SB_LUT4 mult_17_i404_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3715[5] ), 
            .I2(GND_net), .I3(GND_net), .O(n600_adj_5516));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i404_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6394_14_lut (.I0(GND_net), .I1(n18971[11]), .I2(n980), 
            .I3(n52496), .O(n18637[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6394_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6394_13_lut (.I0(GND_net), .I1(n18971[10]), .I2(n907), 
            .I3(n52495), .O(n18637[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6394_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6394_13 (.CI(n52495), .I0(n18971[10]), .I1(n907), .CO(n52496));
    SB_LUT4 add_6037_21_lut (.I0(GND_net), .I1(n13158[18]), .I2(GND_net), 
            .I3(n51648), .O(n12096[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6037_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6394_12_lut (.I0(GND_net), .I1(n18971[9]), .I2(n834), 
            .I3(n52494), .O(n18637[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6394_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6478_5_lut (.I0(GND_net), .I1(n19847[2]), .I2(n335), .I3(n51548), 
            .O(n19689[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6478_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6394_12 (.CI(n52494), .I0(n18971[9]), .I1(n834), .CO(n52495));
    SB_CARRY add_6478_5 (.CI(n51548), .I0(n19847[2]), .I1(n335), .CO(n51549));
    SB_CARRY add_6292_9 (.CI(n51431), .I0(n17517[6]), .I1(n606), .CO(n51432));
    SB_LUT4 add_6394_11_lut (.I0(GND_net), .I1(n18971[8]), .I2(n761), 
            .I3(n52493), .O(n18637[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6394_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6292_8_lut (.I0(GND_net), .I1(n17517[5]), .I2(n533), .I3(n51430), 
            .O(n16974[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6292_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_13_add_3_20 (.CI(n51159), .I0(GND_net), .I1(n1[18]), 
            .CO(n51160));
    SB_LUT4 add_18_15_lut (.I0(GND_net), .I1(n257[13]), .I2(n49[13]), 
            .I3(n51084), .O(n352[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6292_8 (.CI(n51430), .I0(n17517[5]), .I1(n533), .CO(n51431));
    SB_CARRY add_6394_11 (.CI(n52493), .I0(n18971[8]), .I1(n761), .CO(n52494));
    SB_LUT4 add_6394_10_lut (.I0(GND_net), .I1(n18971[7]), .I2(n688), 
            .I3(n52492), .O(n18637[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6394_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_13_add_3_19_lut (.I0(GND_net), .I1(GND_net), .I2(n1[17]), 
            .I3(n51158), .O(n182[17])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_18_15 (.CI(n51084), .I0(n257[13]), .I1(n49[13]), .CO(n51085));
    SB_CARRY add_6394_10 (.CI(n52492), .I0(n18971[7]), .I1(n688), .CO(n52493));
    SB_LUT4 add_6394_9_lut (.I0(GND_net), .I1(n18971[6]), .I2(n615), .I3(n52491), 
            .O(n18637[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6394_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_13_add_3_19 (.CI(n51158), .I0(GND_net), .I1(n1[17]), 
            .CO(n51159));
    SB_CARRY add_6394_9 (.CI(n52491), .I0(n18971[6]), .I1(n615), .CO(n52492));
    SB_LUT4 add_6478_4_lut (.I0(GND_net), .I1(n19847[1]), .I2(n262), .I3(n51547), 
            .O(n19689[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6478_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6394_8_lut (.I0(GND_net), .I1(n18971[5]), .I2(n542), .I3(n52490), 
            .O(n18637[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6394_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6394_8 (.CI(n52490), .I0(n18971[5]), .I1(n542), .CO(n52491));
    SB_LUT4 add_6394_7_lut (.I0(GND_net), .I1(n18971[4]), .I2(n469), .I3(n52489), 
            .O(n18637[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6394_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6292_7_lut (.I0(GND_net), .I1(n17517[4]), .I2(n460), .I3(n51429), 
            .O(n16974[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6292_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_i453_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3715[5] ), 
            .I2(GND_net), .I3(GND_net), .O(n673_adj_5515));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i453_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i23360_1_lut (.I0(n376), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n37313));   // verilog/motorControl.v(51[18:38])
    defparam i23360_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_6394_7 (.CI(n52489), .I0(n18971[4]), .I1(n469), .CO(n52490));
    SB_LUT4 add_6394_6_lut (.I0(GND_net), .I1(n18971[3]), .I2(n396), .I3(n52488), 
            .O(n18637[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6394_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6394_6 (.CI(n52488), .I0(n18971[3]), .I1(n396), .CO(n52489));
    SB_LUT4 add_6394_5_lut (.I0(GND_net), .I1(n18971[2]), .I2(n323), .I3(n52487), 
            .O(n18637[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6394_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6394_5 (.CI(n52487), .I0(n18971[2]), .I1(n323), .CO(n52488));
    SB_LUT4 add_6394_4_lut (.I0(GND_net), .I1(n18971[1]), .I2(n250), .I3(n52486), 
            .O(n18637[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6394_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i745_2_lut (.I0(\Kp[15] ), .I1(n55[8]), .I2(GND_net), 
            .I3(GND_net), .O(n1108));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i745_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6394_4 (.CI(n52486), .I0(n18971[1]), .I1(n250), .CO(n52487));
    SB_LUT4 add_6394_3_lut (.I0(GND_net), .I1(n18971[0]), .I2(n177), .I3(n52485), 
            .O(n18637[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6394_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6394_3 (.CI(n52485), .I0(n18971[0]), .I1(n177), .CO(n52486));
    SB_LUT4 add_6394_2_lut (.I0(GND_net), .I1(n35_adj_5270), .I2(n104), 
            .I3(GND_net), .O(n18637[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6394_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6394_2 (.CI(GND_net), .I0(n35_adj_5270), .I1(n104), .CO(n52485));
    SB_LUT4 add_6499_8_lut (.I0(GND_net), .I1(n20004[5]), .I2(n560_adj_5267), 
            .I3(n52484), .O(n19893[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6499_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6499_7_lut (.I0(GND_net), .I1(n20004[4]), .I2(n487_adj_5266), 
            .I3(n52483), .O(n19893[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6499_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6499_7 (.CI(n52483), .I0(n20004[4]), .I1(n487_adj_5266), 
            .CO(n52484));
    SB_LUT4 unary_minus_20_inv_0_i1_1_lut (.I0(deadband[0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5683[0]));   // verilog/motorControl.v(52[43:52])
    defparam unary_minus_20_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_6499_6_lut (.I0(GND_net), .I1(n20004[3]), .I2(n414_adj_5265), 
            .I3(n52482), .O(n19893[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6499_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_i502_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3715[5] ), 
            .I2(GND_net), .I3(GND_net), .O(n746_adj_5512));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i502_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6499_6 (.CI(n52482), .I0(n20004[3]), .I1(n414_adj_5265), 
            .CO(n52483));
    SB_LUT4 mult_17_i551_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3715[5] ), 
            .I2(GND_net), .I3(GND_net), .O(n819_adj_5511));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i551_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6499_5_lut (.I0(GND_net), .I1(n20004[2]), .I2(n341_adj_5264), 
            .I3(n52481), .O(n19893[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6499_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6499_5 (.CI(n52481), .I0(n20004[2]), .I1(n341_adj_5264), 
            .CO(n52482));
    SB_LUT4 add_6499_4_lut (.I0(GND_net), .I1(n20004[1]), .I2(n268_adj_5263), 
            .I3(n52480), .O(n19893[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6499_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6499_4 (.CI(n52480), .I0(n20004[1]), .I1(n268_adj_5263), 
            .CO(n52481));
    SB_LUT4 add_6499_3_lut (.I0(GND_net), .I1(n20004[0]), .I2(n195_adj_5262), 
            .I3(n52479), .O(n19893[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6499_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6499_3 (.CI(n52479), .I0(n20004[0]), .I1(n195_adj_5262), 
            .CO(n52480));
    SB_CARRY add_6037_21 (.CI(n51648), .I0(n13158[18]), .I1(GND_net), 
            .CO(n51649));
    SB_LUT4 add_6499_2_lut (.I0(GND_net), .I1(n53_adj_5261), .I2(n122_adj_5260), 
            .I3(GND_net), .O(n19893[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6499_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6499_2 (.CI(GND_net), .I0(n53_adj_5261), .I1(n122_adj_5260), 
            .CO(n52479));
    SB_LUT4 add_6418_13_lut (.I0(GND_net), .I1(n19255[10]), .I2(n910_adj_5259), 
            .I3(n52478), .O(n18971[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6418_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6418_12_lut (.I0(GND_net), .I1(n19255[9]), .I2(n837_adj_5258), 
            .I3(n52477), .O(n18971[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6418_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_i600_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3715[5] ), 
            .I2(GND_net), .I3(GND_net), .O(n892_adj_5510));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i600_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6418_12 (.CI(n52477), .I0(n19255[9]), .I1(n837_adj_5258), 
            .CO(n52478));
    SB_LUT4 mult_16_i739_2_lut (.I0(\Kp[15] ), .I1(n55[5]), .I2(GND_net), 
            .I3(GND_net), .O(n1099));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i739_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i649_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3715[5] ), 
            .I2(GND_net), .I3(GND_net), .O(n965_adj_5508));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i649_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i698_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3715[5] ), 
            .I2(GND_net), .I3(GND_net), .O(n1038_adj_5507));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i698_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6418_11_lut (.I0(GND_net), .I1(n19255[8]), .I2(n764_adj_5243), 
            .I3(n52476), .O(n18971[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6418_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6418_11 (.CI(n52476), .I0(n19255[8]), .I1(n764_adj_5243), 
            .CO(n52477));
    SB_LUT4 add_6418_10_lut (.I0(GND_net), .I1(n19255[7]), .I2(n691_adj_5242), 
            .I3(n52475), .O(n18971[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6418_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6418_10 (.CI(n52475), .I0(n19255[7]), .I1(n691_adj_5242), 
            .CO(n52476));
    SB_LUT4 mult_17_i747_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3715[5] ), 
            .I2(GND_net), .I3(GND_net), .O(n1111_adj_5506));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i747_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_20_inv_0_i2_1_lut (.I0(deadband[1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5683[1]));   // verilog/motorControl.v(52[43:52])
    defparam unary_minus_20_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_6418_9_lut (.I0(GND_net), .I1(n19255[6]), .I2(n618_adj_5241), 
            .I3(n52474), .O(n18971[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6418_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6418_9 (.CI(n52474), .I0(n19255[6]), .I1(n618_adj_5241), 
            .CO(n52475));
    SB_LUT4 add_6418_8_lut (.I0(GND_net), .I1(n19255[5]), .I2(n545_adj_5240), 
            .I3(n52473), .O(n18971[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6418_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6418_8 (.CI(n52473), .I0(n19255[5]), .I1(n545_adj_5240), 
            .CO(n52474));
    SB_LUT4 add_6418_7_lut (.I0(GND_net), .I1(n19255[4]), .I2(n472_adj_5239), 
            .I3(n52472), .O(n18971[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6418_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6418_7 (.CI(n52472), .I0(n19255[4]), .I1(n472_adj_5239), 
            .CO(n52473));
    SB_LUT4 add_6418_6_lut (.I0(GND_net), .I1(n19255[3]), .I2(n399_adj_5238), 
            .I3(n52471), .O(n18971[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6418_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6418_6 (.CI(n52471), .I0(n19255[3]), .I1(n399_adj_5238), 
            .CO(n52472));
    SB_LUT4 add_6418_5_lut (.I0(GND_net), .I1(n19255[2]), .I2(n326_adj_5237), 
            .I3(n52470), .O(n18971[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6418_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6292_7 (.CI(n51429), .I0(n17517[4]), .I1(n460), .CO(n51430));
    SB_CARRY add_6418_5 (.CI(n52470), .I0(n19255[2]), .I1(n326_adj_5237), 
            .CO(n52471));
    SB_LUT4 add_6418_4_lut (.I0(GND_net), .I1(n19255[1]), .I2(n253_adj_5236), 
            .I3(n52469), .O(n18971[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6418_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6418_4 (.CI(n52469), .I0(n19255[1]), .I1(n253_adj_5236), 
            .CO(n52470));
    SB_LUT4 add_6418_3_lut (.I0(GND_net), .I1(n19255[0]), .I2(n180_adj_5235), 
            .I3(n52468), .O(n18971[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6418_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6418_3 (.CI(n52468), .I0(n19255[0]), .I1(n180_adj_5235), 
            .CO(n52469));
    SB_LUT4 add_6418_2_lut (.I0(GND_net), .I1(n38), .I2(n107_adj_5234), 
            .I3(GND_net), .O(n18971[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6418_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6418_2 (.CI(GND_net), .I0(n38), .I1(n107_adj_5234), .CO(n52468));
    SB_LUT4 add_6440_12_lut (.I0(GND_net), .I1(n19493[9]), .I2(n840_adj_5233), 
            .I3(n52467), .O(n19255[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6440_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6440_11_lut (.I0(GND_net), .I1(n19493[8]), .I2(n767_adj_5231), 
            .I3(n52466), .O(n19255[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6440_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6440_11 (.CI(n52466), .I0(n19493[8]), .I1(n767_adj_5231), 
            .CO(n52467));
    SB_LUT4 add_6440_10_lut (.I0(GND_net), .I1(n19493[7]), .I2(n694_adj_5230), 
            .I3(n52465), .O(n19255[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6440_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6440_10 (.CI(n52465), .I0(n19493[7]), .I1(n694_adj_5230), 
            .CO(n52466));
    SB_LUT4 add_6440_9_lut (.I0(GND_net), .I1(n19493[6]), .I2(n621_adj_5229), 
            .I3(n52464), .O(n19255[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6440_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6440_9 (.CI(n52464), .I0(n19493[6]), .I1(n621_adj_5229), 
            .CO(n52465));
    SB_LUT4 add_6292_6_lut (.I0(GND_net), .I1(n17517[3]), .I2(n387), .I3(n51428), 
            .O(n16974[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6292_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6440_8_lut (.I0(GND_net), .I1(n19493[5]), .I2(n548_adj_5228), 
            .I3(n52463), .O(n19255[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6440_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6440_8 (.CI(n52463), .I0(n19493[5]), .I1(n548_adj_5228), 
            .CO(n52464));
    SB_LUT4 add_6440_7_lut (.I0(GND_net), .I1(n19493[4]), .I2(n475_adj_5227), 
            .I3(n52462), .O(n19255[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6440_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6440_7 (.CI(n52462), .I0(n19493[4]), .I1(n475_adj_5227), 
            .CO(n52463));
    SB_LUT4 add_6440_6_lut (.I0(GND_net), .I1(n19493[3]), .I2(n402_adj_5226), 
            .I3(n52461), .O(n19255[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6440_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6440_6 (.CI(n52461), .I0(n19493[3]), .I1(n402_adj_5226), 
            .CO(n52462));
    SB_LUT4 add_6440_5_lut (.I0(GND_net), .I1(n19493[2]), .I2(n329_adj_5225), 
            .I3(n52460), .O(n19255[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6440_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6037_20_lut (.I0(GND_net), .I1(n13158[17]), .I2(GND_net), 
            .I3(n51647), .O(n12096[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6037_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6440_5 (.CI(n52460), .I0(n19493[2]), .I1(n329_adj_5225), 
            .CO(n52461));
    SB_LUT4 add_6440_4_lut (.I0(GND_net), .I1(n19493[1]), .I2(n256_adj_5223), 
            .I3(n52459), .O(n19255[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6440_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6440_4 (.CI(n52459), .I0(n19493[1]), .I1(n256_adj_5223), 
            .CO(n52460));
    SB_LUT4 add_6440_3_lut (.I0(GND_net), .I1(n19493[0]), .I2(n183_adj_5222), 
            .I3(n52458), .O(n19255[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6440_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i77_2_lut (.I0(\Kp[1] ), .I1(n55[17]), .I2(GND_net), 
            .I3(GND_net), .O(n113_adj_5503));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i77_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6440_3 (.CI(n52458), .I0(n19493[0]), .I1(n183_adj_5222), 
            .CO(n52459));
    SB_LUT4 add_6440_2_lut (.I0(GND_net), .I1(n41_adj_5221), .I2(n110), 
            .I3(GND_net), .O(n19255[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6440_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6440_2 (.CI(GND_net), .I0(n41_adj_5221), .I1(n110), .CO(n52458));
    SB_LUT4 mult_16_i30_2_lut (.I0(\Kp[0] ), .I1(n55[18]), .I2(GND_net), 
            .I3(GND_net), .O(n44_adj_5502));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i30_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6037_20 (.CI(n51647), .I0(n13158[17]), .I1(GND_net), 
            .CO(n51648));
    SB_CARRY add_6478_4 (.CI(n51547), .I0(n19847[1]), .I1(n262), .CO(n51548));
    SB_LUT4 mult_16_i126_2_lut (.I0(\Kp[2] ), .I1(n55[17]), .I2(GND_net), 
            .I3(GND_net), .O(n186_adj_5501));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i126_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i175_2_lut (.I0(\Kp[3] ), .I1(n55[17]), .I2(GND_net), 
            .I3(GND_net), .O(n259_adj_5500));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i175_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i224_2_lut (.I0(\Kp[4] ), .I1(n55[17]), .I2(GND_net), 
            .I3(GND_net), .O(n332_adj_5498));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i224_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_18_14_lut (.I0(GND_net), .I1(n257[12]), .I2(n49[12]), 
            .I3(n51083), .O(n352[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6037_19_lut (.I0(GND_net), .I1(n13158[16]), .I2(GND_net), 
            .I3(n51646), .O(n12096[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6037_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i273_2_lut (.I0(\Kp[5] ), .I1(n55[17]), .I2(GND_net), 
            .I3(GND_net), .O(n405_adj_5497));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i273_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6292_6 (.CI(n51428), .I0(n17517[3]), .I1(n387), .CO(n51429));
    SB_LUT4 add_6478_3_lut (.I0(GND_net), .I1(n19847[0]), .I2(n189), .I3(n51546), 
            .O(n19689[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6478_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6037_19 (.CI(n51646), .I0(n13158[16]), .I1(GND_net), 
            .CO(n51647));
    SB_LUT4 unary_minus_20_inv_0_i3_1_lut (.I0(deadband[2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5683[2]));   // verilog/motorControl.v(52[43:52])
    defparam unary_minus_20_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_16_i322_2_lut (.I0(\Kp[6] ), .I1(n55[17]), .I2(GND_net), 
            .I3(GND_net), .O(n478_adj_5495));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i322_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i371_2_lut (.I0(\Kp[7] ), .I1(n55[17]), .I2(GND_net), 
            .I3(GND_net), .O(n551_adj_5494));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i371_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i420_2_lut (.I0(\Kp[8] ), .I1(n55[17]), .I2(GND_net), 
            .I3(GND_net), .O(n624_adj_5493));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i420_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6292_5_lut (.I0(GND_net), .I1(n17517[2]), .I2(n314), .I3(n51427), 
            .O(n16974[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6292_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i469_2_lut (.I0(\Kp[9] ), .I1(n55[17]), .I2(GND_net), 
            .I3(GND_net), .O(n697_adj_5492));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i469_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i518_2_lut (.I0(\Kp[10] ), .I1(n55[17]), .I2(GND_net), 
            .I3(GND_net), .O(n770_adj_5491));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i518_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i59_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3715[4] ), 
            .I2(GND_net), .I3(GND_net), .O(n86_adj_5490));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i59_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i12_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3715[5] ), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_5489));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i12_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i108_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3715[4] ), 
            .I2(GND_net), .I3(GND_net), .O(n159_adj_5488));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i108_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i51502_3_lut_4_lut (.I0(n130[3]), .I1(n182[3]), .I2(n182[2]), 
            .I3(n130[2]), .O(n67196));   // verilog/motorControl.v(48[21:44])
    defparam i51502_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 LessThan_12_i6_3_lut_3_lut (.I0(n130[3]), .I1(n182[3]), .I2(n182[2]), 
            .I3(GND_net), .O(n6_c));   // verilog/motorControl.v(48[21:44])
    defparam LessThan_12_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 mult_17_i157_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3715[4] ), 
            .I2(GND_net), .I3(GND_net), .O(n232_adj_5487));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i157_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i206_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3715[4] ), 
            .I2(GND_net), .I3(GND_net), .O(n305_adj_5486));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i206_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_20_inv_0_i4_1_lut (.I0(deadband[3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5683[3]));   // verilog/motorControl.v(52[43:52])
    defparam unary_minus_20_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_17_i255_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3715[4] ), 
            .I2(GND_net), .I3(GND_net), .O(n378_adj_5483));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i255_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_20_inv_0_i5_1_lut (.I0(deadband[4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5683[4]));   // verilog/motorControl.v(52[43:52])
    defparam unary_minus_20_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_20_inv_0_i6_1_lut (.I0(deadband[5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5683[5]));   // verilog/motorControl.v(52[43:52])
    defparam unary_minus_20_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_20_inv_0_i7_1_lut (.I0(deadband[6]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5683[6]));   // verilog/motorControl.v(52[43:52])
    defparam unary_minus_20_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_20_inv_0_i8_1_lut (.I0(deadband[7]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5683[7]));   // verilog/motorControl.v(52[43:52])
    defparam unary_minus_20_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_16_i57_2_lut (.I0(\Kp[1] ), .I1(n55[7]), .I2(GND_net), 
            .I3(GND_net), .O(n83_adj_5476));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i57_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i10_2_lut (.I0(\Kp[0] ), .I1(n55[8]), .I2(GND_net), 
            .I3(GND_net), .O(n14_adj_5475));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i10_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i304_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3715[4] ), 
            .I2(GND_net), .I3(GND_net), .O(n451_adj_5474));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i304_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_20_inv_0_i9_1_lut (.I0(deadband[8]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5683[8]));   // verilog/motorControl.v(52[43:52])
    defparam unary_minus_20_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_17_i353_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3715[4] ), 
            .I2(GND_net), .I3(GND_net), .O(n524_adj_5472));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i353_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_20_inv_0_i10_1_lut (.I0(deadband[9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5683[9]));   // verilog/motorControl.v(52[43:52])
    defparam unary_minus_20_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_17_i402_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3715[4] ), 
            .I2(GND_net), .I3(GND_net), .O(n597_adj_5469));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i402_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i106_2_lut (.I0(\Kp[2] ), .I1(n55[7]), .I2(GND_net), 
            .I3(GND_net), .O(n156_adj_5468));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i106_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i155_2_lut (.I0(\Kp[3] ), .I1(n55[7]), .I2(GND_net), 
            .I3(GND_net), .O(n229_adj_5467));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i155_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i52258_2_lut_4_lut (.I0(deadband[21]), .I1(n352[21]), .I2(deadband[9]), 
            .I3(n367), .O(n67952));
    defparam i52258_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 mult_17_i451_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3715[4] ), 
            .I2(GND_net), .I3(GND_net), .O(n670_adj_5466));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i451_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i204_2_lut (.I0(\Kp[4] ), .I1(n55[7]), .I2(GND_net), 
            .I3(GND_net), .O(n302_adj_5465));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i204_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_20_inv_0_i11_1_lut (.I0(deadband[10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5683[10]));   // verilog/motorControl.v(52[43:52])
    defparam unary_minus_20_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_17_i500_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3715[4] ), 
            .I2(GND_net), .I3(GND_net), .O(n743_adj_5463));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i500_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i549_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3715[4] ), 
            .I2(GND_net), .I3(GND_net), .O(n816_adj_5462));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i549_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i253_2_lut (.I0(\Kp[5] ), .I1(n55[7]), .I2(GND_net), 
            .I3(GND_net), .O(n375_adj_5461));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i253_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_20_inv_0_i12_1_lut (.I0(deadband[11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5683[11]));   // verilog/motorControl.v(52[43:52])
    defparam unary_minus_20_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_17_i598_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3715[4] ), 
            .I2(GND_net), .I3(GND_net), .O(n889_adj_5459));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i598_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_20_inv_0_i13_1_lut (.I0(deadband[12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5683[12]));   // verilog/motorControl.v(52[43:52])
    defparam unary_minus_20_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_16_i302_2_lut (.I0(\Kp[6] ), .I1(n55[7]), .I2(GND_net), 
            .I3(GND_net), .O(n448_adj_5456));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i302_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i647_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3715[4] ), 
            .I2(GND_net), .I3(GND_net), .O(n962_adj_5455));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i647_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i52268_2_lut_4_lut (.I0(deadband[16]), .I1(n352[16]), .I2(deadband[7]), 
            .I3(n352[7]), .O(n67962));
    defparam i52268_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 mult_16_i63_2_lut (.I0(\Kp[1] ), .I1(n55[10]), .I2(GND_net), 
            .I3(GND_net), .O(n92));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i63_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i16_2_lut (.I0(\Kp[0] ), .I1(n55[11]), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_5454));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i16_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i351_2_lut (.I0(\Kp[7] ), .I1(n55[7]), .I2(GND_net), 
            .I3(GND_net), .O(n521_adj_5453));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i351_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i696_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3715[4] ), 
            .I2(GND_net), .I3(GND_net), .O(n1035_adj_5452));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i696_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i400_2_lut (.I0(\Kp[8] ), .I1(n55[7]), .I2(GND_net), 
            .I3(GND_net), .O(n594_adj_5451));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i400_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i745_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3715[4] ), 
            .I2(GND_net), .I3(GND_net), .O(n1108_adj_5450));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i745_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i112_2_lut (.I0(\Kp[2] ), .I1(n55[10]), .I2(GND_net), 
            .I3(GND_net), .O(n165_adj_5449));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i112_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_20_inv_0_i14_1_lut (.I0(deadband[13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5683[13]));   // verilog/motorControl.v(52[43:52])
    defparam unary_minus_20_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_16_i449_2_lut (.I0(\Kp[9] ), .I1(n55[7]), .I2(GND_net), 
            .I3(GND_net), .O(n667_adj_5447));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i449_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i161_2_lut (.I0(\Kp[3] ), .I1(n55[10]), .I2(GND_net), 
            .I3(GND_net), .O(n238));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i161_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i498_2_lut (.I0(\Kp[10] ), .I1(n55[7]), .I2(GND_net), 
            .I3(GND_net), .O(n740_adj_5446));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i498_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i547_2_lut (.I0(\Kp[11] ), .I1(n55[7]), .I2(GND_net), 
            .I3(GND_net), .O(n813_adj_5445));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i547_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i57_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3715[3] ), 
            .I2(GND_net), .I3(GND_net), .O(n83));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i57_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i10_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3715[4] ), 
            .I2(GND_net), .I3(GND_net), .O(n14_adj_5444));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i10_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i51800_3_lut_4_lut (.I0(IntegralLimit[3]), .I1(n130[3]), .I2(n130[2]), 
            .I3(IntegralLimit[2]), .O(n67494));   // verilog/motorControl.v(46[12:34])
    defparam i51800_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 mult_16_i596_2_lut (.I0(\Kp[12] ), .I1(n55[7]), .I2(GND_net), 
            .I3(GND_net), .O(n886_adj_5443));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i596_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_10_i6_3_lut_3_lut (.I0(IntegralLimit[3]), .I1(n130[3]), 
            .I2(n130[2]), .I3(GND_net), .O(n6_adj_5564));   // verilog/motorControl.v(46[12:34])
    defparam LessThan_10_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 mult_17_i106_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3715[3] ), 
            .I2(GND_net), .I3(GND_net), .O(n156_adj_5442));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i106_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i210_2_lut (.I0(\Kp[4] ), .I1(n55[10]), .I2(GND_net), 
            .I3(GND_net), .O(n311));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i210_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i37005_2_lut_3_lut_4_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3715[21] ), 
            .I2(\PID_CONTROLLER.integral_23__N_3715[20] ), .I3(\Ki[1] ), 
            .O(n20207[0]));   // verilog/motorControl.v(51[27:38])
    defparam i37005_2_lut_3_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 mult_17_i155_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3715[3] ), 
            .I2(GND_net), .I3(GND_net), .O(n229));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i155_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_20_inv_0_i15_1_lut (.I0(deadband[14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5683[14]));   // verilog/motorControl.v(52[43:52])
    defparam unary_minus_20_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i37007_2_lut_3_lut_4_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3715[21] ), 
            .I2(\PID_CONTROLLER.integral_23__N_3715[20] ), .I3(\Ki[1] ), 
            .O(n50890));   // verilog/motorControl.v(51[27:38])
    defparam i37007_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 mult_17_i204_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3715[3] ), 
            .I2(GND_net), .I3(GND_net), .O(n302));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i204_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i253_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3715[3] ), 
            .I2(GND_net), .I3(GND_net), .O(n375_adj_5440));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i253_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i302_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3715[3] ), 
            .I2(GND_net), .I3(GND_net), .O(n448_adj_5439));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i302_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i259_2_lut (.I0(\Kp[5] ), .I1(n55[10]), .I2(GND_net), 
            .I3(GND_net), .O(n384_adj_5438));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i259_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_20_inv_0_i16_1_lut (.I0(deadband[15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5683[15]));   // verilog/motorControl.v(52[43:52])
    defparam unary_minus_20_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_16_i69_2_lut (.I0(\Kp[1] ), .I1(n55[13]), .I2(GND_net), 
            .I3(GND_net), .O(n101));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i69_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i22_2_lut (.I0(\Kp[0] ), .I1(n55[14]), .I2(GND_net), 
            .I3(GND_net), .O(n32_adj_5275));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i22_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i5954_2_lut_4_lut (.I0(control_update), .I1(n69824), .I2(PWMLimit[23]), 
            .I3(n352[23]), .O(n11595));
    defparam i5954_2_lut_4_lut.LUT_INIT = 16'h2a02;
    SB_LUT4 unary_minus_20_inv_0_i17_1_lut (.I0(deadband[16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5683[16]));   // verilog/motorControl.v(52[43:52])
    defparam unary_minus_20_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_16_i645_2_lut (.I0(\Kp[13] ), .I1(n55[7]), .I2(GND_net), 
            .I3(GND_net), .O(n959_adj_5434));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i645_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i351_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3715[3] ), 
            .I2(GND_net), .I3(GND_net), .O(n521));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i351_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i400_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3715[3] ), 
            .I2(GND_net), .I3(GND_net), .O(n594));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i400_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i443_2_lut (.I0(\Kp[9] ), .I1(n55[4]), .I2(GND_net), 
            .I3(GND_net), .O(n658));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i443_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i52191_2_lut_4_lut (.I0(PWMLimit[16]), .I1(n352[16]), .I2(PWMLimit[12]), 
            .I3(n352[12]), .O(n67885));
    defparam i52191_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 mult_16_i308_2_lut (.I0(\Kp[6] ), .I1(n55[10]), .I2(GND_net), 
            .I3(GND_net), .O(n457));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i308_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i449_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3715[3] ), 
            .I2(GND_net), .I3(GND_net), .O(n667));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i449_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i52197_2_lut_4_lut (.I0(PWMLimit[14]), .I1(n352[14]), .I2(PWMLimit[13]), 
            .I3(n352[13]), .O(n67891));
    defparam i52197_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i29534_4_lut (.I0(PWMLimit[1]), .I1(n61943), .I2(n37330), 
            .I3(n11595), .O(n51[1]));   // verilog/motorControl.v(41[14] 62[8])
    defparam i29534_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 LessThan_25_i6_3_lut_3_lut (.I0(n352[3]), .I1(n432[3]), .I2(n432[2]), 
            .I3(GND_net), .O(n6_adj_5565));   // verilog/motorControl.v(55[23:39])
    defparam LessThan_25_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 i52177_3_lut_4_lut (.I0(n352[3]), .I1(n432[3]), .I2(n432[2]), 
            .I3(n352[2]), .O(n67871));   // verilog/motorControl.v(55[23:39])
    defparam i52177_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 mult_16_i492_2_lut (.I0(\Kp[10] ), .I1(n55[4]), .I2(GND_net), 
            .I3(GND_net), .O(n731));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i492_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i694_2_lut (.I0(\Kp[14] ), .I1(n55[7]), .I2(GND_net), 
            .I3(GND_net), .O(n1032_adj_5433));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i694_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i357_2_lut (.I0(\Kp[7] ), .I1(n55[10]), .I2(GND_net), 
            .I3(GND_net), .O(n530));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i357_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i118_2_lut (.I0(\Kp[2] ), .I1(n55[13]), .I2(GND_net), 
            .I3(GND_net), .O(n174));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i118_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i498_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3715[3] ), 
            .I2(GND_net), .I3(GND_net), .O(n740));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i498_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_20_inv_0_i18_1_lut (.I0(deadband[17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5683[17]));   // verilog/motorControl.v(52[43:52])
    defparam unary_minus_20_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_17_i547_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3715[3] ), 
            .I2(GND_net), .I3(GND_net), .O(n813));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i547_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_20_inv_0_i19_1_lut (.I0(deadband[18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5683[18]));   // verilog/motorControl.v(52[43:52])
    defparam unary_minus_20_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i13829_3_lut (.I0(n352[2]), .I1(n432[2]), .I2(n11597), .I3(GND_net), 
            .O(n27827));   // verilog/motorControl.v(41[14] 62[8])
    defparam i13829_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29533_4_lut (.I0(PWMLimit[2]), .I1(n61943), .I2(n27827), 
            .I3(n11595), .O(n51[2]));   // verilog/motorControl.v(41[14] 62[8])
    defparam i29533_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 i13824_3_lut (.I0(n352[3]), .I1(n432[3]), .I2(n11597), .I3(GND_net), 
            .O(n27822));   // verilog/motorControl.v(41[14] 62[8])
    defparam i13824_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_17_i596_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3715[3] ), 
            .I2(GND_net), .I3(GND_net), .O(n886));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i596_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_20_inv_0_i20_1_lut (.I0(deadband[19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5683[19]));   // verilog/motorControl.v(52[43:52])
    defparam unary_minus_20_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_17_i645_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3715[3] ), 
            .I2(GND_net), .I3(GND_net), .O(n959));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i645_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i29532_4_lut (.I0(PWMLimit[3]), .I1(n61943), .I2(n27822), 
            .I3(n11595), .O(n51[3]));   // verilog/motorControl.v(41[14] 62[8])
    defparam i29532_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 i23363_3_lut_4_lut (.I0(n376), .I1(n456), .I2(n455), .I3(n375), 
            .O(n4_adj_5566));   // verilog/motorControl.v(51[18:38])
    defparam i23363_3_lut_4_lut.LUT_INIT = 16'h40f4;
    SB_LUT4 i13819_3_lut (.I0(n352[4]), .I1(n432[4]), .I2(n11597), .I3(GND_net), 
            .O(n27817));   // verilog/motorControl.v(41[14] 62[8])
    defparam i13819_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29531_4_lut (.I0(PWMLimit[4]), .I1(n61943), .I2(n27817), 
            .I3(n11595), .O(n51[4]));   // verilog/motorControl.v(41[14] 62[8])
    defparam i29531_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 mult_16_i71_2_lut (.I0(\Kp[1] ), .I1(n55[14]), .I2(GND_net), 
            .I3(GND_net), .O(n104_adj_5428));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i71_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i24_2_lut (.I0(\Kp[0] ), .I1(n55[15]), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_5427));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i24_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i120_2_lut (.I0(\Kp[2] ), .I1(n55[14]), .I2(GND_net), 
            .I3(GND_net), .O(n177_adj_5426));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i120_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_20_inv_0_i21_1_lut (.I0(deadband[20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5683[20]));   // verilog/motorControl.v(52[43:52])
    defparam unary_minus_20_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_16_i406_2_lut (.I0(\Kp[8] ), .I1(n55[10]), .I2(GND_net), 
            .I3(GND_net), .O(n603));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i406_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i36916_2_lut_3_lut (.I0(\Kp[1] ), .I1(n55[22]), .I2(n62), 
            .I3(GND_net), .O(n20087[0]));   // verilog/motorControl.v(51[18:24])
    defparam i36916_2_lut_3_lut.LUT_INIT = 16'h7878;
    SB_LUT4 i1_3_lut_4_lut (.I0(\Kp[1] ), .I1(n55[22]), .I2(n62), .I3(n63605), 
            .O(n20087[1]));   // verilog/motorControl.v(51[18:24])
    defparam i1_3_lut_4_lut.LUT_INIT = 16'h7f80;
    SB_LUT4 i37041_3_lut_4_lut (.I0(n62_adj_5567), .I1(n131), .I2(n204), 
            .I3(n20207[0]), .O(n4_adj_30));   // verilog/motorControl.v(51[27:38])
    defparam i37041_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 unary_minus_20_inv_0_i22_1_lut (.I0(deadband[21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5683[21]));   // verilog/motorControl.v(52[43:52])
    defparam unary_minus_20_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_3_lut_4_lut_adj_1723 (.I0(n62_adj_5567), .I1(n131), .I2(n204), 
            .I3(n20207[0]), .O(n20182));   // verilog/motorControl.v(51[27:38])
    defparam i1_3_lut_4_lut_adj_1723.LUT_INIT = 16'h8778;
    SB_LUT4 mult_16_i169_2_lut (.I0(\Kp[3] ), .I1(n55[14]), .I2(GND_net), 
            .I3(GND_net), .O(n250_adj_5421));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i169_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i218_2_lut (.I0(\Kp[4] ), .I1(n55[14]), .I2(GND_net), 
            .I3(GND_net), .O(n323_adj_5420));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i218_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i455_2_lut (.I0(\Kp[9] ), .I1(n55[10]), .I2(GND_net), 
            .I3(GND_net), .O(n676));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i455_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i743_2_lut (.I0(\Kp[15] ), .I1(n55[7]), .I2(GND_net), 
            .I3(GND_net), .O(n1105_adj_5419));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i743_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i52213_3_lut_4_lut (.I0(PWMLimit[3]), .I1(n352[3]), .I2(n352[2]), 
            .I3(PWMLimit[2]), .O(n67907));   // verilog/motorControl.v(53[14:29])
    defparam i52213_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 unary_minus_20_inv_0_i23_1_lut (.I0(deadband[22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5683[22]));   // verilog/motorControl.v(52[43:52])
    defparam unary_minus_20_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_13_inv_0_i15_1_lut (.I0(IntegralLimit[14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[14]));   // verilog/motorControl.v(49[22:36])
    defparam unary_minus_13_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i13814_3_lut (.I0(n352[5]), .I1(n432[5]), .I2(n11597), .I3(GND_net), 
            .O(n27812));   // verilog/motorControl.v(41[14] 62[8])
    defparam i13814_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29530_4_lut (.I0(PWMLimit[5]), .I1(n61943), .I2(n27812), 
            .I3(n11595), .O(n51[5]));   // verilog/motorControl.v(41[14] 62[8])
    defparam i29530_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 i13809_3_lut (.I0(n352[6]), .I1(n432[6]), .I2(n11597), .I3(GND_net), 
            .O(n27807));   // verilog/motorControl.v(41[14] 62[8])
    defparam i13809_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29529_4_lut (.I0(PWMLimit[6]), .I1(n61943), .I2(n27807), 
            .I3(n11595), .O(n51[6]));   // verilog/motorControl.v(41[14] 62[8])
    defparam i29529_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 LessThan_23_i6_3_lut_3_lut (.I0(PWMLimit[3]), .I1(n352[3]), 
            .I2(n352[2]), .I3(GND_net), .O(n6_adj_5195));   // verilog/motorControl.v(53[14:29])
    defparam LessThan_23_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 unary_minus_20_inv_0_i24_1_lut (.I0(deadband[23]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5683[23]));   // verilog/motorControl.v(52[43:52])
    defparam unary_minus_20_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_16_i267_2_lut (.I0(\Kp[5] ), .I1(n55[14]), .I2(GND_net), 
            .I3(GND_net), .O(n396_adj_5415));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i267_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i13804_3_lut (.I0(n352[7]), .I1(n432[7]), .I2(n11597), .I3(GND_net), 
            .O(n27802));   // verilog/motorControl.v(41[14] 62[8])
    defparam i13804_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29528_4_lut (.I0(PWMLimit[7]), .I1(n61943), .I2(n27802), 
            .I3(n11595), .O(n51[7]));   // verilog/motorControl.v(41[14] 62[8])
    defparam i29528_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 mult_17_i694_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3715[3] ), 
            .I2(GND_net), .I3(GND_net), .O(n1032));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i694_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_19_i41_2_lut (.I0(deadband[20]), .I1(n352[20]), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_5571));   // verilog/motorControl.v(52[12:29])
    defparam LessThan_19_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_19_i39_2_lut (.I0(deadband[19]), .I1(n352[19]), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_5572));   // verilog/motorControl.v(52[12:29])
    defparam LessThan_19_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_16_i504_2_lut (.I0(\Kp[10] ), .I1(n55[10]), .I2(GND_net), 
            .I3(GND_net), .O(n749));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i504_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i52318_3_lut_4_lut (.I0(deadband[3]), .I1(n352[3]), .I2(n352[2]), 
            .I3(deadband[2]), .O(n68012));   // verilog/motorControl.v(52[12:29])
    defparam i52318_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 LessThan_19_i45_2_lut (.I0(deadband[22]), .I1(n352[22]), .I2(GND_net), 
            .I3(GND_net), .O(n45_adj_5573));   // verilog/motorControl.v(52[12:29])
    defparam LessThan_19_i45_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_19_i43_2_lut (.I0(deadband[21]), .I1(n352[21]), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_5574));   // verilog/motorControl.v(52[12:29])
    defparam LessThan_19_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_19_i37_2_lut (.I0(deadband[18]), .I1(n352[18]), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_5575));   // verilog/motorControl.v(52[12:29])
    defparam LessThan_19_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_17_i77_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3715[13] ), 
            .I2(GND_net), .I3(GND_net), .O(n113_adj_5414));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i77_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_19_i6_3_lut_3_lut (.I0(deadband[3]), .I1(n352[3]), 
            .I2(n352[2]), .I3(GND_net), .O(n6_adj_5576));   // verilog/motorControl.v(52[12:29])
    defparam LessThan_19_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 LessThan_19_i29_2_lut (.I0(deadband[14]), .I1(n352[14]), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_5577));   // verilog/motorControl.v(52[12:29])
    defparam LessThan_19_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_19_i31_2_lut (.I0(deadband[15]), .I1(n361), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_5578));   // verilog/motorControl.v(52[12:29])
    defparam LessThan_19_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_19_i21_2_lut (.I0(deadband[10]), .I1(n352[10]), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_5579));   // verilog/motorControl.v(52[12:29])
    defparam LessThan_19_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_19_i23_2_lut (.I0(deadband[11]), .I1(n352[11]), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_5580));   // verilog/motorControl.v(52[12:29])
    defparam LessThan_19_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_17_i30_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3715[14] ), 
            .I2(GND_net), .I3(GND_net), .O(n44_adj_5413));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i30_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_19_i25_2_lut (.I0(deadband[12]), .I1(n352[12]), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_5581));   // verilog/motorControl.v(52[12:29])
    defparam LessThan_19_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_19_i17_2_lut (.I0(deadband[8]), .I1(n352[8]), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_5582));   // verilog/motorControl.v(52[12:29])
    defparam LessThan_19_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_19_i9_2_lut (.I0(deadband[4]), .I1(n352[4]), .I2(GND_net), 
            .I3(GND_net), .O(n9_adj_5583));   // verilog/motorControl.v(52[12:29])
    defparam LessThan_19_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 unary_minus_26_inv_0_i1_1_lut (.I0(PWMLimit[0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5682[0]));   // verilog/motorControl.v(56[22:31])
    defparam unary_minus_26_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 LessThan_19_i35_2_lut (.I0(deadband[17]), .I1(n352[17]), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_5584));   // verilog/motorControl.v(52[12:29])
    defparam LessThan_19_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_19_i33_2_lut (.I0(deadband[16]), .I1(n352[16]), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_5585));   // verilog/motorControl.v(52[12:29])
    defparam LessThan_19_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_19_i11_2_lut (.I0(deadband[5]), .I1(n352[5]), .I2(GND_net), 
            .I3(GND_net), .O(n11_adj_5586));   // verilog/motorControl.v(52[12:29])
    defparam LessThan_19_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_19_i13_2_lut (.I0(deadband[6]), .I1(n352[6]), .I2(GND_net), 
            .I3(GND_net), .O(n13_adj_5587));   // verilog/motorControl.v(52[12:29])
    defparam LessThan_19_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_19_i15_2_lut (.I0(deadband[7]), .I1(n352[7]), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_5588));   // verilog/motorControl.v(52[12:29])
    defparam LessThan_19_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_19_i27_2_lut (.I0(deadband[13]), .I1(n352[13]), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_5589));   // verilog/motorControl.v(52[12:29])
    defparam LessThan_19_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_23_i41_2_lut (.I0(PWMLimit[20]), .I1(n352[20]), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_5590));   // verilog/motorControl.v(53[14:29])
    defparam LessThan_23_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_17_i743_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3715[3] ), 
            .I2(GND_net), .I3(GND_net), .O(n1105));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i743_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_23_i37_2_lut (.I0(PWMLimit[18]), .I1(n352[18]), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_5591));   // verilog/motorControl.v(53[14:29])
    defparam LessThan_23_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_23_i39_2_lut (.I0(PWMLimit[19]), .I1(n352[19]), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_5592));   // verilog/motorControl.v(53[14:29])
    defparam LessThan_23_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_23_i35_2_lut (.I0(PWMLimit[17]), .I1(n352[17]), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_5593));   // verilog/motorControl.v(53[14:29])
    defparam LessThan_23_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_23_i23_2_lut (.I0(PWMLimit[11]), .I1(n352[11]), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_5594));   // verilog/motorControl.v(53[14:29])
    defparam LessThan_23_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_23_i21_2_lut (.I0(PWMLimit[10]), .I1(n352[10]), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_5595));   // verilog/motorControl.v(53[14:29])
    defparam LessThan_23_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i52199_4_lut (.I0(n27_adj_5183), .I1(n25_adj_5199), .I2(n23_adj_5594), 
            .I3(n21_adj_5595), .O(n67893));
    defparam i52199_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 mux_14_i24_3_lut (.I0(n130[23]), .I1(n182[23]), .I2(n181), 
            .I3(GND_net), .O(n207[23]));   // verilog/motorControl.v(48[18] 50[12])
    defparam mux_14_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_16_i316_2_lut (.I0(\Kp[6] ), .I1(n55[14]), .I2(GND_net), 
            .I3(GND_net), .O(n469_adj_5410));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i316_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_15_i24_3_lut (.I0(n207[23]), .I1(IntegralLimit[23]), .I2(n155), 
            .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3715[23] ));   // verilog/motorControl.v(48[18] 50[12])
    defparam mux_15_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_26_inv_0_i2_1_lut (.I0(PWMLimit[1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5682[1]));   // verilog/motorControl.v(56[22:31])
    defparam unary_minus_26_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i52193_4_lut (.I0(n33_adj_5200), .I1(n31), .I2(n29_adj_5184), 
            .I3(n67893), .O(n67887));
    defparam i52193_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 LessThan_23_i26_3_lut (.I0(n352[13]), .I1(n352[14]), .I2(n29_adj_5184), 
            .I3(GND_net), .O(n26_adj_5597));   // verilog/motorControl.v(53[14:29])
    defparam LessThan_23_i26_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_14_i23_3_lut (.I0(n130[22]), .I1(n182[22]), .I2(n181), 
            .I3(GND_net), .O(n207[22]));   // verilog/motorControl.v(48[18] 50[12])
    defparam mux_14_i23_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_15_i23_3_lut (.I0(n207[22]), .I1(IntegralLimit[22]), .I2(n155), 
            .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3715[22] ));   // verilog/motorControl.v(48[18] 50[12])
    defparam mux_15_i23_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_16_i365_2_lut (.I0(\Kp[7] ), .I1(n55[14]), .I2(GND_net), 
            .I3(GND_net), .O(n542_adj_5408));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i365_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_14_i22_3_lut (.I0(n130[21]), .I1(n182[21]), .I2(n181), 
            .I3(GND_net), .O(n207[21]));   // verilog/motorControl.v(48[18] 50[12])
    defparam mux_14_i22_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_23_i28_3_lut (.I0(n26_adj_5597), .I1(n361), .I2(n31), 
            .I3(GND_net), .O(n28_adj_5598));   // verilog/motorControl.v(53[14:29])
    defparam LessThan_23_i28_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_23_i24_3_lut (.I0(n352[12]), .I1(n352[16]), .I2(n33_adj_5200), 
            .I3(GND_net), .O(n24_adj_5599));   // verilog/motorControl.v(53[14:29])
    defparam LessThan_23_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_23_i22_3_lut (.I0(n352[10]), .I1(n352[11]), .I2(n23_adj_5594), 
            .I3(GND_net), .O(n22_adj_5600));   // verilog/motorControl.v(53[14:29])
    defparam LessThan_23_i22_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_15_i22_3_lut (.I0(n207[21]), .I1(IntegralLimit[21]), .I2(n155), 
            .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3715[21] ));   // verilog/motorControl.v(48[18] 50[12])
    defparam mux_15_i22_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_23_i32_3_lut (.I0(n24_adj_5599), .I1(n352[17]), .I2(n35_adj_5593), 
            .I3(GND_net), .O(n32_adj_5601));   // verilog/motorControl.v(53[14:29])
    defparam LessThan_23_i32_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i54042_4_lut (.I0(n32_adj_5601), .I1(n22_adj_5600), .I2(n35_adj_5593), 
            .I3(n67885), .O(n69736));   // verilog/motorControl.v(53[14:29])
    defparam i54042_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i54043_3_lut (.I0(n69736), .I1(n352[18]), .I2(n37_adj_5591), 
            .I3(GND_net), .O(n69737));   // verilog/motorControl.v(53[14:29])
    defparam i54043_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53934_3_lut (.I0(n69737), .I1(n352[19]), .I2(n39_adj_5592), 
            .I3(GND_net), .O(n69628));   // verilog/motorControl.v(53[14:29])
    defparam i53934_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_14_i21_3_lut (.I0(n130[20]), .I1(n182[20]), .I2(n181), 
            .I3(GND_net), .O(n207[20]));   // verilog/motorControl.v(48[18] 50[12])
    defparam mux_14_i21_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53778_4_lut (.I0(n39_adj_5592), .I1(n37_adj_5591), .I2(n35_adj_5593), 
            .I3(n67887), .O(n69472));
    defparam i53778_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i54133_4_lut (.I0(n28_adj_5598), .I1(n20_adj_31), .I2(n31), 
            .I3(n67891), .O(n69827));   // verilog/motorControl.v(53[14:29])
    defparam i54133_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 mux_15_i21_3_lut (.I0(n207[20]), .I1(IntegralLimit[20]), .I2(n155), 
            .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3715[20] ));   // verilog/motorControl.v(48[18] 50[12])
    defparam mux_15_i21_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52599_3_lut (.I0(n69628), .I1(n352[20]), .I2(n41_adj_5590), 
            .I3(GND_net), .O(n68293));   // verilog/motorControl.v(53[14:29])
    defparam i52599_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_16_i553_2_lut (.I0(\Kp[11] ), .I1(n55[10]), .I2(GND_net), 
            .I3(GND_net), .O(n822));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i553_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i54212_4_lut (.I0(n68293), .I1(n69827), .I2(n41_adj_5590), 
            .I3(n69472), .O(n69906));   // verilog/motorControl.v(53[14:29])
    defparam i54212_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 mux_14_i20_3_lut (.I0(n130[19]), .I1(n182[19]), .I2(n181), 
            .I3(GND_net), .O(n212));   // verilog/motorControl.v(48[18] 50[12])
    defparam mux_14_i20_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i54213_3_lut (.I0(n69906), .I1(n352[21]), .I2(PWMLimit[21]), 
            .I3(GND_net), .O(n69907));   // verilog/motorControl.v(53[14:29])
    defparam i54213_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 mux_14_i19_3_lut (.I0(n130[18]), .I1(n182[18]), .I2(n181), 
            .I3(GND_net), .O(n213));   // verilog/motorControl.v(48[18] 50[12])
    defparam mux_14_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i54130_3_lut (.I0(n69907), .I1(n352[22]), .I2(PWMLimit[22]), 
            .I3(GND_net), .O(n69824));   // verilog/motorControl.v(53[14:29])
    defparam i54130_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 mult_17_i55_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3715[2] ), 
            .I2(GND_net), .I3(GND_net), .O(n80_adj_5407));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i55_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i54101_3_lut (.I0(n69824), .I1(PWMLimit[23]), .I2(n352[23]), 
            .I3(GND_net), .O(n405_adj_5603));   // verilog/motorControl.v(53[14:29])
    defparam i54101_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 mult_17_i8_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3715[3] ), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_5406));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i8_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i52252_4_lut (.I0(n352[6]), .I1(n352[5]), .I2(n59[6]), .I3(n59[5]), 
            .O(n67946));
    defparam i52252_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 i53104_3_lut (.I0(n352[7]), .I1(n67946), .I2(n59[7]), .I3(GND_net), 
            .O(n68798));
    defparam i53104_3_lut.LUT_INIT = 16'hdede;
    SB_LUT4 mult_17_i104_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3715[2] ), 
            .I2(GND_net), .I3(GND_net), .O(n153_adj_5405));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i104_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_14_i14_3_lut (.I0(n130[13]), .I1(n182[13]), .I2(n181), 
            .I3(GND_net), .O(n207[13]));   // verilog/motorControl.v(48[18] 50[12])
    defparam mux_14_i14_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_21_i27_rep_73_2_lut (.I0(n352[13]), .I1(n59[13]), .I2(GND_net), 
            .I3(GND_net), .O(n71315));   // verilog/motorControl.v(52[33:53])
    defparam LessThan_21_i27_rep_73_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mux_15_i14_3_lut (.I0(n207[13]), .I1(IntegralLimit[13]), .I2(n155), 
            .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3715[13] ));   // verilog/motorControl.v(48[18] 50[12])
    defparam mux_15_i14_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53092_4_lut (.I0(n352[14]), .I1(n71315), .I2(n59[14]), .I3(n68798), 
            .O(n68786));
    defparam i53092_4_lut.LUT_INIT = 16'hdeff;
    SB_LUT4 LessThan_21_i31_rep_67_2_lut (.I0(n361), .I1(n59[15]), .I2(GND_net), 
            .I3(GND_net), .O(n71309));   // verilog/motorControl.v(52[33:53])
    defparam LessThan_21_i31_rep_67_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_17_i153_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3715[2] ), 
            .I2(GND_net), .I3(GND_net), .O(n226_adj_5404));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i153_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_14_i13_3_lut (.I0(n130[12]), .I1(n182[12]), .I2(n181), 
            .I3(GND_net), .O(n219));   // verilog/motorControl.v(48[18] 50[12])
    defparam mux_14_i13_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52248_4_lut (.I0(n352[8]), .I1(n352[4]), .I2(n59[8]), .I3(n59[4]), 
            .O(n67942));
    defparam i52248_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 i53100_3_lut (.I0(n367), .I1(n67942), .I2(n59[9]), .I3(GND_net), 
            .O(n68794));
    defparam i53100_3_lut.LUT_INIT = 16'hdede;
    SB_LUT4 mult_17_i126_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3715[13] ), 
            .I2(GND_net), .I3(GND_net), .O(n186_adj_5403));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i126_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i541_2_lut (.I0(\Kp[11] ), .I1(n55[4]), .I2(GND_net), 
            .I3(GND_net), .O(n804_adj_5273));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i541_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i202_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3715[2] ), 
            .I2(GND_net), .I3(GND_net), .O(n299_adj_5402));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i202_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_14_i12_3_lut (.I0(n130[11]), .I1(n182[11]), .I2(n181), 
            .I3(GND_net), .O(n207[11]));   // verilog/motorControl.v(48[18] 50[12])
    defparam mux_14_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_21_i21_rep_88_2_lut (.I0(n352[10]), .I1(n59[10]), .I2(GND_net), 
            .I3(GND_net), .O(n71330));   // verilog/motorControl.v(52[33:53])
    defparam LessThan_21_i21_rep_88_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mux_15_i12_3_lut (.I0(n207[11]), .I1(IntegralLimit[11]), .I2(n155), 
            .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3715[11] ));   // verilog/motorControl.v(48[18] 50[12])
    defparam mux_15_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53098_4_lut (.I0(n352[11]), .I1(n71330), .I2(n59[11]), .I3(n68794), 
            .O(n68792));
    defparam i53098_4_lut.LUT_INIT = 16'hdeff;
    SB_LUT4 mult_17_i251_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3715[2] ), 
            .I2(GND_net), .I3(GND_net), .O(n372_adj_5401));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i251_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_14_i11_3_lut (.I0(n130[10]), .I1(n182[10]), .I2(n181), 
            .I3(GND_net), .O(n207[10]));   // verilog/motorControl.v(48[18] 50[12])
    defparam mux_14_i11_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_15_i11_3_lut (.I0(n207[10]), .I1(IntegralLimit[10]), .I2(n155), 
            .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3715[10] ));   // verilog/motorControl.v(48[18] 50[12])
    defparam mux_15_i11_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_14_i10_3_lut (.I0(n130[9]), .I1(n182[9]), .I2(n181), .I3(GND_net), 
            .O(n207[9]));   // verilog/motorControl.v(48[18] 50[12])
    defparam mux_14_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_15_i10_3_lut (.I0(n207[9]), .I1(IntegralLimit[9]), .I2(n155), 
            .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3715[9] ));   // verilog/motorControl.v(48[18] 50[12])
    defparam mux_15_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_21_i25_rep_83_2_lut (.I0(n352[12]), .I1(n59[12]), .I2(GND_net), 
            .I3(GND_net), .O(n71325));   // verilog/motorControl.v(52[33:53])
    defparam LessThan_21_i25_rep_83_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_21_i16_3_lut (.I0(n59[9]), .I1(n59[21]), .I2(n352[21]), 
            .I3(GND_net), .O(n16_adj_5605));   // verilog/motorControl.v(52[33:53])
    defparam LessThan_21_i16_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i52215_4_lut (.I0(n352[21]), .I1(n367), .I2(n59[21]), .I3(n59[9]), 
            .O(n67909));
    defparam i52215_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 mult_17_i300_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3715[2] ), 
            .I2(GND_net), .I3(GND_net), .O(n445_adj_5400));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i300_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i175_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3715[13] ), 
            .I2(GND_net), .I3(GND_net), .O(n259));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i175_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_14_i9_3_lut (.I0(n130[8]), .I1(n182[8]), .I2(n181), .I3(GND_net), 
            .O(n207[8]));   // verilog/motorControl.v(48[18] 50[12])
    defparam mux_14_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_15_i9_3_lut (.I0(n207[8]), .I1(IntegralLimit[8]), .I2(n155), 
            .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3715[8] ));   // verilog/motorControl.v(48[18] 50[12])
    defparam mux_15_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_21_i8_3_lut (.I0(n59[4]), .I1(n59[8]), .I2(n352[8]), 
            .I3(GND_net), .O(n8_adj_5607));   // verilog/motorControl.v(52[33:53])
    defparam LessThan_21_i8_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 mult_17_i349_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3715[2] ), 
            .I2(GND_net), .I3(GND_net), .O(n518_adj_5399));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i349_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_14_i8_3_lut (.I0(n130[7]), .I1(n182[7]), .I2(n181), .I3(GND_net), 
            .O(n207[7]));   // verilog/motorControl.v(48[18] 50[12])
    defparam mux_14_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_15_i8_3_lut (.I0(n207[7]), .I1(IntegralLimit[7]), .I2(n155), 
            .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3715[7] ));   // verilog/motorControl.v(48[18] 50[12])
    defparam mux_15_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_21_i24_3_lut (.I0(n16_adj_5605), .I1(n59[22]), .I2(n352[22]), 
            .I3(GND_net), .O(n24_adj_5608));   // verilog/motorControl.v(52[33:53])
    defparam LessThan_21_i24_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 mult_17_i398_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3715[2] ), 
            .I2(GND_net), .I3(GND_net), .O(n591_adj_5398));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i398_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_14_i7_3_lut (.I0(n130[6]), .I1(n182[6]), .I2(n181), .I3(GND_net), 
            .O(n207[6]));   // verilog/motorControl.v(48[18] 50[12])
    defparam mux_14_i7_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_15_i7_3_lut (.I0(n207[6]), .I1(IntegralLimit[6]), .I2(n155), 
            .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3715[6] ));   // verilog/motorControl.v(48[18] 50[12])
    defparam mux_15_i7_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_16_i414_2_lut (.I0(\Kp[8] ), .I1(n55[14]), .I2(GND_net), 
            .I3(GND_net), .O(n615_adj_5397));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i414_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_14_i6_3_lut (.I0(n130[5]), .I1(n182[5]), .I2(n181), .I3(GND_net), 
            .O(n207[5]));   // verilog/motorControl.v(48[18] 50[12])
    defparam mux_14_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_15_i6_3_lut (.I0(n207[5]), .I1(IntegralLimit[5]), .I2(n155), 
            .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3715[5] ));   // verilog/motorControl.v(48[18] 50[12])
    defparam mux_15_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52256_4_lut (.I0(n352[3]), .I1(n352[2]), .I2(n59[3]), .I3(n59[2]), 
            .O(n67950));
    defparam i52256_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 mult_17_i447_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3715[2] ), 
            .I2(GND_net), .I3(GND_net), .O(n664_adj_5396));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i447_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_14_i5_3_lut (.I0(n130[4]), .I1(n182[4]), .I2(n181), .I3(GND_net), 
            .O(n207[4]));   // verilog/motorControl.v(48[18] 50[12])
    defparam mux_14_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_17_i496_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3715[2] ), 
            .I2(GND_net), .I3(GND_net), .O(n737_adj_5395));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i496_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_21_i9_rep_81_2_lut (.I0(n352[4]), .I1(n59[4]), .I2(GND_net), 
            .I3(GND_net), .O(n71323));   // verilog/motorControl.v(52[33:53])
    defparam LessThan_21_i9_rep_81_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mux_15_i5_3_lut (.I0(n207[4]), .I1(IntegralLimit[4]), .I2(n155), 
            .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3715[4] ));   // verilog/motorControl.v(48[18] 50[12])
    defparam mux_15_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_17_i545_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3715[2] ), 
            .I2(GND_net), .I3(GND_net), .O(n810_adj_5394));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i545_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i52254_4_lut (.I0(n352[5]), .I1(n71323), .I2(n59[5]), .I3(n67950), 
            .O(n67948));
    defparam i52254_4_lut.LUT_INIT = 16'h5a7b;
    SB_LUT4 unary_minus_26_inv_0_i3_1_lut (.I0(PWMLimit[2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5682[2]));   // verilog/motorControl.v(56[22:31])
    defparam unary_minus_26_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_16_i602_2_lut (.I0(\Kp[12] ), .I1(n55[10]), .I2(GND_net), 
            .I3(GND_net), .O(n895));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i602_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_21_i13_rep_109_2_lut (.I0(n352[6]), .I1(n59[6]), .I2(GND_net), 
            .I3(GND_net), .O(n71351));   // verilog/motorControl.v(52[33:53])
    defparam LessThan_21_i13_rep_109_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mux_14_i4_3_lut (.I0(n130[3]), .I1(n182[3]), .I2(n181), .I3(GND_net), 
            .O(n207[3]));   // verilog/motorControl.v(48[18] 50[12])
    defparam mux_14_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53481_4_lut (.I0(n352[7]), .I1(n71351), .I2(n59[7]), .I3(n67948), 
            .O(n69175));
    defparam i53481_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 mult_16_i463_2_lut (.I0(\Kp[9] ), .I1(n55[14]), .I2(GND_net), 
            .I3(GND_net), .O(n688_adj_5391));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i463_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i594_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3715[2] ), 
            .I2(GND_net), .I3(GND_net), .O(n883_adj_5390));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i594_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_15_i4_3_lut (.I0(n207[3]), .I1(IntegralLimit[3]), .I2(n155), 
            .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3715[3] ));   // verilog/motorControl.v(48[18] 50[12])
    defparam mux_15_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_14_i3_3_lut (.I0(n130[2]), .I1(n182[2]), .I2(n181), .I3(GND_net), 
            .O(n207[2]));   // verilog/motorControl.v(48[18] 50[12])
    defparam mux_14_i3_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_17_i643_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3715[2] ), 
            .I2(GND_net), .I3(GND_net), .O(n956_adj_5389));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i643_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_15_i3_3_lut (.I0(n207[2]), .I1(IntegralLimit[2]), .I2(n155), 
            .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3715[2] ));   // verilog/motorControl.v(48[18] 50[12])
    defparam mux_15_i3_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_14_i2_3_lut (.I0(n130[1]), .I1(n182[1]), .I2(n181), .I3(GND_net), 
            .O(n230));   // verilog/motorControl.v(48[18] 50[12])
    defparam mux_14_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_21_i17_rep_106_2_lut (.I0(n352[8]), .I1(n59[8]), .I2(GND_net), 
            .I3(GND_net), .O(n71348));   // verilog/motorControl.v(52[33:53])
    defparam LessThan_21_i17_rep_106_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i53102_4_lut (.I0(n367), .I1(n71348), .I2(n59[9]), .I3(n69175), 
            .O(n68796));
    defparam i53102_4_lut.LUT_INIT = 16'hdeff;
    SB_LUT4 mult_16_i651_2_lut (.I0(\Kp[13] ), .I1(n55[10]), .I2(GND_net), 
            .I3(GND_net), .O(n968));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i651_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i692_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3715[2] ), 
            .I2(GND_net), .I3(GND_net), .O(n1029_adj_5388));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i692_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i13799_3_lut (.I0(n352[8]), .I1(n432[8]), .I2(n11597), .I3(GND_net), 
            .O(n27797));   // verilog/motorControl.v(41[14] 62[8])
    defparam i13799_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53784_4_lut (.I0(n352[11]), .I1(n71330), .I2(n59[11]), .I3(n68796), 
            .O(n69478));
    defparam i53784_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 i29527_4_lut (.I0(PWMLimit[8]), .I1(n61943), .I2(n27797), 
            .I3(n11595), .O(n51[8]));   // verilog/motorControl.v(41[14] 62[8])
    defparam i29527_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 i52239_4_lut (.I0(n352[13]), .I1(n71325), .I2(n59[13]), .I3(n69478), 
            .O(n67933));
    defparam i52239_4_lut.LUT_INIT = 16'h5a7b;
    SB_LUT4 i13794_3_lut (.I0(n367), .I1(n432[9]), .I2(n11597), .I3(GND_net), 
            .O(n27792));   // verilog/motorControl.v(41[14] 62[8])
    defparam i13794_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_21_i29_rep_71_2_lut (.I0(n352[14]), .I1(n59[14]), .I2(GND_net), 
            .I3(GND_net), .O(n71313));   // verilog/motorControl.v(52[33:53])
    defparam LessThan_21_i29_rep_71_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i29526_4_lut (.I0(PWMLimit[9]), .I1(n61943), .I2(n27792), 
            .I3(n11595), .O(n51[9]));   // verilog/motorControl.v(41[14] 62[8])
    defparam i29526_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 i53475_4_lut (.I0(n361), .I1(n71313), .I2(n59[15]), .I3(n67933), 
            .O(n69169));
    defparam i53475_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 unary_minus_26_inv_0_i4_1_lut (.I0(PWMLimit[3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5682[3]));   // verilog/motorControl.v(56[22:31])
    defparam unary_minus_26_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_17_i741_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3715[2] ), 
            .I2(GND_net), .I3(GND_net), .O(n1102_adj_5386));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i741_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i13789_3_lut (.I0(n352[10]), .I1(n432[10]), .I2(n11597), .I3(GND_net), 
            .O(n27787));   // verilog/motorControl.v(41[14] 62[8])
    defparam i13789_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29525_4_lut (.I0(PWMLimit[10]), .I1(n61943), .I2(n27787), 
            .I3(n11595), .O(n51[10]));   // verilog/motorControl.v(41[14] 62[8])
    defparam i29525_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 unary_minus_26_inv_0_i5_1_lut (.I0(PWMLimit[4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5682[4]));   // verilog/motorControl.v(56[22:31])
    defparam unary_minus_26_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 LessThan_21_i33_rep_99_2_lut (.I0(n352[16]), .I1(n59[16]), .I2(GND_net), 
            .I3(GND_net), .O(n71341));   // verilog/motorControl.v(52[33:53])
    defparam LessThan_21_i33_rep_99_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i54030_4_lut (.I0(n352[17]), .I1(n71341), .I2(n59[17]), .I3(n69169), 
            .O(n69724));
    defparam i54030_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 LessThan_21_i37_rep_62_2_lut (.I0(n352[18]), .I1(n59[18]), .I2(GND_net), 
            .I3(GND_net), .O(n71304));   // verilog/motorControl.v(52[33:53])
    defparam LessThan_21_i37_rep_62_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i54245_4_lut (.I0(n352[19]), .I1(n71304), .I2(n59[19]), .I3(n69724), 
            .O(n69939));
    defparam i54245_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 LessThan_21_i41_rep_59_2_lut (.I0(n352[20]), .I1(n59[20]), .I2(GND_net), 
            .I3(GND_net), .O(n71301));   // verilog/motorControl.v(52[33:53])
    defparam LessThan_21_i41_rep_59_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i52284_4_lut (.I0(n27_adj_5589), .I1(n15_adj_5588), .I2(n13_adj_5587), 
            .I3(n11_adj_5586), .O(n67978));
    defparam i52284_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 mult_16_i512_2_lut (.I0(\Kp[10] ), .I1(n55[14]), .I2(GND_net), 
            .I3(GND_net), .O(n761_adj_5384));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i512_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i561_2_lut (.I0(\Kp[11] ), .I1(n55[14]), .I2(GND_net), 
            .I3(GND_net), .O(n834_adj_5383));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i561_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_19_i12_3_lut (.I0(n352[7]), .I1(n352[16]), .I2(n33_adj_5585), 
            .I3(GND_net), .O(n12_adj_5611));   // verilog/motorControl.v(52[12:29])
    defparam LessThan_19_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_19_i10_3_lut (.I0(n352[5]), .I1(n352[6]), .I2(n13_adj_5587), 
            .I3(GND_net), .O(n10_adj_5612));   // verilog/motorControl.v(52[12:29])
    defparam LessThan_19_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_19_i30_3_lut (.I0(n12_adj_5611), .I1(n352[17]), .I2(n35_adj_5584), 
            .I3(GND_net), .O(n30_adj_5613));   // verilog/motorControl.v(52[12:29])
    defparam LessThan_19_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53138_4_lut (.I0(n13_adj_5587), .I1(n11_adj_5586), .I2(n9_adj_5583), 
            .I3(n68012), .O(n68832));
    defparam i53138_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i53134_4_lut (.I0(n19), .I1(n17_adj_5582), .I2(n15_adj_5588), 
            .I3(n68832), .O(n68828));
    defparam i53134_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 mult_16_i700_2_lut (.I0(\Kp[14] ), .I1(n55[10]), .I2(GND_net), 
            .I3(GND_net), .O(n1041));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i700_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i54076_4_lut (.I0(n25_adj_5581), .I1(n23_adj_5580), .I2(n21_adj_5579), 
            .I3(n68828), .O(n69770));
    defparam i54076_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i53497_4_lut (.I0(n31_adj_5578), .I1(n29_adj_5577), .I2(n27_adj_5589), 
            .I3(n69770), .O(n69191));
    defparam i53497_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i54157_4_lut (.I0(n37_adj_5575), .I1(n35_adj_5584), .I2(n33_adj_5585), 
            .I3(n69191), .O(n69851));
    defparam i54157_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 unary_minus_26_inv_0_i6_1_lut (.I0(PWMLimit[5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5682[5]));   // verilog/motorControl.v(56[22:31])
    defparam unary_minus_26_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_17_i224_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3715[13] ), 
            .I2(GND_net), .I3(GND_net), .O(n332_adj_5380));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i224_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i53649_3_lut (.I0(n6_adj_5576), .I1(n352[10]), .I2(n21_adj_5579), 
            .I3(GND_net), .O(n69343));   // verilog/motorControl.v(52[12:29])
    defparam i53649_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_17_i53_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3715[1] ), 
            .I2(GND_net), .I3(GND_net), .O(n77_adj_5379));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i53_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i6_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3715[2] ), 
            .I2(GND_net), .I3(GND_net), .O(n8_adj_5378));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i6_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i610_2_lut (.I0(\Kp[12] ), .I1(n55[14]), .I2(GND_net), 
            .I3(GND_net), .O(n907_adj_5376));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i610_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_19_i16_3_lut (.I0(n367), .I1(n352[21]), .I2(n43_adj_5574), 
            .I3(GND_net), .O(n16_adj_5615));   // verilog/motorControl.v(52[12:29])
    defparam LessThan_19_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_16_i749_2_lut (.I0(\Kp[15] ), .I1(n55[10]), .I2(GND_net), 
            .I3(GND_net), .O(n1114));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i749_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_26_inv_0_i7_1_lut (.I0(PWMLimit[6]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5682[6]));   // verilog/motorControl.v(56[22:31])
    defparam unary_minus_26_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_17_i102_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3715[1] ), 
            .I2(GND_net), .I3(GND_net), .O(n150_adj_5374));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i102_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i151_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3715[1] ), 
            .I2(GND_net), .I3(GND_net), .O(n223_adj_5372));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i151_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_19_i8_3_lut (.I0(n352[4]), .I1(n352[8]), .I2(n17_adj_5582), 
            .I3(GND_net), .O(n8_adj_5616));   // verilog/motorControl.v(52[12:29])
    defparam LessThan_19_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_19_i24_3_lut (.I0(n16_adj_5615), .I1(n352[22]), .I2(n45_adj_5573), 
            .I3(GND_net), .O(n24_adj_5617));   // verilog/motorControl.v(52[12:29])
    defparam LessThan_19_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_26_inv_0_i8_1_lut (.I0(PWMLimit[7]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5682[7]));   // verilog/motorControl.v(56[22:31])
    defparam unary_minus_26_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i52290_4_lut (.I0(n21_adj_5579), .I1(n19), .I2(n17_adj_5582), 
            .I3(n9_adj_5583), .O(n67984));
    defparam i52290_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i53650_3_lut (.I0(n69343), .I1(n352[11]), .I2(n23_adj_5580), 
            .I3(GND_net), .O(n69344));   // verilog/motorControl.v(52[12:29])
    defparam i53650_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52260_4_lut (.I0(n43_adj_5574), .I1(n25_adj_5581), .I2(n23_adj_5580), 
            .I3(n67984), .O(n67954));
    defparam i52260_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i53561_4_lut (.I0(n24_adj_5617), .I1(n8_adj_5616), .I2(n45_adj_5573), 
            .I3(n67952), .O(n69255));   // verilog/motorControl.v(52[12:29])
    defparam i53561_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i52575_3_lut (.I0(n69344), .I1(n352[12]), .I2(n25_adj_5581), 
            .I3(GND_net), .O(n68269));   // verilog/motorControl.v(52[12:29])
    defparam i52575_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_16_i659_2_lut (.I0(\Kp[13] ), .I1(n55[14]), .I2(GND_net), 
            .I3(GND_net), .O(n980_adj_5370));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i659_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i200_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3715[1] ), 
            .I2(GND_net), .I3(GND_net), .O(n296_adj_5369));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i200_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i273_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3715[13] ), 
            .I2(GND_net), .I3(GND_net), .O(n405));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i273_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_21_i12_3_lut (.I0(n59[7]), .I1(n59[16]), .I2(n352[16]), 
            .I3(GND_net), .O(n12_adj_5618));   // verilog/motorControl.v(52[33:53])
    defparam LessThan_21_i12_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 mult_17_i322_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3715[13] ), 
            .I2(GND_net), .I3(GND_net), .O(n478));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i322_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_26_inv_0_i9_1_lut (.I0(PWMLimit[8]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5682[8]));   // verilog/motorControl.v(56[22:31])
    defparam unary_minus_26_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i53635_3_lut (.I0(n4_adj_32), .I1(n59[13]), .I2(n352[13]), 
            .I3(GND_net), .O(n69329));   // verilog/motorControl.v(52[33:53])
    defparam i53635_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i53636_3_lut (.I0(n69329), .I1(n59[14]), .I2(n352[14]), .I3(GND_net), 
            .O(n69330));   // verilog/motorControl.v(52[33:53])
    defparam i53636_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i13784_3_lut (.I0(n352[11]), .I1(n432[11]), .I2(n11597), .I3(GND_net), 
            .O(n27782));   // verilog/motorControl.v(41[14] 62[8])
    defparam i13784_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29524_4_lut (.I0(PWMLimit[11]), .I1(n61943), .I2(n27782), 
            .I3(n11595), .O(n51[11]));   // verilog/motorControl.v(41[14] 62[8])
    defparam i29524_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 i13779_3_lut (.I0(n352[12]), .I1(n432[12]), .I2(n11597), .I3(GND_net), 
            .O(n27777));   // verilog/motorControl.v(41[14] 62[8])
    defparam i13779_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52227_4_lut (.I0(n352[16]), .I1(n352[7]), .I2(n59[16]), .I3(n59[7]), 
            .O(n67921));
    defparam i52227_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 LessThan_21_i35_rep_94_2_lut (.I0(n352[17]), .I1(n59[17]), .I2(GND_net), 
            .I3(GND_net), .O(n71336));   // verilog/motorControl.v(52[33:53])
    defparam LessThan_21_i35_rep_94_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_21_i10_3_lut (.I0(n59[5]), .I1(n59[6]), .I2(n352[6]), 
            .I3(GND_net), .O(n10_adj_5620));   // verilog/motorControl.v(52[33:53])
    defparam LessThan_21_i10_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i29523_4_lut (.I0(PWMLimit[12]), .I1(n61943), .I2(n27777), 
            .I3(n11595), .O(n51[12]));   // verilog/motorControl.v(41[14] 62[8])
    defparam i29523_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 LessThan_21_i30_3_lut (.I0(n12_adj_5618), .I1(n59[17]), .I2(n352[17]), 
            .I3(GND_net), .O(n30_adj_5621));   // verilog/motorControl.v(52[33:53])
    defparam LessThan_21_i30_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i52229_4_lut (.I0(n352[16]), .I1(n71309), .I2(n59[16]), .I3(n68786), 
            .O(n67923));
    defparam i52229_4_lut.LUT_INIT = 16'h5a7b;
    SB_LUT4 i54040_4_lut (.I0(n30_adj_5621), .I1(n10_adj_5620), .I2(n71336), 
            .I3(n67921), .O(n69734));   // verilog/motorControl.v(52[33:53])
    defparam i54040_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i52587_3_lut (.I0(n69330), .I1(n59[15]), .I2(n361), .I3(GND_net), 
            .O(n68281));   // verilog/motorControl.v(52[33:53])
    defparam i52587_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i54232_4_lut (.I0(n68281), .I1(n69734), .I2(n71336), .I3(n67923), 
            .O(n69926));   // verilog/motorControl.v(52[33:53])
    defparam i54232_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i54233_3_lut (.I0(n69926), .I1(n59[18]), .I2(n352[18]), .I3(GND_net), 
            .O(n69927));   // verilog/motorControl.v(52[33:53])
    defparam i54233_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 LessThan_21_i6_3_lut (.I0(n59[2]), .I1(n59[3]), .I2(n352[3]), 
            .I3(GND_net), .O(n6_adj_5622));   // verilog/motorControl.v(52[33:53])
    defparam LessThan_21_i6_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i53639_3_lut (.I0(n6_adj_5622), .I1(n59[10]), .I2(n352[10]), 
            .I3(GND_net), .O(n69333));   // verilog/motorControl.v(52[33:53])
    defparam i53639_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i53640_3_lut (.I0(n69333), .I1(n59[11]), .I2(n352[11]), .I3(GND_net), 
            .O(n69334));   // verilog/motorControl.v(52[33:53])
    defparam i53640_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i13774_3_lut (.I0(n352[13]), .I1(n432[13]), .I2(n11597), .I3(GND_net), 
            .O(n27772));   // verilog/motorControl.v(41[14] 62[8])
    defparam i13774_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29522_4_lut (.I0(PWMLimit[13]), .I1(n61943), .I2(n27772), 
            .I3(n11595), .O(n51[13]));   // verilog/motorControl.v(41[14] 62[8])
    defparam i29522_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 unary_minus_26_inv_0_i10_1_lut (.I0(PWMLimit[9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5682[9]));   // verilog/motorControl.v(56[22:31])
    defparam unary_minus_26_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i52219_4_lut (.I0(n352[21]), .I1(n71325), .I2(n59[21]), .I3(n68792), 
            .O(n67913));
    defparam i52219_4_lut.LUT_INIT = 16'h5a7b;
    SB_LUT4 mult_17_i371_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3715[13] ), 
            .I2(GND_net), .I3(GND_net), .O(n551));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i371_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i249_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3715[1] ), 
            .I2(GND_net), .I3(GND_net), .O(n369_adj_5363));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i249_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_21_i45_rep_56_2_lut (.I0(n352[22]), .I1(n59[22]), .I2(GND_net), 
            .I3(GND_net), .O(n71298));   // verilog/motorControl.v(52[33:53])
    defparam LessThan_21_i45_rep_56_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i53563_4_lut (.I0(n24_adj_5608), .I1(n8_adj_5607), .I2(n71298), 
            .I3(n67909), .O(n69257));   // verilog/motorControl.v(52[33:53])
    defparam i53563_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 unary_minus_26_inv_0_i11_1_lut (.I0(PWMLimit[10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5682[10]));   // verilog/motorControl.v(56[22:31])
    defparam unary_minus_26_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_17_i298_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3715[1] ), 
            .I2(GND_net), .I3(GND_net), .O(n442_adj_5361));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i298_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i420_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3715[13] ), 
            .I2(GND_net), .I3(GND_net), .O(n624));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i420_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i52585_3_lut (.I0(n69334), .I1(n59[12]), .I2(n352[12]), .I3(GND_net), 
            .O(n68279));   // verilog/motorControl.v(52[33:53])
    defparam i52585_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i13769_3_lut (.I0(n352[14]), .I1(n432[14]), .I2(n11597), .I3(GND_net), 
            .O(n27767));   // verilog/motorControl.v(41[14] 62[8])
    defparam i13769_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i54190_3_lut (.I0(n69927), .I1(n59[19]), .I2(n352[19]), .I3(GND_net), 
            .O(n69884));   // verilog/motorControl.v(52[33:53])
    defparam i54190_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i29521_4_lut (.I0(PWMLimit[14]), .I1(n61943), .I2(n27767), 
            .I3(n11595), .O(n51[14]));   // verilog/motorControl.v(41[14] 62[8])
    defparam i29521_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 i52221_4_lut (.I0(n352[21]), .I1(n71301), .I2(n59[21]), .I3(n69939), 
            .O(n67915));
    defparam i52221_4_lut.LUT_INIT = 16'h5a7b;
    SB_LUT4 mult_17_i347_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3715[1] ), 
            .I2(GND_net), .I3(GND_net), .O(n515_adj_5357));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i347_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i396_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3715[1] ), 
            .I2(GND_net), .I3(GND_net), .O(n588_adj_5356));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i396_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i13764_3_lut (.I0(n361), .I1(n432[15]), .I2(n11597), .I3(GND_net), 
            .O(n27762));   // verilog/motorControl.v(41[14] 62[8])
    defparam i13764_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53893_4_lut (.I0(n68279), .I1(n69257), .I2(n71298), .I3(n67913), 
            .O(n69587));   // verilog/motorControl.v(52[33:53])
    defparam i53893_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i29520_4_lut (.I0(PWMLimit[15]), .I1(n61943), .I2(n27762), 
            .I3(n11595), .O(n51[15]));   // verilog/motorControl.v(41[14] 62[8])
    defparam i29520_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 i13759_3_lut (.I0(n352[16]), .I1(n432[16]), .I2(n11597), .I3(GND_net), 
            .O(n27757));   // verilog/motorControl.v(41[14] 62[8])
    defparam i13759_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_26_inv_0_i12_1_lut (.I0(PWMLimit[11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5682[11]));   // verilog/motorControl.v(56[22:31])
    defparam unary_minus_26_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i29519_4_lut (.I0(PWMLimit[16]), .I1(n61943), .I2(n27757), 
            .I3(n11595), .O(n51[16]));   // verilog/motorControl.v(41[14] 62[8])
    defparam i29519_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 i13754_3_lut (.I0(n352[17]), .I1(n432[17]), .I2(n11597), .I3(GND_net), 
            .O(n27752));   // verilog/motorControl.v(41[14] 62[8])
    defparam i13754_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29518_4_lut (.I0(PWMLimit[17]), .I1(n61943), .I2(n27752), 
            .I3(n11595), .O(n51[17]));   // verilog/motorControl.v(41[14] 62[8])
    defparam i29518_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 i52593_3_lut (.I0(n69884), .I1(n59[20]), .I2(n352[20]), .I3(GND_net), 
            .O(n68287));   // verilog/motorControl.v(52[33:53])
    defparam i52593_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 LessThan_19_i4_4_lut (.I0(deadband[0]), .I1(n375), .I2(deadband[1]), 
            .I3(n376), .O(n4_adj_5623));   // verilog/motorControl.v(52[12:29])
    defparam LessThan_19_i4_4_lut.LUT_INIT = 16'h4d0c;
    SB_LUT4 i53645_3_lut (.I0(n4_adj_5623), .I1(n352[13]), .I2(n27_adj_5589), 
            .I3(GND_net), .O(n69339));   // verilog/motorControl.v(52[12:29])
    defparam i53645_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53646_3_lut (.I0(n69339), .I1(n352[14]), .I2(n29_adj_5577), 
            .I3(GND_net), .O(n69340));   // verilog/motorControl.v(52[12:29])
    defparam i53646_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_17_i445_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3715[1] ), 
            .I2(GND_net), .I3(GND_net), .O(n661_adj_5353));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i445_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i13749_3_lut (.I0(n352[18]), .I1(n432[18]), .I2(n11597), .I3(GND_net), 
            .O(n27747));   // verilog/motorControl.v(41[14] 62[8])
    defparam i13749_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29517_4_lut (.I0(PWMLimit[18]), .I1(n61943), .I2(n27747), 
            .I3(n11595), .O(n51[18]));   // verilog/motorControl.v(41[14] 62[8])
    defparam i29517_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 i52275_4_lut (.I0(n33_adj_5585), .I1(n31_adj_5578), .I2(n29_adj_5577), 
            .I3(n67978), .O(n67969));
    defparam i52275_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i54038_4_lut (.I0(n30_adj_5613), .I1(n10_adj_5612), .I2(n35_adj_5584), 
            .I3(n67962), .O(n69732));   // verilog/motorControl.v(52[12:29])
    defparam i54038_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i52577_3_lut (.I0(n69340), .I1(n361), .I2(n31_adj_5578), .I3(GND_net), 
            .O(n68271));   // verilog/motorControl.v(52[12:29])
    defparam i52577_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i54230_4_lut (.I0(n68271), .I1(n69732), .I2(n35_adj_5584), 
            .I3(n67969), .O(n69924));   // verilog/motorControl.v(52[12:29])
    defparam i54230_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 unary_minus_26_inv_0_i13_1_lut (.I0(PWMLimit[12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5682[12]));   // verilog/motorControl.v(56[22:31])
    defparam unary_minus_26_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i54231_3_lut (.I0(n69924), .I1(n352[18]), .I2(n37_adj_5575), 
            .I3(GND_net), .O(n69925));   // verilog/motorControl.v(52[12:29])
    defparam i54231_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i54192_3_lut (.I0(n69925), .I1(n352[19]), .I2(n39_adj_5572), 
            .I3(GND_net), .O(n69886));   // verilog/motorControl.v(52[12:29])
    defparam i54192_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52262_4_lut (.I0(n43_adj_5574), .I1(n41_adj_5571), .I2(n39_adj_5572), 
            .I3(n69851), .O(n67956));
    defparam i52262_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i53891_4_lut (.I0(n68269), .I1(n69255), .I2(n45_adj_5573), 
            .I3(n67954), .O(n69585));   // verilog/motorControl.v(52[12:29])
    defparam i53891_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i13744_3_lut (.I0(n352[19]), .I1(n432[19]), .I2(n11597), .I3(GND_net), 
            .O(n27742));   // verilog/motorControl.v(41[14] 62[8])
    defparam i13744_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52583_3_lut (.I0(n69886), .I1(n352[20]), .I2(n41_adj_5571), 
            .I3(GND_net), .O(n68277));   // verilog/motorControl.v(52[12:29])
    defparam i52583_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i54096_4_lut (.I0(n68277), .I1(n69585), .I2(n45_adj_5573), 
            .I3(n67956), .O(n69790));   // verilog/motorControl.v(52[12:29])
    defparam i54096_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 mult_17_i469_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3715[13] ), 
            .I2(GND_net), .I3(GND_net), .O(n697));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i469_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i29516_4_lut (.I0(PWMLimit[19]), .I1(n61943), .I2(n27742), 
            .I3(n11595), .O(n51[19]));   // verilog/motorControl.v(41[14] 62[8])
    defparam i29516_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 i54098_4_lut (.I0(n68287), .I1(n69587), .I2(n71298), .I3(n67915), 
            .O(n69792));   // verilog/motorControl.v(52[33:53])
    defparam i54098_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 mult_17_i494_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3715[1] ), 
            .I2(GND_net), .I3(GND_net), .O(n734_adj_5351));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i494_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i518_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3715[13] ), 
            .I2(GND_net), .I3(GND_net), .O(n770));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i518_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i13739_3_lut (.I0(n352[20]), .I1(n432[20]), .I2(n11597), .I3(GND_net), 
            .O(n27737));   // verilog/motorControl.v(41[14] 62[8])
    defparam i13739_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1724 (.I0(n69790), .I1(control_update), .I2(deadband[23]), 
            .I3(n352[23]), .O(n63567));
    defparam i1_4_lut_adj_1724.LUT_INIT = 16'h4c04;
    SB_LUT4 i29515_4_lut (.I0(PWMLimit[20]), .I1(n61943), .I2(n27737), 
            .I3(n11595), .O(n51[20]));   // verilog/motorControl.v(41[14] 62[8])
    defparam i29515_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 i1_4_lut_adj_1725 (.I0(n63567), .I1(n69792), .I2(n352[23]), 
            .I3(n47_adj_5416), .O(n61943));
    defparam i1_4_lut_adj_1725.LUT_INIT = 16'h0a22;
    SB_LUT4 i13734_3_lut (.I0(n352[21]), .I1(n432[21]), .I2(n11597), .I3(GND_net), 
            .O(n27732));   // verilog/motorControl.v(41[14] 62[8])
    defparam i13734_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29514_4_lut (.I0(PWMLimit[21]), .I1(n61943), .I2(n27732), 
            .I3(n11595), .O(n51[21]));   // verilog/motorControl.v(41[14] 62[8])
    defparam i29514_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 mult_17_i543_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3715[1] ), 
            .I2(GND_net), .I3(GND_net), .O(n807_adj_5349));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i543_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i81_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3715[15] ), 
            .I2(GND_net), .I3(GND_net), .O(n119_adj_5348));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i81_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i13729_3_lut (.I0(n352[22]), .I1(n432[22]), .I2(n11597), .I3(GND_net), 
            .O(n27727));   // verilog/motorControl.v(41[14] 62[8])
    defparam i13729_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29513_4_lut (.I0(PWMLimit[22]), .I1(n61943), .I2(n27727), 
            .I3(n11595), .O(n51[22]));   // verilog/motorControl.v(41[14] 62[8])
    defparam i29513_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 mult_17_i34_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3715[16] ), 
            .I2(GND_net), .I3(GND_net), .O(n50_adj_5347));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i34_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i592_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3715[1] ), 
            .I2(GND_net), .I3(GND_net), .O(n880_adj_5346));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i592_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i13724_3_lut (.I0(n352[23]), .I1(n432[23]), .I2(n11597), .I3(GND_net), 
            .O(n27722));   // verilog/motorControl.v(41[14] 62[8])
    defparam i13724_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29512_4_lut (.I0(PWMLimit[23]), .I1(n61943), .I2(n27722), 
            .I3(n11595), .O(n51[23]));   // verilog/motorControl.v(41[14] 62[8])
    defparam i29512_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 mult_17_i641_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3715[1] ), 
            .I2(GND_net), .I3(GND_net), .O(n953_adj_5345));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i641_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_26_inv_0_i14_1_lut (.I0(PWMLimit[13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5682[13]));   // verilog/motorControl.v(56[22:31])
    defparam unary_minus_26_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_16_i51_2_lut (.I0(\Kp[1] ), .I1(n55[4]), .I2(GND_net), 
            .I3(GND_net), .O(n74_adj_5343));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i51_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i4_2_lut (.I0(\Kp[0] ), .I1(n55[5]), .I2(GND_net), 
            .I3(GND_net), .O(n5_adj_5342));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i4_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i690_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3715[1] ), 
            .I2(GND_net), .I3(GND_net), .O(n1026_adj_5341));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i690_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_26_inv_0_i15_1_lut (.I0(PWMLimit[14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5682[14]));   // verilog/motorControl.v(56[22:31])
    defparam unary_minus_26_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_17_i739_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3715[1] ), 
            .I2(GND_net), .I3(GND_net), .O(n1099_adj_5338));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i739_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut_adj_1726 (.I0(n20181), .I1(n6), .I2(n36845), .I3(\Ki[4] ), 
            .O(n20133[3]));   // verilog/motorControl.v(51[27:38])
    defparam i1_4_lut_adj_1726.LUT_INIT = 16'h9666;
    SB_LUT4 LessThan_25_i39_2_lut (.I0(n352[19]), .I1(n432[19]), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_5625));   // verilog/motorControl.v(55[23:39])
    defparam LessThan_25_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_25_i41_2_lut (.I0(n352[20]), .I1(n432[20]), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_5626));   // verilog/motorControl.v(55[23:39])
    defparam LessThan_25_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1727 (.I0(n20216[0]), .I1(n50890), .I2(\Ki[2] ), 
            .I3(\PID_CONTROLLER.integral_23__N_3715[20] ), .O(n20209));   // verilog/motorControl.v(51[27:38])
    defparam i1_4_lut_adj_1727.LUT_INIT = 16'h9666;
    SB_LUT4 LessThan_25_i45_2_lut (.I0(n352[22]), .I1(n432[22]), .I2(GND_net), 
            .I3(GND_net), .O(n45_adj_5627));   // verilog/motorControl.v(55[23:39])
    defparam LessThan_25_i45_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_25_i43_2_lut (.I0(n352[21]), .I1(n432[21]), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_5628));   // verilog/motorControl.v(55[23:39])
    defparam LessThan_25_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_25_i37_2_lut (.I0(n352[18]), .I1(n432[18]), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_5629));   // verilog/motorControl.v(55[23:39])
    defparam LessThan_25_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_17_i42_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3715[20] ), 
            .I2(GND_net), .I3(GND_net), .O(n62_adj_5567));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i42_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_25_i23_2_lut (.I0(n352[11]), .I1(n432[11]), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_5630));   // verilog/motorControl.v(55[23:39])
    defparam LessThan_25_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_25_i25_2_lut (.I0(n352[12]), .I1(n432[12]), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_5631));   // verilog/motorControl.v(55[23:39])
    defparam LessThan_25_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_25_i29_2_lut (.I0(n352[14]), .I1(n432[14]), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_5632));   // verilog/motorControl.v(55[23:39])
    defparam LessThan_25_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_25_i31_2_lut (.I0(n361), .I1(n432[15]), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_5633));   // verilog/motorControl.v(55[23:39])
    defparam LessThan_25_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_25_i35_2_lut (.I0(n352[17]), .I1(n432[17]), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_5634));   // verilog/motorControl.v(55[23:39])
    defparam LessThan_25_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_25_i11_2_lut (.I0(n352[5]), .I1(n432[5]), .I2(GND_net), 
            .I3(GND_net), .O(n11_adj_5635));   // verilog/motorControl.v(55[23:39])
    defparam LessThan_25_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_25_i13_2_lut (.I0(n352[6]), .I1(n432[6]), .I2(GND_net), 
            .I3(GND_net), .O(n13_adj_5636));   // verilog/motorControl.v(55[23:39])
    defparam LessThan_25_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i36955_4_lut (.I0(\Ki[0] ), .I1(\Ki[1] ), .I2(\PID_CONTROLLER.integral_23__N_3715[22] ), 
            .I3(\PID_CONTROLLER.integral_23__N_3715[21] ), .O(n20216[0]));   // verilog/motorControl.v(51[27:38])
    defparam i36955_4_lut.LUT_INIT = 16'h6ca0;
    SB_LUT4 LessThan_25_i27_2_lut (.I0(n352[13]), .I1(n432[13]), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_5637));   // verilog/motorControl.v(55[23:39])
    defparam LessThan_25_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_25_i15_2_lut (.I0(n352[7]), .I1(n432[7]), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_5638));   // verilog/motorControl.v(55[23:39])
    defparam LessThan_25_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_25_i33_2_lut (.I0(n352[16]), .I1(n432[16]), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_5639));   // verilog/motorControl.v(55[23:39])
    defparam LessThan_25_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_25_i9_2_lut (.I0(n352[4]), .I1(n432[4]), .I2(GND_net), 
            .I3(GND_net), .O(n9_adj_5640));   // verilog/motorControl.v(55[23:39])
    defparam LessThan_25_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_25_i17_2_lut (.I0(n352[8]), .I1(n432[8]), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_5641));   // verilog/motorControl.v(55[23:39])
    defparam LessThan_25_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_17_i95_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3715[22] ), 
            .I2(GND_net), .I3(GND_net), .O(n140_adj_5642));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i95_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut_adj_1728 (.I0(n36845), .I1(\Ki[2] ), .I2(\Ki[5] ), 
            .I3(\PID_CONTROLLER.integral_23__N_3715[21] ), .O(n63559));   // verilog/motorControl.v(51[27:38])
    defparam i1_4_lut_adj_1728.LUT_INIT = 16'h6ca0;
    SB_LUT4 LessThan_25_i19_2_lut (.I0(n367), .I1(n432[9]), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_5643));   // verilog/motorControl.v(55[23:39])
    defparam LessThan_25_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1729 (.I0(n36816), .I1(\Ki[3] ), .I2(\Ki[4] ), 
            .I3(\PID_CONTROLLER.integral_23__N_3715[20] ), .O(n63581));   // verilog/motorControl.v(51[27:38])
    defparam i1_4_lut_adj_1729.LUT_INIT = 16'h6ca0;
    SB_LUT4 LessThan_25_i21_2_lut (.I0(n352[10]), .I1(n432[10]), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_5644));   // verilog/motorControl.v(55[23:39])
    defparam LessThan_25_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i52164_4_lut (.I0(n21_adj_5644), .I1(n19_adj_5643), .I2(n17_adj_5641), 
            .I3(n9_adj_5640), .O(n67858));
    defparam i52164_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i37018_4_lut (.I0(n20216[0]), .I1(\Ki[2] ), .I2(n50890), .I3(\PID_CONTROLLER.integral_23__N_3715[20] ), 
            .O(n4_adj_5645));   // verilog/motorControl.v(51[27:38])
    defparam i37018_4_lut.LUT_INIT = 16'he8a0;
    SB_LUT4 i36957_4_lut (.I0(\Ki[0] ), .I1(\Ki[1] ), .I2(\PID_CONTROLLER.integral_23__N_3715[22] ), 
            .I3(\PID_CONTROLLER.integral_23__N_3715[21] ), .O(n50839));   // verilog/motorControl.v(51[27:38])
    defparam i36957_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i52156_4_lut (.I0(n27_adj_5637), .I1(n15_adj_5638), .I2(n13_adj_5636), 
            .I3(n11_adj_5635), .O(n67850));
    defparam i52156_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 LessThan_25_i12_3_lut (.I0(n432[7]), .I1(n432[16]), .I2(n33_adj_5639), 
            .I3(GND_net), .O(n12_adj_5646));   // verilog/motorControl.v(55[23:39])
    defparam LessThan_25_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1730 (.I0(n63559), .I1(\Ki[0] ), .I2(n140_adj_5642), 
            .I3(\PID_CONTROLLER.integral_23__N_3715[23] ), .O(n63561));   // verilog/motorControl.v(51[27:38])
    defparam i1_4_lut_adj_1730.LUT_INIT = 16'h695a;
    SB_LUT4 LessThan_25_i10_3_lut (.I0(n432[5]), .I1(n432[6]), .I2(n13_adj_5636), 
            .I3(GND_net), .O(n10_adj_5647));   // verilog/motorControl.v(55[23:39])
    defparam LessThan_25_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut_adj_1731 (.I0(n50839), .I1(n4_adj_5645), .I2(n63581), 
            .I3(GND_net), .O(n61017));   // verilog/motorControl.v(51[27:38])
    defparam i1_3_lut_adj_1731.LUT_INIT = 16'h9696;
    SB_LUT4 LessThan_25_i30_3_lut (.I0(n12_adj_5646), .I1(n432[17]), .I2(n35_adj_5634), 
            .I3(GND_net), .O(n30_adj_5648));   // verilog/motorControl.v(55[23:39])
    defparam LessThan_25_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53042_4_lut (.I0(n13_adj_5636), .I1(n11_adj_5635), .I2(n9_adj_5640), 
            .I3(n67871), .O(n68736));
    defparam i53042_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i53038_4_lut (.I0(n19_adj_5643), .I1(n17_adj_5641), .I2(n15_adj_5638), 
            .I3(n68736), .O(n68732));
    defparam i53038_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i54006_4_lut (.I0(n25_adj_5631), .I1(n23_adj_5630), .I2(n21_adj_5644), 
            .I3(n68732), .O(n69700));
    defparam i54006_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i53447_4_lut (.I0(n31_adj_5633), .I1(n29_adj_5632), .I2(n27_adj_5637), 
            .I3(n69700), .O(n69141));
    defparam i53447_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i54125_4_lut (.I0(n37_adj_5629), .I1(n35_adj_5634), .I2(n33_adj_5639), 
            .I3(n69141), .O(n69819));
    defparam i54125_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i36850_4_lut (.I0(n20181), .I1(n36845), .I2(n6), .I3(\Ki[4] ), 
            .O(n8_adj_5649));   // verilog/motorControl.v(51[27:38])
    defparam i36850_4_lut.LUT_INIT = 16'he8a0;
    SB_LUT4 i1_4_lut_adj_1732 (.I0(n6_adj_33), .I1(n8_adj_5649), .I2(n61017), 
            .I3(n63561), .O(n61429));   // verilog/motorControl.v(51[27:38])
    defparam i1_4_lut_adj_1732.LUT_INIT = 16'h6996;
    SB_LUT4 i53625_3_lut (.I0(n6_adj_5565), .I1(n432[10]), .I2(n21_adj_5644), 
            .I3(GND_net), .O(n69319));   // verilog/motorControl.v(55[23:39])
    defparam i53625_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_25_i16_3_lut (.I0(n432[9]), .I1(n432[21]), .I2(n43_adj_5628), 
            .I3(GND_net), .O(n16_adj_5651));   // verilog/motorControl.v(55[23:39])
    defparam LessThan_25_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_25_i8_3_lut (.I0(n432[4]), .I1(n432[8]), .I2(n17_adj_5641), 
            .I3(GND_net), .O(n8_adj_5652));   // verilog/motorControl.v(55[23:39])
    defparam LessThan_25_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_25_i24_3_lut (.I0(n16_adj_5651), .I1(n432[22]), .I2(n45_adj_5627), 
            .I3(GND_net), .O(n24_adj_5653));   // verilog/motorControl.v(55[23:39])
    defparam LessThan_25_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53626_3_lut (.I0(n69319), .I1(n432[11]), .I2(n23_adj_5630), 
            .I3(GND_net), .O(n69320));   // verilog/motorControl.v(55[23:39])
    defparam i53626_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52140_4_lut (.I0(n43_adj_5628), .I1(n25_adj_5631), .I2(n23_adj_5630), 
            .I3(n67858), .O(n67834));
    defparam i52140_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i53569_4_lut (.I0(n24_adj_5653), .I1(n8_adj_5652), .I2(n45_adj_5627), 
            .I3(n67830), .O(n69263));   // verilog/motorControl.v(55[23:39])
    defparam i53569_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i52601_3_lut (.I0(n69320), .I1(n432[12]), .I2(n25_adj_5631), 
            .I3(GND_net), .O(n68295));   // verilog/motorControl.v(55[23:39])
    defparam i52601_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53623_3_lut (.I0(n4_adj_5566), .I1(n432[13]), .I2(n27_adj_5637), 
            .I3(GND_net), .O(n69317));   // verilog/motorControl.v(55[23:39])
    defparam i53623_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53624_3_lut (.I0(n69317), .I1(n432[14]), .I2(n29_adj_5632), 
            .I3(GND_net), .O(n69318));   // verilog/motorControl.v(55[23:39])
    defparam i53624_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52152_4_lut (.I0(n33_adj_5639), .I1(n31_adj_5633), .I2(n29_adj_5632), 
            .I3(n67850), .O(n67846));
    defparam i52152_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i54044_4_lut (.I0(n30_adj_5648), .I1(n10_adj_5647), .I2(n35_adj_5634), 
            .I3(n67844), .O(n69738));   // verilog/motorControl.v(55[23:39])
    defparam i54044_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i52603_3_lut (.I0(n69318), .I1(n432[15]), .I2(n31_adj_5633), 
            .I3(GND_net), .O(n68297));   // verilog/motorControl.v(55[23:39])
    defparam i52603_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i54234_4_lut (.I0(n68297), .I1(n69738), .I2(n35_adj_5634), 
            .I3(n67846), .O(n69928));   // verilog/motorControl.v(55[23:39])
    defparam i54234_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i54235_3_lut (.I0(n69928), .I1(n432[18]), .I2(n37_adj_5629), 
            .I3(GND_net), .O(n69929));   // verilog/motorControl.v(55[23:39])
    defparam i54235_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i54186_3_lut (.I0(n69929), .I1(n432[19]), .I2(n39_adj_5625), 
            .I3(GND_net), .O(n69880));   // verilog/motorControl.v(55[23:39])
    defparam i54186_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52142_4_lut (.I0(n43_adj_5628), .I1(n41_adj_5626), .I2(n39_adj_5625), 
            .I3(n69819), .O(n67836));
    defparam i52142_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i53897_4_lut (.I0(n68295), .I1(n69263), .I2(n45_adj_5627), 
            .I3(n67834), .O(n69591));   // verilog/motorControl.v(55[23:39])
    defparam i53897_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i52609_3_lut (.I0(n69880), .I1(n432[20]), .I2(n41_adj_5626), 
            .I3(GND_net), .O(n68303));   // verilog/motorControl.v(55[23:39])
    defparam i52609_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i54102_4_lut (.I0(n68303), .I1(n69591), .I2(n45_adj_5627), 
            .I3(n67836), .O(n69796));   // verilog/motorControl.v(55[23:39])
    defparam i54102_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i54103_3_lut (.I0(n69796), .I1(n352[23]), .I2(n432[23]), .I3(GND_net), 
            .O(n69797));   // verilog/motorControl.v(55[23:39])
    defparam i54103_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i5956_3_lut (.I0(control_update), .I1(n405_adj_5603), .I2(n69797), 
            .I3(GND_net), .O(n11597));   // verilog/motorControl.v(20[7:21])
    defparam i5956_3_lut.LUT_INIT = 16'ha8a8;
    SB_LUT4 i29066_4_lut (.I0(PWMLimit[0]), .I1(n61943), .I2(n27629), 
            .I3(n11595), .O(n51[0]));   // verilog/motorControl.v(41[14] 62[8])
    defparam i29066_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 LessThan_10_i41_2_lut (.I0(IntegralLimit[20]), .I1(n130[20]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_5654));   // verilog/motorControl.v(46[12:34])
    defparam LessThan_10_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_10_i39_2_lut (.I0(IntegralLimit[19]), .I1(n130[19]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_5655));   // verilog/motorControl.v(46[12:34])
    defparam LessThan_10_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_10_i45_2_lut (.I0(IntegralLimit[22]), .I1(n130[22]), 
            .I2(GND_net), .I3(GND_net), .O(n45_adj_5656));   // verilog/motorControl.v(46[12:34])
    defparam LessThan_10_i45_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_10_i43_2_lut (.I0(IntegralLimit[21]), .I1(n130[21]), 
            .I2(GND_net), .I3(GND_net), .O(n43_adj_5657));   // verilog/motorControl.v(46[12:34])
    defparam LessThan_10_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i36878_2_lut_3_lut (.I0(\Kp[0] ), .I1(n55[23]), .I2(\Kp[1] ), 
            .I3(GND_net), .O(n50749));   // verilog/motorControl.v(51[18:24])
    defparam i36878_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 mult_17_i130_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3715[15] ), 
            .I2(GND_net), .I3(GND_net), .O(n192_adj_5335));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i130_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_2_lut_3_lut (.I0(\Kp[2] ), .I1(\Kp[0] ), .I2(\Kp[1] ), 
            .I3(GND_net), .O(n61580));
    defparam i2_2_lut_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 LessThan_10_i29_2_lut (.I0(IntegralLimit[14]), .I1(n130[14]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_5658));   // verilog/motorControl.v(46[12:34])
    defparam LessThan_10_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_10_i31_2_lut (.I0(IntegralLimit[15]), .I1(n130[15]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_5659));   // verilog/motorControl.v(46[12:34])
    defparam LessThan_10_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_10_i23_2_lut (.I0(IntegralLimit[11]), .I1(n130[11]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_5660));   // verilog/motorControl.v(46[12:34])
    defparam LessThan_10_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_10_i25_2_lut (.I0(IntegralLimit[12]), .I1(n130[12]), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_5661));   // verilog/motorControl.v(46[12:34])
    defparam LessThan_10_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_10_i37_2_lut (.I0(IntegralLimit[18]), .I1(n130[18]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_5662));   // verilog/motorControl.v(46[12:34])
    defparam LessThan_10_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 unary_minus_26_inv_0_i16_1_lut (.I0(PWMLimit[15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5682[15]));   // verilog/motorControl.v(56[22:31])
    defparam unary_minus_26_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 LessThan_10_i35_2_lut (.I0(IntegralLimit[17]), .I1(n130[17]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_5663));   // verilog/motorControl.v(46[12:34])
    defparam LessThan_10_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_10_i33_2_lut (.I0(IntegralLimit[16]), .I1(n130[16]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_5664));   // verilog/motorControl.v(46[12:34])
    defparam LessThan_10_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_10_i9_2_lut (.I0(IntegralLimit[4]), .I1(n130[4]), .I2(GND_net), 
            .I3(GND_net), .O(n9_adj_5665));   // verilog/motorControl.v(46[12:34])
    defparam LessThan_10_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_10_i17_2_lut (.I0(IntegralLimit[8]), .I1(n130[8]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_5666));   // verilog/motorControl.v(46[12:34])
    defparam LessThan_10_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_10_i19_2_lut (.I0(IntegralLimit[9]), .I1(n130[9]), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_5667));   // verilog/motorControl.v(46[12:34])
    defparam LessThan_10_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_10_i21_2_lut (.I0(IntegralLimit[10]), .I1(n130[10]), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_5668));   // verilog/motorControl.v(46[12:34])
    defparam LessThan_10_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_10_i11_2_lut (.I0(IntegralLimit[5]), .I1(n130[5]), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_5669));   // verilog/motorControl.v(46[12:34])
    defparam LessThan_10_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_10_i13_2_lut (.I0(IntegralLimit[6]), .I1(n130[6]), 
            .I2(GND_net), .I3(GND_net), .O(n13_adj_5670));   // verilog/motorControl.v(46[12:34])
    defparam LessThan_10_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_10_i15_2_lut (.I0(IntegralLimit[7]), .I1(n130[7]), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_5671));   // verilog/motorControl.v(46[12:34])
    defparam LessThan_10_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_10_i27_2_lut (.I0(IntegralLimit[13]), .I1(n130[13]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_5672));   // verilog/motorControl.v(46[12:34])
    defparam LessThan_10_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i51764_4_lut (.I0(n21_adj_5668), .I1(n19_adj_5667), .I2(n17_adj_5666), 
            .I3(n9_adj_5665), .O(n67458));
    defparam i51764_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i51751_4_lut (.I0(n27_adj_5672), .I1(n15_adj_5671), .I2(n13_adj_5670), 
            .I3(n11_adj_5669), .O(n67445));
    defparam i51751_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 LessThan_10_i12_3_lut (.I0(n130[7]), .I1(n130[16]), .I2(n33_adj_5664), 
            .I3(GND_net), .O(n12_adj_5673));   // verilog/motorControl.v(46[12:34])
    defparam LessThan_10_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_10_i10_3_lut (.I0(n130[5]), .I1(n130[6]), .I2(n13_adj_5670), 
            .I3(GND_net), .O(n10_adj_5674));   // verilog/motorControl.v(46[12:34])
    defparam LessThan_10_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_10_i30_3_lut (.I0(n12_adj_5673), .I1(n130[17]), .I2(n35_adj_5663), 
            .I3(GND_net), .O(n30_adj_5675));   // verilog/motorControl.v(46[12:34])
    defparam LessThan_10_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52694_4_lut (.I0(n13_adj_5670), .I1(n11_adj_5669), .I2(n9_adj_5665), 
            .I3(n67494), .O(n68388));
    defparam i52694_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i52682_4_lut (.I0(n19_adj_5667), .I1(n17_adj_5666), .I2(n15_adj_5671), 
            .I3(n68388), .O(n68376));
    defparam i52682_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i53919_4_lut (.I0(n25_adj_5661), .I1(n23_adj_5660), .I2(n21_adj_5668), 
            .I3(n68376), .O(n69613));
    defparam i53919_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i53270_4_lut (.I0(n31_adj_5659), .I1(n29_adj_5658), .I2(n27_adj_5672), 
            .I3(n69613), .O(n68964));
    defparam i53270_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i54104_4_lut (.I0(n37_adj_5662), .I1(n35_adj_5663), .I2(n33_adj_5664), 
            .I3(n68964), .O(n69798));
    defparam i54104_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 LessThan_10_i16_3_lut (.I0(n130[9]), .I1(n130[21]), .I2(n43_adj_5657), 
            .I3(GND_net), .O(n16_adj_5676));   // verilog/motorControl.v(46[12:34])
    defparam LessThan_10_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53557_3_lut (.I0(n6_adj_5564), .I1(n130[10]), .I2(n21_adj_5668), 
            .I3(GND_net), .O(n69251));   // verilog/motorControl.v(46[12:34])
    defparam i53557_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53558_3_lut (.I0(n69251), .I1(n130[11]), .I2(n23_adj_5660), 
            .I3(GND_net), .O(n69252));   // verilog/motorControl.v(46[12:34])
    defparam i53558_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_10_i8_3_lut (.I0(n130[4]), .I1(n130[8]), .I2(n17_adj_5666), 
            .I3(GND_net), .O(n8_adj_5677));   // verilog/motorControl.v(46[12:34])
    defparam LessThan_10_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_10_i24_3_lut (.I0(n16_adj_5676), .I1(n130[22]), .I2(n45_adj_5656), 
            .I3(GND_net), .O(n24_adj_5678));   // verilog/motorControl.v(46[12:34])
    defparam LessThan_10_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51540_4_lut (.I0(n43_adj_5657), .I1(n25_adj_5661), .I2(n23_adj_5660), 
            .I3(n67458), .O(n67234));
    defparam i51540_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i53246_4_lut (.I0(n24_adj_5678), .I1(n8_adj_5677), .I2(n45_adj_5656), 
            .I3(n67202), .O(n68940));   // verilog/motorControl.v(46[12:34])
    defparam i53246_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i52561_3_lut (.I0(n69252), .I1(n130[12]), .I2(n25_adj_5661), 
            .I3(GND_net), .O(n68255));   // verilog/motorControl.v(46[12:34])
    defparam i52561_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_10_i4_4_lut (.I0(n130[0]), .I1(n130[1]), .I2(IntegralLimit[1]), 
            .I3(IntegralLimit[0]), .O(n4_adj_5679));   // verilog/motorControl.v(46[12:34])
    defparam LessThan_10_i4_4_lut.LUT_INIT = 16'h0c8e;
    SB_LUT4 i53343_3_lut (.I0(n4_adj_5679), .I1(n130[13]), .I2(n27_adj_5672), 
            .I3(GND_net), .O(n69037));   // verilog/motorControl.v(46[12:34])
    defparam i53343_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53344_3_lut (.I0(n69037), .I1(n130[14]), .I2(n29_adj_5658), 
            .I3(GND_net), .O(n69038));   // verilog/motorControl.v(46[12:34])
    defparam i53344_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51737_4_lut (.I0(n33_adj_5664), .I1(n31_adj_5659), .I2(n29_adj_5658), 
            .I3(n67445), .O(n67431));
    defparam i51737_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i54131_4_lut (.I0(n30_adj_5675), .I1(n10_adj_5674), .I2(n35_adj_5663), 
            .I3(n67423), .O(n69825));   // verilog/motorControl.v(46[12:34])
    defparam i54131_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i52563_3_lut (.I0(n69038), .I1(n130[15]), .I2(n31_adj_5659), 
            .I3(GND_net), .O(n68257));   // verilog/motorControl.v(46[12:34])
    defparam i52563_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i54272_4_lut (.I0(n68257), .I1(n69825), .I2(n35_adj_5663), 
            .I3(n67431), .O(n69966));   // verilog/motorControl.v(46[12:34])
    defparam i54272_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i54273_3_lut (.I0(n69966), .I1(n130[18]), .I2(n37_adj_5662), 
            .I3(GND_net), .O(n69967));   // verilog/motorControl.v(46[12:34])
    defparam i54273_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i54239_3_lut (.I0(n69967), .I1(n130[19]), .I2(n39_adj_5655), 
            .I3(GND_net), .O(n69933));   // verilog/motorControl.v(46[12:34])
    defparam i54239_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51587_4_lut (.I0(n43_adj_5657), .I1(n41_adj_5654), .I2(n39_adj_5655), 
            .I3(n69798), .O(n67281));
    defparam i51587_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i53885_4_lut (.I0(n68255), .I1(n68940), .I2(n45_adj_5656), 
            .I3(n67234), .O(n69579));   // verilog/motorControl.v(46[12:34])
    defparam i53885_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i54174_3_lut (.I0(n69933), .I1(n130[20]), .I2(n41_adj_5654), 
            .I3(GND_net), .O(n40_adj_5680));   // verilog/motorControl.v(46[12:34])
    defparam i54174_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_16_i100_2_lut (.I0(\Kp[2] ), .I1(n55[4]), .I2(GND_net), 
            .I3(GND_net), .O(n147_adj_5333));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i100_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i53887_4_lut (.I0(n40_adj_5680), .I1(n69579), .I2(n45_adj_5656), 
            .I3(n67281), .O(n69581));   // verilog/motorControl.v(46[12:34])
    defparam i53887_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 unary_minus_26_inv_0_i17_1_lut (.I0(PWMLimit[16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5682[16]));   // verilog/motorControl.v(56[22:31])
    defparam unary_minus_26_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_17_i179_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3715[15] ), 
            .I2(GND_net), .I3(GND_net), .O(n265_adj_5331));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i179_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i51_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3715[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n74));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i51_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i4_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3715[1] ), 
            .I2(GND_net), .I3(GND_net), .O(n5_adj_5329));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i4_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i149_2_lut (.I0(\Kp[3] ), .I1(n55[4]), .I2(GND_net), 
            .I3(GND_net), .O(n220_adj_5328));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i149_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i167_2_lut (.I0(\Kp[3] ), .I1(n55[13]), .I2(GND_net), 
            .I3(GND_net), .O(n247));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i167_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i100_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3715[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n147_adj_5327));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i100_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i149_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3715[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n220));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i149_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i198_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3715[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n293_adj_5326));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i198_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i247_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3715[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n366_adj_5325));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i247_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i296_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3715[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n439_adj_5324));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i296_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i53888_3_lut (.I0(n69581), .I1(IntegralLimit[23]), .I2(n130[23]), 
            .I3(GND_net), .O(n155));   // verilog/motorControl.v(46[12:34])
    defparam i53888_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 mult_17_i345_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3715[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n512_adj_5323));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i345_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i394_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3715[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n585_adj_5322));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i394_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i590_2_lut (.I0(\Kp[12] ), .I1(n55[4]), .I2(GND_net), 
            .I3(GND_net), .O(n877_adj_5211));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i590_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_12_i41_2_lut (.I0(n130[20]), .I1(n182[20]), .I2(GND_net), 
            .I3(GND_net), .O(n41));   // verilog/motorControl.v(48[21:44])
    defparam LessThan_12_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 unary_minus_26_inv_0_i18_1_lut (.I0(PWMLimit[17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5682[17]));   // verilog/motorControl.v(56[22:31])
    defparam unary_minus_26_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_16_i216_2_lut (.I0(\Kp[4] ), .I1(n55[13]), .I2(GND_net), 
            .I3(GND_net), .O(n320));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i216_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_12_i39_2_lut (.I0(n130[19]), .I1(n182[19]), .I2(GND_net), 
            .I3(GND_net), .O(n39));   // verilog/motorControl.v(48[21:44])
    defparam LessThan_12_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_12_i45_2_lut (.I0(n130[22]), .I1(n182[22]), .I2(GND_net), 
            .I3(GND_net), .O(n45));   // verilog/motorControl.v(48[21:44])
    defparam LessThan_12_i45_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_17_i443_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3715[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n658_adj_5319));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i443_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_12_i43_2_lut (.I0(n130[21]), .I1(n182[21]), .I2(GND_net), 
            .I3(GND_net), .O(n43));   // verilog/motorControl.v(48[21:44])
    defparam LessThan_12_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_12_i37_2_lut (.I0(n130[18]), .I1(n182[18]), .I2(GND_net), 
            .I3(GND_net), .O(n37));   // verilog/motorControl.v(48[21:44])
    defparam LessThan_12_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_12_i29_2_lut (.I0(n130[14]), .I1(n182[14]), .I2(GND_net), 
            .I3(GND_net), .O(n29));   // verilog/motorControl.v(48[21:44])
    defparam LessThan_12_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_17_i492_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3715[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n731_adj_5318));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i492_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_12_i31_2_lut (.I0(n130[15]), .I1(n182[15]), .I2(GND_net), 
            .I3(GND_net), .O(n31_c));   // verilog/motorControl.v(48[21:44])
    defparam LessThan_12_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_12_i23_2_lut (.I0(n130[11]), .I1(n182[11]), .I2(GND_net), 
            .I3(GND_net), .O(n23));   // verilog/motorControl.v(48[21:44])
    defparam LessThan_12_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_12_i25_2_lut (.I0(n130[12]), .I1(n182[12]), .I2(GND_net), 
            .I3(GND_net), .O(n25));   // verilog/motorControl.v(48[21:44])
    defparam LessThan_12_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_12_i35_2_lut (.I0(n130[17]), .I1(n182[17]), .I2(GND_net), 
            .I3(GND_net), .O(n35));   // verilog/motorControl.v(48[21:44])
    defparam LessThan_12_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_12_i33_2_lut (.I0(n130[16]), .I1(n182[16]), .I2(GND_net), 
            .I3(GND_net), .O(n33_c));   // verilog/motorControl.v(48[21:44])
    defparam LessThan_12_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_12_i11_2_lut (.I0(n130[5]), .I1(n182[5]), .I2(GND_net), 
            .I3(GND_net), .O(n11));   // verilog/motorControl.v(48[21:44])
    defparam LessThan_12_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_12_i13_2_lut (.I0(n130[6]), .I1(n182[6]), .I2(GND_net), 
            .I3(GND_net), .O(n13));   // verilog/motorControl.v(48[21:44])
    defparam LessThan_12_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_12_i15_2_lut (.I0(n130[7]), .I1(n182[7]), .I2(GND_net), 
            .I3(GND_net), .O(n15));   // verilog/motorControl.v(48[21:44])
    defparam LessThan_12_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_12_i27_2_lut (.I0(n130[13]), .I1(n182[13]), .I2(GND_net), 
            .I3(GND_net), .O(n27));   // verilog/motorControl.v(48[21:44])
    defparam LessThan_12_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_12_i9_2_lut (.I0(n130[4]), .I1(n182[4]), .I2(GND_net), 
            .I3(GND_net), .O(n9));   // verilog/motorControl.v(48[21:44])
    defparam LessThan_12_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_12_i17_2_lut (.I0(n130[8]), .I1(n182[8]), .I2(GND_net), 
            .I3(GND_net), .O(n17));   // verilog/motorControl.v(48[21:44])
    defparam LessThan_12_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_12_i19_2_lut (.I0(n130[9]), .I1(n182[9]), .I2(GND_net), 
            .I3(GND_net), .O(n19_c));   // verilog/motorControl.v(48[21:44])
    defparam LessThan_12_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_12_i21_2_lut (.I0(n130[10]), .I1(n182[10]), .I2(GND_net), 
            .I3(GND_net), .O(n21));   // verilog/motorControl.v(48[21:44])
    defparam LessThan_12_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i52402_4_lut (.I0(n21), .I1(n19_c), .I2(n17), .I3(n9), .O(n68096));
    defparam i52402_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i52376_4_lut (.I0(n27), .I1(n15), .I2(n13), .I3(n11), .O(n68070));
    defparam i52376_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 mult_16_i265_2_lut (.I0(\Kp[5] ), .I1(n55[13]), .I2(GND_net), 
            .I3(GND_net), .O(n393));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i265_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i314_2_lut (.I0(\Kp[6] ), .I1(n55[13]), .I2(GND_net), 
            .I3(GND_net), .O(n466));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i314_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_12_i12_3_lut (.I0(n182[7]), .I1(n182[16]), .I2(n33_c), 
            .I3(GND_net), .O(n12_adj_5681));   // verilog/motorControl.v(48[21:44])
    defparam LessThan_12_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_12_i10_3_lut (.I0(n182[5]), .I1(n182[6]), .I2(n13), 
            .I3(GND_net), .O(n10_adj_5147));   // verilog/motorControl.v(48[21:44])
    defparam LessThan_12_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_12_i30_3_lut (.I0(n12_adj_5681), .I1(n182[17]), .I2(n35), 
            .I3(GND_net), .O(n30_adj_5146));   // verilog/motorControl.v(48[21:44])
    defparam LessThan_12_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52330_2_lut_4_lut (.I0(n130[21]), .I1(n182[21]), .I2(n130[9]), 
            .I3(n182[9]), .O(n68024));
    defparam i52330_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    
endmodule
//
// Verilog Description of module \quadrature_decoder(0) 
//

module \quadrature_decoder(0)  (ENCODER1_B_N_keep, n1779, ENCODER1_A_N_keep, 
            n1786, GND_net, n1788, n1790, n1792, n1794, n1796, 
            \encoder1_position[25] , \encoder1_position[24] , \encoder1_position[23] , 
            \encoder1_position[22] , \encoder1_position[21] , \encoder1_position[20] , 
            b_prev, \a_new[1] , \encoder1_position[19] , \encoder1_position[18] , 
            \encoder1_position[17] , \encoder1_position[16] , \encoder1_position[15] , 
            \encoder1_position[14] , \encoder1_position[13] , \encoder1_position[12] , 
            \encoder1_position[11] , \encoder1_position[10] , \encoder1_position[9] , 
            \encoder1_position[8] , \encoder1_position[7] , \encoder1_position[6] , 
            \encoder1_position[5] , \encoder1_position[4] , \encoder1_position[3] , 
            \encoder1_position[2] , n1822, n1824, VCC_net, n29649, 
            a_prev, n29614, n1784, position_31__N_3836, \b_new[1] , 
            n29402, debounce_cnt_N_3833) /* synthesis lattice_noprune=1 */ ;
    input ENCODER1_B_N_keep;
    input n1779;
    input ENCODER1_A_N_keep;
    output n1786;
    input GND_net;
    output n1788;
    output n1790;
    output n1792;
    output n1794;
    output n1796;
    output \encoder1_position[25] ;
    output \encoder1_position[24] ;
    output \encoder1_position[23] ;
    output \encoder1_position[22] ;
    output \encoder1_position[21] ;
    output \encoder1_position[20] ;
    output b_prev;
    output \a_new[1] ;
    output \encoder1_position[19] ;
    output \encoder1_position[18] ;
    output \encoder1_position[17] ;
    output \encoder1_position[16] ;
    output \encoder1_position[15] ;
    output \encoder1_position[14] ;
    output \encoder1_position[13] ;
    output \encoder1_position[12] ;
    output \encoder1_position[11] ;
    output \encoder1_position[10] ;
    output \encoder1_position[9] ;
    output \encoder1_position[8] ;
    output \encoder1_position[7] ;
    output \encoder1_position[6] ;
    output \encoder1_position[5] ;
    output \encoder1_position[4] ;
    output \encoder1_position[3] ;
    output \encoder1_position[2] ;
    output n1822;
    output n1824;
    input VCC_net;
    input n29649;
    output a_prev;
    input n29614;
    output n1784;
    output position_31__N_3836;
    output \b_new[1] ;
    input n29402;
    output debounce_cnt_N_3833;
    
    wire [1:0]b_new;   // vhdl/quadrature_decoder.vhd(40[9:14])
    wire [1:0]a_new;   // vhdl/quadrature_decoder.vhd(39[9:14])
    wire [31:0]n133;
    
    wire direction_N_3840, n52362, n52361, n52360, n52359, n52358, 
        n52357, n52356, n52355, n52354, n52353, n52352, n52351, 
        n52350, n52349, n52348, n52347, n52346, n52345, n52344, 
        n52343, n52342, n52341, n52340, n52339, n52338, n52337, 
        n52336, n52335, n52334, n52333, n52332;
    
    SB_DFF b_new_i0 (.Q(b_new[0]), .C(n1779), .D(ENCODER1_B_N_keep));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_DFF a_new_i0 (.Q(a_new[0]), .C(n1779), .D(ENCODER1_A_N_keep));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_LUT4 position_1940_add_4_33_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(n1786), .I3(n52362), .O(n133[31])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1940_add_4_33_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 position_1940_add_4_32_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(n1788), .I3(n52361), .O(n133[30])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1940_add_4_32_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1940_add_4_32 (.CI(n52361), .I0(direction_N_3840), 
            .I1(n1788), .CO(n52362));
    SB_LUT4 position_1940_add_4_31_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(n1790), .I3(n52360), .O(n133[29])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1940_add_4_31_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1940_add_4_31 (.CI(n52360), .I0(direction_N_3840), 
            .I1(n1790), .CO(n52361));
    SB_LUT4 position_1940_add_4_30_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(n1792), .I3(n52359), .O(n133[28])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1940_add_4_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1940_add_4_30 (.CI(n52359), .I0(direction_N_3840), 
            .I1(n1792), .CO(n52360));
    SB_LUT4 position_1940_add_4_29_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(n1794), .I3(n52358), .O(n133[27])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1940_add_4_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1940_add_4_29 (.CI(n52358), .I0(direction_N_3840), 
            .I1(n1794), .CO(n52359));
    SB_LUT4 position_1940_add_4_28_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(n1796), .I3(n52357), .O(n133[26])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1940_add_4_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1940_add_4_28 (.CI(n52357), .I0(direction_N_3840), 
            .I1(n1796), .CO(n52358));
    SB_LUT4 position_1940_add_4_27_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder1_position[25] ), .I3(n52356), .O(n133[25])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1940_add_4_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1940_add_4_27 (.CI(n52356), .I0(direction_N_3840), 
            .I1(\encoder1_position[25] ), .CO(n52357));
    SB_LUT4 position_1940_add_4_26_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder1_position[24] ), .I3(n52355), .O(n133[24])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1940_add_4_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1940_add_4_26 (.CI(n52355), .I0(direction_N_3840), 
            .I1(\encoder1_position[24] ), .CO(n52356));
    SB_LUT4 position_1940_add_4_25_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder1_position[23] ), .I3(n52354), .O(n133[23])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1940_add_4_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1940_add_4_25 (.CI(n52354), .I0(direction_N_3840), 
            .I1(\encoder1_position[23] ), .CO(n52355));
    SB_LUT4 position_1940_add_4_24_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder1_position[22] ), .I3(n52353), .O(n133[22])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1940_add_4_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1940_add_4_24 (.CI(n52353), .I0(direction_N_3840), 
            .I1(\encoder1_position[22] ), .CO(n52354));
    SB_LUT4 position_1940_add_4_23_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder1_position[21] ), .I3(n52352), .O(n133[21])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1940_add_4_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1940_add_4_23 (.CI(n52352), .I0(direction_N_3840), 
            .I1(\encoder1_position[21] ), .CO(n52353));
    SB_LUT4 position_1940_add_4_22_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder1_position[20] ), .I3(n52351), .O(n133[20])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1940_add_4_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 b_prev_I_0_48_2_lut (.I0(b_prev), .I1(\a_new[1] ), .I2(GND_net), 
            .I3(GND_net), .O(direction_N_3840));   // vhdl/quadrature_decoder.vhd(64[18:37])
    defparam b_prev_I_0_48_2_lut.LUT_INIT = 16'h9999;
    SB_CARRY position_1940_add_4_22 (.CI(n52351), .I0(direction_N_3840), 
            .I1(\encoder1_position[20] ), .CO(n52352));
    SB_LUT4 position_1940_add_4_21_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder1_position[19] ), .I3(n52350), .O(n133[19])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1940_add_4_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1940_add_4_21 (.CI(n52350), .I0(direction_N_3840), 
            .I1(\encoder1_position[19] ), .CO(n52351));
    SB_LUT4 position_1940_add_4_20_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder1_position[18] ), .I3(n52349), .O(n133[18])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1940_add_4_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1940_add_4_20 (.CI(n52349), .I0(direction_N_3840), 
            .I1(\encoder1_position[18] ), .CO(n52350));
    SB_LUT4 position_1940_add_4_19_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder1_position[17] ), .I3(n52348), .O(n133[17])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1940_add_4_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1940_add_4_19 (.CI(n52348), .I0(direction_N_3840), 
            .I1(\encoder1_position[17] ), .CO(n52349));
    SB_LUT4 position_1940_add_4_18_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder1_position[16] ), .I3(n52347), .O(n133[16])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1940_add_4_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1940_add_4_18 (.CI(n52347), .I0(direction_N_3840), 
            .I1(\encoder1_position[16] ), .CO(n52348));
    SB_LUT4 position_1940_add_4_17_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder1_position[15] ), .I3(n52346), .O(n133[15])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1940_add_4_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1940_add_4_17 (.CI(n52346), .I0(direction_N_3840), 
            .I1(\encoder1_position[15] ), .CO(n52347));
    SB_LUT4 position_1940_add_4_16_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder1_position[14] ), .I3(n52345), .O(n133[14])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1940_add_4_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1940_add_4_16 (.CI(n52345), .I0(direction_N_3840), 
            .I1(\encoder1_position[14] ), .CO(n52346));
    SB_LUT4 position_1940_add_4_15_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder1_position[13] ), .I3(n52344), .O(n133[13])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1940_add_4_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1940_add_4_15 (.CI(n52344), .I0(direction_N_3840), 
            .I1(\encoder1_position[13] ), .CO(n52345));
    SB_LUT4 position_1940_add_4_14_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder1_position[12] ), .I3(n52343), .O(n133[12])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1940_add_4_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1940_add_4_14 (.CI(n52343), .I0(direction_N_3840), 
            .I1(\encoder1_position[12] ), .CO(n52344));
    SB_LUT4 position_1940_add_4_13_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder1_position[11] ), .I3(n52342), .O(n133[11])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1940_add_4_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1940_add_4_13 (.CI(n52342), .I0(direction_N_3840), 
            .I1(\encoder1_position[11] ), .CO(n52343));
    SB_LUT4 position_1940_add_4_12_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder1_position[10] ), .I3(n52341), .O(n133[10])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1940_add_4_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1940_add_4_12 (.CI(n52341), .I0(direction_N_3840), 
            .I1(\encoder1_position[10] ), .CO(n52342));
    SB_LUT4 position_1940_add_4_11_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder1_position[9] ), .I3(n52340), .O(n133[9])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1940_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1940_add_4_11 (.CI(n52340), .I0(direction_N_3840), 
            .I1(\encoder1_position[9] ), .CO(n52341));
    SB_LUT4 position_1940_add_4_10_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder1_position[8] ), .I3(n52339), .O(n133[8])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1940_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1940_add_4_10 (.CI(n52339), .I0(direction_N_3840), 
            .I1(\encoder1_position[8] ), .CO(n52340));
    SB_LUT4 position_1940_add_4_9_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder1_position[7] ), .I3(n52338), .O(n133[7])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1940_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1940_add_4_9 (.CI(n52338), .I0(direction_N_3840), 
            .I1(\encoder1_position[7] ), .CO(n52339));
    SB_LUT4 position_1940_add_4_8_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder1_position[6] ), .I3(n52337), .O(n133[6])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1940_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1940_add_4_8 (.CI(n52337), .I0(direction_N_3840), 
            .I1(\encoder1_position[6] ), .CO(n52338));
    SB_LUT4 position_1940_add_4_7_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder1_position[5] ), .I3(n52336), .O(n133[5])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1940_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1940_add_4_7 (.CI(n52336), .I0(direction_N_3840), 
            .I1(\encoder1_position[5] ), .CO(n52337));
    SB_LUT4 position_1940_add_4_6_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder1_position[4] ), .I3(n52335), .O(n133[4])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1940_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1940_add_4_6 (.CI(n52335), .I0(direction_N_3840), 
            .I1(\encoder1_position[4] ), .CO(n52336));
    SB_LUT4 position_1940_add_4_5_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder1_position[3] ), .I3(n52334), .O(n133[3])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1940_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1940_add_4_5 (.CI(n52334), .I0(direction_N_3840), 
            .I1(\encoder1_position[3] ), .CO(n52335));
    SB_LUT4 position_1940_add_4_4_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder1_position[2] ), .I3(n52333), .O(n133[2])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1940_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1940_add_4_4 (.CI(n52333), .I0(direction_N_3840), 
            .I1(\encoder1_position[2] ), .CO(n52334));
    SB_LUT4 position_1940_add_4_3_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(n1822), .I3(n52332), .O(n133[1])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1940_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1940_add_4_3 (.CI(n52332), .I0(direction_N_3840), 
            .I1(n1822), .CO(n52333));
    SB_LUT4 position_1940_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(n1824), 
            .I3(VCC_net), .O(n133[0])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1940_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1940_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(n1824), 
            .CO(n52332));
    SB_DFF a_prev_40 (.Q(a_prev), .C(n1779), .D(n29649));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_DFF direction_42 (.Q(n1784), .C(n1779), .D(n29614));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_DFFE position_1940__i0 (.Q(n1824), .C(n1779), .E(position_31__N_3836), 
            .D(n133[0]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1940__i31 (.Q(n1786), .C(n1779), .E(position_31__N_3836), 
            .D(n133[31]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1940__i30 (.Q(n1788), .C(n1779), .E(position_31__N_3836), 
            .D(n133[30]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1940__i29 (.Q(n1790), .C(n1779), .E(position_31__N_3836), 
            .D(n133[29]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1940__i28 (.Q(n1792), .C(n1779), .E(position_31__N_3836), 
            .D(n133[28]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1940__i27 (.Q(n1794), .C(n1779), .E(position_31__N_3836), 
            .D(n133[27]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1940__i26 (.Q(n1796), .C(n1779), .E(position_31__N_3836), 
            .D(n133[26]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1940__i25 (.Q(\encoder1_position[25] ), .C(n1779), 
            .E(position_31__N_3836), .D(n133[25]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1940__i24 (.Q(\encoder1_position[24] ), .C(n1779), 
            .E(position_31__N_3836), .D(n133[24]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1940__i23 (.Q(\encoder1_position[23] ), .C(n1779), 
            .E(position_31__N_3836), .D(n133[23]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1940__i22 (.Q(\encoder1_position[22] ), .C(n1779), 
            .E(position_31__N_3836), .D(n133[22]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1940__i21 (.Q(\encoder1_position[21] ), .C(n1779), 
            .E(position_31__N_3836), .D(n133[21]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1940__i20 (.Q(\encoder1_position[20] ), .C(n1779), 
            .E(position_31__N_3836), .D(n133[20]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1940__i19 (.Q(\encoder1_position[19] ), .C(n1779), 
            .E(position_31__N_3836), .D(n133[19]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1940__i18 (.Q(\encoder1_position[18] ), .C(n1779), 
            .E(position_31__N_3836), .D(n133[18]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1940__i17 (.Q(\encoder1_position[17] ), .C(n1779), 
            .E(position_31__N_3836), .D(n133[17]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1940__i16 (.Q(\encoder1_position[16] ), .C(n1779), 
            .E(position_31__N_3836), .D(n133[16]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1940__i15 (.Q(\encoder1_position[15] ), .C(n1779), 
            .E(position_31__N_3836), .D(n133[15]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1940__i14 (.Q(\encoder1_position[14] ), .C(n1779), 
            .E(position_31__N_3836), .D(n133[14]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1940__i13 (.Q(\encoder1_position[13] ), .C(n1779), 
            .E(position_31__N_3836), .D(n133[13]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1940__i12 (.Q(\encoder1_position[12] ), .C(n1779), 
            .E(position_31__N_3836), .D(n133[12]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1940__i11 (.Q(\encoder1_position[11] ), .C(n1779), 
            .E(position_31__N_3836), .D(n133[11]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1940__i10 (.Q(\encoder1_position[10] ), .C(n1779), 
            .E(position_31__N_3836), .D(n133[10]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1940__i9 (.Q(\encoder1_position[9] ), .C(n1779), .E(position_31__N_3836), 
            .D(n133[9]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1940__i8 (.Q(\encoder1_position[8] ), .C(n1779), .E(position_31__N_3836), 
            .D(n133[8]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1940__i7 (.Q(\encoder1_position[7] ), .C(n1779), .E(position_31__N_3836), 
            .D(n133[7]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1940__i6 (.Q(\encoder1_position[6] ), .C(n1779), .E(position_31__N_3836), 
            .D(n133[6]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1940__i5 (.Q(\encoder1_position[5] ), .C(n1779), .E(position_31__N_3836), 
            .D(n133[5]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1940__i4 (.Q(\encoder1_position[4] ), .C(n1779), .E(position_31__N_3836), 
            .D(n133[4]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1940__i3 (.Q(\encoder1_position[3] ), .C(n1779), .E(position_31__N_3836), 
            .D(n133[3]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1940__i2 (.Q(\encoder1_position[2] ), .C(n1779), .E(position_31__N_3836), 
            .D(n133[2]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1940__i1 (.Q(n1822), .C(n1779), .E(position_31__N_3836), 
            .D(n133[1]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFF a_new_i1 (.Q(\a_new[1] ), .C(n1779), .D(a_new[0]));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_DFF b_new_i1 (.Q(\b_new[1] ), .C(n1779), .D(b_new[0]));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_DFF b_prev_41 (.Q(b_prev), .C(n1779), .D(n29402));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_LUT4 position_31__I_938_4_lut (.I0(a_prev), .I1(b_prev), .I2(\a_new[1] ), 
            .I3(\b_new[1] ), .O(position_31__N_3836));   // vhdl/quadrature_decoder.vhd(63[11:57])
    defparam position_31__I_938_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 debounce_cnt_I_937_4_lut (.I0(a_new[0]), .I1(b_new[0]), .I2(\a_new[1] ), 
            .I3(\b_new[1] ), .O(debounce_cnt_N_3833));   // vhdl/quadrature_decoder.vhd(53[8:58])
    defparam debounce_cnt_I_937_4_lut.LUT_INIT = 16'h7bde;
    
endmodule
//
// Verilog Description of module coms
//

module coms (n29895, VCC_net, \data_in_frame[5] , clk16MHz, GND_net, 
            n29892, \data_out_frame[6] , \data_out_frame[5] , \data_out_frame[4] , 
            \Ki[7] , n2873, \data_out_frame[8] , n58623, n58622, n29583, 
            \data_in_frame[21] , \data_out_frame[18] , \FRAME_MATCHER.i_31__N_2509 , 
            displacement, \Ki[6] , \FRAME_MATCHER.state[3] , \data_out_frame[25] , 
            n8, \data_out_frame[22] , \Ki[5] , \data_out_frame[23] , 
            n59477, \data_out_frame[19] , n53457, n58957, \Ki[4] , 
            n59223, \data_out_frame[16] , \data_out_frame[24] , n59452, 
            n59455, n58938, n29890, n25, n30, n26, n54456, n53546, 
            \data_out_frame[21] , \Ki[3] , \Ki[2] , \data_out_frame[20] , 
            \data_out_frame[17] , pwm_setpoint, n59241, n59406, n58978, 
            n29885, n29881, n29878, \data_in_frame[4] , n57914, n57916, 
            n57918, \Ki[1] , n29861, n29858, n29855, \Kp[15] , \Kp[14] , 
            n29851, \data_in_frame[3][6] , \data_in_frame[3][5] , \Kp[13] , 
            \Kp[12] , \Kp[11] , \Kp[10] , encoder0_position_scaled, 
            \Kp[9] , \data_out_frame[15] , n59124, \Kp[8] , n58621, 
            \data_out_frame[12] , \Kp[7] , \data_out_frame[13] , n59274, 
            n58620, \Kp[6] , \data_out_frame[14] , \Kp[5] , \Kp[4] , 
            n58671, \Kp[3] , \Kp[2] , n70020, reset, setpoint, \Kp[1] , 
            n2076, n25764, \data_in_frame[11] , IntegralLimit, n58619, 
            n54490, \data_out_frame[9] , n58495, n2217, n58618, n58617, 
            n58616, n58615, n58614, n58613, n58612, \data_out_frame[10] , 
            n58611, n58610, n58609, n58608, n58607, n58606, n58605, 
            n58604, \data_out_frame[11] , n58603, n58602, n58601, 
            n58600, n58599, n58598, n58597, n58596, n58595, n58594, 
            n58593, n58592, n58591, n58590, n58589, n58588, \data_in_frame[12] , 
            n30494, n28975, \byte_transmit_counter[2] , n58587, \data_in_frame[16] , 
            deadband, n58586, \byte_transmit_counter[1] , \byte_transmit_counter[0] , 
            n58585, n58887, \data_out_frame[7] , n36, n26143, n26376, 
            n58584, n58583, n58582, n58581, n58580, n58579, n58578, 
            n58577, n58576, n58575, n58574, n58573, n30510, n28959, 
            \data_in_frame[1] , n26210, n29786, \data_in_frame[23] , 
            n53515, n54620, n29771, \data_in_frame[0] , n29639, n29650, 
            \data_in_frame[0][3] , n29765, n29764, n57968, n29668, 
            n29674, n29756, \data_in_frame[0][6] , n59055, \FRAME_MATCHER.i[0] , 
            n43501, n163, rx_data, n59027, n22, neopxl_color, n7, 
            encoder1_position_scaled, n15, n15_adj_11, n19, \data_out_frame[1][1] , 
            \data_out_frame[3][1] , PWMLimit, n28, n375, n376, n4, 
            n58572, n58571, n58570, n58569, n58568, \data_in_frame[6] , 
            \data_in_frame[8] , n58567, n58566, n58565, n58564, n58496, 
            n58499, \data_out_frame[0][3] , \data_out_frame[1][3] , n28947, 
            \data_out_frame[3][3] , n58500, n28945, n58501, n58503, 
            \Ki[8] , \Ki[9] , \Ki[10] , \Ki[11] , \Ki[12] , \Ki[13] , 
            n58505, \Ki[14] , \Ki[15] , n58507, n58508, n58509, 
            n58510, n58511, n58512, n58513, n71165, n71003, n58514, 
            n58515, n58493, n58516, n58517, n28929, n28928, n58518, 
            n58519, n58520, \data_out_frame[1][6] , \data_out_frame[3][6] , 
            n29643, \FRAME_MATCHER.rx_data_ready_prev , n29642, n61932, 
            n29638, \data_out_frame[1][7] , \data_out_frame[3][7] , n29637, 
            current_limit, n29636, control_mode, n29635, n29634, n29633, 
            n29632, n29631, n29630, n29629, n29627, n29626, n29625, 
            n29624, n29623, n58521, \data_out_frame[1][0] , n58522, 
            n58523, n29621, n71225, n70991, \FRAME_MATCHER.i[3] , 
            \FRAME_MATCHER.i[4] , n8_adj_12, n29618, n29617, n29616, 
            n29615, n29613, n29612, n29608, n29607, n29606, n29605, 
            n29604, n29582, n29574, n29558, n29557, n29556, \Ki[0] , 
            \Kp[0] , n28921, n58524, n58525, n58526, n58527, n58528, 
            n58529, n58530, n58531, n58532, n58533, n58534, n58535, 
            n58536, n58492, n58537, n58538, n58539, n28903, n58540, 
            n58541, n58494, n58542, n58543, n58544, \FRAME_MATCHER.i[5] , 
            tx_active, n58545, n28895, n28894, n58546, \data_out_frame[0][4] , 
            n22734, \data_out_frame[3][4] , ID, \data_out_frame[0][2] , 
            n58670, n58669, n58668, n58667, n59299, \data_out_frame[26][2] , 
            n30439, n30438, n30437, n30421, \data_in_frame[0][0] , 
            n30391, n30305, n30273, n29898, n29901, n57890, n57886, 
            n30255, n29417, n29420, n29423, n29426, n57882, n29432, 
            n57878, \data_in_frame[17] , n57876, n57874, n57872, n57868, 
            n57864, n57860, n57856, n57852, \data_in_frame[18] , n57850, 
            n29930, \data_in_frame[7] , n30218, n29934, n29937, n29940, 
            n58666, n29943, n29946, n57846, n29955, n29958, n29961, 
            n29964, n30205, n29970, n29973, n29976, n30199, n30198, 
            n30030, n58665, n58106, n58108, n58060, n30043, n30046, 
            n30049, n30053, n30056, n30059, n30062, n57932, n57936, 
            n30072, n30169, n30075, n30079, n57996, n30110, n30154, 
            n29468, \data_out_frame[1][5] , n58664, n57842, n29474, 
            n57838, n57834, n58663, n57986, \data_in_frame[20] , n57980, 
            n29520, n29523, n57974, n29535, n29539, n29542, n29551, 
            \data_out_frame[27][2] , n29570, n58662, n58661, n58660, 
            n58659, n58658, n29575, n58657, n58506, n58656, n58655, 
            n58654, n58653, n58652, n58651, n58650, n58649, n58648, 
            n58647, n29578, n58646, n58645, n58644, n58643, n58642, 
            n58641, n58640, n58639, n58638, n58637, n58636, n58635, 
            n58634, n58633, n58632, n29410, n160, n58547, n29405, 
            n29403, n70997, n159, n58548, n58549, n58550, n58551, 
            n58552, n58553, n58504, n58498, n58554, n58555, n58556, 
            n58557, n58558, n58497, n58502, n58559, n58631, n58630, 
            n58629, n58628, n58560, n58561, n58562, n58563, LED_c, 
            DE_c, n58627, n58626, n58625, n58624, \pwm_counter[22] , 
            n45, \pwm_counter[21] , n43, n8_adj_13, n59638, \duty[3] , 
            \duty[0] , n260, n7_adj_14, n54113, n8_adj_15, n59430, 
            n40820, n455, n11597, n37330, n26282, n59007, n59215, 
            n58805, n59153, n25700, n58928, n87, n75, n33697, 
            n98, rx_data_ready, Kp_23__N_748, n28309, n28311, n367, 
            n19_adj_16, n361, n31, n28313, n43503, n18, n20, n230, 
            n155, \PID_CONTROLLER.integral_23__N_3715[1] , n161, n58418, 
            n59644, n33, n401, n4_adj_17, n26372, n28307, \current[7] , 
            \current[6] , \current[5] , \current[4] , \current[3] , 
            \current[2] , \current[1] , \current[0] , \current[15] , 
            n456, n27629, \current[11] , \current[10] , \current[9] , 
            \current[8] , n63789, n63793, n67140, n7_adj_18, n28385, 
            n70919, r_SM_Main, tx_o, r_Clock_Count, n4938, n29, 
            n23, \o_Rx_DV_N_3488[12] , \o_Rx_DV_N_3488[24] , n27, n29581, 
            \r_SM_Main_2__N_3536[1] , n59648, n60274, n6, tx_enable, 
            baudrate, r_Clock_Count_adj_29, \o_Rx_DV_N_3488[2] , \o_Rx_DV_N_3488[1] , 
            \o_Rx_DV_N_3488[3] , \o_Rx_DV_N_3488[4] , \o_Rx_DV_N_3488[5] , 
            \o_Rx_DV_N_3488[6] , \o_Rx_DV_N_3488[8] , \o_Rx_DV_N_3488[7] , 
            \r_Bit_Index[0] , n61449, n62163, \r_SM_Main_2__N_3446[1] , 
            r_Rx_Data, \r_SM_Main[1]_adj_27 , \r_SM_Main[2]_adj_28 , RX_N_2, 
            n25515, n62091, n60815, n62089, \o_Rx_DV_N_3488[0] , n4935, 
            n27901, n59702, n62513, n62417, n62465, n62401, n30420, 
            n54640, n30416, n62433, n30126, n30125, n30124, n30123, 
            n30122, n30121, n30120, n62481, n58684, n62497, n62449, 
            n27661) /* synthesis syn_module_defined=1 */ ;
    input n29895;
    input VCC_net;
    output [7:0]\data_in_frame[5] ;
    input clk16MHz;
    input GND_net;
    input n29892;
    output [7:0]\data_out_frame[6] ;
    output [7:0]\data_out_frame[5] ;
    output [7:0]\data_out_frame[4] ;
    output \Ki[7] ;
    input n2873;
    output [7:0]\data_out_frame[8] ;
    input n58623;
    input n58622;
    input n29583;
    output [7:0]\data_in_frame[21] ;
    output [7:0]\data_out_frame[18] ;
    output \FRAME_MATCHER.i_31__N_2509 ;
    input [23:0]displacement;
    output \Ki[6] ;
    output \FRAME_MATCHER.state[3] ;
    output [7:0]\data_out_frame[25] ;
    input n8;
    output [7:0]\data_out_frame[22] ;
    output \Ki[5] ;
    output [7:0]\data_out_frame[23] ;
    output n59477;
    output [7:0]\data_out_frame[19] ;
    input n53457;
    output n58957;
    output \Ki[4] ;
    output n59223;
    output [7:0]\data_out_frame[16] ;
    output [7:0]\data_out_frame[24] ;
    output n59452;
    input n59455;
    input n58938;
    input n29890;
    input n25;
    input n30;
    input n26;
    input n54456;
    output n53546;
    output [7:0]\data_out_frame[21] ;
    output \Ki[3] ;
    output \Ki[2] ;
    output [7:0]\data_out_frame[20] ;
    output [7:0]\data_out_frame[17] ;
    input [23:0]pwm_setpoint;
    input n59241;
    input n59406;
    input n58978;
    input n29885;
    input n29881;
    input n29878;
    output [7:0]\data_in_frame[4] ;
    input n57914;
    input n57916;
    input n57918;
    output \Ki[1] ;
    input n29861;
    input n29858;
    input n29855;
    output \Kp[15] ;
    output \Kp[14] ;
    input n29851;
    output \data_in_frame[3][6] ;
    output \data_in_frame[3][5] ;
    output \Kp[13] ;
    output \Kp[12] ;
    output \Kp[11] ;
    output \Kp[10] ;
    input [23:0]encoder0_position_scaled;
    output \Kp[9] ;
    output [7:0]\data_out_frame[15] ;
    output n59124;
    output \Kp[8] ;
    input n58621;
    output [7:0]\data_out_frame[12] ;
    output \Kp[7] ;
    output [7:0]\data_out_frame[13] ;
    output n59274;
    input n58620;
    output \Kp[6] ;
    output [7:0]\data_out_frame[14] ;
    output \Kp[5] ;
    output \Kp[4] ;
    input n58671;
    output \Kp[3] ;
    output \Kp[2] ;
    output n70020;
    input reset;
    output [23:0]setpoint;
    output \Kp[1] ;
    input n2076;
    input n25764;
    output [7:0]\data_in_frame[11] ;
    output [23:0]IntegralLimit;
    input n58619;
    output n54490;
    output [7:0]\data_out_frame[9] ;
    input n58495;
    input n2217;
    input n58618;
    input n58617;
    input n58616;
    input n58615;
    input n58614;
    input n58613;
    input n58612;
    output [7:0]\data_out_frame[10] ;
    input n58611;
    input n58610;
    input n58609;
    input n58608;
    input n58607;
    input n58606;
    input n58605;
    input n58604;
    output [7:0]\data_out_frame[11] ;
    input n58603;
    input n58602;
    input n58601;
    input n58600;
    input n58599;
    input n58598;
    input n58597;
    input n58596;
    input n58595;
    input n58594;
    input n58593;
    input n58592;
    input n58591;
    input n58590;
    input n58589;
    input n58588;
    output [7:0]\data_in_frame[12] ;
    input n30494;
    input n28975;
    output \byte_transmit_counter[2] ;
    input n58587;
    output [7:0]\data_in_frame[16] ;
    output [23:0]deadband;
    input n58586;
    output \byte_transmit_counter[1] ;
    output \byte_transmit_counter[0] ;
    input n58585;
    output n58887;
    output [7:0]\data_out_frame[7] ;
    output n36;
    output n26143;
    output n26376;
    input n58584;
    input n58583;
    input n58582;
    input n58581;
    input n58580;
    input n58579;
    input n58578;
    input n58577;
    input n58576;
    input n58575;
    input n58574;
    input n58573;
    input n30510;
    input n28959;
    output [7:0]\data_in_frame[1] ;
    input n26210;
    input n29786;
    output [7:0]\data_in_frame[23] ;
    output n53515;
    output n54620;
    input n29771;
    output [7:0]\data_in_frame[0] ;
    input n29639;
    input n29650;
    output \data_in_frame[0][3] ;
    input n29765;
    input n29764;
    input n57968;
    input n29668;
    input n29674;
    input n29756;
    output \data_in_frame[0][6] ;
    output n59055;
    output \FRAME_MATCHER.i[0] ;
    output n43501;
    output n163;
    output [7:0]rx_data;
    input n59027;
    output n22;
    output [23:0]neopxl_color;
    output n7;
    input [23:0]encoder1_position_scaled;
    input n15;
    input n15_adj_11;
    output n19;
    output \data_out_frame[1][1] ;
    output \data_out_frame[3][1] ;
    output [23:0]PWMLimit;
    input n28;
    input n375;
    input n376;
    output n4;
    input n58572;
    input n58571;
    input n58570;
    input n58569;
    input n58568;
    output [7:0]\data_in_frame[6] ;
    output [7:0]\data_in_frame[8] ;
    input n58567;
    input n58566;
    input n58565;
    input n58564;
    input n58496;
    input n58499;
    output \data_out_frame[0][3] ;
    output \data_out_frame[1][3] ;
    input n28947;
    output \data_out_frame[3][3] ;
    input n58500;
    input n28945;
    input n58501;
    input n58503;
    output \Ki[8] ;
    output \Ki[9] ;
    output \Ki[10] ;
    output \Ki[11] ;
    output \Ki[12] ;
    output \Ki[13] ;
    input n58505;
    output \Ki[14] ;
    output \Ki[15] ;
    input n58507;
    input n58508;
    input n58509;
    input n58510;
    input n58511;
    input n58512;
    input n58513;
    input n71165;
    input n71003;
    input n58514;
    input n58515;
    input n58493;
    input n58516;
    input n58517;
    input n28929;
    input n28928;
    input n58518;
    input n58519;
    input n58520;
    output \data_out_frame[1][6] ;
    output \data_out_frame[3][6] ;
    input n29643;
    output \FRAME_MATCHER.rx_data_ready_prev ;
    input n29642;
    output n61932;
    input n29638;
    output \data_out_frame[1][7] ;
    output \data_out_frame[3][7] ;
    input n29637;
    output [15:0]current_limit;
    input n29636;
    output [7:0]control_mode;
    input n29635;
    input n29634;
    input n29633;
    input n29632;
    input n29631;
    input n29630;
    input n29629;
    input n29627;
    input n29626;
    input n29625;
    input n29624;
    input n29623;
    input n58521;
    output \data_out_frame[1][0] ;
    input n58522;
    input n58523;
    input n29621;
    input n71225;
    input n70991;
    output \FRAME_MATCHER.i[3] ;
    output \FRAME_MATCHER.i[4] ;
    output n8_adj_12;
    input n29618;
    input n29617;
    input n29616;
    input n29615;
    input n29613;
    input n29612;
    input n29608;
    input n29607;
    input n29606;
    input n29605;
    input n29604;
    input n29582;
    input n29574;
    input n29558;
    input n29557;
    input n29556;
    output \Ki[0] ;
    output \Kp[0] ;
    input n28921;
    input n58524;
    input n58525;
    input n58526;
    input n58527;
    input n58528;
    input n58529;
    input n58530;
    input n58531;
    input n58532;
    input n58533;
    input n58534;
    input n58535;
    input n58536;
    input n58492;
    input n58537;
    input n58538;
    input n58539;
    input n28903;
    input n58540;
    input n58541;
    input n58494;
    input n58542;
    input n58543;
    input n58544;
    output \FRAME_MATCHER.i[5] ;
    output tx_active;
    input n58545;
    input n28895;
    input n28894;
    input n58546;
    output \data_out_frame[0][4] ;
    output n22734;
    output \data_out_frame[3][4] ;
    input [7:0]ID;
    output \data_out_frame[0][2] ;
    input n58670;
    input n58669;
    input n58668;
    input n58667;
    output n59299;
    output \data_out_frame[26][2] ;
    input n30439;
    input n30438;
    input n30437;
    input n30421;
    output \data_in_frame[0][0] ;
    input n30391;
    input n30305;
    input n30273;
    input n29898;
    input n29901;
    input n57890;
    input n57886;
    input n30255;
    input n29417;
    input n29420;
    input n29423;
    input n29426;
    input n57882;
    input n29432;
    input n57878;
    output [7:0]\data_in_frame[17] ;
    input n57876;
    input n57874;
    input n57872;
    input n57868;
    input n57864;
    input n57860;
    input n57856;
    input n57852;
    output [7:0]\data_in_frame[18] ;
    input n57850;
    input n29930;
    output [7:0]\data_in_frame[7] ;
    input n30218;
    input n29934;
    input n29937;
    input n29940;
    input n58666;
    input n29943;
    input n29946;
    input n57846;
    input n29955;
    input n29958;
    input n29961;
    input n29964;
    input n30205;
    input n29970;
    input n29973;
    input n29976;
    input n30199;
    input n30198;
    input n30030;
    input n58665;
    input n58106;
    input n58108;
    input n58060;
    input n30043;
    input n30046;
    input n30049;
    input n30053;
    input n30056;
    input n30059;
    input n30062;
    input n57932;
    input n57936;
    input n30072;
    input n30169;
    input n30075;
    input n30079;
    input n57996;
    input n30110;
    input n30154;
    input n29468;
    output \data_out_frame[1][5] ;
    input n58664;
    input n57842;
    input n29474;
    input n57838;
    input n57834;
    input n58663;
    input n57986;
    output [7:0]\data_in_frame[20] ;
    input n57980;
    input n29520;
    input n29523;
    input n57974;
    input n29535;
    input n29539;
    input n29542;
    input n29551;
    output \data_out_frame[27][2] ;
    input n29570;
    input n58662;
    input n58661;
    input n58660;
    input n58659;
    input n58658;
    input n29575;
    input n58657;
    input n58506;
    input n58656;
    input n58655;
    input n58654;
    input n58653;
    input n58652;
    input n58651;
    input n58650;
    input n58649;
    input n58648;
    input n58647;
    input n29578;
    input n58646;
    input n58645;
    input n58644;
    input n58643;
    input n58642;
    input n58641;
    input n58640;
    input n58639;
    input n58638;
    input n58637;
    input n58636;
    input n58635;
    input n58634;
    input n58633;
    input n58632;
    input n29410;
    input n160;
    input n58547;
    input n29405;
    input n29403;
    input n70997;
    output n159;
    input n58548;
    input n58549;
    input n58550;
    input n58551;
    input n58552;
    input n58553;
    input n58504;
    input n58498;
    input n58554;
    input n58555;
    input n58556;
    input n58557;
    input n58558;
    input n58497;
    input n58502;
    input n58559;
    input n58631;
    input n58630;
    input n58629;
    input n58628;
    input n58560;
    input n58561;
    input n58562;
    input n58563;
    output LED_c;
    output DE_c;
    input n58627;
    input n58626;
    input n58625;
    input n58624;
    input \pwm_counter[22] ;
    output n45;
    input \pwm_counter[21] ;
    output n43;
    output n8_adj_13;
    output n59638;
    input \duty[3] ;
    input \duty[0] ;
    input n260;
    output n7_adj_14;
    input n54113;
    output n8_adj_15;
    input n59430;
    output n40820;
    input n455;
    input n11597;
    output n37330;
    output n26282;
    output n59007;
    output n59215;
    output n58805;
    output n59153;
    output n25700;
    output n58928;
    input n87;
    output n75;
    output n33697;
    output n98;
    output rx_data_ready;
    output Kp_23__N_748;
    output n28309;
    output n28311;
    input n367;
    output n19_adj_16;
    input n361;
    output n31;
    output n28313;
    output n43503;
    input n18;
    output n20;
    input n230;
    input n155;
    output \PID_CONTROLLER.integral_23__N_3715[1] ;
    output n161;
    output n58418;
    output n59644;
    input n33;
    input n401;
    output n4_adj_17;
    input n26372;
    output n28307;
    input \current[7] ;
    input \current[6] ;
    input \current[5] ;
    input \current[4] ;
    input \current[3] ;
    input \current[2] ;
    input \current[1] ;
    input \current[0] ;
    input \current[15] ;
    input n456;
    output n27629;
    input \current[11] ;
    input \current[10] ;
    input \current[9] ;
    input \current[8] ;
    input n63789;
    output n63793;
    input n67140;
    output n7_adj_18;
    output n28385;
    output n70919;
    output [2:0]r_SM_Main;
    output tx_o;
    output [8:0]r_Clock_Count;
    input n4938;
    output n29;
    output n23;
    output \o_Rx_DV_N_3488[12] ;
    output \o_Rx_DV_N_3488[24] ;
    output n27;
    input n29581;
    input \r_SM_Main_2__N_3536[1] ;
    input n59648;
    input n60274;
    output n6;
    output tx_enable;
    input [31:0]baudrate;
    output [7:0]r_Clock_Count_adj_29;
    output \o_Rx_DV_N_3488[2] ;
    output \o_Rx_DV_N_3488[1] ;
    output \o_Rx_DV_N_3488[3] ;
    output \o_Rx_DV_N_3488[4] ;
    output \o_Rx_DV_N_3488[5] ;
    output \o_Rx_DV_N_3488[6] ;
    output \o_Rx_DV_N_3488[8] ;
    output \o_Rx_DV_N_3488[7] ;
    output \r_Bit_Index[0] ;
    output n61449;
    input n62163;
    input \r_SM_Main_2__N_3446[1] ;
    output r_Rx_Data;
    output \r_SM_Main[1]_adj_27 ;
    output \r_SM_Main[2]_adj_28 ;
    input RX_N_2;
    output n25515;
    input n62091;
    output n60815;
    output n62089;
    output \o_Rx_DV_N_3488[0] ;
    input n4935;
    output n27901;
    output n59702;
    output n62513;
    output n62417;
    output n62465;
    output n62401;
    input n30420;
    input n54640;
    input n30416;
    output n62433;
    input n30126;
    input n30125;
    input n30124;
    input n30123;
    input n30122;
    input n30121;
    input n30120;
    output n62481;
    input n58684;
    output n62497;
    output n62449;
    output n27661;
    
    wire clk16MHz /* synthesis SET_AS_NETWORK=clk16MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    
    wire n58673;
    wire [7:0]byte_transmit_counter;   // verilog/coms.v(105[12:33])
    
    wire n51015, n58672, n59281, Kp_23__N_1748, n37, n29688, n2, 
        n2_adj_4733;
    wire [31:0]\FRAME_MATCHER.state_31__N_2612 ;
    
    wire n2_adj_4734, n29689, n26327, n59212, n3, n59197, n58994, 
        n60824, n3_adj_4735, n53491, n3_adj_4736, n3_adj_4737, n29690, 
        n59382, n3_adj_4738, n53466, n59052, n3_adj_4739, n60844, 
        n54479, n25678, n54450, n10, n59490, n59074, n6_c, n29691, 
        n54114, n14, n10_adj_4740, n60980, n59332, n12, n54566, 
        n59149, n59353, n10_adj_4741, n26225, n59421;
    wire [31:0]\FRAME_MATCHER.i ;   // verilog/coms.v(118[11:12])
    
    wire n40660, n59448, n59484, n10_adj_4742, n3_adj_4743, n61721, 
        n6_adj_4744, n59356, n3_adj_4745, n26168, n58953, n59424, 
        n12_adj_4746, n8_adj_4747, n2_adj_4748, n29692, n29693, n59400, 
        n28_c, n2_adj_4749, n32, n59162, n30_adj_4750, n2_adj_4751, 
        n59030, n54525, n31_c, n2_adj_4752, n53928, n58987, n53717, 
        n29_c, n29586;
    wire [7:0]\data_in_frame[22] ;   // verilog/coms.v(99[12:25])
    
    wire n2_adj_4753, n60591, n29877, n29589, n2_adj_4754, n8_adj_4755, 
        n3_adj_4756, n2_adj_4757, n29592, n29694, n54570, n61136, 
        n3_adj_4758;
    wire [7:0]\data_in_frame[2] ;   // verilog/coms.v(99[12:25])
    
    wire n29695, n29696, n2_adj_4759, n6_adj_4760, n3_adj_4761, n29596, 
        n58126;
    wire [7:0]\data_in_frame[3] ;   // verilog/coms.v(99[12:25])
    
    wire n29845, n29599, n29841, n29838, n6_adj_4762, n25142, n3_adj_4763, 
        n54397, n58990, n8_adj_4764, n53626, n59218, n3_adj_4765, 
        n53644, n60897, n59403, n58893, n53735, n54568, n59344, 
        n59040, n12_adj_4766, n26180, n54552, n53897, n29697, n29698, 
        n29699, n6_adj_4767, n29700, n2_adj_4768, n29701, n54415, 
        n54529, n26739, n54220, n60541, n58809, n2_adj_4769, n2_adj_4770, 
        n26585, n6_adj_4771, n2_adj_4772, n53610, n59186, n53707, 
        n25650, n58944, n2_adj_4773, n2_adj_4774, n29702, n2_adj_4775, 
        n58975, n2_adj_4776, n2107, n59021, n10_adj_4777, n1673, 
        n58782, n59287, n18_c, n59112, n59442, n17, n29703, n59335, 
        n59012, n19_c, n25052, n10_adj_4778, n59171, n1510, n26049, 
        n14_adj_4779, n2_adj_4780, n1513, n2_adj_4781, n70022, n54413, 
        n2_adj_4782, n26206, n59089, n2_adj_4783, n29704, n26350, 
        n58680, n51014, n29705, n29706, n29835, n2_adj_4784, n29707, 
        n24, n29708, n26817, n14_adj_4785, n59308, n59024, n15_c, 
        n2_adj_4786, n2068;
    wire [23:0]n4760;
    
    wire n27674, n29832, n29709, n61441, n58679, n51013, n59329, 
        n22_c, n58935, n18_adj_4787, n26_adj_4788, n59168, n70024, 
        n2_adj_4789, n29710, n29711, n58678, n51012, n29712, n60743, 
        n2_adj_4790, n29713, n6_adj_4791, n23650, n2_adj_4792, n2_adj_4793, 
        n2_adj_4794, n2_adj_4795, n29829, n29714, n26849, n25872, 
        n12_adj_4796, n54432, n8_adj_4797, n59189, n71081, n66954, 
        n71150, n29826, n53640, n7_c, n23652, n14_adj_4798, n7_adj_4799;
    wire [7:0]tx_data;   // verilog/coms.v(108[13:20])
    
    wire n2_adj_4800, n6_adj_4801, n53933, n54434, n6_adj_4802, n16, 
        n17_adj_4803, n61261, n29715, n53583, n58984, n2_adj_4804, 
        n2_adj_4805, n2_adj_4806, n2_adj_4807, n2_adj_4808, n2_adj_4809, 
        n2_adj_4810, n2_adj_4811, n2_adj_4812, n2_adj_4813, n2_adj_4814, 
        n2_adj_4815, n2_adj_4816, n2_adj_4817, n2_adj_4818, n2_adj_4819, 
        n59338, n10_adj_4820, n3_adj_4821, n29716, n59384, n6_adj_4822, 
        n53449, n58677, n51011, n2_adj_4823, n2_adj_4824, n2_adj_4825, 
        n2_adj_4826, n2_adj_4827, n2_adj_4828, n2_adj_4829, n2_adj_4830, 
        n2_adj_4831, n2_adj_4832, n29717, n2_adj_4833, n2_adj_4834, 
        n2_adj_4835, n2_adj_4836, n2_adj_4837, n29718, n29719, n2_adj_4838, 
        n58676, n51010, n29823, n2_adj_4839, n29720, n29750, n2_adj_4840, 
        n58675, n51009, n58674, tx_transmit_N_3416, n29753, n2_adj_4841, 
        n29820, n29752, n26618, n1169, n12_adj_4842, n59296, n29749, 
        n6_adj_4843;
    wire [7:0]\data_in_frame[15] ;   // verilog/coms.v(99[12:25])
    
    wire n29748, n26_adj_4844, n29817, n29747, n29746, n29609, n25682, 
        n25611, n58867, n42, n26046, n58931, n40, n29813, n29810, 
        n71138, n2_adj_4845, n71141, n2_adj_4846, n2_adj_4847, n58864, 
        n41, n2_adj_4848, n58858, n59229, n39, n29745, n26563, 
        n1130, n44, n48, n29744, n29743, n29742, n58861, n58821, 
        n43_c, n8_adj_4849, n7_adj_4850, n4_c, n2_adj_4851, n2_adj_4852, 
        n29741, n8_adj_4853, n12_adj_4854, n2_adj_4855, n58873, n29807;
    wire [7:0]\data_in_frame[14] ;   // verilog/coms.v(99[12:25])
    
    wire n29740, n2_adj_4856, n2_adj_4857, n2_adj_4858, n58910, n6_adj_4859, 
        n26347, n1699, n29739, n2_adj_4860, n53470, n54430, n29751, 
        n29755, n26483, n29804, n26039, n2_adj_4861, n2_adj_4862;
    wire [7:0]\data_in_frame[19] ;   // verilog/coms.v(99[12:25])
    
    wire n58897, n26298, n29801, n29754, n8_adj_4863, n7_adj_4864, 
        n29798, n1312, n26022, n59350, n26649, n1835, n29738, 
        n29737, n29795, n6_adj_4865, n29736, n25614, n54458, n59067, 
        n54516, n58969, n58771, n59323, n29792, n10_adj_4866, n58941, 
        n59326, n14_adj_4867, n59436, n29735, n58972, n1191, n14_adj_4868, 
        n10_adj_4869, n29789, n59462, n1720, n53638, n36_adj_4870, 
        n58855, n25640, n59268, n34, n26_adj_4871, n40_adj_4872, 
        n58833, n38, n39_adj_4873, n29734, n59418, n59305, n37_adj_4874, 
        n29783, n29780, n59481, n29733, n29777, n29774, n58785, 
        n53489, n59244, n6_adj_4875, n64430, n64431, n71078, n58138;
    wire [7:0]\data_in_frame[0]_c ;   // verilog/coms.v(99[12:25])
    
    wire n29653, n29656, n59415, n58140, n58132, n64482, n64481, 
        n58830, n6_adj_4876, n59265, n58950, n10_adj_4877, n14_adj_4878, 
        n13, n15_adj_4879;
    wire [7:0]\data_in_frame[13] ;   // verilog/coms.v(99[12:25])
    
    wire n29732, n58802, n29731, n58883, n29730, n25685, n6_adj_4880, 
        n58880, n29729, n29728, n6_adj_4881, n12_adj_4882, n10_adj_4883, 
        n59253, n26716, n10_adj_4884, n10_adj_4885, \FRAME_MATCHER.i_31__N_2511 , 
        n29727, n29726, n132, n10_adj_4886, n67115, n40681, n3_adj_4887, 
        n29725, n161_c, n3468, n40817, n58720, n2_adj_4889, n2_adj_4890, 
        n2_adj_4891, n2_adj_4892, n2_adj_4893, n29724, n2_adj_4895, 
        n2_adj_4896, n28051, n64422, n64423, n64421, n64064, n29723, 
        n29722, n70895, n14_adj_4902, n2_adj_4903, n29721, n2_adj_4904, 
        n2_adj_4905, Kp_23__N_878, n58818, n7_adj_4906, n2_adj_4907, 
        n2_adj_4908, n2_adj_4909, n2_adj_4910, n1, n2_adj_4911, n64382, 
        n58731, n58752, n30145, n64472, n2_adj_4912, n29687, n64473, 
        n2_adj_4913, n2_adj_4914, n29686, n29685, n64458, n29684, 
        n29683, n29682, n2_adj_4915, n64457, n64484, n64485, n29681, 
        n2_adj_4916, n2_adj_4917, n2_adj_4918, n64401, n64400, n29680, 
        n2_adj_4919, n64487, n64488, n30102, n64368, n2_adj_4920, 
        n64367, n69187, n2_adj_4921, n2_adj_4922, n2_adj_4923, n2_adj_4924, 
        n2_adj_4925, n2_adj_4926, n2_adj_4927, n2_adj_4928, n2_adj_4929, 
        n2_adj_4930, n28045, n30099, n64404, n64405, n30095, n64403, 
        n2_adj_4931, n70961, n67143, n2_adj_4932, n71207, n70955, 
        n69199, n28043, n64395, n2_adj_4933, n2_adj_4934, n64396, 
        n64394, n2_adj_4935, n2_adj_4936, n64547, n64548, n2_adj_4937, 
        n30092, n2_adj_4938, n64554, n64553, n70967, n66934, n2_adj_4939, 
        n2_adj_4940, n2_adj_4941, n64529, n64530, n64437, n2_adj_4942, 
        n2_adj_4943, n64436, n2_adj_4944, n64419, n28104, n64420, 
        n64418, n2_adj_4945, n30089, n2_adj_4946, n2_adj_4947, n2_adj_4948, 
        n30085, n70973, n67162, n69121, n70907, n69122, n70883, 
        n71219, n69205, n70925, n30082, \FRAME_MATCHER.i_31__N_2514 , 
        n1951, n60750, n4452, n8_adj_4949, n22687, n63955, n26967, 
        n3303, \FRAME_MATCHER.i_31__N_2512 , n2060, n1954, n1957, 
        n63978, n61412, n57728, n1955, n25463, n20350, n2049, 
        n771, \FRAME_MATCHER.i_31__N_2508 , n2048, n8_adj_4950, n29504, 
        n6_adj_4951, n29501, n25388, n25474, \FRAME_MATCHER.i_31__N_2507 , 
        n27541, n60982, n25468, n26964;
    wire [7:0]\data_in[2] ;   // verilog/coms.v(98[12:19])
    wire [7:0]\data_in[1] ;   // verilog/coms.v(98[12:19])
    
    wire n25538;
    wire [7:0]\data_in[3] ;   // verilog/coms.v(98[12:19])
    
    wire n18_adj_4953, n29569;
    wire [7:0]\data_in[0] ;   // verilog/coms.v(98[12:19])
    
    wire n20_c, n29559, n29555, n29554, n29498, n29534, n15_adj_4954, 
        n2_adj_4955, n25380, n10_adj_4956, n64186, n9, n25493, n2_adj_4957, 
        n2_adj_4958, n2_adj_4959, n2_adj_4960, n2_adj_4961, n2_adj_4962, 
        n2_adj_4963, n2_adj_4964, n2_adj_4965, n2_adj_4966, n2_adj_4967, 
        n2_adj_4968, n2_adj_4969, n2_adj_4970, n2_adj_4971, n2_adj_4972, 
        n2_adj_4973, n2_adj_4974, n2_adj_4975, n29495, n2_adj_4976, 
        n2_adj_4977, n2_adj_4978, n2_adj_4979, n2_adj_4980, n10_adj_4981, 
        n14_adj_4982, n25487, n16_adj_4983, n22_adj_4984, n29492, 
        n20_adj_4985, n29489, n24_adj_4986, n16_adj_4987, n17_adj_4988, 
        n16_adj_4989, n17_adj_4990, n27978, \FRAME_MATCHER.i_31__N_2513 , 
        n33690, n29486, n10_adj_4991;
    wire [2:0]r_SM_Main_2__N_3545;
    
    wire n43563, n1_adj_4992, n61225, n42843, n6_adj_4993, n2_adj_4994, 
        n71283, n2_adj_4995, n29483, n28830, n2_adj_4996, n2_adj_4997, 
        n67065, n2_adj_4998, n67066, n27980, n27982, n2_adj_4999, 
        n59010, n27984, n27986, n27988, n27990, n27992, n27994, 
        n27996, n27998, n28000, n28002, n28004, n28006, n28008, 
        n28010, n28012, n28014, n28016, n28018, n28020, n28022, 
        n28024, n28026, n28028, n28030, n28032, n28034, n28036, 
        n28038, n28040, n2_adj_5000, n2_adj_5001, n2_adj_5002, n2_adj_5003, 
        n2_adj_5004, n2_adj_5005, n2_adj_5006, n2_adj_5007, n53570, 
        n25906, n54511, n2_adj_5008, n2_adj_5009, n2_adj_5010, n2_adj_5011;
    wire [7:0]\data_out_frame[26] ;   // verilog/coms.v(100[12:26])
    
    wire n58467, n35423, n6_adj_5012, n59003, n58472, n58473, n58470, 
        n58474, n30436, n30435, n30434, n29369, n30432, n30428, 
        n30427, n29372, n29375, n29378, n22_adj_5013, n29384, n29387, 
        n29390, n30396, n29393, n30394, n30393, n29396, n30390, 
        n30389, n30388, n29399, n30373, n30349, n30322, n30321, 
        n30320, n30314, n30307, n30306, n30304, n30303, n30302, 
        n30301, n30300, n30299, n30298, n30297, n30296, n30295, 
        n30294, n30293, n30292, n30291, n30290, n30289, n30288, 
        n30287, n30286, n30285, n30284, n30283, n30282, n30281, 
        n30280, n30279, n30278, n30277, n30276, n30275, n30274, 
        n29407, n30271, n30268, n30265, n30264, n29904, n29908, 
        n30260, n30257, n29911, n29914, n29918, n30227, n29921, 
        n29924, n29927, n2_adj_5014, n58092;
    wire [7:0]\data_in_frame[7]_c ;   // verilog/coms.v(99[12:25])
    
    wire n58086, n29979;
    wire [7:0]\data_in_frame[9] ;   // verilog/coms.v(99[12:25])
    
    wire n29982, n29985, n29989, n29992, n29995, n29998, n30001, 
        n30004;
    wire [7:0]\data_in_frame[10] ;   // verilog/coms.v(99[12:25])
    
    wire n30007, n30010, n30013, n30017, n30020, n30023, n30027, 
        n2_adj_5015, n2_adj_5016, n2_adj_5017, n30106, n30098, n71039, 
        n67165, n71042, n4_adj_5018, n4_adj_5019, n58468, n58475, 
        n58000, n58476;
    wire [7:0]\data_out_frame[27] ;   // verilog/coms.v(100[12:26])
    
    wire n58477, n58478, n58479, n2_adj_5020, n70913, n67141, n58471, 
        n71189, n70931, n69115, n2_adj_5021, n64466, n58480, n64467, 
        n58469, n58481, n64494, n64493, n67049, n64413, n2_adj_5022, 
        n2_adj_5023, n2_adj_5024, n64414, n2_adj_5025, n64412, n58482, 
        n2_adj_5026, n70871, n70859, n14_adj_5027, n7_adj_5028, n71036, 
        n71030, n9_adj_5029, n28337, n40663, n29406, n92, n40696, 
        n40711, n7_adj_5030, n7_adj_5031, n7_adj_5032, n7_adj_5033, 
        n64407, n64408, n64406, n3_adj_5034, n1_adj_5035, n1_adj_5036, 
        n1_adj_5037, n1_adj_5038, n1_adj_5039, n1_adj_5040, n1_adj_5041, 
        n28833, n5, n28832, n26865, n71255, n70889, n1_adj_5042, 
        n2_adj_5043, n2_adj_5044, n70901, n2_adj_5045, n2_adj_5046, 
        n28304, n52300, n67044, n52299, n67043, n52298, n67042, 
        n52297, n67037, n52296, n67036, n52295, n67028, n52294, 
        n67003, n52293, n66999, n52292, n66998, n52291, n66997, 
        n52290, n66993, n52289, n66992, n52288, n66973, n52287, 
        n66972, n52286, n66967, n52285, n66966, n52284, n66962, 
        n52283, n66959, n52282, n66955, n52281, n66953, n52280, 
        n66952, n52279, n66951, n52278, n66944, n52277, n66942, 
        n52276, n66941, n52275, n66940, n52274, n66939, n52273, 
        n66938, n52272, n66937, n52271, n66936, n52270, n66935;
    wire [31:0]n133;
    
    wire n4_adj_5048, n5_adj_5049, n71024, n25815, n71027, n54460, 
        n54116, n54572, n26689, n59226, n63809, n59232, n59380, 
        n54447, n63815, n61135, n59183, n61398, n47954, n59235, 
        n59379, n54411, n63951, n63743, n59341, n61410, n53713, 
        Kp_23__N_1551, n59409, n59284, n53503, n59427, n10_adj_5050, 
        n26239, n25744, n53442, n8_adj_5051, n58760, n25979, n7_adj_5053, 
        n26435, n59368, n59083, n25112, n54513, n54630, n7_adj_5054, 
        n59046, n58812, n59259, n25843, n59371, n59018, n22_adj_5055, 
        n28_adj_5056, n53511, n26_adj_5057, n54588, n27_c, n59092, 
        n58981, n25_adj_5058, n26605, n25853, n26359, n54527, n59459, 
        n59097, n14_adj_5059, n9_adj_5060, n59374, n59134, n53460, 
        n59206, n63675, n63677, n59174, n59060, n59146, Kp_23__N_1389, 
        n63687, n59137, n63689, n58960, n63695, n61382, n54155, 
        n59439, n63701, n59471, n63707, n26755, n25724, n10_adj_5061, 
        n58851, n26639, n61117, n59165, n60961, n54033, n10_adj_5062, 
        n54475, Kp_23__N_1607, n58925, n6_adj_5063, n59033, n26085, 
        n59106, n5_adj_5064, n54473, n26134, n54452, n59143, n6_adj_5065, 
        n26438, n59199, n59194, n6_adj_5066, n54518, n54417, n5_adj_5067, 
        n59080, n61279, n10_adj_5068, n59100, n54520, n63929, n59109, 
        n63935, n59256, n58894, n59412, n63939, n70018, n26633, 
        n63945, n63897, n63899, n140, n59121, n63903, n59064, 
        n58792, n63909, n59474, n59397, n63915, n54468, n59316, 
        n6_adj_5070, Kp_23__N_1271, n25925, n25807, n4_adj_5072, n59177, 
        n10_adj_5073, n59180, n63857, n63859, Kp_23__N_669, n63863, 
        n59468, n59391, n63869, n58914, n25818, n63875, n61424, 
        n63881, n54436, n63749, n58870, n53832, n25987, n6_adj_5074, 
        n59278, n63629, n59156, n63635, n58947, n59271, n6_adj_5075, 
        n59000, n10_adj_5076, n59320, n58799, n58836, n26774, n54002, 
        n3_adj_5077, n59394, n10_adj_5078, n14_adj_5079, n10_adj_5080, 
        n25661, n26411, n59140, n6_adj_5081, n59362, n23833, n25751, 
        n58901, n6_adj_5082, n26608, n23922, n70014, n63647, n59487, 
        n26680, n63653, n26426, n54404, n61299, n26219, Kp_23__N_1080, 
        n59302, n59247, n10_adj_5083, n6_adj_5084, n58848, n59103, 
        n10_adj_5085, n60903, n59086, n10_adj_5086, n53031, n64050, 
        n26288, n23926, n25758, n63719, n59077, n61271, n8_adj_5087, 
        n63723, n63725, n6_adj_5088, n25953, n63727, n8_adj_5089, 
        n63729, n63731, n63837, n5_adj_5090, n63825, n58789, n58815, 
        n58876, n64048, n63831, n61285, n63733, n63801, n63807, 
        n63843, n61908, n63739, n25786, n26251, n59290, n10_adj_5091, 
        n26316, n58824, n25860, n26343, Kp_23__N_974, n25869, n58827, 
        n12_adj_5092, n58922, n6_adj_5093, n25878, Kp_23__N_993, n7_adj_5094, 
        n6_adj_5095, n59202, n26544, n58997, n63755, n8_adj_5096, 
        n58755, n59365, n6_adj_5097, n10_adj_5098, n64040, n25892, 
        n64182, n26_adj_5099, n64184, n54308, n25_adj_5100, n25455, 
        n67106, n12_adj_5101, n10_adj_5102, n11, n9_adj_5103, n6_adj_5104, 
        n22_adj_5105, n70026, n1_adj_5106, n27_adj_5107, n67093, n26_adj_5108, 
        n17_adj_5109, n63981, n27_adj_5110, n44_adj_5111, n42_adj_5112, 
        n29_adj_5113, n43_adj_5114, n41_adj_5115, n23_c, n40_adj_5116, 
        n39_adj_5117, n50, n45_adj_5118, n71258, n64471, n71018, 
        n71252, n71246, n64383, n64480, n71240, n70943, n71012, 
        n71015, n71234, n71006, n71009, n71228, n70949, n71216, 
        n59250, n58842, n71204, n70970, n26368, n70964, n70958, 
        n71198, n70937, n70952, n71186, n70946, n70940, n70934, 
        n33_adj_5126, n33693, n70928, n70922, n70916, n70910, n70904, 
        n70898, n70892, n70886, n70880, n70868, n70856, n27233;
    
    SB_DFFE data_in_frame_0___i46 (.Q(\data_in_frame[5] [5]), .C(clk16MHz), 
            .E(VCC_net), .D(n29895));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 add_1097_9_lut (.I0(n58672), .I1(byte_transmit_counter[7]), 
            .I2(GND_net), .I3(n51015), .O(n58673)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1097_9_lut.LUT_INIT = 16'h8228;
    SB_DFFE data_in_frame_0___i45 (.Q(\data_in_frame[5] [4]), .C(clk16MHz), 
            .E(VCC_net), .D(n29892));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i3_4_lut_3_lut_4_lut (.I0(\data_out_frame[6] [2]), .I1(\data_out_frame[5] [7]), 
            .I2(\data_out_frame[6] [3]), .I3(\data_out_frame[4] [2]), .O(n59281));   // verilog/coms.v(77[16:43])
    defparam i3_4_lut_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i15682_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n37), .I2(\data_in_frame[5] [7]), 
            .I3(\Ki[7] ), .O(n29688));   // verilog/coms.v(148[4] 304[11])
    defparam i15682_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFFESS data_out_frame_0___i67 (.Q(\data_out_frame[8] [2]), .C(clk16MHz), 
            .E(n2873), .D(n2), .S(n58623));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i68 (.Q(\data_out_frame[8] [3]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4733), .S(n58622));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i176 (.Q(\data_in_frame[21] [7]), .C(clk16MHz), 
           .D(n29583));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_775_Select_145_i2_4_lut (.I0(\data_out_frame[18] [1]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[17]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4734));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_145_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i15683_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n37), .I2(\data_in_frame[5] [6]), 
            .I3(\Ki[6] ), .O(n29689));   // verilog/coms.v(148[4] 304[11])
    defparam i15683_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 select_775_Select_223_i3_4_lut (.I0(n26327), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(n59212), .I3(\data_out_frame[25] [6]), .O(n3));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_223_i3_4_lut.LUT_INIT = 16'h8448;
    SB_LUT4 i1_2_lut (.I0(\data_out_frame[25] [5]), .I1(n59197), .I2(GND_net), 
            .I3(GND_net), .O(n59212));
    defparam i1_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 select_775_Select_222_i3_4_lut (.I0(n58994), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(n59212), .I3(n60824), .O(n3_adj_4735));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_222_i3_4_lut.LUT_INIT = 16'h8448;
    SB_LUT4 select_775_Select_221_i3_3_lut (.I0(n53491), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(n58994), .I3(GND_net), .O(n3_adj_4736));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_221_i3_3_lut.LUT_INIT = 16'h8484;
    SB_LUT4 select_775_Select_220_i3_4_lut (.I0(n53491), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(n8), .I3(\data_out_frame[22] [6]), .O(n3_adj_4737));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_220_i3_4_lut.LUT_INIT = 16'h8448;
    SB_LUT4 i15684_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n37), .I2(\data_in_frame[5] [5]), 
            .I3(\Ki[5] ), .O(n29690));   // verilog/coms.v(148[4] 304[11])
    defparam i15684_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 select_775_Select_219_i3_2_lut (.I0(n59382), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4738));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_219_i3_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 select_775_Select_218_i3_4_lut (.I0(n53466), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(n59052), .I3(\data_out_frame[23] [0]), .O(n3_adj_4739));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_218_i3_4_lut.LUT_INIT = 16'h8448;
    SB_LUT4 i4_4_lut (.I0(n60844), .I1(n54479), .I2(n25678), .I3(n54450), 
            .O(n10));
    defparam i4_4_lut.LUT_INIT = 16'h9669;
    SB_LUT4 i5_3_lut (.I0(n59477), .I1(n10), .I2(\data_out_frame[19] [0]), 
            .I3(GND_net), .O(n59490));
    defparam i5_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i4_4_lut_adj_1057 (.I0(n53457), .I1(n59074), .I2(n59490), 
            .I3(n6_c), .O(n58957));
    defparam i4_4_lut_adj_1057.LUT_INIT = 16'h6996;
    SB_LUT4 i15685_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n37), .I2(\data_in_frame[5] [4]), 
            .I3(\Ki[4] ), .O(n29691));   // verilog/coms.v(148[4] 304[11])
    defparam i15685_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i6_4_lut (.I0(n59490), .I1(n54114), .I2(n59223), .I3(\data_out_frame[16] [4]), 
            .O(n14));
    defparam i6_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut (.I0(\data_out_frame[18] [5]), .I1(n14), .I2(n10_adj_4740), 
            .I3(n60980), .O(n53466));
    defparam i7_4_lut.LUT_INIT = 16'h9669;
    SB_LUT4 i5_4_lut (.I0(\data_out_frame[23] [1]), .I1(n59332), .I2(\data_out_frame[24] [7]), 
            .I3(n53466), .O(n12));
    defparam i5_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1058 (.I0(n54566), .I1(n12), .I2(n58957), .I3(n59149), 
            .O(n59382));
    defparam i6_4_lut_adj_1058.LUT_INIT = 16'h9669;
    SB_LUT4 i4_4_lut_adj_1059 (.I0(n59452), .I1(n59353), .I2(\data_out_frame[16] [5]), 
            .I3(n59455), .O(n10_adj_4741));
    defparam i4_4_lut_adj_1059.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut (.I0(n26225), .I1(n59421), .I2(n10_adj_4741), .I3(n58938), 
            .O(n59477));
    defparam i1_4_lut.LUT_INIT = 16'h9669;
    SB_DFFE data_in_frame_0___i44 (.Q(\data_in_frame[5] [3]), .C(clk16MHz), 
            .E(VCC_net), .D(n29890));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_adj_1060 (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(GND_net), .I3(GND_net), .O(n40660));
    defparam i1_2_lut_adj_1060.LUT_INIT = 16'hbbbb;
    SB_LUT4 i1_4_lut_adj_1061 (.I0(\data_out_frame[25] [3]), .I1(n25), .I2(n30), 
            .I3(n26), .O(n53491));
    defparam i1_4_lut_adj_1061.LUT_INIT = 16'h9669;
    SB_LUT4 i4_4_lut_adj_1062 (.I0(n59448), .I1(n53491), .I2(n59197), 
            .I3(n59484), .O(n10_adj_4742));
    defparam i4_4_lut_adj_1062.LUT_INIT = 16'h9669;
    SB_LUT4 select_775_Select_217_i3_4_lut (.I0(n59382), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(n10_adj_4742), .I3(n54456), .O(n3_adj_4743));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_217_i3_4_lut.LUT_INIT = 16'h8448;
    SB_LUT4 i3_4_lut (.I0(\data_out_frame[24] [6]), .I1(\data_out_frame[25] [0]), 
            .I2(\data_out_frame[25] [1]), .I3(n61721), .O(n59052));
    defparam i3_4_lut.LUT_INIT = 16'h9669;
    SB_LUT4 i2_2_lut (.I0(n59448), .I1(n59052), .I2(GND_net), .I3(GND_net), 
            .O(n6_adj_4744));
    defparam i2_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 select_775_Select_216_i3_4_lut (.I0(\data_out_frame[25] [2]), 
            .I1(\FRAME_MATCHER.state[3] ), .I2(n6_adj_4744), .I3(n59356), 
            .O(n3_adj_4745));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_216_i3_4_lut.LUT_INIT = 16'h8448;
    SB_LUT4 i12_2_lut (.I0(\data_out_frame[23] [1]), .I1(\data_out_frame[23] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n26168));   // verilog/coms.v(100[12:26])
    defparam i12_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i5_4_lut_adj_1063 (.I0(n58953), .I1(n59424), .I2(n53546), 
            .I3(\data_out_frame[19] [0]), .O(n12_adj_4746));
    defparam i5_4_lut_adj_1063.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1064 (.I0(\data_out_frame[23] [3]), .I1(\data_out_frame[21] [1]), 
            .I2(n12_adj_4746), .I3(n8_adj_4747), .O(n59197));
    defparam i1_4_lut_adj_1064.LUT_INIT = 16'h9669;
    SB_LUT4 select_775_Select_144_i2_4_lut (.I0(\data_out_frame[18] [0]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[16]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4748));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_144_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i28805_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n37), .I2(\data_in_frame[5] [3]), 
            .I3(\Ki[3] ), .O(n29692));   // verilog/coms.v(148[4] 304[11])
    defparam i28805_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i15687_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n37), .I2(\data_in_frame[5] [2]), 
            .I3(\Ki[2] ), .O(n29693));   // verilog/coms.v(148[4] 304[11])
    defparam i15687_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i10_4_lut (.I0(n26168), .I1(n59400), .I2(n26327), .I3(\data_out_frame[20] [1]), 
            .O(n28_c));
    defparam i10_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 select_775_Select_143_i2_4_lut (.I0(\data_out_frame[17] [7]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[7]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4749));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_143_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i14_3_lut (.I0(\data_out_frame[24] [7]), .I1(n28_c), .I2(\data_out_frame[24] [6]), 
            .I3(GND_net), .O(n32));
    defparam i14_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i12_4_lut (.I0(\data_out_frame[23] [4]), .I1(n59241), .I2(n59406), 
            .I3(n59162), .O(n30_adj_4750));
    defparam i12_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 select_775_Select_142_i2_4_lut (.I0(\data_out_frame[17] [6]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[6]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4751));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_142_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i13_4_lut (.I0(n59030), .I1(n54525), .I2(n58978), .I3(\data_out_frame[23] [7]), 
            .O(n31_c));
    defparam i13_4_lut.LUT_INIT = 16'h9669;
    SB_LUT4 select_775_Select_141_i2_4_lut (.I0(\data_out_frame[17] [5]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[5]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4752));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_141_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFFE data_in_frame_0___i43 (.Q(\data_in_frame[5] [2]), .C(clk16MHz), 
            .E(VCC_net), .D(n29885));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i11_4_lut (.I0(n53928), .I1(n58987), .I2(n59197), .I3(n53717), 
            .O(n29_c));
    defparam i11_4_lut.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0___i177 (.Q(\data_in_frame[22] [0]), .C(clk16MHz), 
           .D(n29586));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_775_Select_140_i2_4_lut (.I0(\data_out_frame[17] [4]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[4]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4753));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_140_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFFE data_in_frame_0___i42 (.Q(\data_in_frame[5] [1]), .C(clk16MHz), 
            .E(VCC_net), .D(n29881));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i41 (.Q(\data_in_frame[5] [0]), .C(clk16MHz), 
            .E(VCC_net), .D(n29878));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i17_4_lut (.I0(n29_c), .I1(n31_c), .I2(n30_adj_4750), .I3(n32), 
            .O(n60591));
    defparam i17_4_lut.LUT_INIT = 16'h6996;
    SB_DFFE data_in_frame_0___i40 (.Q(\data_in_frame[4] [7]), .C(clk16MHz), 
            .E(VCC_net), .D(n29877));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i3_4_lut_adj_1065 (.I0(n60591), .I1(\data_out_frame[25] [6]), 
            .I2(\data_out_frame[25] [4]), .I3(\data_out_frame[25] [5]), 
            .O(n59484));
    defparam i3_4_lut_adj_1065.LUT_INIT = 16'h9669;
    SB_DFF data_in_frame_0___i178 (.Q(\data_in_frame[22] [1]), .C(clk16MHz), 
           .D(n29589));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_adj_1066 (.I0(\data_out_frame[25] [3]), .I1(n59484), 
            .I2(GND_net), .I3(GND_net), .O(n59356));
    defparam i1_2_lut_adj_1066.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1067 (.I0(\data_out_frame[25] [2]), .I1(\data_out_frame[25] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n59149));
    defparam i1_2_lut_adj_1067.LUT_INIT = 16'h6666;
    SB_DFFE data_in_frame_0___i39 (.Q(\data_in_frame[4] [6]), .C(clk16MHz), 
            .E(VCC_net), .D(n57914));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i38 (.Q(\data_in_frame[4] [5]), .C(clk16MHz), 
            .E(VCC_net), .D(n57916));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_775_Select_139_i2_4_lut (.I0(\data_out_frame[17] [3]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[3]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4754));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_139_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFFE data_in_frame_0___i37 (.Q(\data_in_frame[4] [4]), .C(clk16MHz), 
            .E(VCC_net), .D(n57918));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_775_Select_215_i3_4_lut (.I0(\data_out_frame[25] [0]), 
            .I1(\FRAME_MATCHER.state[3] ), .I2(n8_adj_4755), .I3(n59149), 
            .O(n3_adj_4756));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_215_i3_4_lut.LUT_INIT = 16'h8448;
    SB_LUT4 i1_2_lut_adj_1068 (.I0(\data_out_frame[24] [5]), .I1(\data_out_frame[24] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n59030));
    defparam i1_2_lut_adj_1068.LUT_INIT = 16'h6666;
    SB_LUT4 select_775_Select_138_i2_4_lut (.I0(\data_out_frame[17] [2]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[2]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4757));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_138_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFF data_in_frame_0___i179 (.Q(\data_in_frame[22] [2]), .C(clk16MHz), 
           .D(n29592));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i15688_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n37), .I2(\data_in_frame[5] [1]), 
            .I3(\Ki[1] ), .O(n29694));   // verilog/coms.v(148[4] 304[11])
    defparam i15688_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFFE data_in_frame_0___i36 (.Q(\data_in_frame[4] [3]), .C(clk16MHz), 
            .E(VCC_net), .D(n29861));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i35 (.Q(\data_in_frame[4] [2]), .C(clk16MHz), 
            .E(VCC_net), .D(n29858));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_775_Select_214_i3_4_lut (.I0(n54570), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(n59030), .I3(n61136), .O(n3_adj_4758));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_214_i3_4_lut.LUT_INIT = 16'h4884;
    SB_DFFE data_in_frame_0___i34 (.Q(\data_in_frame[4] [1]), .C(clk16MHz), 
            .E(VCC_net), .D(n29855));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i15689_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n37), .I2(\data_in_frame[2] [7]), 
            .I3(\Kp[15] ), .O(n29695));   // verilog/coms.v(148[4] 304[11])
    defparam i15689_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i15690_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n37), .I2(\data_in_frame[2] [6]), 
            .I3(\Kp[14] ), .O(n29696));   // verilog/coms.v(148[4] 304[11])
    defparam i15690_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 select_775_Select_137_i2_4_lut (.I0(\data_out_frame[17] [1]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[1]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4759));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_137_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_775_Select_213_i3_4_lut (.I0(\data_out_frame[24] [4]), 
            .I1(\FRAME_MATCHER.state[3] ), .I2(n6_adj_4760), .I3(\data_out_frame[24] [3]), 
            .O(n3_adj_4761));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_213_i3_4_lut.LUT_INIT = 16'h4884;
    SB_DFF data_in_frame_0___i180 (.Q(\data_in_frame[22] [3]), .C(clk16MHz), 
           .D(n29596));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i33 (.Q(\data_in_frame[4] [0]), .C(clk16MHz), 
            .E(VCC_net), .D(n29851));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i32 (.Q(\data_in_frame[3] [7]), .C(clk16MHz), 
            .E(VCC_net), .D(n58126));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i31 (.Q(\data_in_frame[3][6] ), .C(clk16MHz), 
            .E(VCC_net), .D(n29845));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i181 (.Q(\data_in_frame[22] [4]), .C(clk16MHz), 
           .D(n29599));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i30 (.Q(\data_in_frame[3][5] ), .C(clk16MHz), 
            .E(VCC_net), .D(n29841));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i29 (.Q(\data_in_frame[3] [4]), .C(clk16MHz), 
            .E(VCC_net), .D(n29838));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_775_Select_211_i3_4_lut (.I0(\data_out_frame[24] [1]), 
            .I1(\FRAME_MATCHER.state[3] ), .I2(n6_adj_4762), .I3(n25142), 
            .O(n3_adj_4763));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_211_i3_4_lut.LUT_INIT = 16'h4884;
    SB_LUT4 i2_3_lut (.I0(n54397), .I1(n58990), .I2(\data_out_frame[24] [1]), 
            .I3(GND_net), .O(n59400));
    defparam i2_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i3_3_lut (.I0(\data_out_frame[24] [0]), .I1(\data_out_frame[23] [6]), 
            .I2(n59400), .I3(GND_net), .O(n8_adj_4764));
    defparam i3_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 select_775_Select_210_i3_4_lut (.I0(n53626), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(n8_adj_4764), .I3(n59218), .O(n3_adj_4765));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_210_i3_4_lut.LUT_INIT = 16'h8448;
    SB_LUT4 i2_3_lut_adj_1069 (.I0(n53644), .I1(n54397), .I2(n60897), 
            .I3(GND_net), .O(n53717));
    defparam i2_3_lut_adj_1069.LUT_INIT = 16'h6969;
    SB_LUT4 i2_3_lut_adj_1070 (.I0(\data_out_frame[21] [7]), .I1(n59403), 
            .I2(n53717), .I3(GND_net), .O(n59218));
    defparam i2_3_lut_adj_1070.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1071 (.I0(n58893), .I1(\data_out_frame[22] [4]), 
            .I2(n54566), .I3(GND_net), .O(n61721));
    defparam i2_3_lut_adj_1071.LUT_INIT = 16'h6969;
    SB_LUT4 i2_3_lut_adj_1072 (.I0(n53735), .I1(n59218), .I2(\data_out_frame[23] [7]), 
            .I3(GND_net), .O(n54568));
    defparam i2_3_lut_adj_1072.LUT_INIT = 16'h9696;
    SB_LUT4 i5_4_lut_adj_1073 (.I0(\data_out_frame[21] [7]), .I1(n58893), 
            .I2(n59344), .I3(n59040), .O(n12_adj_4766));
    defparam i5_4_lut_adj_1073.LUT_INIT = 16'h9669;
    SB_LUT4 i6_4_lut_adj_1074 (.I0(n26180), .I1(n12_adj_4766), .I2(n59332), 
            .I3(n54552), .O(n58987));
    defparam i6_4_lut_adj_1074.LUT_INIT = 16'h9669;
    SB_LUT4 i2_3_lut_adj_1075 (.I0(\data_out_frame[22] [4]), .I1(\data_out_frame[22] [3]), 
            .I2(n53897), .I3(GND_net), .O(n54525));
    defparam i2_3_lut_adj_1075.LUT_INIT = 16'h9696;
    SB_LUT4 i15691_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n37), .I2(\data_in_frame[2] [5]), 
            .I3(\Kp[13] ), .O(n29697));   // verilog/coms.v(148[4] 304[11])
    defparam i15691_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i15692_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n37), .I2(\data_in_frame[2] [4]), 
            .I3(\Kp[12] ), .O(n29698));   // verilog/coms.v(148[4] 304[11])
    defparam i15692_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_2_lut_adj_1076 (.I0(\data_out_frame[22] [5]), .I1(n53928), 
            .I2(GND_net), .I3(GND_net), .O(n54566));
    defparam i1_2_lut_adj_1076.LUT_INIT = 16'h6666;
    SB_LUT4 i15693_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n37), .I2(\data_in_frame[2] [3]), 
            .I3(\Kp[11] ), .O(n29699));   // verilog/coms.v(148[4] 304[11])
    defparam i15693_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4_4_lut_adj_1077 (.I0(\data_out_frame[20] [0]), .I1(\data_out_frame[22] [2]), 
            .I2(\data_out_frame[17] [6]), .I3(n6_adj_4767), .O(n59040));
    defparam i4_4_lut_adj_1077.LUT_INIT = 16'h6996;
    SB_LUT4 i15694_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n37), .I2(\data_in_frame[2] [2]), 
            .I3(\Kp[10] ), .O(n29700));   // verilog/coms.v(148[4] 304[11])
    defparam i15694_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_4_lut_adj_1078 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[8] [6]), 
            .I2(encoder0_position_scaled[6]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4768));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1078.LUT_INIT = 16'ha088;
    SB_LUT4 i15695_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n37), .I2(\data_in_frame[2] [1]), 
            .I3(\Kp[9] ), .O(n29701));   // verilog/coms.v(148[4] 304[11])
    defparam i15695_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_2_lut_adj_1079 (.I0(\data_out_frame[20] [2]), .I1(n54415), 
            .I2(GND_net), .I3(GND_net), .O(n54529));
    defparam i1_2_lut_adj_1079.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1080 (.I0(n26739), .I1(n54220), .I2(\data_out_frame[15] [6]), 
            .I3(GND_net), .O(n60541));
    defparam i2_3_lut_adj_1080.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_1081 (.I0(\data_out_frame[17] [7]), .I1(n58809), 
            .I2(\data_out_frame[19] [7]), .I3(n60541), .O(n53897));
    defparam i3_4_lut_adj_1081.LUT_INIT = 16'h9669;
    SB_LUT4 select_775_Select_136_i2_4_lut (.I0(\data_out_frame[17] [0]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[0]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4769));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_136_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i2_3_lut_adj_1082 (.I0(\data_out_frame[21] [6]), .I1(n60897), 
            .I2(n53735), .I3(GND_net), .O(n58990));
    defparam i2_3_lut_adj_1082.LUT_INIT = 16'h6969;
    SB_LUT4 select_775_Select_135_i2_4_lut (.I0(\data_out_frame[16] [7]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[15]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4770));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_135_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i4_4_lut_adj_1083 (.I0(\data_out_frame[18] [0]), .I1(n60541), 
            .I2(n26585), .I3(n6_adj_4771), .O(n54415));
    defparam i4_4_lut_adj_1083.LUT_INIT = 16'h9669;
    SB_LUT4 select_775_Select_134_i2_4_lut (.I0(\data_out_frame[16] [6]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[14]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4772));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_134_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i2_3_lut_adj_1084 (.I0(\data_out_frame[22] [0]), .I1(\data_out_frame[19] [6]), 
            .I2(n53610), .I3(GND_net), .O(n53644));
    defparam i2_3_lut_adj_1084.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_1085 (.I0(\data_out_frame[16] [3]), .I1(n59186), 
            .I2(n59124), .I3(\data_out_frame[16] [2]), .O(n53707));   // verilog/coms.v(88[17:70])
    defparam i3_4_lut_adj_1085.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1086 (.I0(n25650), .I1(n58944), .I2(\data_out_frame[17] [4]), 
            .I3(GND_net), .O(n53610));
    defparam i2_3_lut_adj_1086.LUT_INIT = 16'h9696;
    SB_LUT4 select_775_Select_133_i2_4_lut (.I0(\data_out_frame[16] [5]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[13]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4773));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_133_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_4_lut_adj_1087 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[16] [4]), 
            .I2(pwm_setpoint[12]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4774));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1087.LUT_INIT = 16'ha088;
    SB_LUT4 i15696_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n37), .I2(\data_in_frame[2] [0]), 
            .I3(\Kp[8] ), .O(n29702));   // verilog/coms.v(148[4] 304[11])
    defparam i15696_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 select_775_Select_131_i2_4_lut (.I0(\data_out_frame[16] [3]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[11]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4775));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_131_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_adj_1088 (.I0(\data_out_frame[20] [6]), .I1(\data_out_frame[20] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n26180));
    defparam i1_2_lut_adj_1088.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1089 (.I0(\data_out_frame[15] [1]), .I1(\data_out_frame[19] [5]), 
            .I2(n58975), .I3(n53610), .O(n54397));
    defparam i1_4_lut_adj_1089.LUT_INIT = 16'h9669;
    SB_DFFESS data_out_frame_0___i69 (.Q(\data_out_frame[8] [4]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4776), .S(n58621));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_adj_1090 (.I0(\data_out_frame[19] [0]), .I1(\data_out_frame[19] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n59421));
    defparam i1_2_lut_adj_1090.LUT_INIT = 16'h6666;
    SB_LUT4 i13_2_lut (.I0(\data_out_frame[19] [7]), .I1(\data_out_frame[19] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n2107));   // verilog/coms.v(100[12:26])
    defparam i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1091 (.I0(\data_out_frame[12] [4]), .I1(\data_out_frame[12] [7]), 
            .I2(\data_out_frame[12] [2]), .I3(n59021), .O(n10_adj_4777));   // verilog/coms.v(88[17:28])
    defparam i4_4_lut_adj_1091.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_1092 (.I0(\data_out_frame[12] [1]), .I1(n10_adj_4777), 
            .I2(\data_out_frame[12] [3]), .I3(GND_net), .O(n1673));   // verilog/coms.v(88[17:28])
    defparam i5_3_lut_adj_1092.LUT_INIT = 16'h9696;
    SB_LUT4 i7_4_lut_adj_1093 (.I0(\data_out_frame[8] [2]), .I1(n58782), 
            .I2(n59287), .I3(n1673), .O(n18_c));
    defparam i7_4_lut_adj_1093.LUT_INIT = 16'h6996;
    SB_LUT4 i6_3_lut (.I0(\data_out_frame[12] [0]), .I1(n59112), .I2(n59442), 
            .I3(GND_net), .O(n17));
    defparam i6_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i21810_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n37), .I2(\data_in_frame[3] [7]), 
            .I3(\Kp[7] ), .O(n29703));   // verilog/coms.v(148[4] 304[11])
    defparam i21810_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i8_4_lut (.I0(n59335), .I1(n59012), .I2(n59281), .I3(\data_out_frame[6] [1]), 
            .O(n19_c));
    defparam i8_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i2_4_lut (.I0(n19_c), .I1(n25052), .I2(n17), .I3(n18_c), 
            .O(n10_adj_4778));
    defparam i2_4_lut.LUT_INIT = 16'h9669;
    SB_LUT4 i6_4_lut_adj_1094 (.I0(n59171), .I1(n1510), .I2(n26049), .I3(\data_out_frame[13] [7]), 
            .O(n14_adj_4779));
    defparam i6_4_lut_adj_1094.LUT_INIT = 16'h6996;
    SB_LUT4 select_775_Select_130_i2_4_lut (.I0(\data_out_frame[16] [2]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[10]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4780));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_130_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i7_4_lut_adj_1095 (.I0(n1513), .I1(n14_adj_4779), .I2(n10_adj_4778), 
            .I3(n1673), .O(n60980));
    defparam i7_4_lut_adj_1095.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1096 (.I0(\data_out_frame[18] [6]), .I1(n60980), 
            .I2(GND_net), .I3(GND_net), .O(n59274));
    defparam i1_2_lut_adj_1096.LUT_INIT = 16'h9999;
    SB_DFFESS data_out_frame_0___i70 (.Q(\data_out_frame[8] [5]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4781), .S(n58620));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i3_4_lut_adj_1097 (.I0(\data_out_frame[18] [5]), .I1(n59274), 
            .I2(n70022), .I3(n54413), .O(n59424));
    defparam i3_4_lut_adj_1097.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1098 (.I0(\data_out_frame[17] [7]), .I1(\data_out_frame[17] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n26585));
    defparam i1_2_lut_adj_1098.LUT_INIT = 16'h6666;
    SB_LUT4 select_775_Select_129_i2_4_lut (.I0(\data_out_frame[16] [1]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[9]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4782));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_129_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i3_4_lut_adj_1099 (.I0(n25650), .I1(n26206), .I2(\data_out_frame[15] [3]), 
            .I3(\data_out_frame[17] [5]), .O(n59089));
    defparam i3_4_lut_adj_1099.LUT_INIT = 16'h6996;
    SB_LUT4 select_775_Select_128_i2_4_lut (.I0(\data_out_frame[16] [0]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[8]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4783));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_128_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i15698_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n37), .I2(\data_in_frame[3][6] ), 
            .I3(\Kp[6] ), .O(n29704));   // verilog/coms.v(148[4] 304[11])
    defparam i15698_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_2_lut_adj_1100 (.I0(\data_out_frame[16] [3]), .I1(\data_out_frame[14] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n26350));
    defparam i1_2_lut_adj_1100.LUT_INIT = 16'h6666;
    SB_LUT4 add_1097_8_lut (.I0(n58672), .I1(byte_transmit_counter[6]), 
            .I2(GND_net), .I3(n51014), .O(n58680)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1097_8_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i15699_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n37), .I2(\data_in_frame[3][5] ), 
            .I3(\Kp[5] ), .O(n29705));   // verilog/coms.v(148[4] 304[11])
    defparam i15699_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i15700_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n37), .I2(\data_in_frame[3] [4]), 
            .I3(\Kp[4] ), .O(n29706));   // verilog/coms.v(148[4] 304[11])
    defparam i15700_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2_3_lut_adj_1101 (.I0(n54552), .I1(n59089), .I2(\data_out_frame[18] [0]), 
            .I3(GND_net), .O(n58809));
    defparam i2_3_lut_adj_1101.LUT_INIT = 16'h6969;
    SB_DFFE data_in_frame_0___i28 (.Q(\data_in_frame[3] [3]), .C(clk16MHz), 
            .E(VCC_net), .D(n29835));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i71 (.Q(\data_out_frame[8] [6]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4768), .S(n58671));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_775_Select_127_i2_4_lut (.I0(\data_out_frame[15] [7]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[23]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4784));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_127_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i15701_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n37), .I2(\data_in_frame[3] [3]), 
            .I3(\Kp[3] ), .O(n29707));   // verilog/coms.v(148[4] 304[11])
    defparam i15701_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i10_4_lut_adj_1102 (.I0(n58953), .I1(n53735), .I2(n58809), 
            .I3(n26350), .O(n24));
    defparam i10_4_lut_adj_1102.LUT_INIT = 16'h6996;
    SB_LUT4 i15702_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n37), .I2(\data_in_frame[3] [2]), 
            .I3(\Kp[2] ), .O(n29708));   // verilog/coms.v(148[4] 304[11])
    defparam i15702_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5_3_lut_adj_1103 (.I0(n70020), .I1(\data_out_frame[17] [5]), 
            .I2(n26817), .I3(GND_net), .O(n14_adj_4785));
    defparam i5_3_lut_adj_1103.LUT_INIT = 16'h6969;
    SB_LUT4 i6_4_lut_adj_1104 (.I0(n59308), .I1(\data_out_frame[17] [3]), 
            .I2(n26585), .I3(n59024), .O(n15_c));
    defparam i6_4_lut_adj_1104.LUT_INIT = 16'h6996;
    SB_LUT4 select_775_Select_126_i2_4_lut (.I0(\data_out_frame[15] [6]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[22]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4786));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_126_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFFR \FRAME_MATCHER.state_FSM_i1  (.Q(Kp_23__N_1748), .C(clk16MHz), 
            .D(n2068), .R(reset));   // verilog/coms.v(148[4] 304[11])
    SB_CARRY add_1097_8 (.CI(n51014), .I0(byte_transmit_counter[6]), .I1(GND_net), 
            .CO(n51015));
    SB_DFFER setpoint_i0_i0 (.Q(setpoint[0]), .C(clk16MHz), .E(n27674), 
            .D(n4760[0]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i27 (.Q(\data_in_frame[3] [2]), .C(clk16MHz), 
            .E(VCC_net), .D(n29832));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i15703_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n37), .I2(\data_in_frame[3] [1]), 
            .I3(\Kp[1] ), .O(n29709));   // verilog/coms.v(148[4] 304[11])
    defparam i15703_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 select_775_Select_69_i2_4_lut (.I0(\data_out_frame[8] [5]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder0_position_scaled[5]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4781));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_69_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i8_4_lut_adj_1105 (.I0(n15_c), .I1(\data_out_frame[16] [5]), 
            .I2(n14_adj_4785), .I3(\data_out_frame[17] [4]), .O(n61441));
    defparam i8_4_lut_adj_1105.LUT_INIT = 16'h6996;
    SB_LUT4 add_1097_7_lut (.I0(n58672), .I1(byte_transmit_counter[5]), 
            .I2(GND_net), .I3(n51013), .O(n58679)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1097_7_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i8_4_lut_adj_1106 (.I0(n59329), .I1(\data_out_frame[18] [1]), 
            .I2(\data_out_frame[19] [3]), .I3(n2076), .O(n22_c));
    defparam i8_4_lut_adj_1106.LUT_INIT = 16'h6996;
    SB_LUT4 i12_4_lut_adj_1107 (.I0(n58935), .I1(n24), .I2(n18_adj_4787), 
            .I3(n25764), .O(n26_adj_4788));
    defparam i12_4_lut_adj_1107.LUT_INIT = 16'h6996;
    SB_LUT4 i54330_4_lut (.I0(n61441), .I1(\data_out_frame[14] [4]), .I2(n59168), 
            .I3(\data_out_frame[18] [5]), .O(n70024));
    defparam i54330_4_lut.LUT_INIT = 16'h9669;
    SB_LUT4 select_775_Select_125_i2_4_lut (.I0(\data_out_frame[15] [5]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[21]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4789));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_125_i2_4_lut.LUT_INIT = 16'hc088;
    SB_CARRY add_1097_7 (.CI(n51013), .I0(byte_transmit_counter[5]), .I1(GND_net), 
            .CO(n51014));
    SB_LUT4 i15704_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n37), .I2(\data_in_frame[11] [7]), 
            .I3(IntegralLimit[23]), .O(n29710));   // verilog/coms.v(148[4] 304[11])
    defparam i15704_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i15705_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n37), .I2(\data_in_frame[11] [6]), 
            .I3(IntegralLimit[22]), .O(n29711));   // verilog/coms.v(148[4] 304[11])
    defparam i15705_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 add_1097_6_lut (.I0(n58672), .I1(byte_transmit_counter[4]), 
            .I2(GND_net), .I3(n51012), .O(n58678)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1097_6_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i15706_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n37), .I2(\data_in_frame[11] [5]), 
            .I3(IntegralLimit[21]), .O(n29712));   // verilog/coms.v(148[4] 304[11])
    defparam i15706_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i13_4_lut_adj_1108 (.I0(n70024), .I1(n26_adj_4788), .I2(n22_c), 
            .I3(n2107), .O(n60743));
    defparam i13_4_lut_adj_1108.LUT_INIT = 16'h9669;
    SB_LUT4 select_775_Select_124_i2_4_lut (.I0(\data_out_frame[15] [4]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[20]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4790));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_124_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i15707_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n37), .I2(\data_in_frame[11] [4]), 
            .I3(IntegralLimit[20]), .O(n29713));   // verilog/coms.v(148[4] 304[11])
    defparam i15707_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4_4_lut_adj_1109 (.I0(\data_out_frame[19] [5]), .I1(n60743), 
            .I2(n59421), .I3(n6_adj_4791), .O(n23650));
    defparam i4_4_lut_adj_1109.LUT_INIT = 16'h6996;
    SB_LUT4 select_775_Select_123_i2_4_lut (.I0(\data_out_frame[15] [3]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[19]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4792));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_123_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_adj_1110 (.I0(\data_out_frame[16] [0]), .I1(\data_out_frame[18] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n59168));
    defparam i1_2_lut_adj_1110.LUT_INIT = 16'h6666;
    SB_LUT4 select_775_Select_122_i2_4_lut (.I0(\data_out_frame[15] [2]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[18]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4793));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_122_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_775_Select_121_i2_4_lut (.I0(\data_out_frame[15] [1]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[17]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4794));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_121_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFFESS data_out_frame_0___i72 (.Q(\data_out_frame[8] [7]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4795), .S(n58619));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i26 (.Q(\data_in_frame[3] [1]), .C(clk16MHz), 
            .E(VCC_net), .D(n29829));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i22866_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n37), .I2(\data_in_frame[11] [3]), 
            .I3(IntegralLimit[19]), .O(n29714));   // verilog/coms.v(148[4] 304[11])
    defparam i22866_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5_4_lut_adj_1111 (.I0(n26849), .I1(n26739), .I2(\data_out_frame[17] [7]), 
            .I3(n25872), .O(n12_adj_4796));
    defparam i5_4_lut_adj_1111.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1112 (.I0(\data_out_frame[18] [1]), .I1(n54432), 
            .I2(n12_adj_4796), .I3(n8_adj_4797), .O(n59189));
    defparam i1_4_lut_adj_1112.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_55442 (.I0(byte_transmit_counter[3]), 
            .I1(n71081), .I2(n66954), .I3(byte_transmit_counter[4]), .O(n71150));
    defparam byte_transmit_counter_3__bdd_4_lut_55442.LUT_INIT = 16'he4aa;
    SB_DFFE data_in_frame_0___i25 (.Q(\data_in_frame[3] [0]), .C(clk16MHz), 
            .E(VCC_net), .D(n29826));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i2_3_lut_adj_1113 (.I0(\data_out_frame[15] [7]), .I1(\data_out_frame[13] [7]), 
            .I2(n53640), .I3(GND_net), .O(n54490));
    defparam i2_3_lut_adj_1113.LUT_INIT = 16'h9696;
    SB_LUT4 i4_4_lut_adj_1114 (.I0(n7_c), .I1(n54432), .I2(n54490), .I3(n59189), 
            .O(n23652));
    defparam i4_4_lut_adj_1114.LUT_INIT = 16'h6996;
    SB_LUT4 n71150_bdd_4_lut (.I0(n71150), .I1(n14_adj_4798), .I2(n7_adj_4799), 
            .I3(byte_transmit_counter[4]), .O(tx_data[5]));
    defparam n71150_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFFESS data_out_frame_0___i73 (.Q(\data_out_frame[9] [0]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4800), .S(n58495));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_adj_1115 (.I0(\data_out_frame[22] [1]), .I1(n23650), 
            .I2(GND_net), .I3(GND_net), .O(n59344));
    defparam i1_2_lut_adj_1115.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1116 (.I0(n2217), .I1(n54397), .I2(n23650), .I3(n6_adj_4801), 
            .O(n53933));
    defparam i4_4_lut_adj_1116.LUT_INIT = 16'h6996;
    SB_LUT4 select_775_Select_68_i2_4_lut (.I0(\data_out_frame[8] [4]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder0_position_scaled[4]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4776));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_68_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i4_4_lut_adj_1117 (.I0(\data_out_frame[16] [2]), .I1(n54432), 
            .I2(n54434), .I3(n6_adj_4802), .O(n60844));
    defparam i4_4_lut_adj_1117.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1118 (.I0(n54415), .I1(n2217), .I2(n58990), .I3(n53897), 
            .O(n16));
    defparam i6_4_lut_adj_1118.LUT_INIT = 16'h9669;
    SB_LUT4 i7_4_lut_adj_1119 (.I0(n60844), .I1(n53933), .I2(n59344), 
            .I3(n23652), .O(n17_adj_4803));
    defparam i7_4_lut_adj_1119.LUT_INIT = 16'h9669;
    SB_LUT4 i9_4_lut (.I0(n17_adj_4803), .I1(n53644), .I2(n16), .I3(n61261), 
            .O(n25142));
    defparam i9_4_lut.LUT_INIT = 16'h9669;
    SB_LUT4 i22897_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n37), .I2(\data_in_frame[11] [2]), 
            .I3(IntegralLimit[18]), .O(n29715));   // verilog/coms.v(148[4] 304[11])
    defparam i22897_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i3_4_lut_adj_1120 (.I0(n54529), .I1(n59040), .I2(n54552), 
            .I3(\data_out_frame[22] [3]), .O(n54570));
    defparam i3_4_lut_adj_1120.LUT_INIT = 16'h9669;
    SB_LUT4 i2_3_lut_adj_1121 (.I0(n53626), .I1(n53583), .I2(\data_out_frame[23] [5]), 
            .I3(GND_net), .O(n26327));
    defparam i2_3_lut_adj_1121.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1122 (.I0(n61136), .I1(n59448), .I2(GND_net), 
            .I3(GND_net), .O(n58984));
    defparam i1_2_lut_adj_1122.LUT_INIT = 16'h9999;
    SB_DFFESS data_out_frame_0___i74 (.Q(\data_out_frame[9] [1]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4804), .S(n58618));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i75 (.Q(\data_out_frame[9] [2]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4805), .S(n58617));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i76 (.Q(\data_out_frame[9] [3]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4806), .S(n58616));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i77 (.Q(\data_out_frame[9] [4]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4807), .S(n58615));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i78 (.Q(\data_out_frame[9] [5]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4808), .S(n58614));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i79 (.Q(\data_out_frame[9] [6]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4809), .S(n58613));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i80 (.Q(\data_out_frame[9] [7]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4810), .S(n58612));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i81 (.Q(\data_out_frame[10] [0]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4811), .S(n58611));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i82 (.Q(\data_out_frame[10] [1]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4812), .S(n58610));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i83 (.Q(\data_out_frame[10] [2]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4813), .S(n58609));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i84 (.Q(\data_out_frame[10] [3]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4814), .S(n58608));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i85 (.Q(\data_out_frame[10] [4]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4815), .S(n58607));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i86 (.Q(\data_out_frame[10] [5]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4816), .S(n58606));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i87 (.Q(\data_out_frame[10] [6]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4817), .S(n58605));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i88 (.Q(\data_out_frame[10] [7]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4818), .S(n58604));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i89 (.Q(\data_out_frame[11] [0]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4819), .S(n58603));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i4_4_lut_adj_1123 (.I0(n58984), .I1(n26327), .I2(n54570), 
            .I3(n59338), .O(n10_adj_4820));
    defparam i4_4_lut_adj_1123.LUT_INIT = 16'h9669;
    SB_LUT4 select_775_Select_209_i3_4_lut (.I0(n54568), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(n10_adj_4820), .I3(n61721), .O(n3_adj_4821));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_209_i3_4_lut.LUT_INIT = 16'h8448;
    SB_LUT4 i22935_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n37), .I2(\data_in_frame[11] [1]), 
            .I3(IntegralLimit[17]), .O(n29716));   // verilog/coms.v(148[4] 304[11])
    defparam i22935_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4_4_lut_adj_1124 (.I0(\data_out_frame[12] [7]), .I1(\data_out_frame[10] [5]), 
            .I2(n59384), .I3(n6_adj_4822), .O(n26206));   // verilog/coms.v(77[16:27])
    defparam i4_4_lut_adj_1124.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1125 (.I0(\data_out_frame[15] [2]), .I1(n26206), 
            .I2(n53449), .I3(\data_out_frame[17] [3]), .O(n58975));
    defparam i3_4_lut_adj_1125.LUT_INIT = 16'h6996;
    SB_CARRY add_1097_6 (.CI(n51012), .I0(byte_transmit_counter[4]), .I1(GND_net), 
            .CO(n51013));
    SB_LUT4 add_1097_5_lut (.I0(n58672), .I1(byte_transmit_counter[3]), 
            .I2(GND_net), .I3(n51011), .O(n58677)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1097_5_lut.LUT_INIT = 16'h8228;
    SB_DFFESS data_out_frame_0___i90 (.Q(\data_out_frame[11] [1]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4823), .S(n58602));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i91 (.Q(\data_out_frame[11] [2]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4824), .S(n58601));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i92 (.Q(\data_out_frame[11] [3]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4825), .S(n58600));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i93 (.Q(\data_out_frame[11] [4]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4826), .S(n58599));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i94 (.Q(\data_out_frame[11] [5]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4827), .S(n58598));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i95 (.Q(\data_out_frame[11] [6]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4828), .S(n58597));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i96 (.Q(\data_out_frame[11] [7]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4829), .S(n58596));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i97 (.Q(\data_out_frame[12] [0]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4830), .S(n58595));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i98 (.Q(\data_out_frame[12] [1]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4831), .S(n58594));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i99 (.Q(\data_out_frame[12] [2]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4832), .S(n58593));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i15711_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n37), .I2(\data_in_frame[11] [0]), 
            .I3(IntegralLimit[16]), .O(n29717));   // verilog/coms.v(148[4] 304[11])
    defparam i15711_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFFESS data_out_frame_0___i100 (.Q(\data_out_frame[12] [3]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4833), .S(n58592));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i101 (.Q(\data_out_frame[12] [4]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4834), .S(n58591));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i102 (.Q(\data_out_frame[12] [5]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4835), .S(n58590));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i103 (.Q(\data_out_frame[12] [6]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4836), .S(n58589));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i104 (.Q(\data_out_frame[12] [7]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4837), .S(n58588));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i15712_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n37), .I2(\data_in_frame[12] [7]), 
            .I3(IntegralLimit[15]), .O(n29718));   // verilog/coms.v(148[4] 304[11])
    defparam i15712_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i15713_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n37), .I2(\data_in_frame[12] [6]), 
            .I3(IntegralLimit[14]), .O(n29719));   // verilog/coms.v(148[4] 304[11])
    defparam i15713_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFFESS data_out_frame_0___i105 (.Q(\data_out_frame[13] [0]), .C(clk16MHz), 
            .E(n30494), .D(n2_adj_4838), .S(n28975));   // verilog/coms.v(130[12] 305[6])
    SB_CARRY add_1097_5 (.CI(n51011), .I0(byte_transmit_counter[3]), .I1(GND_net), 
            .CO(n51012));
    SB_LUT4 add_1097_4_lut (.I0(n58672), .I1(\byte_transmit_counter[2] ), 
            .I2(GND_net), .I3(n51010), .O(n58676)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1097_4_lut.LUT_INIT = 16'h8228;
    SB_DFFE data_in_frame_0___i24 (.Q(\data_in_frame[2] [7]), .C(clk16MHz), 
            .E(VCC_net), .D(n29823));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i106 (.Q(\data_out_frame[13] [1]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4839), .S(n58587));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_adj_1126 (.I0(\data_out_frame[12] [1]), .I1(n25052), 
            .I2(GND_net), .I3(GND_net), .O(n58935));
    defparam i1_2_lut_adj_1126.LUT_INIT = 16'h6666;
    SB_LUT4 i15714_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n37), .I2(\data_in_frame[12] [5]), 
            .I3(IntegralLimit[13]), .O(n29720));   // verilog/coms.v(148[4] 304[11])
    defparam i15714_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i15744_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n37), .I2(\data_in_frame[16] [6]), 
            .I3(deadband[6]), .O(n29750));   // verilog/coms.v(148[4] 304[11])
    defparam i15744_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_CARRY add_1097_4 (.CI(n51010), .I0(\byte_transmit_counter[2] ), .I1(GND_net), 
            .CO(n51011));
    SB_DFFESS data_out_frame_0___i107 (.Q(\data_out_frame[13] [2]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4840), .S(n58586));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 add_1097_3_lut (.I0(n58672), .I1(\byte_transmit_counter[1] ), 
            .I2(GND_net), .I3(n51009), .O(n58675)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1097_3_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_1097_3 (.CI(n51009), .I0(\byte_transmit_counter[1] ), .I1(GND_net), 
            .CO(n51010));
    SB_LUT4 i2_3_lut_adj_1127 (.I0(\data_out_frame[16] [5]), .I1(n58953), 
            .I2(\data_out_frame[16] [3]), .I3(GND_net), .O(n25872));   // verilog/coms.v(88[17:28])
    defparam i2_3_lut_adj_1127.LUT_INIT = 16'h9696;
    SB_LUT4 add_1097_2_lut (.I0(n58672), .I1(\byte_transmit_counter[0] ), 
            .I2(tx_transmit_N_3416), .I3(GND_net), .O(n58674)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1097_2_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i15747_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n37), .I2(\data_in_frame[16] [3]), 
            .I3(deadband[3]), .O(n29753));   // verilog/coms.v(148[4] 304[11])
    defparam i15747_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_2_lut_adj_1128 (.I0(\data_out_frame[14] [3]), .I1(n54114), 
            .I2(GND_net), .I3(GND_net), .O(n54413));
    defparam i1_2_lut_adj_1128.LUT_INIT = 16'h6666;
    SB_DFFESS data_out_frame_0___i108 (.Q(\data_out_frame[13] [3]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4841), .S(n58585));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i23 (.Q(\data_in_frame[2] [6]), .C(clk16MHz), 
            .E(VCC_net), .D(n29820));   // verilog/coms.v(130[12] 305[6])
    SB_CARRY add_1097_2 (.CI(GND_net), .I0(\byte_transmit_counter[0] ), 
            .I1(tx_transmit_N_3416), .CO(n51009));
    SB_LUT4 i15746_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n37), .I2(\data_in_frame[16] [4]), 
            .I3(deadband[4]), .O(n29752));   // verilog/coms.v(148[4] 304[11])
    defparam i15746_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_2_lut_adj_1129 (.I0(\data_out_frame[11] [3]), .I1(\data_out_frame[11] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n26618));   // verilog/coms.v(88[17:70])
    defparam i1_2_lut_adj_1129.LUT_INIT = 16'h6666;
    SB_LUT4 i5_4_lut_adj_1130 (.I0(n1169), .I1(n58887), .I2(\data_out_frame[13] [4]), 
            .I3(\data_out_frame[7] [1]), .O(n12_adj_4842));
    defparam i5_4_lut_adj_1130.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1131 (.I0(n26618), .I1(n12_adj_4842), .I2(n59296), 
            .I3(n36), .O(n54220));
    defparam i6_4_lut_adj_1131.LUT_INIT = 16'h6996;
    SB_LUT4 i15743_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n37), .I2(\data_in_frame[16] [7]), 
            .I3(deadband[7]), .O(n29749));   // verilog/coms.v(148[4] 304[11])
    defparam i15743_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_2_lut_adj_1132 (.I0(\data_out_frame[10] [6]), .I1(\data_out_frame[10] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_4843));   // verilog/coms.v(88[17:63])
    defparam i1_2_lut_adj_1132.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1133 (.I0(\data_out_frame[10] [3]), .I1(\data_out_frame[10] [7]), 
            .I2(\data_out_frame[10] [2]), .I3(n6_adj_4843), .O(n58782));   // verilog/coms.v(88[17:63])
    defparam i4_4_lut_adj_1133.LUT_INIT = 16'h6996;
    SB_LUT4 i15742_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n37), .I2(\data_in_frame[15] [0]), 
            .I3(deadband[8]), .O(n29748));   // verilog/coms.v(148[4] 304[11])
    defparam i15742_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_2_lut_adj_1134 (.I0(\data_out_frame[9] [0]), .I1(\data_out_frame[9] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n59296));
    defparam i1_2_lut_adj_1134.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1135 (.I0(\data_out_frame[9] [1]), .I1(\data_out_frame[6] [6]), 
            .I2(\data_out_frame[4] [4]), .I3(n26143), .O(n26_adj_4844));
    defparam i1_4_lut_adj_1135.LUT_INIT = 16'h6996;
    SB_DFFE data_in_frame_0___i22 (.Q(\data_in_frame[2] [5]), .C(clk16MHz), 
            .E(VCC_net), .D(n29817));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i23663_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n37), .I2(\data_in_frame[15] [1]), 
            .I3(deadband[9]), .O(n29747));   // verilog/coms.v(148[4] 304[11])
    defparam i23663_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i15740_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n37), .I2(\data_in_frame[15] [2]), 
            .I3(deadband[10]), .O(n29746));   // verilog/coms.v(148[4] 304[11])
    defparam i15740_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF data_in_frame_0___i182 (.Q(\data_in_frame[22] [5]), .C(clk16MHz), 
           .D(n29609));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i17_4_lut_adj_1136 (.I0(n25682), .I1(n25611), .I2(\data_out_frame[7] [2]), 
            .I3(n58867), .O(n42));
    defparam i17_4_lut_adj_1136.LUT_INIT = 16'h6996;
    SB_LUT4 i15_4_lut (.I0(\data_out_frame[9] [6]), .I1(n26046), .I2(n26376), 
            .I3(n58931), .O(n40));
    defparam i15_4_lut.LUT_INIT = 16'h6996;
    SB_DFFE data_in_frame_0___i21 (.Q(\data_in_frame[2] [4]), .C(clk16MHz), 
            .E(VCC_net), .D(n29813));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i20 (.Q(\data_in_frame[2] [3]), .C(clk16MHz), 
            .E(VCC_net), .D(n29810));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_55412 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[10] [1]), .I2(\data_out_frame[11] [1]), 
            .I3(\byte_transmit_counter[1] ), .O(n71138));
    defparam byte_transmit_counter_0__bdd_4_lut_55412.LUT_INIT = 16'he4aa;
    SB_DFFESS data_out_frame_0___i109 (.Q(\data_out_frame[13] [4]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4845), .S(n58584));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 n71138_bdd_4_lut (.I0(n71138), .I1(\data_out_frame[9] [1]), 
            .I2(\data_out_frame[8] [1]), .I3(\byte_transmit_counter[1] ), 
            .O(n71141));
    defparam n71138_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFFESS data_out_frame_0___i110 (.Q(\data_out_frame[13] [5]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4846), .S(n58583));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i111 (.Q(\data_out_frame[13] [6]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4847), .S(n58582));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i16_4_lut (.I0(\data_out_frame[6] [3]), .I1(n58864), .I2(\data_out_frame[7] [1]), 
            .I3(\data_out_frame[8] [7]), .O(n41));
    defparam i16_4_lut.LUT_INIT = 16'h6996;
    SB_DFFESS data_out_frame_0___i112 (.Q(\data_out_frame[13] [7]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4848), .S(n58581));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i14_4_lut (.I0(n59296), .I1(\data_out_frame[9] [5]), .I2(n58858), 
            .I3(n59229), .O(n39));
    defparam i14_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i15739_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n37), .I2(\data_in_frame[15] [3]), 
            .I3(deadband[11]), .O(n29745));   // verilog/coms.v(148[4] 304[11])
    defparam i15739_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i19_4_lut (.I0(\data_out_frame[4] [6]), .I1(n26563), .I2(n1130), 
            .I3(n26_adj_4844), .O(n44));
    defparam i19_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i23_4_lut (.I0(n39), .I1(n41), .I2(n40), .I3(n42), .O(n48));
    defparam i23_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i15738_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n37), .I2(\data_in_frame[15] [4]), 
            .I3(deadband[12]), .O(n29744));   // verilog/coms.v(148[4] 304[11])
    defparam i15738_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i15737_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n37), .I2(\data_in_frame[15] [5]), 
            .I3(deadband[13]), .O(n29743));   // verilog/coms.v(148[4] 304[11])
    defparam i15737_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i15736_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n37), .I2(\data_in_frame[15] [6]), 
            .I3(deadband[14]), .O(n29742));   // verilog/coms.v(148[4] 304[11])
    defparam i15736_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i18_4_lut (.I0(n58861), .I1(\data_out_frame[7] [0]), .I2(n58821), 
            .I3(\data_out_frame[4] [5]), .O(n43_c));
    defparam i18_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i2_2_lut_adj_1137 (.I0(\data_out_frame[10] [0]), .I1(\data_out_frame[11] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n8_adj_4849));
    defparam i2_2_lut_adj_1137.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1138 (.I0(\data_out_frame[11] [4]), .I1(n43_c), 
            .I2(n48), .I3(n44), .O(n7_adj_4850));
    defparam i1_4_lut_adj_1138.LUT_INIT = 16'h9669;
    SB_LUT4 i5_4_lut_adj_1139 (.I0(n26618), .I1(n7_adj_4850), .I2(n26376), 
            .I3(n8_adj_4849), .O(n59442));
    defparam i5_4_lut_adj_1139.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1140 (.I0(n4_c), .I1(\data_out_frame[15] [2]), 
            .I2(\data_out_frame[15] [3]), .I3(GND_net), .O(n58944));
    defparam i2_3_lut_adj_1140.LUT_INIT = 16'h9696;
    SB_DFFESS data_out_frame_0___i113 (.Q(\data_out_frame[14] [0]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4851), .S(n58580));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i114 (.Q(\data_out_frame[14] [1]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4852), .S(n58579));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i15735_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n37), .I2(\data_in_frame[15] [7]), 
            .I3(deadband[15]), .O(n29741));   // verilog/coms.v(148[4] 304[11])
    defparam i15735_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_2_lut_adj_1141 (.I0(n59384), .I1(\data_out_frame[11] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n8_adj_4853));   // verilog/coms.v(88[17:63])
    defparam i1_2_lut_adj_1141.LUT_INIT = 16'h6666;
    SB_LUT4 i5_4_lut_adj_1142 (.I0(\data_out_frame[10] [4]), .I1(\data_out_frame[11] [6]), 
            .I2(n59442), .I3(\data_out_frame[11] [5]), .O(n12_adj_4854));   // verilog/coms.v(88[17:63])
    defparam i5_4_lut_adj_1142.LUT_INIT = 16'h6996;
    SB_DFFESS data_out_frame_0___i115 (.Q(\data_out_frame[14] [2]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4855), .S(n58578));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_4_lut_adj_1143 (.I0(\data_out_frame[14] [1]), .I1(n58782), 
            .I2(n12_adj_4854), .I3(n8_adj_4853), .O(n59171));
    defparam i1_4_lut_adj_1143.LUT_INIT = 16'h9669;
    SB_LUT4 i2_3_lut_adj_1144 (.I0(n58873), .I1(\data_out_frame[8] [4]), 
            .I2(\data_out_frame[6] [1]), .I3(GND_net), .O(n58861));   // verilog/coms.v(77[16:43])
    defparam i2_3_lut_adj_1144.LUT_INIT = 16'h9696;
    SB_DFFE data_in_frame_0___i19 (.Q(\data_in_frame[2] [2]), .C(clk16MHz), 
            .E(VCC_net), .D(n29807));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i15734_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n37), .I2(\data_in_frame[14] [0]), 
            .I3(deadband[16]), .O(n29740));   // verilog/coms.v(148[4] 304[11])
    defparam i15734_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFFESS data_out_frame_0___i116 (.Q(\data_out_frame[14] [3]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4856), .S(n58577));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i117 (.Q(\data_out_frame[14] [4]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4857), .S(n58576));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i118 (.Q(\data_out_frame[14] [5]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4858), .S(n58575));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i4_4_lut_adj_1145 (.I0(n26143), .I1(\data_out_frame[9] [2]), 
            .I2(n58910), .I3(n6_adj_4859), .O(n26347));   // verilog/coms.v(100[12:26])
    defparam i4_4_lut_adj_1145.LUT_INIT = 16'h6996;
    SB_LUT4 i911_2_lut (.I0(\data_out_frame[13] [7]), .I1(\data_out_frame[13] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n1699));   // verilog/coms.v(74[16:27])
    defparam i911_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i15733_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n37), .I2(\data_in_frame[14] [1]), 
            .I3(deadband[17]), .O(n29739));   // verilog/coms.v(148[4] 304[11])
    defparam i15733_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFFESS data_out_frame_0___i119 (.Q(\data_out_frame[14] [6]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4860), .S(n58574));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_adj_1146 (.I0(\data_out_frame[6] [0]), .I1(\data_out_frame[5] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n25682));   // verilog/coms.v(75[16:27])
    defparam i1_2_lut_adj_1146.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1147 (.I0(n26347), .I1(n53470), .I2(GND_net), 
            .I3(GND_net), .O(n54430));
    defparam i1_2_lut_adj_1147.LUT_INIT = 16'h6666;
    SB_LUT4 i15745_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n37), .I2(\data_in_frame[16] [5]), 
            .I3(deadband[5]), .O(n29751));   // verilog/coms.v(148[4] 304[11])
    defparam i15745_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i23371_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n37), .I2(\data_in_frame[16] [1]), 
            .I3(deadband[1]), .O(n29755));   // verilog/coms.v(148[4] 304[11])
    defparam i23371_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_2_lut_adj_1148 (.I0(\data_out_frame[9] [3]), .I1(\data_out_frame[9] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n26046));
    defparam i1_2_lut_adj_1148.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1149 (.I0(n1169), .I1(n26143), .I2(n26483), .I3(n26046), 
            .O(n59112));
    defparam i3_4_lut_adj_1149.LUT_INIT = 16'h6996;
    SB_DFFE data_in_frame_0___i18 (.Q(\data_in_frame[2] [1]), .C(clk16MHz), 
            .E(VCC_net), .D(n29804));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_adj_1150 (.I0(\data_out_frame[7] [1]), .I1(n26039), 
            .I2(GND_net), .I3(GND_net), .O(n26483));
    defparam i1_2_lut_adj_1150.LUT_INIT = 16'h6666;
    SB_DFFESS data_out_frame_0___i120 (.Q(\data_out_frame[14] [7]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4861), .S(n58573));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i121 (.Q(\data_out_frame[15] [0]), .C(clk16MHz), 
            .E(n30510), .D(n2_adj_4862), .S(n28959));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 mux_1052_i1_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n37), .I2(\data_in_frame[3] [0]), 
            .I3(\data_in_frame[19] [0]), .O(n4760[0]));   // verilog/coms.v(148[4] 304[11])
    defparam mux_1052_i1_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 i1_2_lut_adj_1151 (.I0(\data_out_frame[4] [7]), .I1(n58897), 
            .I2(GND_net), .I3(GND_net), .O(n1169));   // verilog/coms.v(74[16:62])
    defparam i1_2_lut_adj_1151.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1152 (.I0(n26298), .I1(\data_out_frame[11] [4]), 
            .I2(\data_out_frame[9] [3]), .I3(GND_net), .O(n58910));
    defparam i2_3_lut_adj_1152.LUT_INIT = 16'h9696;
    SB_DFFE data_in_frame_0___i17 (.Q(\data_in_frame[2] [0]), .C(clk16MHz), 
            .E(VCC_net), .D(n29801));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i15748_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n37), .I2(\data_in_frame[16] [2]), 
            .I3(deadband[2]), .O(n29754));   // verilog/coms.v(148[4] 304[11])
    defparam i15748_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2_2_lut_adj_1153 (.I0(\data_out_frame[11] [3]), .I1(\data_out_frame[9] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n8_adj_4863));
    defparam i2_2_lut_adj_1153.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1154 (.I0(n58910), .I1(n26563), .I2(\data_out_frame[8] [7]), 
            .I3(n1169), .O(n7_adj_4864));
    defparam i1_4_lut_adj_1154.LUT_INIT = 16'h6996;
    SB_DFFE data_in_frame_0___i16 (.Q(\data_in_frame[1] [7]), .C(clk16MHz), 
            .E(VCC_net), .D(n29798));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i5_4_lut_adj_1155 (.I0(n26483), .I1(n7_adj_4864), .I2(\data_out_frame[13] [5]), 
            .I3(n8_adj_4863), .O(n26739));
    defparam i5_4_lut_adj_1155.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1156 (.I0(n1312), .I1(n59112), .I2(\data_out_frame[11] [5]), 
            .I3(GND_net), .O(n53470));
    defparam i2_3_lut_adj_1156.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1157 (.I0(n26022), .I1(n59350), .I2(\data_out_frame[14] [0]), 
            .I3(GND_net), .O(n26649));
    defparam i2_3_lut_adj_1157.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1158 (.I0(n26649), .I1(n53470), .I2(n26739), 
            .I3(GND_net), .O(n53640));
    defparam i2_3_lut_adj_1158.LUT_INIT = 16'h9696;
    SB_LUT4 i1047_2_lut (.I0(\data_out_frame[15] [7]), .I1(\data_out_frame[15] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n1835));   // verilog/coms.v(74[16:27])
    defparam i1047_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i15732_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n37), .I2(\data_in_frame[14] [2]), 
            .I3(deadband[18]), .O(n29738));   // verilog/coms.v(148[4] 304[11])
    defparam i15732_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i15731_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n37), .I2(\data_in_frame[14] [3]), 
            .I3(deadband[19]), .O(n29737));   // verilog/coms.v(148[4] 304[11])
    defparam i15731_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFFE data_in_frame_0___i15 (.Q(\data_in_frame[1] [6]), .C(clk16MHz), 
            .E(VCC_net), .D(n29795));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i2_3_lut_adj_1159 (.I0(\data_out_frame[4] [4]), .I1(\data_out_frame[4] [3]), 
            .I2(\data_out_frame[6] [5]), .I3(GND_net), .O(n26563));
    defparam i2_3_lut_adj_1159.LUT_INIT = 16'h9696;
    SB_LUT4 i4_4_lut_adj_1160 (.I0(\data_out_frame[9] [5]), .I1(\data_out_frame[7] [4]), 
            .I2(\data_out_frame[5] [1]), .I3(n6_adj_4865), .O(n26022));   // verilog/coms.v(76[16:34])
    defparam i4_4_lut_adj_1160.LUT_INIT = 16'h6996;
    SB_LUT4 i15730_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n37), .I2(\data_in_frame[14] [4]), 
            .I3(deadband[20]), .O(n29736));   // verilog/coms.v(148[4] 304[11])
    defparam i15730_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_2_lut_adj_1161 (.I0(\data_out_frame[4] [7]), .I1(\data_out_frame[7] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n58931));
    defparam i1_2_lut_adj_1161.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1162 (.I0(n25614), .I1(n58931), .I2(n26039), 
            .I3(GND_net), .O(n1312));
    defparam i2_3_lut_adj_1162.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1163 (.I0(\data_out_frame[9] [4]), .I1(n59012), 
            .I2(GND_net), .I3(GND_net), .O(n59350));
    defparam i1_2_lut_adj_1163.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_4_lut_4_lut (.I0(n54458), .I1(n59067), .I2(n54516), 
            .I3(n58969), .O(n58771));
    defparam i1_2_lut_4_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1164 (.I0(\data_out_frame[9] [7]), .I1(\data_out_frame[10] [0]), 
            .I2(n25611), .I3(n26022), .O(n59323));   // verilog/coms.v(79[16:43])
    defparam i3_4_lut_adj_1164.LUT_INIT = 16'h6996;
    SB_DFFE data_in_frame_0___i14 (.Q(\data_in_frame[1] [5]), .C(clk16MHz), 
            .E(VCC_net), .D(n29792));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i2_2_lut_adj_1165 (.I0(\data_out_frame[7] [4]), .I1(n59323), 
            .I2(GND_net), .I3(GND_net), .O(n10_adj_4866));   // verilog/coms.v(77[16:27])
    defparam i2_2_lut_adj_1165.LUT_INIT = 16'h6666;
    SB_LUT4 i6_4_lut_adj_1166 (.I0(\data_out_frame[12] [1]), .I1(n58941), 
            .I2(n59326), .I3(\data_out_frame[12] [0]), .O(n14_adj_4867));   // verilog/coms.v(77[16:27])
    defparam i6_4_lut_adj_1166.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1167 (.I0(\data_out_frame[14] [2]), .I1(n14_adj_4867), 
            .I2(n10_adj_4866), .I3(n59350), .O(n59124));   // verilog/coms.v(77[16:27])
    defparam i7_4_lut_adj_1167.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1168 (.I0(\data_out_frame[11] [0]), .I1(\data_out_frame[11] [1]), 
            .I2(\data_out_frame[8] [4]), .I3(GND_net), .O(n59287));   // verilog/coms.v(77[16:43])
    defparam i2_3_lut_adj_1168.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1169 (.I0(\data_out_frame[8] [5]), .I1(\data_out_frame[8] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n59436));   // verilog/coms.v(77[16:43])
    defparam i1_2_lut_adj_1169.LUT_INIT = 16'h6666;
    SB_LUT4 i15729_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n37), .I2(\data_in_frame[14] [5]), 
            .I3(deadband[21]), .O(n29735));   // verilog/coms.v(148[4] 304[11])
    defparam i15729_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i342_2_lut (.I0(\data_out_frame[4] [5]), .I1(\data_out_frame[4] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n1130));   // verilog/coms.v(79[16:27])
    defparam i342_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1170 (.I0(\data_out_frame[5] [2]), .I1(\data_out_frame[5] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n25614));   // verilog/coms.v(76[16:34])
    defparam i1_2_lut_adj_1170.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1171 (.I0(\data_out_frame[5] [3]), .I1(\data_out_frame[5] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n25611));   // verilog/coms.v(74[16:62])
    defparam i1_2_lut_adj_1171.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1172 (.I0(\data_out_frame[6] [4]), .I1(\data_out_frame[8] [6]), 
            .I2(\data_out_frame[4] [2]), .I3(GND_net), .O(n58821));   // verilog/coms.v(77[16:27])
    defparam i2_3_lut_adj_1172.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_1173 (.I0(\data_out_frame[8] [5]), .I1(n58972), 
            .I2(\data_out_frame[6] [3]), .I3(\data_out_frame[4] [1]), .O(n26376));   // verilog/coms.v(78[16:43])
    defparam i3_4_lut_adj_1173.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1174 (.I0(n25611), .I1(n25614), .I2(n1191), .I3(\data_out_frame[5] [4]), 
            .O(n58897));   // verilog/coms.v(74[16:62])
    defparam i3_4_lut_adj_1174.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1175 (.I0(\data_out_frame[4] [5]), .I1(n58897), 
            .I2(\data_out_frame[5] [0]), .I3(\data_out_frame[6] [7]), .O(n26143));   // verilog/coms.v(74[16:62])
    defparam i3_4_lut_adj_1175.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1176 (.I0(\data_out_frame[8] [7]), .I1(n26298), 
            .I2(GND_net), .I3(GND_net), .O(n58887));
    defparam i1_2_lut_adj_1176.LUT_INIT = 16'h6666;
    SB_LUT4 i6_4_lut_adj_1177 (.I0(n59436), .I1(\data_out_frame[8] [7]), 
            .I2(n59287), .I3(\data_out_frame[10] [6]), .O(n14_adj_4868));   // verilog/coms.v(77[16:43])
    defparam i6_4_lut_adj_1177.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1178 (.I0(\data_out_frame[13] [2]), .I1(n14_adj_4868), 
            .I2(n10_adj_4869), .I3(n58873), .O(n25650));   // verilog/coms.v(77[16:43])
    defparam i7_4_lut_adj_1178.LUT_INIT = 16'h6996;
    SB_DFFE data_in_frame_0___i13 (.Q(\data_in_frame[1] [4]), .C(clk16MHz), 
            .E(VCC_net), .D(n29789));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_adj_1179 (.I0(\data_out_frame[13] [1]), .I1(n26563), 
            .I2(GND_net), .I3(GND_net), .O(n59462));   // verilog/coms.v(77[16:27])
    defparam i1_2_lut_adj_1179.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1180 (.I0(n25650), .I1(n26210), .I2(GND_net), 
            .I3(GND_net), .O(n1720));   // verilog/coms.v(77[16:43])
    defparam i1_2_lut_adj_1180.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1181 (.I0(\data_out_frame[14] [4]), .I1(n59124), 
            .I2(GND_net), .I3(GND_net), .O(n53638));
    defparam i1_2_lut_adj_1181.LUT_INIT = 16'h6666;
    SB_LUT4 i14_4_lut_adj_1182 (.I0(\data_out_frame[10] [7]), .I1(n53638), 
            .I2(n1720), .I3(n59462), .O(n36_adj_4870));
    defparam i14_4_lut_adj_1182.LUT_INIT = 16'h6996;
    SB_DFFE data_in_frame_0___i190 (.Q(\data_in_frame[23] [5]), .C(clk16MHz), 
            .E(VCC_net), .D(n29786));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i12_4_lut_adj_1183 (.I0(n58855), .I1(n25640), .I2(n59436), 
            .I3(n59268), .O(n34));
    defparam i12_4_lut_adj_1183.LUT_INIT = 16'h6996;
    SB_LUT4 i18_4_lut_adj_1184 (.I0(\data_out_frame[8] [1]), .I1(n36_adj_4870), 
            .I2(n26_adj_4871), .I3(n1835), .O(n40_adj_4872));
    defparam i18_4_lut_adj_1184.LUT_INIT = 16'h6996;
    SB_LUT4 i16_4_lut_adj_1185 (.I0(n58833), .I1(n54430), .I2(n25682), 
            .I3(n1699), .O(n38));
    defparam i16_4_lut_adj_1185.LUT_INIT = 16'h9669;
    SB_LUT4 i17_3_lut (.I0(n53640), .I1(n34), .I2(\data_out_frame[14] [3]), 
            .I3(GND_net), .O(n39_adj_4873));
    defparam i17_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i15728_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n37), .I2(\data_in_frame[14] [6]), 
            .I3(deadband[22]), .O(n29734));   // verilog/coms.v(148[4] 304[11])
    defparam i15728_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i15_4_lut_adj_1186 (.I0(n59418), .I1(n59171), .I2(n59305), 
            .I3(n58944), .O(n37_adj_4874));
    defparam i15_4_lut_adj_1186.LUT_INIT = 16'h6996;
    SB_DFFE data_in_frame_0___i12 (.Q(\data_in_frame[1] [3]), .C(clk16MHz), 
            .E(VCC_net), .D(n29783));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i21_4_lut (.I0(n37_adj_4874), .I1(n39_adj_4873), .I2(n38), 
            .I3(n40_adj_4872), .O(n53515));
    defparam i21_4_lut.LUT_INIT = 16'h6996;
    SB_DFFE data_in_frame_0___i11 (.Q(\data_in_frame[1] [2]), .C(clk16MHz), 
            .E(VCC_net), .D(n29780));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_adj_1187 (.I0(n70020), .I1(n54620), .I2(GND_net), 
            .I3(GND_net), .O(n59481));
    defparam i1_2_lut_adj_1187.LUT_INIT = 16'h6666;
    SB_LUT4 i15727_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n37), .I2(\data_in_frame[14] [7]), 
            .I3(deadband[23]), .O(n29733));   // verilog/coms.v(148[4] 304[11])
    defparam i15727_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFFE data_in_frame_0___i10 (.Q(\data_in_frame[1] [1]), .C(clk16MHz), 
            .E(VCC_net), .D(n29777));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i9 (.Q(\data_in_frame[1] [0]), .C(clk16MHz), 
            .E(VCC_net), .D(n29774));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i2_3_lut_adj_1188 (.I0(\data_out_frame[16] [3]), .I1(n59455), 
            .I2(\data_out_frame[16] [4]), .I3(GND_net), .O(n58785));
    defparam i2_3_lut_adj_1188.LUT_INIT = 16'h9696;
    SB_DFFE data_in_frame_0___i8 (.Q(\data_in_frame[0] [7]), .C(clk16MHz), 
            .E(VCC_net), .D(n29771));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_adj_1189 (.I0(n53489), .I1(n59244), .I2(GND_net), 
            .I3(GND_net), .O(n6_adj_4875));
    defparam i1_2_lut_adj_1189.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1190 (.I0(\data_out_frame[21] [3]), .I1(\data_out_frame[17] [1]), 
            .I2(n26225), .I3(n6_adj_4875), .O(n53583));
    defparam i4_4_lut_adj_1190.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1191 (.I0(\data_out_frame[21] [2]), .I1(n54479), 
            .I2(\data_out_frame[19] [0]), .I3(n54450), .O(n53546));
    defparam i3_4_lut_adj_1191.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut (.I0(\byte_transmit_counter[1] ), 
            .I1(n64430), .I2(n64431), .I3(\byte_transmit_counter[2] ), 
            .O(n71078));
    defparam byte_transmit_counter_1__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_DFF data_in_frame_0___i2 (.Q(\data_in_frame[0] [1]), .C(clk16MHz), 
           .D(n29639));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i3 (.Q(\data_in_frame[0]_c [2]), .C(clk16MHz), 
           .D(n58138));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i4 (.Q(\data_in_frame[0][3] ), .C(clk16MHz), 
           .D(n29650));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i183 (.Q(\data_in_frame[22] [6]), .C(clk16MHz), 
           .D(n29653));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i184 (.Q(\data_in_frame[22] [7]), .C(clk16MHz), 
           .D(n29656));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i2_3_lut_adj_1192 (.I0(n53546), .I1(n53583), .I2(\data_out_frame[23] [4]), 
            .I3(GND_net), .O(n60824));
    defparam i2_3_lut_adj_1192.LUT_INIT = 16'h9696;
    SB_DFF data_in_frame_0___i185 (.Q(\data_in_frame[23] [0]), .C(clk16MHz), 
           .D(n29765));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_adj_1193 (.I0(\data_out_frame[6] [2]), .I1(\data_out_frame[10] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n59415));   // verilog/coms.v(75[16:27])
    defparam i1_2_lut_adj_1193.LUT_INIT = 16'h6666;
    SB_DFF data_in_frame_0___i186 (.Q(\data_in_frame[23] [1]), .C(clk16MHz), 
           .D(n29764));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i187 (.Q(\data_in_frame[23] [2]), .C(clk16MHz), 
           .D(n57968));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i188 (.Q(\data_in_frame[23] [3]), .C(clk16MHz), 
           .D(n29668));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i5 (.Q(\data_in_frame[0]_c [4]), .C(clk16MHz), 
           .D(n58140));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i189 (.Q(\data_in_frame[23] [4]), .C(clk16MHz), 
           .D(n29674));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i6 (.Q(\data_in_frame[0]_c [5]), .C(clk16MHz), 
           .D(n58132));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 n71078_bdd_4_lut (.I0(n71078), .I1(n64482), .I2(n64481), .I3(\byte_transmit_counter[2] ), 
            .O(n71081));
    defparam n71078_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_adj_1194 (.I0(n58830), .I1(n59415), .I2(GND_net), 
            .I3(GND_net), .O(n6_adj_4876));   // verilog/coms.v(75[16:27])
    defparam i1_2_lut_adj_1194.LUT_INIT = 16'h6666;
    SB_DFFE data_in_frame_0___i7 (.Q(\data_in_frame[0][6] ), .C(clk16MHz), 
            .E(VCC_net), .D(n29756));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i4_4_lut_adj_1195 (.I0(\data_out_frame[8] [3]), .I1(\data_out_frame[10] [2]), 
            .I2(n59265), .I3(n6_adj_4876), .O(n26049));   // verilog/coms.v(75[16:27])
    defparam i4_4_lut_adj_1195.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1196 (.I0(\data_out_frame[12] [5]), .I1(\data_out_frame[14] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n58833));   // verilog/coms.v(88[17:63])
    defparam i1_2_lut_adj_1196.LUT_INIT = 16'h6666;
    SB_DFFR deadband_i0_i1 (.Q(deadband[1]), .C(clk16MHz), .D(n29755), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i2_3_lut_adj_1197 (.I0(\data_out_frame[8] [0]), .I1(\data_out_frame[7] [4]), 
            .I2(\data_out_frame[7] [7]), .I3(GND_net), .O(n58867));   // verilog/coms.v(77[16:27])
    defparam i2_3_lut_adj_1197.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1198 (.I0(\data_out_frame[9] [6]), .I1(\data_out_frame[5] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n59326));   // verilog/coms.v(77[16:27])
    defparam i1_2_lut_adj_1198.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1199 (.I0(\data_out_frame[7] [6]), .I1(\data_out_frame[7] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n58950));   // verilog/coms.v(78[16:27])
    defparam i1_2_lut_adj_1199.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1200 (.I0(n58950), .I1(\data_out_frame[10] [1]), 
            .I2(\data_out_frame[5] [6]), .I3(n59326), .O(n10_adj_4877));   // verilog/coms.v(77[16:27])
    defparam i4_4_lut_adj_1200.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_1201 (.I0(n58867), .I1(n10_adj_4877), .I2(\data_out_frame[10] [0]), 
            .I3(GND_net), .O(n1510));   // verilog/coms.v(77[16:27])
    defparam i5_3_lut_adj_1201.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1202 (.I0(\data_out_frame[12] [2]), .I1(n1510), 
            .I2(GND_net), .I3(GND_net), .O(n25640));   // verilog/coms.v(77[16:43])
    defparam i1_2_lut_adj_1202.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1203 (.I0(\data_out_frame[17] [0]), .I1(n59055), 
            .I2(\data_out_frame[14] [4]), .I3(GND_net), .O(n26817));   // verilog/coms.v(77[16:43])
    defparam i2_3_lut_adj_1203.LUT_INIT = 16'h9696;
    SB_LUT4 i375_2_lut (.I0(\data_out_frame[5] [7]), .I1(\data_out_frame[5] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n1191));   // verilog/coms.v(74[16:27])
    defparam i375_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1204 (.I0(\data_out_frame[4] [3]), .I1(\data_out_frame[6] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n58972));   // verilog/coms.v(78[16:43])
    defparam i1_2_lut_adj_1204.LUT_INIT = 16'h6666;
    SB_LUT4 i5_3_lut_adj_1205 (.I0(\data_out_frame[10] [6]), .I1(\data_out_frame[10] [4]), 
            .I2(n58864), .I3(GND_net), .O(n14_adj_4878));   // verilog/coms.v(88[17:28])
    defparam i5_3_lut_adj_1205.LUT_INIT = 16'h9696;
    SB_LUT4 i4_2_lut (.I0(\data_out_frame[12] [6]), .I1(\data_out_frame[8] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n13));   // verilog/coms.v(88[17:28])
    defparam i4_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i6_4_lut_adj_1206 (.I0(n59335), .I1(\data_out_frame[12] [7]), 
            .I2(\data_out_frame[4] [2]), .I3(n58972), .O(n15_adj_4879));   // verilog/coms.v(88[17:28])
    defparam i6_4_lut_adj_1206.LUT_INIT = 16'h6996;
    SB_DFFR deadband_i0_i2 (.Q(deadband[2]), .C(clk16MHz), .D(n29754), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_4_lut_adj_1207 (.I0(n15_adj_4879), .I1(\data_out_frame[13] [0]), 
            .I2(n13), .I3(n14_adj_4878), .O(n4_c));
    defparam i1_4_lut_adj_1207.LUT_INIT = 16'h6996;
    SB_DFFR deadband_i0_i3 (.Q(deadband[3]), .C(clk16MHz), .D(n29753), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i22329_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n37), .I2(\data_in_frame[13] [1]), 
            .I3(IntegralLimit[1]), .O(n29732));   // verilog/coms.v(148[4] 304[11])
    defparam i22329_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFFR deadband_i0_i4 (.Q(deadband[4]), .C(clk16MHz), .D(n29752), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_adj_1208 (.I0(\data_out_frame[15] [0]), .I1(\data_out_frame[15] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n58855));
    defparam i1_2_lut_adj_1208.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1209 (.I0(\data_out_frame[16] [7]), .I1(\data_out_frame[19] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n26225));   // verilog/coms.v(79[16:43])
    defparam i1_2_lut_adj_1209.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1210 (.I0(\data_out_frame[16] [6]), .I1(n26817), 
            .I2(GND_net), .I3(GND_net), .O(n58802));   // verilog/coms.v(88[17:28])
    defparam i1_2_lut_adj_1210.LUT_INIT = 16'h6666;
    SB_LUT4 i15725_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n37), .I2(\data_in_frame[13] [2]), 
            .I3(IntegralLimit[2]), .O(n29731));   // verilog/coms.v(148[4] 304[11])
    defparam i15725_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_2_lut_adj_1211 (.I0(\data_out_frame[6] [3]), .I1(\data_out_frame[4] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n58883));   // verilog/coms.v(77[16:43])
    defparam i1_2_lut_adj_1211.LUT_INIT = 16'h6666;
    SB_LUT4 i15724_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n37), .I2(\data_in_frame[13] [3]), 
            .I3(IntegralLimit[3]), .O(n29730));   // verilog/coms.v(148[4] 304[11])
    defparam i15724_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i3_4_lut_adj_1212 (.I0(\data_out_frame[7] [7]), .I1(n58883), 
            .I2(\data_out_frame[10] [5]), .I3(\data_out_frame[14] [7]), 
            .O(n59418));   // verilog/coms.v(75[16:27])
    defparam i3_4_lut_adj_1212.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1213 (.I0(\data_out_frame[8] [1]), .I1(\data_out_frame[7] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n58858));   // verilog/coms.v(78[16:27])
    defparam i1_2_lut_adj_1213.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1214 (.I0(\data_out_frame[5] [3]), .I1(\data_out_frame[7] [5]), 
            .I2(\data_out_frame[9] [7]), .I3(GND_net), .O(n59229));
    defparam i2_3_lut_adj_1214.LUT_INIT = 16'h9696;
    SB_LUT4 i4_4_lut_adj_1215 (.I0(n25685), .I1(\data_out_frame[5] [7]), 
            .I2(n58858), .I3(n6_adj_4880), .O(n1513));   // verilog/coms.v(78[16:27])
    defparam i4_4_lut_adj_1215.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1216 (.I0(\data_out_frame[8] [3]), .I1(\data_out_frame[8] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n58880));   // verilog/coms.v(75[16:27])
    defparam i1_2_lut_adj_1216.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1217 (.I0(\data_out_frame[4] [1]), .I1(\data_out_frame[5] [5]), 
            .I2(\data_out_frame[8] [1]), .I3(GND_net), .O(n59265));   // verilog/coms.v(75[16:27])
    defparam i2_3_lut_adj_1217.LUT_INIT = 16'h9696;
    SB_DFFR deadband_i0_i5 (.Q(deadband[5]), .C(clk16MHz), .D(n29751), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_adj_1218 (.I0(\data_out_frame[12] [5]), .I1(\data_out_frame[12] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n59021));   // verilog/coms.v(88[17:28])
    defparam i1_2_lut_adj_1218.LUT_INIT = 16'h6666;
    SB_DFFR deadband_i0_i6 (.Q(deadband[6]), .C(clk16MHz), .D(n29750), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i7 (.Q(deadband[7]), .C(clk16MHz), .D(n29749), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i8 (.Q(deadband[8]), .C(clk16MHz), .D(n29748), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_adj_1219 (.I0(\data_out_frame[5] [4]), .I1(\data_out_frame[7] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n58941));   // verilog/coms.v(77[16:27])
    defparam i1_2_lut_adj_1219.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1220 (.I0(\data_out_frame[10] [3]), .I1(\data_out_frame[6] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n59268));   // verilog/coms.v(88[17:70])
    defparam i1_2_lut_adj_1220.LUT_INIT = 16'h6666;
    SB_LUT4 i15723_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n37), .I2(\data_in_frame[13] [4]), 
            .I3(IntegralLimit[4]), .O(n29729));   // verilog/coms.v(148[4] 304[11])
    defparam i15723_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFFR deadband_i0_i9 (.Q(deadband[9]), .C(clk16MHz), .D(n29747), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i10 (.Q(deadband[10]), .C(clk16MHz), .D(n29746), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i11 (.Q(deadband[11]), .C(clk16MHz), .D(n29745), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i12 (.Q(deadband[12]), .C(clk16MHz), .D(n29744), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i15722_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n37), .I2(\data_in_frame[13] [5]), 
            .I3(IntegralLimit[5]), .O(n29728));   // verilog/coms.v(148[4] 304[11])
    defparam i15722_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2_3_lut_adj_1221 (.I0(\data_out_frame[6] [0]), .I1(\data_out_frame[10] [2]), 
            .I2(\data_out_frame[7] [7]), .I3(GND_net), .O(n25685));   // verilog/coms.v(88[17:70])
    defparam i2_3_lut_adj_1221.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_1222 (.I0(\data_out_frame[8] [2]), .I1(n58941), 
            .I2(\data_out_frame[4] [0]), .I3(\data_out_frame[8] [0]), .O(n58830));   // verilog/coms.v(75[16:27])
    defparam i3_4_lut_adj_1222.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1223 (.I0(\data_out_frame[14] [5]), .I1(\data_out_frame[12] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_4881));   // verilog/coms.v(88[17:70])
    defparam i1_2_lut_adj_1223.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1224 (.I0(n58830), .I1(n25685), .I2(n59268), 
            .I3(n6_adj_4881), .O(n59329));   // verilog/coms.v(88[17:70])
    defparam i4_4_lut_adj_1224.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut_adj_1225 (.I0(n59021), .I1(n59265), .I2(\data_out_frame[10] [3]), 
            .I3(n58880), .O(n12_adj_4882));   // verilog/coms.v(75[16:27])
    defparam i5_4_lut_adj_1225.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1226 (.I0(\data_out_frame[5] [6]), .I1(n12_adj_4882), 
            .I2(n59418), .I3(\data_out_frame[8] [4]), .O(n53449));   // verilog/coms.v(75[16:27])
    defparam i6_4_lut_adj_1226.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1227 (.I0(\data_out_frame[17] [2]), .I1(\data_out_frame[17] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n59024));
    defparam i1_2_lut_adj_1227.LUT_INIT = 16'h6666;
    SB_DFFR deadband_i0_i13 (.Q(deadband[13]), .C(clk16MHz), .D(n29743), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i3_4_lut_adj_1228 (.I0(\data_out_frame[16] [7]), .I1(n26849), 
            .I2(n53449), .I3(\data_out_frame[15] [0]), .O(n53489));
    defparam i3_4_lut_adj_1228.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1229 (.I0(\data_out_frame[21] [5]), .I1(n53489), 
            .I2(\data_out_frame[19] [3]), .I3(n59024), .O(n10_adj_4883));
    defparam i4_4_lut_adj_1229.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_1230 (.I0(n59253), .I1(n10_adj_4883), .I2(n26716), 
            .I3(GND_net), .O(n59403));
    defparam i5_3_lut_adj_1230.LUT_INIT = 16'h9696;
    SB_LUT4 i4_4_lut_adj_1231 (.I0(n58802), .I1(n26225), .I2(\data_out_frame[21] [4]), 
            .I3(n59253), .O(n10_adj_4884));   // verilog/coms.v(79[16:43])
    defparam i4_4_lut_adj_1231.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_1232 (.I0(\data_out_frame[19] [3]), .I1(n10_adj_4884), 
            .I2(\data_out_frame[17] [2]), .I3(GND_net), .O(n53626));   // verilog/coms.v(79[16:43])
    defparam i5_3_lut_adj_1232.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_4_lut (.I0(\data_out_frame[20] [3]), .I1(\data_out_frame[20] [1]), 
            .I2(\data_out_frame[20] [2]), .I3(\data_out_frame[18] [3]), 
            .O(n6_c));
    defparam i1_2_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1233 (.I0(\data_out_frame[19] [4]), .I1(n4_c), 
            .I2(\data_out_frame[15] [0]), .I3(\data_out_frame[17] [2]), 
            .O(n10_adj_4885));
    defparam i4_4_lut_adj_1233.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_1234 (.I0(n58975), .I1(n10_adj_4885), .I2(n26716), 
            .I3(GND_net), .O(n60897));
    defparam i5_3_lut_adj_1234.LUT_INIT = 16'h9696;
    SB_DFFR deadband_i0_i14 (.Q(deadband[14]), .C(clk16MHz), .D(n29742), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_adj_1235 (.I0(reset), .I1(\FRAME_MATCHER.i_31__N_2511 ), 
            .I2(GND_net), .I3(GND_net), .O(n58672));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_adj_1235.LUT_INIT = 16'h4444;
    SB_DFFR deadband_i0_i15 (.Q(deadband[15]), .C(clk16MHz), .D(n29741), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i15721_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n37), .I2(\data_in_frame[13] [6]), 
            .I3(IntegralLimit[6]), .O(n29727));   // verilog/coms.v(148[4] 304[11])
    defparam i15721_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i15720_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n37), .I2(\data_in_frame[13] [7]), 
            .I3(IntegralLimit[7]), .O(n29726));   // verilog/coms.v(148[4] 304[11])
    defparam i15720_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFFR deadband_i0_i16 (.Q(deadband[16]), .C(clk16MHz), .D(n29740), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i3_4_lut_adj_1236 (.I0(\FRAME_MATCHER.i[0] ), .I1(n43501), .I2(\FRAME_MATCHER.i [2]), 
            .I3(\FRAME_MATCHER.i [1]), .O(n132));
    defparam i3_4_lut_adj_1236.LUT_INIT = 16'h0040;
    SB_LUT4 i4_4_lut_adj_1237 (.I0(n60897), .I1(n53626), .I2(\data_out_frame[25] [6]), 
            .I3(n59162), .O(n10_adj_4886));
    defparam i4_4_lut_adj_1237.LUT_INIT = 16'h9669;
    SB_DFFR deadband_i0_i17 (.Q(deadband[17]), .C(clk16MHz), .D(n29739), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i18 (.Q(deadband[18]), .C(clk16MHz), .D(n29738), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i26750_4_lut (.I0(n163), .I1(n67115), .I2(rx_data[7]), .I3(\data_in_frame[4] [7]), 
            .O(n40681));   // verilog/coms.v(94[13:20])
    defparam i26750_4_lut.LUT_INIT = 16'hfac0;
    SB_LUT4 i26751_3_lut (.I0(n40681), .I1(\data_in_frame[4] [7]), .I2(reset), 
            .I3(GND_net), .O(n29877));   // verilog/TinyFPGA_B.v(47[5:10])
    defparam i26751_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 select_775_Select_208_i3_4_lut (.I0(\data_out_frame[25] [7]), 
            .I1(\FRAME_MATCHER.state[3] ), .I2(n10_adj_4886), .I3(n60824), 
            .O(n3_adj_4887));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_208_i3_4_lut.LUT_INIT = 16'h8448;
    SB_DFFR deadband_i0_i19 (.Q(deadband[19]), .C(clk16MHz), .D(n29737), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i15719_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n37), .I2(\data_in_frame[12] [0]), 
            .I3(IntegralLimit[8]), .O(n29725));   // verilog/coms.v(148[4] 304[11])
    defparam i15719_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i6_2_lut_4_lut (.I0(\data_out_frame[20] [3]), .I1(\data_out_frame[20] [1]), 
            .I2(\data_out_frame[20] [2]), .I3(n59027), .O(n22));
    defparam i6_2_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1238 (.I0(n161_c), .I1(n3468), .I2(reset), .I3(n40817), 
            .O(n58720));
    defparam i3_4_lut_adj_1238.LUT_INIT = 16'hf7ff;
    SB_LUT4 select_775_Select_207_i2_4_lut (.I0(\data_out_frame[25] [7]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[7]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4889));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_207_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_775_Select_206_i2_4_lut (.I0(\data_out_frame[25] [6]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[6]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4890));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_206_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFFR deadband_i0_i20 (.Q(deadband[20]), .C(clk16MHz), .D(n29736), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i21 (.Q(deadband[21]), .C(clk16MHz), .D(n29735), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_775_Select_205_i2_4_lut (.I0(\data_out_frame[25] [5]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[5]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4891));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_205_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFFR deadband_i0_i22 (.Q(deadband[22]), .C(clk16MHz), .D(n29734), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_4_lut_adj_1239 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[25] [4]), 
            .I2(neopxl_color[4]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4892));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1239.LUT_INIT = 16'ha088;
    SB_DFFR deadband_i0_i23 (.Q(deadband[23]), .C(clk16MHz), .D(n29733), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFS IntegralLimit_i0_i1 (.Q(IntegralLimit[1]), .C(clk16MHz), .D(n29732), 
            .S(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i2 (.Q(IntegralLimit[2]), .C(clk16MHz), .D(n29731), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_775_Select_61_i2_4_lut (.I0(\data_out_frame[7] [5]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder0_position_scaled[13]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4893));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_61_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i48787_3_lut (.I0(\data_out_frame[16] [5]), .I1(\data_out_frame[17] [5]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n64481));
    defparam i48787_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48788_3_lut (.I0(\data_out_frame[18] [5]), .I1(\data_out_frame[19] [5]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n64482));
    defparam i48788_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i54315_3_lut (.I0(rx_data[5]), .I1(\data_in_frame[0]_c [5]), 
            .I2(n7), .I3(GND_net), .O(n58132));   // verilog/coms.v(94[13:20])
    defparam i54315_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFR IntegralLimit_i0_i3 (.Q(IntegralLimit[3]), .C(clk16MHz), .D(n29730), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i15718_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n37), .I2(\data_in_frame[12] [1]), 
            .I3(IntegralLimit[9]), .O(n29724));   // verilog/coms.v(148[4] 304[11])
    defparam i15718_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 select_775_Select_60_i2_4_lut (.I0(\data_out_frame[7] [4]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder0_position_scaled[12]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4895));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_60_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_775_Select_59_i2_4_lut (.I0(\data_out_frame[7] [3]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder0_position_scaled[11]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4896));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_59_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i20_4_lut (.I0(encoder1_position_scaled[16]), .I1(displacement[16]), 
            .I2(n15), .I3(n15_adj_11), .O(n19));
    defparam i20_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i54317_3_lut (.I0(rx_data[4]), .I1(\data_in_frame[0]_c [4]), 
            .I2(n7), .I3(GND_net), .O(n58140));   // verilog/coms.v(94[13:20])
    defparam i54317_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFS IntegralLimit_i0_i4 (.Q(IntegralLimit[4]), .C(clk16MHz), .D(n29729), 
            .S(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFS IntegralLimit_i0_i5 (.Q(IntegralLimit[5]), .C(clk16MHz), .D(n29728), 
            .S(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i6 (.Q(IntegralLimit[6]), .C(clk16MHz), .D(n29727), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i7 (.Q(IntegralLimit[7]), .C(clk16MHz), .D(n29726), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i8 (.Q(IntegralLimit[8]), .C(clk16MHz), .D(n29725), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i14045_3_lut (.I0(\data_out_frame[1][1] ), .I1(\data_out_frame[3][1] ), 
            .I2(\byte_transmit_counter[1] ), .I3(GND_net), .O(n28051));   // verilog/coms.v(109[34:55])
    defparam i14045_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48728_3_lut (.I0(\data_out_frame[6] [1]), .I1(\data_out_frame[7] [1]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n64422));
    defparam i48728_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48729_4_lut (.I0(n64422), .I1(n28051), .I2(\byte_transmit_counter[2] ), 
            .I3(\byte_transmit_counter[0] ), .O(n64423));
    defparam i48729_4_lut.LUT_INIT = 16'haca0;
    SB_DFFR IntegralLimit_i0_i9 (.Q(IntegralLimit[9]), .C(clk16MHz), .D(n29724), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i48727_3_lut (.I0(\data_out_frame[4] [1]), .I1(\data_out_frame[5] [1]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n64421));
    defparam i48727_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48379_2_lut (.I0(PWMLimit[1]), .I1(PWMLimit[0]), .I2(GND_net), 
            .I3(GND_net), .O(n64064));
    defparam i48379_2_lut.LUT_INIT = 16'heeee;
    SB_DFFR IntegralLimit_i0_i10 (.Q(IntegralLimit[10]), .C(clk16MHz), .D(n29723), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i11 (.Q(IntegralLimit[11]), .C(clk16MHz), .D(n29722), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i23357_4_lut (.I0(n64064), .I1(n28), .I2(n375), .I3(n376), 
            .O(n4));
    defparam i23357_4_lut.LUT_INIT = 16'h3530;
    SB_LUT4 i30053106_i1_3_lut (.I0(n71141), .I1(n70895), .I2(\byte_transmit_counter[2] ), 
            .I3(GND_net), .O(n14_adj_4902));
    defparam i30053106_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 select_775_Select_58_i2_4_lut (.I0(\data_out_frame[7] [2]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder0_position_scaled[10]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4903));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_58_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFFR IntegralLimit_i0_i12 (.Q(IntegralLimit[12]), .C(clk16MHz), .D(n29721), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i13 (.Q(IntegralLimit[13]), .C(clk16MHz), .D(n29720), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i14 (.Q(IntegralLimit[14]), .C(clk16MHz), .D(n29719), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i15 (.Q(IntegralLimit[15]), .C(clk16MHz), .D(n29718), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i16 (.Q(IntegralLimit[16]), .C(clk16MHz), .D(n29717), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i17 (.Q(IntegralLimit[17]), .C(clk16MHz), .D(n29716), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i18 (.Q(IntegralLimit[18]), .C(clk16MHz), .D(n29715), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i19 (.Q(IntegralLimit[19]), .C(clk16MHz), .D(n29714), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i22584_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n37), .I2(\data_in_frame[12] [4]), 
            .I3(IntegralLimit[12]), .O(n29721));   // verilog/coms.v(148[4] 304[11])
    defparam i22584_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFFR IntegralLimit_i0_i20 (.Q(IntegralLimit[20]), .C(clk16MHz), .D(n29713), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i22583_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n37), .I2(\data_in_frame[12] [3]), 
            .I3(IntegralLimit[11]), .O(n29722));   // verilog/coms.v(148[4] 304[11])
    defparam i22583_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFFR IntegralLimit_i0_i21 (.Q(IntegralLimit[21]), .C(clk16MHz), .D(n29712), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i22 (.Q(IntegralLimit[22]), .C(clk16MHz), .D(n29711), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i23 (.Q(IntegralLimit[23]), .C(clk16MHz), .D(n29710), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFS Kp_i1 (.Q(\Kp[1] ), .C(clk16MHz), .D(n29709), .S(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Kp_i2 (.Q(\Kp[2] ), .C(clk16MHz), .D(n29708), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i54316_3_lut (.I0(rx_data[2]), .I1(\data_in_frame[0]_c [2]), 
            .I2(n7), .I3(GND_net), .O(n58138));   // verilog/coms.v(94[13:20])
    defparam i54316_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFS Kp_i3 (.Q(\Kp[3] ), .C(clk16MHz), .D(n29707), .S(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i122 (.Q(\data_out_frame[15] [1]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4794), .S(n58572));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i123 (.Q(\data_out_frame[15] [2]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4793), .S(n58571));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Kp_i4 (.Q(\Kp[4] ), .C(clk16MHz), .D(n29706), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i124 (.Q(\data_out_frame[15] [3]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4792), .S(n58570));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i125 (.Q(\data_out_frame[15] [4]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4790), .S(n58569));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Kp_i5 (.Q(\Kp[5] ), .C(clk16MHz), .D(n29705), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_775_Select_203_i2_4_lut (.I0(\data_out_frame[25] [3]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[3]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4904));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_203_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i48737_3_lut (.I0(\data_out_frame[22] [5]), .I1(\data_out_frame[23] [5]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n64431));
    defparam i48737_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48736_3_lut (.I0(\data_out_frame[20] [5]), .I1(\data_out_frame[21] [5]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n64430));
    defparam i48736_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1240 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[25] [2]), 
            .I2(neopxl_color[2]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4905));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1240.LUT_INIT = 16'ha088;
    SB_DFFR Kp_i6 (.Q(\Kp[6] ), .C(clk16MHz), .D(n29704), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Kp_i7 (.Q(\Kp[7] ), .C(clk16MHz), .D(n29703), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i15717_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n37), .I2(\data_in_frame[12] [2]), 
            .I3(IntegralLimit[10]), .O(n29723));   // verilog/coms.v(148[4] 304[11])
    defparam i15717_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFFR Kp_i8 (.Q(\Kp[8] ), .C(clk16MHz), .D(n29702), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i126 (.Q(\data_out_frame[15] [5]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4789), .S(n58568));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 equal_1931_i7_2_lut_4_lut (.I0(\data_in_frame[6] [5]), .I1(Kp_23__N_878), 
            .I2(n58818), .I3(\data_in_frame[8] [6]), .O(n7_adj_4906));   // verilog/coms.v(239[9:81])
    defparam equal_1931_i7_2_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 select_775_Select_201_i2_4_lut (.I0(\data_out_frame[25] [1]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[1]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4907));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_201_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFFESS data_out_frame_0___i127 (.Q(\data_out_frame[15] [6]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4786), .S(n58567));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Kp_i9 (.Q(\Kp[9] ), .C(clk16MHz), .D(n29701), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i128 (.Q(\data_out_frame[15] [7]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4784), .S(n58566));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i129 (.Q(\data_out_frame[16] [0]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4783), .S(n58565));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i130 (.Q(\data_out_frame[16] [1]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4782), .S(n58564));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Kp_i10 (.Q(\Kp[10] ), .C(clk16MHz), .D(n29700), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_775_Select_200_i2_4_lut (.I0(\data_out_frame[25] [0]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[0]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4908));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_200_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFFR Kp_i11 (.Q(\Kp[11] ), .C(clk16MHz), .D(n29699), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Kp_i12 (.Q(\Kp[12] ), .C(clk16MHz), .D(n29698), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Kp_i13 (.Q(\Kp[13] ), .C(clk16MHz), .D(n29697), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_775_Select_199_i2_4_lut (.I0(\data_out_frame[24] [7]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[15]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4909));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_199_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFFR Kp_i14 (.Q(\Kp[14] ), .C(clk16MHz), .D(n29696), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i131 (.Q(\data_out_frame[16] [2]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4780), .S(n58496));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_775_Select_198_i2_4_lut (.I0(\data_out_frame[24] [6]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[14]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4910));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_198_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFFR Kp_i15 (.Q(\Kp[15] ), .C(clk16MHz), .D(n29695), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i132 (.Q(\data_out_frame[16] [3]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4775), .S(n58499));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Ki_i1 (.Q(\Ki[1] ), .C(clk16MHz), .D(n29694), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_3_i1_3_lut (.I0(\data_out_frame[0][3] ), 
            .I1(\data_out_frame[1][3] ), .I2(\byte_transmit_counter[0] ), 
            .I3(GND_net), .O(n1));   // verilog/coms.v(109[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_3_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 select_775_Select_197_i2_4_lut (.I0(\data_out_frame[24] [5]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[13]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4911));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_197_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFFR Ki_i2 (.Q(\Ki[2] ), .C(clk16MHz), .D(n29693), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Ki_i3 (.Q(\Ki[3] ), .C(clk16MHz), .D(n29692), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Ki_i4 (.Q(\Ki[4] ), .C(clk16MHz), .D(n29691), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Ki_i5 (.Q(\Ki[5] ), .C(clk16MHz), .D(n29690), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Ki_i6 (.Q(\Ki[6] ), .C(clk16MHz), .D(n29689), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i133 (.Q(\data_out_frame[16] [4]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4774), .S(n28947));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i48688_4_lut (.I0(n1), .I1(\data_out_frame[3][3] ), .I2(\byte_transmit_counter[1] ), 
            .I3(\byte_transmit_counter[0] ), .O(n64382));
    defparam i48688_4_lut.LUT_INIT = 16'hca0a;
    SB_LUT4 i16139_3_lut_4_lut (.I0(n58731), .I1(n58752), .I2(rx_data[7]), 
            .I3(\data_in_frame[13] [7]), .O(n30145));
    defparam i16139_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i48778_3_lut (.I0(\data_out_frame[8] [4]), .I1(\data_out_frame[9] [4]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n64472));
    defparam i48778_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFR Ki_i7 (.Q(\Ki[7] ), .C(clk16MHz), .D(n29688), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i134 (.Q(\data_out_frame[16] [5]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4773), .S(n58500));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_775_Select_196_i2_4_lut (.I0(\data_out_frame[24] [4]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[12]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4912));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_196_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFFESS data_out_frame_0___i135 (.Q(\data_out_frame[16] [6]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4772), .S(n28945));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i136 (.Q(\data_out_frame[16] [7]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4770), .S(n58501));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i137 (.Q(\data_out_frame[17] [0]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4769), .S(n58503));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Ki_i8 (.Q(\Ki[8] ), .C(clk16MHz), .D(n29687), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i48779_3_lut (.I0(\data_out_frame[10] [4]), .I1(\data_out_frame[11] [4]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n64473));
    defparam i48779_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1241 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[24] [3]), 
            .I2(neopxl_color[11]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4913));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1241.LUT_INIT = 16'ha088;
    SB_LUT4 select_775_Select_194_i2_4_lut (.I0(\data_out_frame[24] [2]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[10]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4914));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_194_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFFR Ki_i9 (.Q(\Ki[9] ), .C(clk16MHz), .D(n29686), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Ki_i10 (.Q(\Ki[10] ), .C(clk16MHz), .D(n29685), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i48764_3_lut (.I0(\data_out_frame[14] [4]), .I1(\data_out_frame[15] [4]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n64458));
    defparam i48764_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFR Ki_i11 (.Q(\Ki[11] ), .C(clk16MHz), .D(n29684), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Ki_i12 (.Q(\Ki[12] ), .C(clk16MHz), .D(n29683), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Ki_i13 (.Q(\Ki[13] ), .C(clk16MHz), .D(n29682), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_775_Select_193_i2_4_lut (.I0(\data_out_frame[24] [1]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[9]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4915));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_193_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i48763_3_lut (.I0(\data_out_frame[12] [4]), .I1(\data_out_frame[13] [4]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n64457));
    defparam i48763_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48790_3_lut (.I0(\data_out_frame[8] [0]), .I1(\data_out_frame[9] [0]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n64484));
    defparam i48790_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48791_3_lut (.I0(\data_out_frame[10] [0]), .I1(\data_out_frame[11] [0]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n64485));
    defparam i48791_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFESS data_out_frame_0___i138 (.Q(\data_out_frame[17] [1]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4759), .S(n58505));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Ki_i14 (.Q(\Ki[14] ), .C(clk16MHz), .D(n29681), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_775_Select_192_i2_4_lut (.I0(\data_out_frame[24] [0]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[8]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4916));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_192_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_775_Select_191_i2_4_lut (.I0(\data_out_frame[23] [7]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[23]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4917));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_191_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_775_Select_190_i2_4_lut (.I0(\data_out_frame[23] [6]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[22]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4918));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_190_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i48707_3_lut (.I0(\data_out_frame[14] [0]), .I1(\data_out_frame[15] [0]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n64401));
    defparam i48707_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48706_3_lut (.I0(\data_out_frame[12] [0]), .I1(\data_out_frame[13] [0]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n64400));
    defparam i48706_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFR Ki_i15 (.Q(\Ki[15] ), .C(clk16MHz), .D(n29680), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i139 (.Q(\data_out_frame[17] [2]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4757), .S(n58507));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_775_Select_189_i2_4_lut (.I0(\data_out_frame[23] [5]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[21]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4919));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_189_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i48793_3_lut (.I0(\data_out_frame[8] [6]), .I1(\data_out_frame[9] [6]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n64487));
    defparam i48793_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFESS data_out_frame_0___i140 (.Q(\data_out_frame[17] [3]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4754), .S(n58508));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i141 (.Q(\data_out_frame[17] [4]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4753), .S(n58509));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i142 (.Q(\data_out_frame[17] [5]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4752), .S(n58510));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i143 (.Q(\data_out_frame[17] [6]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4751), .S(n58511));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i144 (.Q(\data_out_frame[17] [7]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4749), .S(n58512));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i48794_3_lut (.I0(\data_out_frame[10] [6]), .I1(\data_out_frame[11] [6]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n64488));
    defparam i48794_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16096_3_lut_4_lut (.I0(n58731), .I1(n58752), .I2(rx_data[6]), 
            .I3(\data_in_frame[13] [6]), .O(n30102));
    defparam i16096_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i48674_3_lut (.I0(\data_out_frame[14] [6]), .I1(\data_out_frame[15] [6]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n64368));
    defparam i48674_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 select_775_Select_188_i2_4_lut (.I0(\data_out_frame[23] [4]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[20]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4920));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_188_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i48673_3_lut (.I0(\data_out_frame[12] [6]), .I1(\data_out_frame[13] [6]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n64367));
    defparam i48673_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFESS data_out_frame_0___i145 (.Q(\data_out_frame[18] [0]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4748), .S(n58513));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i53493_3_lut (.I0(n71165), .I1(n71003), .I2(\byte_transmit_counter[2] ), 
            .I3(GND_net), .O(n69187));
    defparam i53493_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFESS data_out_frame_0___i146 (.Q(\data_out_frame[18] [1]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4734), .S(n58514));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i147 (.Q(\data_out_frame[18] [2]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4921), .S(n58515));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i148 (.Q(\data_out_frame[18] [3]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4922), .S(n58493));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i149 (.Q(\data_out_frame[18] [4]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4923), .S(n58516));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i150 (.Q(\data_out_frame[18] [5]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4924), .S(n58517));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i151 (.Q(\data_out_frame[18] [6]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4925), .S(n28929));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i152 (.Q(\data_out_frame[18] [7]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4926), .S(n28928));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i153 (.Q(\data_out_frame[19] [0]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4927), .S(n58518));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_775_Select_187_i2_4_lut (.I0(\data_out_frame[23] [3]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[19]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4928));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_187_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFFESS data_out_frame_0___i154 (.Q(\data_out_frame[19] [1]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4929), .S(n58519));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i155 (.Q(\data_out_frame[19] [2]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4930), .S(n58520));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i3_4_lut_adj_1242 (.I0(reset), .I1(\FRAME_MATCHER.i[0] ), .I2(n40660), 
            .I3(n161_c), .O(n58752));
    defparam i3_4_lut_adj_1242.LUT_INIT = 16'hfbff;
    SB_LUT4 i14039_3_lut (.I0(\data_out_frame[1][6] ), .I1(\data_out_frame[3][6] ), 
            .I2(\byte_transmit_counter[1] ), .I3(GND_net), .O(n28045));   // verilog/coms.v(109[34:55])
    defparam i14039_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF \FRAME_MATCHER.rx_data_ready_prev_4012  (.Q(\FRAME_MATCHER.rx_data_ready_prev ), 
           .C(clk16MHz), .D(n29643));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i16093_3_lut_4_lut (.I0(n58731), .I1(n58752), .I2(rx_data[5]), 
            .I3(\data_in_frame[13] [5]), .O(n30099));
    defparam i16093_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF neopxl_color_i0_i1 (.Q(neopxl_color[1]), .C(clk16MHz), .D(n29642));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i2_3_lut_adj_1243 (.I0(n3468), .I1(n58752), .I2(n40817), .I3(GND_net), 
            .O(n61932));
    defparam i2_3_lut_adj_1243.LUT_INIT = 16'hdfdf;
    SB_LUT4 i48710_3_lut (.I0(\data_out_frame[6] [6]), .I1(\data_out_frame[7] [6]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n64404));
    defparam i48710_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48711_4_lut (.I0(n64404), .I1(n28045), .I2(\byte_transmit_counter[2] ), 
            .I3(\byte_transmit_counter[0] ), .O(n64405));
    defparam i48711_4_lut.LUT_INIT = 16'haca0;
    SB_LUT4 i16089_3_lut_4_lut (.I0(n58731), .I1(n58752), .I2(rx_data[4]), 
            .I3(\data_in_frame[13] [4]), .O(n30095));
    defparam i16089_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i48709_3_lut (.I0(\data_out_frame[4] [6]), .I1(\data_out_frame[5] [6]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n64403));
    defparam i48709_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 select_775_Select_57_i2_4_lut (.I0(\data_out_frame[7] [1]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder0_position_scaled[9]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4931));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_57_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i51953_2_lut (.I0(n70961), .I1(\byte_transmit_counter[2] ), 
            .I2(GND_net), .I3(GND_net), .O(n67143));
    defparam i51953_2_lut.LUT_INIT = 16'h2222;
    SB_DFF neopxl_color_i0_i14 (.Q(neopxl_color[14]), .C(clk16MHz), .D(n29638));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_775_Select_56_i2_4_lut (.I0(\data_out_frame[7] [0]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder0_position_scaled[8]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4932));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_56_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i53505_3_lut (.I0(n71207), .I1(n70955), .I2(\byte_transmit_counter[2] ), 
            .I3(GND_net), .O(n69199));
    defparam i53505_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14037_3_lut (.I0(\data_out_frame[1][7] ), .I1(\data_out_frame[3][7] ), 
            .I2(\byte_transmit_counter[1] ), .I3(GND_net), .O(n28043));   // verilog/coms.v(109[34:55])
    defparam i14037_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48701_3_lut (.I0(\data_out_frame[6] [7]), .I1(\data_out_frame[7] [7]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n64395));
    defparam i48701_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1244 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[6] [7]), 
            .I2(encoder0_position_scaled[23]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4933));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1244.LUT_INIT = 16'ha088;
    SB_LUT4 i1_4_lut_adj_1245 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[6] [6]), 
            .I2(encoder0_position_scaled[22]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4934));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1245.LUT_INIT = 16'ha088;
    SB_LUT4 i48702_4_lut (.I0(n64395), .I1(n28043), .I2(\byte_transmit_counter[2] ), 
            .I3(\byte_transmit_counter[0] ), .O(n64396));
    defparam i48702_4_lut.LUT_INIT = 16'haca0;
    SB_LUT4 i48700_3_lut (.I0(\data_out_frame[4] [7]), .I1(\data_out_frame[5] [7]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n64394));
    defparam i48700_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_adj_1246 (.I0(\data_out_frame[20] [3]), .I1(\data_out_frame[20] [1]), 
            .I2(\data_out_frame[20] [2]), .I3(\data_out_frame[20] [5]), 
            .O(n59223));
    defparam i1_2_lut_4_lut_adj_1246.LUT_INIT = 16'h6996;
    SB_LUT4 select_775_Select_53_i2_4_lut (.I0(\data_out_frame[6] [5]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder0_position_scaled[21]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4935));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_53_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_775_Select_67_i2_4_lut (.I0(\data_out_frame[8] [3]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder0_position_scaled[3]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4733));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_67_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFF current_limit_i0_i7 (.Q(current_limit[7]), .C(clk16MHz), .D(n29637));   // verilog/coms.v(130[12] 305[6])
    SB_DFF control_mode_i0_i4 (.Q(control_mode[4]), .C(clk16MHz), .D(n29636));   // verilog/coms.v(130[12] 305[6])
    SB_DFF control_mode_i0_i3 (.Q(control_mode[3]), .C(clk16MHz), .D(n29635));   // verilog/coms.v(130[12] 305[6])
    SB_DFF control_mode_i0_i2 (.Q(control_mode[2]), .C(clk16MHz), .D(n29634));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_775_Select_52_i2_4_lut (.I0(\data_out_frame[6] [4]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder0_position_scaled[20]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4936));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_52_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFF control_mode_i0_i1 (.Q(control_mode[1]), .C(clk16MHz), .D(n29633));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i23 (.Q(neopxl_color[23]), .C(clk16MHz), .D(n29632));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i22 (.Q(neopxl_color[22]), .C(clk16MHz), .D(n29631));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i48853_3_lut (.I0(\data_out_frame[8] [7]), .I1(\data_out_frame[9] [7]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n64547));
    defparam i48853_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF neopxl_color_i0_i21 (.Q(neopxl_color[21]), .C(clk16MHz), .D(n29630));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i48854_3_lut (.I0(\data_out_frame[10] [7]), .I1(\data_out_frame[11] [7]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n64548));
    defparam i48854_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF neopxl_color_i0_i20 (.Q(neopxl_color[20]), .C(clk16MHz), .D(n29629));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_775_Select_51_i2_4_lut (.I0(\data_out_frame[6] [3]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder0_position_scaled[19]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4937));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_51_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFF neopxl_color_i0_i19 (.Q(neopxl_color[19]), .C(clk16MHz), .D(n29627));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i18 (.Q(neopxl_color[18]), .C(clk16MHz), .D(n29626));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i17 (.Q(neopxl_color[17]), .C(clk16MHz), .D(n29625));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i16 (.Q(neopxl_color[16]), .C(clk16MHz), .D(n29624));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i15 (.Q(neopxl_color[15]), .C(clk16MHz), .D(n29623));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i16086_3_lut_4_lut (.I0(n58731), .I1(n58752), .I2(rx_data[3]), 
            .I3(\data_in_frame[13] [3]), .O(n30092));
    defparam i16086_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 select_775_Select_50_i2_4_lut (.I0(\data_out_frame[6] [2]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder0_position_scaled[18]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4938));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_50_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i48860_3_lut (.I0(\data_out_frame[14] [7]), .I1(\data_out_frame[15] [7]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n64554));
    defparam i48860_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48859_3_lut (.I0(\data_out_frame[12] [7]), .I1(\data_out_frame[13] [7]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n64553));
    defparam i48859_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51563_2_lut (.I0(n70967), .I1(\byte_transmit_counter[2] ), 
            .I2(GND_net), .I3(GND_net), .O(n66934));
    defparam i51563_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 select_775_Select_49_i2_4_lut (.I0(\data_out_frame[6] [1]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder0_position_scaled[17]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4939));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_49_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFFESS data_out_frame_0___i156 (.Q(\data_out_frame[19] [3]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4940), .S(n58521));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_775_Select_48_i2_4_lut (.I0(\data_out_frame[6] [0]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder0_position_scaled[16]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4941));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_48_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i48835_3_lut (.I0(\data_out_frame[16] [7]), .I1(\data_out_frame[17] [7]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n64529));
    defparam i48835_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48836_3_lut (.I0(\data_out_frame[18] [7]), .I1(\data_out_frame[19] [7]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n64530));
    defparam i48836_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48743_3_lut (.I0(\data_out_frame[22] [7]), .I1(\data_out_frame[23] [7]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n64437));
    defparam i48743_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 select_775_Select_47_i2_4_lut (.I0(\data_out_frame[5] [7]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(control_mode[7]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4942));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_47_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_775_Select_46_i2_4_lut (.I0(\data_out_frame[5] [6]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(control_mode[6]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4943));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_46_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i48742_3_lut (.I0(\data_out_frame[20] [7]), .I1(\data_out_frame[21] [7]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n64436));
    defparam i48742_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 select_775_Select_45_i2_4_lut (.I0(\data_out_frame[5] [5]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(control_mode[5]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4944));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_45_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i48725_3_lut (.I0(\data_out_frame[6] [0]), .I1(\data_out_frame[7] [0]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n64419));
    defparam i48725_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48726_4_lut (.I0(n64419), .I1(n28104), .I2(\byte_transmit_counter[2] ), 
            .I3(\data_out_frame[1][0] ), .O(n64420));
    defparam i48726_4_lut.LUT_INIT = 16'ha3a0;
    SB_LUT4 i48724_3_lut (.I0(\data_out_frame[4] [0]), .I1(\data_out_frame[5] [0]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n64418));
    defparam i48724_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 select_775_Select_44_i2_4_lut (.I0(\data_out_frame[5] [4]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(control_mode[4]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4945));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_44_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i16083_3_lut_4_lut (.I0(n58731), .I1(n58752), .I2(rx_data[2]), 
            .I3(\data_in_frame[13] [2]), .O(n30089));
    defparam i16083_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 select_775_Select_43_i2_4_lut (.I0(\data_out_frame[5] [3]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(control_mode[3]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4946));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_43_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFFESS data_out_frame_0___i157 (.Q(\data_out_frame[19] [4]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4947), .S(n58522));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i158 (.Q(\data_out_frame[19] [5]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4948), .S(n58523));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i2 (.Q(neopxl_color[2]), .C(clk16MHz), .D(n29621));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i16079_3_lut_4_lut (.I0(n58731), .I1(n58752), .I2(rx_data[1]), 
            .I3(\data_in_frame[13] [1]), .O(n30085));
    defparam i16079_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i52408_2_lut (.I0(n70973), .I1(\byte_transmit_counter[2] ), 
            .I2(GND_net), .I3(GND_net), .O(n67162));
    defparam i52408_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i53427_3_lut (.I0(n71225), .I1(n70991), .I2(\byte_transmit_counter[2] ), 
            .I3(GND_net), .O(n69121));
    defparam i53427_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53428_4_lut (.I0(n69121), .I1(n70907), .I2(byte_transmit_counter[3]), 
            .I3(\byte_transmit_counter[2] ), .O(n69122));
    defparam i53428_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i53511_3_lut (.I0(n70883), .I1(n71219), .I2(\byte_transmit_counter[2] ), 
            .I3(GND_net), .O(n69205));
    defparam i53511_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48678_3_lut (.I0(n70925), .I1(n69122), .I2(byte_transmit_counter[4]), 
            .I3(GND_net), .O(tx_data[3]));
    defparam i48678_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16076_3_lut_4_lut (.I0(n58731), .I1(n58752), .I2(rx_data[0]), 
            .I3(\data_in_frame[13] [0]), .O(n30082));
    defparam i16076_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_4_lut_adj_1247 (.I0(\FRAME_MATCHER.i_31__N_2514 ), .I1(n1951), 
            .I2(n60750), .I3(n4452), .O(n8_adj_4949));   // verilog/coms.v(118[11:12])
    defparam i1_4_lut_adj_1247.LUT_INIT = 16'ha0a2;
    SB_LUT4 i1_4_lut_adj_1248 (.I0(n8_adj_4949), .I1(n1951), .I2(n22687), 
            .I3(n63955), .O(n26967));   // verilog/coms.v(118[11:12])
    defparam i1_4_lut_adj_1248.LUT_INIT = 16'hbbba;
    SB_LUT4 i456_2_lut (.I0(n3303), .I1(\FRAME_MATCHER.i_31__N_2512 ), .I2(GND_net), 
            .I3(GND_net), .O(n2060));   // verilog/coms.v(148[4] 304[11])
    defparam i456_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_3_lut_4_lut (.I0(\data_out_frame[20] [3]), .I1(n23652), 
            .I2(n60844), .I3(\data_out_frame[20] [4]), .O(n53928));
    defparam i1_2_lut_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i48298_4_lut (.I0(n1951), .I1(n1954), .I2(n3303), .I3(n1957), 
            .O(n63978));   // verilog/coms.v(139[4] 141[7])
    defparam i48298_4_lut.LUT_INIT = 16'h0a02;
    SB_LUT4 i1_4_lut_adj_1249 (.I0(\FRAME_MATCHER.i_31__N_2512 ), .I1(n1954), 
            .I2(n63978), .I3(n61412), .O(n57728));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1249.LUT_INIT = 16'hb3a0;
    SB_LUT4 i6672_4_lut (.I0(n1955), .I1(\FRAME_MATCHER.state[3] ), .I2(n1957), 
            .I3(n25463), .O(n20350));   // verilog/coms.v(148[4] 304[11])
    defparam i6672_4_lut.LUT_INIT = 16'heccc;
    SB_LUT4 i445_2_lut (.I0(\FRAME_MATCHER.state_31__N_2612 [3]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(GND_net), .I3(GND_net), .O(n2049));   // verilog/coms.v(148[4] 304[11])
    defparam i445_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i444_2_lut (.I0(n771), .I1(\FRAME_MATCHER.i_31__N_2508 ), .I2(GND_net), 
            .I3(GND_net), .O(n2048));   // verilog/coms.v(148[4] 304[11])
    defparam i444_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i15498_3_lut_4_lut (.I0(n8_adj_4950), .I1(n58720), .I2(rx_data[7]), 
            .I3(\data_in_frame[19] [7]), .O(n29504));
    defparam i15498_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_adj_1250 (.I0(\FRAME_MATCHER.i[0] ), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [1]), .I3(GND_net), .O(n6_adj_4951));   // verilog/coms.v(118[11:12])
    defparam i2_3_lut_adj_1250.LUT_INIT = 16'hecec;
    SB_LUT4 i15495_3_lut_4_lut (.I0(n8_adj_4950), .I1(n58720), .I2(rx_data[6]), 
            .I3(\data_in_frame[19] [6]), .O(n29501));
    defparam i15495_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i29138_4_lut (.I0(n25388), .I1(\FRAME_MATCHER.i [31]), .I2(n6_adj_4951), 
            .I3(\FRAME_MATCHER.i[3] ), .O(n771));   // verilog/coms.v(160[9:60])
    defparam i29138_4_lut.LUT_INIT = 16'h3332;
    SB_LUT4 i1_2_lut_adj_1251 (.I0(\FRAME_MATCHER.i[4] ), .I1(n25474), .I2(GND_net), 
            .I3(GND_net), .O(n25388));   // verilog/coms.v(157[7:23])
    defparam i1_2_lut_adj_1251.LUT_INIT = 16'heeee;
    SB_LUT4 i29147_4_lut (.I0(n25388), .I1(\FRAME_MATCHER.i [31]), .I2(n8_adj_12), 
            .I3(\FRAME_MATCHER.i[3] ), .O(n3303));   // verilog/coms.v(230[9:54])
    defparam i29147_4_lut.LUT_INIT = 16'h3222;
    SB_LUT4 i2_2_lut_adj_1252 (.I0(n3303), .I1(\FRAME_MATCHER.i_31__N_2512 ), 
            .I2(GND_net), .I3(GND_net), .O(n22687));   // verilog/coms.v(148[4] 304[11])
    defparam i2_2_lut_adj_1252.LUT_INIT = 16'h4444;
    SB_LUT4 i3_2_lut (.I0(n25463), .I1(\FRAME_MATCHER.i_31__N_2507 ), .I2(GND_net), 
            .I3(GND_net), .O(n27541));   // verilog/coms.v(148[4] 304[11])
    defparam i3_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i2_4_lut_adj_1253 (.I0(n4452), .I1(n27541), .I2(\FRAME_MATCHER.i_31__N_2514 ), 
            .I3(n22687), .O(n60982));   // verilog/coms.v(148[4] 304[11])
    defparam i2_4_lut_adj_1253.LUT_INIT = 16'hffdc;
    SB_LUT4 i1_4_lut_adj_1254 (.I0(n25468), .I1(n1957), .I2(n1955), .I3(n60982), 
            .O(n26964));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1254.LUT_INIT = 16'hbaaa;
    SB_DFF current_limit_i0_i8 (.Q(current_limit[8]), .C(clk16MHz), .D(n29618));   // verilog/coms.v(130[12] 305[6])
    SB_DFF current_limit_i0_i9 (.Q(current_limit[9]), .C(clk16MHz), .D(n29617));   // verilog/coms.v(130[12] 305[6])
    SB_DFF current_limit_i0_i10 (.Q(current_limit[10]), .C(clk16MHz), .D(n29616));   // verilog/coms.v(130[12] 305[6])
    SB_DFF current_limit_i0_i11 (.Q(current_limit[11]), .C(clk16MHz), .D(n29615));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i3 (.Q(neopxl_color[3]), .C(clk16MHz), .D(n29613));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i4 (.Q(neopxl_color[4]), .C(clk16MHz), .D(n29612));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i5 (.Q(neopxl_color[5]), .C(clk16MHz), .D(n29608));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i6 (.Q(neopxl_color[6]), .C(clk16MHz), .D(n29607));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i7 (.Q(neopxl_color[7]), .C(clk16MHz), .D(n29606));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i8 (.Q(neopxl_color[8]), .C(clk16MHz), .D(n29605));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i9 (.Q(neopxl_color[9]), .C(clk16MHz), .D(n29604));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i10 (.Q(neopxl_color[10]), .C(clk16MHz), .D(n29582));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i7_4_lut_adj_1255 (.I0(\data_in[2] [6]), .I1(\data_in[1] [2]), 
            .I2(n25538), .I3(\data_in[3] [2]), .O(n18_adj_4953));
    defparam i7_4_lut_adj_1255.LUT_INIT = 16'hfffd;
    SB_DFF current_limit_i0_i12 (.Q(current_limit[12]), .C(clk16MHz), .D(n29574));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i1 (.Q(\data_in[0] [0]), .C(clk16MHz), .D(n29569));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i9_4_lut_adj_1256 (.I0(\data_in[1] [6]), .I1(n18_adj_4953), 
            .I2(\data_in[1] [3]), .I3(\data_in[2] [0]), .O(n20_c));
    defparam i9_4_lut_adj_1256.LUT_INIT = 16'hfffd;
    SB_DFFR PWMLimit_i0_i0 (.Q(PWMLimit[0]), .C(clk16MHz), .D(n29559), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFF current_limit_i0_i0 (.Q(current_limit[0]), .C(clk16MHz), .D(n29558));   // verilog/coms.v(130[12] 305[6])
    SB_DFF control_mode_i0_i0 (.Q(control_mode[0]), .C(clk16MHz), .D(n29557));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i0 (.Q(neopxl_color[0]), .C(clk16MHz), .D(n29556));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Ki_i0 (.Q(\Ki[0] ), .C(clk16MHz), .D(n29555), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Kp_i0 (.Q(\Kp[0] ), .C(clk16MHz), .D(n29554), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i15492_3_lut_4_lut (.I0(n8_adj_4950), .I1(n58720), .I2(rx_data[5]), 
            .I3(\data_in_frame[19] [5]), .O(n29498));
    defparam i15492_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFFR IntegralLimit_i0_i0 (.Q(IntegralLimit[0]), .C(clk16MHz), .D(n29534), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i4_2_lut_adj_1257 (.I0(\data_in[2] [5]), .I1(\data_in[0] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_4954));
    defparam i4_2_lut_adj_1257.LUT_INIT = 16'heeee;
    SB_DFFESS data_out_frame_0___i159 (.Q(\data_out_frame[19] [6]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4955), .S(n28921));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i10_4_lut_adj_1258 (.I0(n15_adj_4954), .I1(n20_c), .I2(\data_in[0] [5]), 
            .I3(\data_in[3] [7]), .O(n25380));
    defparam i10_4_lut_adj_1258.LUT_INIT = 16'hfeff;
    SB_LUT4 i4_4_lut_adj_1259 (.I0(\data_in[1] [7]), .I1(\data_in[0] [0]), 
            .I2(\data_in[1] [1]), .I3(\data_in[0] [4]), .O(n10_adj_4956));
    defparam i4_4_lut_adj_1259.LUT_INIT = 16'hfdff;
    SB_LUT4 i5_3_lut_adj_1260 (.I0(\data_in[3] [4]), .I1(n10_adj_4956), 
            .I2(\data_in[2] [7]), .I3(GND_net), .O(n25538));
    defparam i5_3_lut_adj_1260.LUT_INIT = 16'hdfdf;
    SB_LUT4 i48501_4_lut (.I0(\data_in[1] [5]), .I1(\data_in[0] [3]), .I2(\data_in[2] [2]), 
            .I3(\data_in[1] [0]), .O(n64186));
    defparam i48501_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i1_2_lut_adj_1261 (.I0(\data_in[2] [4]), .I1(\data_in[1] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n9));
    defparam i1_2_lut_adj_1261.LUT_INIT = 16'heeee;
    SB_LUT4 i7_4_lut_adj_1262 (.I0(n9), .I1(n64186), .I2(\data_in[3] [0]), 
            .I3(\data_in[0] [6]), .O(n25493));
    defparam i7_4_lut_adj_1262.LUT_INIT = 16'hffbf;
    SB_DFFESS data_out_frame_0___i160 (.Q(\data_out_frame[19] [7]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4957), .S(n58524));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i161 (.Q(\data_out_frame[20] [0]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4958), .S(n58525));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i162 (.Q(\data_out_frame[20] [1]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4959), .S(n58526));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i163 (.Q(\data_out_frame[20] [2]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4960), .S(n58527));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i164 (.Q(\data_out_frame[20] [3]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4961), .S(n58528));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i165 (.Q(\data_out_frame[20] [4]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4962), .S(n58529));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i166 (.Q(\data_out_frame[20] [5]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4963), .S(n58530));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i167 (.Q(\data_out_frame[20] [6]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4964), .S(n58531));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i168 (.Q(\data_out_frame[20] [7]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4965), .S(n58532));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i169 (.Q(\data_out_frame[21] [0]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4966), .S(n58533));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i170 (.Q(\data_out_frame[21] [1]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4967), .S(n58534));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i171 (.Q(\data_out_frame[21] [2]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4968), .S(n58535));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i172 (.Q(\data_out_frame[21] [3]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4969), .S(n58536));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i173 (.Q(\data_out_frame[21] [4]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4970), .S(n58492));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i174 (.Q(\data_out_frame[21] [5]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4971), .S(n58537));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i175 (.Q(\data_out_frame[21] [6]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4972), .S(n58538));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i176 (.Q(\data_out_frame[21] [7]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4973), .S(n58539));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i177 (.Q(\data_out_frame[22] [0]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4974), .S(n28903));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i178 (.Q(\data_out_frame[22] [1]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4975), .S(n58540));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i15489_3_lut_4_lut (.I0(n8_adj_4950), .I1(n58720), .I2(rx_data[4]), 
            .I3(\data_in_frame[19] [4]), .O(n29495));
    defparam i15489_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFFESS data_out_frame_0___i179 (.Q(\data_out_frame[22] [2]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4976), .S(n58541));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i180 (.Q(\data_out_frame[22] [3]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4977), .S(n58494));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i181 (.Q(\data_out_frame[22] [4]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4978), .S(n58542));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i182 (.Q(\data_out_frame[22] [5]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4979), .S(n58543));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i183 (.Q(\data_out_frame[22] [6]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4980), .S(n58544));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i2_2_lut_adj_1263 (.I0(\data_in[2] [3]), .I1(\data_in[3] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n10_adj_4981));
    defparam i2_2_lut_adj_1263.LUT_INIT = 16'heeee;
    SB_LUT4 i6_4_lut_adj_1264 (.I0(\data_in[0] [2]), .I1(\data_in[3] [3]), 
            .I2(\data_in[3] [1]), .I3(\data_in[0] [7]), .O(n14_adj_4982));
    defparam i6_4_lut_adj_1264.LUT_INIT = 16'hfeff;
    SB_LUT4 i7_4_lut_adj_1265 (.I0(\data_in[3] [6]), .I1(n14_adj_4982), 
            .I2(n10_adj_4981), .I3(\data_in[2] [1]), .O(n25487));
    defparam i7_4_lut_adj_1265.LUT_INIT = 16'hfffd;
    SB_LUT4 i3_2_lut_adj_1266 (.I0(\data_in[1] [3]), .I1(\data_in[1] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n16_adj_4983));
    defparam i3_2_lut_adj_1266.LUT_INIT = 16'hdddd;
    SB_LUT4 i9_4_lut_adj_1267 (.I0(\data_in[3] [7]), .I1(n25487), .I2(\data_in[2] [6]), 
            .I3(\data_in[0] [5]), .O(n22_adj_4984));
    defparam i9_4_lut_adj_1267.LUT_INIT = 16'hfeff;
    SB_LUT4 i15486_3_lut_4_lut (.I0(n8_adj_4950), .I1(n58720), .I2(rx_data[3]), 
            .I3(\data_in_frame[19] [3]), .O(n29492));
    defparam i15486_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i7_3_lut (.I0(\data_in[2] [5]), .I1(\data_in[1] [2]), .I2(n25493), 
            .I3(GND_net), .O(n20_adj_4985));
    defparam i7_3_lut.LUT_INIT = 16'hf7f7;
    SB_LUT4 i15483_3_lut_4_lut (.I0(n8_adj_4950), .I1(n58720), .I2(rx_data[2]), 
            .I3(\data_in_frame[19] [2]), .O(n29489));
    defparam i15483_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11_4_lut_adj_1268 (.I0(n25538), .I1(n22_adj_4984), .I2(n16_adj_4983), 
            .I3(\data_in[0] [1]), .O(n24_adj_4986));
    defparam i11_4_lut_adj_1268.LUT_INIT = 16'hfeff;
    SB_LUT4 i12_4_lut_adj_1269 (.I0(\data_in[2] [0]), .I1(n24_adj_4986), 
            .I2(n20_adj_4985), .I3(\data_in[3] [2]), .O(n1951));
    defparam i12_4_lut_adj_1269.LUT_INIT = 16'hfdff;
    SB_LUT4 i6_4_lut_adj_1270 (.I0(\data_in[2] [2]), .I1(\data_in[1] [0]), 
            .I2(n25487), .I3(\data_in[1] [5]), .O(n16_adj_4987));
    defparam i6_4_lut_adj_1270.LUT_INIT = 16'hfffe;
    SB_LUT4 select_775_Select_120_i2_4_lut (.I0(\data_out_frame[15] [0]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[16]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4862));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_120_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i7_4_lut_adj_1271 (.I0(\data_in[2] [4]), .I1(\data_in[3] [0]), 
            .I2(\data_in[0] [3]), .I3(n25380), .O(n17_adj_4988));
    defparam i7_4_lut_adj_1271.LUT_INIT = 16'hfffd;
    SB_LUT4 i9_4_lut_adj_1272 (.I0(n17_adj_4988), .I1(\data_in[0] [6]), 
            .I2(n16_adj_4987), .I3(\data_in[1] [4]), .O(n1954));
    defparam i9_4_lut_adj_1272.LUT_INIT = 16'hfbff;
    SB_LUT4 i6_4_lut_adj_1273 (.I0(\data_in[3] [6]), .I1(n25493), .I2(\data_in[2] [1]), 
            .I3(n25380), .O(n16_adj_4989));
    defparam i6_4_lut_adj_1273.LUT_INIT = 16'hffef;
    SB_LUT4 i7_4_lut_adj_1274 (.I0(\data_in[0] [7]), .I1(\data_in[2] [3]), 
            .I2(\data_in[0] [2]), .I3(\data_in[3] [1]), .O(n17_adj_4990));
    defparam i7_4_lut_adj_1274.LUT_INIT = 16'hbfff;
    SB_LUT4 i9_4_lut_adj_1275 (.I0(n17_adj_4990), .I1(\data_in[3] [5]), 
            .I2(n16_adj_4989), .I3(\data_in[3] [3]), .O(n1957));
    defparam i9_4_lut_adj_1275.LUT_INIT = 16'hfbff;
    SB_LUT4 select_775_Select_119_i2_4_lut (.I0(\data_out_frame[14] [7]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[7]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4861));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_119_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i362_2_lut (.I0(n1954), .I1(n1951), .I2(GND_net), .I3(GND_net), 
            .O(n1955));   // verilog/coms.v(142[4] 144[7])
    defparam i362_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_775_Select_118_i2_4_lut (.I0(\data_out_frame[14] [6]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[6]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4860));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_118_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFFR \FRAME_MATCHER.i_1938__i0  (.Q(\FRAME_MATCHER.i[0] ), .C(clk16MHz), 
            .D(n27978), .R(reset));   // verilog/coms.v(158[12:15])
    SB_LUT4 select_775_Select_117_i2_4_lut (.I0(\data_out_frame[14] [5]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[5]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4858));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_117_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_adj_1276 (.I0(Kp_23__N_1748), .I1(\FRAME_MATCHER.i_31__N_2513 ), 
            .I2(GND_net), .I3(GND_net), .O(n33690));   // verilog/coms.v(148[4] 304[11])
    defparam i1_2_lut_adj_1276.LUT_INIT = 16'heeee;
    SB_LUT4 i15480_3_lut_4_lut (.I0(n8_adj_4950), .I1(n58720), .I2(rx_data[1]), 
            .I3(\data_in_frame[19] [1]), .O(n29486));
    defparam i15480_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 equal_310_i10_2_lut_3_lut (.I0(\FRAME_MATCHER.i[3] ), .I1(\FRAME_MATCHER.i[4] ), 
            .I2(\FRAME_MATCHER.i[5] ), .I3(GND_net), .O(n10_adj_4991));   // verilog/coms.v(157[7:23])
    defparam equal_310_i10_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 select_775_Select_116_i2_4_lut (.I0(\data_out_frame[14] [4]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[4]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4857));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_116_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_1648_Select_0_i1_2_lut_3_lut_4_lut (.I0(tx_active), .I1(r_SM_Main_2__N_3545[0]), 
            .I2(n43563), .I3(\FRAME_MATCHER.i_31__N_2511 ), .O(n1_adj_4992));   // verilog/coms.v(148[4] 304[11])
    defparam select_1648_Select_0_i1_2_lut_3_lut_4_lut.LUT_INIT = 16'h0100;
    SB_LUT4 i2_4_lut_adj_1277 (.I0(n43563), .I1(n61225), .I2(\FRAME_MATCHER.i_31__N_2511 ), 
            .I3(n42843), .O(n6_adj_4993));   // verilog/coms.v(118[11:12])
    defparam i2_4_lut_adj_1277.LUT_INIT = 16'hccec;
    SB_DFFESS data_out_frame_0___i184 (.Q(\data_out_frame[22] [7]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4994), .S(n58545));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i3_4_lut_adj_1278 (.I0(n33690), .I1(n6_adj_4993), .I2(\FRAME_MATCHER.i_31__N_2509 ), 
            .I3(\FRAME_MATCHER.state_31__N_2612 [3]), .O(n71283));   // verilog/coms.v(118[11:12])
    defparam i3_4_lut_adj_1278.LUT_INIT = 16'heefe;
    SB_LUT4 select_775_Select_115_i2_4_lut (.I0(\data_out_frame[14] [3]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[3]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4856));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_115_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFFESS data_out_frame_0___i185 (.Q(\data_out_frame[23] [0]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4995), .S(n28895));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i15477_3_lut_4_lut (.I0(n8_adj_4950), .I1(n58720), .I2(rx_data[0]), 
            .I3(\data_in_frame[19] [0]), .O(n29483));
    defparam i15477_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1279 (.I0(\data_out_frame[15] [4]), .I1(n25650), 
            .I2(n26210), .I3(n59189), .O(n6_adj_4771));
    defparam i1_2_lut_3_lut_4_lut_adj_1279.LUT_INIT = 16'h6996;
    SB_LUT4 i14824_2_lut_2_lut (.I0(reset), .I1(\FRAME_MATCHER.i_31__N_2508 ), 
            .I2(GND_net), .I3(GND_net), .O(n28830));   // verilog/coms.v(130[12] 305[6])
    defparam i14824_2_lut_2_lut.LUT_INIT = 16'h4444;
    SB_DFFESS data_out_frame_0___i186 (.Q(\data_out_frame[23] [1]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4996), .S(n28894));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i187 (.Q(\data_out_frame[23] [2]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4997), .S(n58546));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_775_Select_114_i2_4_lut (.I0(\data_out_frame[14] [2]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[2]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4855));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_114_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i51556_2_lut (.I0(\data_out_frame[0][4] ), .I1(\byte_transmit_counter[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n67065));
    defparam i51556_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1280 (.I0(\data_out_frame[15] [4]), .I1(n25650), 
            .I2(n26210), .I3(n59089), .O(n53735));
    defparam i1_2_lut_3_lut_4_lut_adj_1280.LUT_INIT = 16'h6996;
    SB_LUT4 select_775_Select_42_i2_4_lut (.I0(\data_out_frame[5] [2]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(control_mode[2]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4998));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_42_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_3_lut_3_lut (.I0(Kp_23__N_1748), .I1(n37), .I2(reset), 
            .I3(GND_net), .O(n22734));   // verilog/coms.v(148[4] 304[11])
    defparam i1_2_lut_3_lut_3_lut.LUT_INIT = 16'h0808;
    SB_LUT4 i51655_2_lut (.I0(\data_out_frame[3][4] ), .I1(\byte_transmit_counter[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n67066));
    defparam i51655_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_775_Select_113_i2_4_lut (.I0(\data_out_frame[14] [1]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[1]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4852));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_113_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFFR \FRAME_MATCHER.i_1938__i31  (.Q(\FRAME_MATCHER.i [31]), .C(clk16MHz), 
            .D(n27980), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_1938__i30  (.Q(\FRAME_MATCHER.i [30]), .C(clk16MHz), 
            .D(n27982), .R(reset));   // verilog/coms.v(158[12:15])
    SB_LUT4 select_775_Select_41_i2_4_lut (.I0(\data_out_frame[5] [1]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(control_mode[1]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4999));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_41_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1281 (.I0(\data_out_frame[16] [6]), .I1(\data_out_frame[16] [4]), 
            .I2(n59010), .I3(\data_out_frame[15] [7]), .O(n8_adj_4797));
    defparam i1_2_lut_3_lut_4_lut_adj_1281.LUT_INIT = 16'h9669;
    SB_LUT4 i1_4_lut_adj_1282 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[14] [0]), 
            .I2(setpoint[0]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4851));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1282.LUT_INIT = 16'ha088;
    SB_DFFR \FRAME_MATCHER.i_1938__i29  (.Q(\FRAME_MATCHER.i [29]), .C(clk16MHz), 
            .D(n27984), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_1938__i28  (.Q(\FRAME_MATCHER.i [28]), .C(clk16MHz), 
            .D(n27986), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_1938__i27  (.Q(\FRAME_MATCHER.i [27]), .C(clk16MHz), 
            .D(n27988), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_1938__i26  (.Q(\FRAME_MATCHER.i [26]), .C(clk16MHz), 
            .D(n27990), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_1938__i25  (.Q(\FRAME_MATCHER.i [25]), .C(clk16MHz), 
            .D(n27992), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_1938__i24  (.Q(\FRAME_MATCHER.i [24]), .C(clk16MHz), 
            .D(n27994), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_1938__i23  (.Q(\FRAME_MATCHER.i [23]), .C(clk16MHz), 
            .D(n27996), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_1938__i22  (.Q(\FRAME_MATCHER.i [22]), .C(clk16MHz), 
            .D(n27998), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_1938__i21  (.Q(\FRAME_MATCHER.i [21]), .C(clk16MHz), 
            .D(n28000), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_1938__i20  (.Q(\FRAME_MATCHER.i [20]), .C(clk16MHz), 
            .D(n28002), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_1938__i19  (.Q(\FRAME_MATCHER.i [19]), .C(clk16MHz), 
            .D(n28004), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_1938__i18  (.Q(\FRAME_MATCHER.i [18]), .C(clk16MHz), 
            .D(n28006), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_1938__i17  (.Q(\FRAME_MATCHER.i [17]), .C(clk16MHz), 
            .D(n28008), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_1938__i16  (.Q(\FRAME_MATCHER.i [16]), .C(clk16MHz), 
            .D(n28010), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_1938__i15  (.Q(\FRAME_MATCHER.i [15]), .C(clk16MHz), 
            .D(n28012), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_1938__i14  (.Q(\FRAME_MATCHER.i [14]), .C(clk16MHz), 
            .D(n28014), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_1938__i13  (.Q(\FRAME_MATCHER.i [13]), .C(clk16MHz), 
            .D(n28016), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_1938__i12  (.Q(\FRAME_MATCHER.i [12]), .C(clk16MHz), 
            .D(n28018), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_1938__i11  (.Q(\FRAME_MATCHER.i [11]), .C(clk16MHz), 
            .D(n28020), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_1938__i10  (.Q(\FRAME_MATCHER.i [10]), .C(clk16MHz), 
            .D(n28022), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_1938__i9  (.Q(\FRAME_MATCHER.i [9]), .C(clk16MHz), 
            .D(n28024), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_1938__i8  (.Q(\FRAME_MATCHER.i [8]), .C(clk16MHz), 
            .D(n28026), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_1938__i7  (.Q(\FRAME_MATCHER.i [7]), .C(clk16MHz), 
            .D(n28028), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_1938__i6  (.Q(\FRAME_MATCHER.i [6]), .C(clk16MHz), 
            .D(n28030), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_1938__i5  (.Q(\FRAME_MATCHER.i[5] ), .C(clk16MHz), 
            .D(n28032), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_1938__i4  (.Q(\FRAME_MATCHER.i[4] ), .C(clk16MHz), 
            .D(n28034), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_1938__i3  (.Q(\FRAME_MATCHER.i[3] ), .C(clk16MHz), 
            .D(n28036), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_1938__i2  (.Q(\FRAME_MATCHER.i [2]), .C(clk16MHz), 
            .D(n28038), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_1938__i1  (.Q(\FRAME_MATCHER.i [1]), .C(clk16MHz), 
            .D(n28040), .R(reset));   // verilog/coms.v(158[12:15])
    SB_LUT4 select_775_Select_40_i2_4_lut (.I0(\data_out_frame[5] [0]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(control_mode[0]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5000));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_40_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_775_Select_39_i2_4_lut (.I0(\data_out_frame[4] [7]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(ID[7]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), .O(n2_adj_5001));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_39_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_775_Select_38_i2_4_lut (.I0(\data_out_frame[4] [6]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(ID[6]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), .O(n2_adj_5002));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_38_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i4_2_lut_3_lut_4_lut (.I0(\data_out_frame[16] [6]), .I1(\data_out_frame[16] [4]), 
            .I2(n59010), .I3(\data_out_frame[19] [4]), .O(n18_adj_4787));
    defparam i4_2_lut_3_lut_4_lut.LUT_INIT = 16'h9669;
    SB_LUT4 select_775_Select_37_i2_4_lut (.I0(\data_out_frame[4] [5]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(ID[5]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), .O(n2_adj_5003));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_37_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_775_Select_36_i2_4_lut (.I0(\data_out_frame[4] [4]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(ID[4]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), .O(n2_adj_5004));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_36_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_775_Select_35_i2_4_lut (.I0(\data_out_frame[4] [3]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(ID[3]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), .O(n2_adj_5005));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_35_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_775_Select_34_i2_4_lut (.I0(\data_out_frame[4] [2]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(ID[2]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), .O(n2_adj_5006));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_34_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_775_Select_111_i2_4_lut (.I0(\data_out_frame[13] [7]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[15]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4848));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_111_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_775_Select_110_i2_4_lut (.I0(\data_out_frame[13] [6]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[14]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4847));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_110_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_775_Select_109_i2_4_lut (.I0(\data_out_frame[13] [5]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[13]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4846));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_109_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_775_Select_33_i2_4_lut (.I0(\data_out_frame[4] [1]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(ID[1]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), .O(n2_adj_5007));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_33_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_775_Select_108_i2_4_lut (.I0(\data_out_frame[13] [4]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[12]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4845));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_108_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1283 (.I0(\data_in_frame[13] [3]), .I1(\data_in_frame[13] [4]), 
            .I2(n53570), .I3(n25906), .O(n54511));   // verilog/coms.v(88[17:63])
    defparam i1_2_lut_3_lut_4_lut_adj_1283.LUT_INIT = 16'h9669;
    SB_DFFESS data_out_frame_0___i3 (.Q(\data_out_frame[0][2] ), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5008), .S(n58670));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i4 (.Q(\data_out_frame[0][3] ), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5009), .S(n58669));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i5 (.Q(\data_out_frame[0][4] ), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5010), .S(n58668));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i9 (.Q(\data_out_frame[1][0] ), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5011), .S(n58667));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1284 (.I0(reset), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[26] [0]), 
            .O(n58467));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1284.LUT_INIT = 16'h5100;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1285 (.I0(\data_in_frame[0]_c [5]), .I1(\data_in_frame[2] [7]), 
            .I2(n35423), .I3(n59299), .O(n6_adj_5012));
    defparam i1_2_lut_3_lut_4_lut_adj_1285.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1286 (.I0(\data_in_frame[0]_c [5]), .I1(\data_in_frame[2] [7]), 
            .I2(n35423), .I3(\data_in_frame[5] [3]), .O(n59003));
    defparam i1_2_lut_3_lut_4_lut_adj_1286.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1287 (.I0(reset), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[26] [1]), 
            .O(n58472));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1287.LUT_INIT = 16'h5100;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1288 (.I0(reset), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[26][2] ), 
            .O(n58473));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1288.LUT_INIT = 16'h5100;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1289 (.I0(reset), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[26] [3]), 
            .O(n58470));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1289.LUT_INIT = 16'h5100;
    SB_DFF current_limit_i0_i13 (.Q(current_limit[13]), .C(clk16MHz), .D(n30439));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1290 (.I0(reset), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[26] [4]), 
            .O(n58474));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1290.LUT_INIT = 16'h5100;
    SB_LUT4 i51913_2_lut_3_lut_4_lut (.I0(\FRAME_MATCHER.i[3] ), .I1(\FRAME_MATCHER.i[4] ), 
            .I2(\FRAME_MATCHER.i[5] ), .I3(n132), .O(n67115));   // verilog/coms.v(94[13:20])
    defparam i51913_2_lut_3_lut_4_lut.LUT_INIT = 16'h0100;
    SB_DFF current_limit_i0_i14 (.Q(current_limit[14]), .C(clk16MHz), .D(n30438));   // verilog/coms.v(130[12] 305[6])
    SB_DFF current_limit_i0_i15 (.Q(current_limit[15]), .C(clk16MHz), .D(n30437));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i1 (.Q(PWMLimit[1]), .C(clk16MHz), .D(n30436), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFS PWMLimit_i0_i2 (.Q(PWMLimit[2]), .C(clk16MHz), .D(n30435), 
            .S(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i3 (.Q(PWMLimit[3]), .C(clk16MHz), .D(n30434), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i117 (.Q(\data_in_frame[14] [4]), .C(clk16MHz), 
           .D(n29369));   // verilog/coms.v(130[12] 305[6])
    SB_DFFS PWMLimit_i0_i4 (.Q(PWMLimit[4]), .C(clk16MHz), .D(n30432), 
            .S(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFS PWMLimit_i0_i5 (.Q(PWMLimit[5]), .C(clk16MHz), .D(n30428), 
            .S(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFS PWMLimit_i0_i6 (.Q(PWMLimit[6]), .C(clk16MHz), .D(n30427), 
            .S(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i118 (.Q(\data_in_frame[14] [5]), .C(clk16MHz), 
           .D(n29372));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i1 (.Q(\data_in_frame[0][0] ), .C(clk16MHz), 
            .E(VCC_net), .D(n30421));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i119 (.Q(\data_in_frame[14] [6]), .C(clk16MHz), 
           .D(n29375));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i120 (.Q(\data_in_frame[14] [7]), .C(clk16MHz), 
           .D(n29378));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i121 (.Q(\data_in_frame[15] [0]), .C(clk16MHz), 
           .D(n22_adj_5013));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i122 (.Q(\data_in_frame[15] [1]), .C(clk16MHz), 
           .D(n29384));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i123 (.Q(\data_in_frame[15] [2]), .C(clk16MHz), 
           .D(n29387));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i124 (.Q(\data_in_frame[15] [3]), .C(clk16MHz), 
           .D(n29390));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i116 (.Q(\data_in_frame[14] [3]), .C(clk16MHz), 
            .E(VCC_net), .D(n30396));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i125 (.Q(\data_in_frame[15] [4]), .C(clk16MHz), 
           .D(n29393));   // verilog/coms.v(130[12] 305[6])
    SB_DFFS PWMLimit_i0_i7 (.Q(PWMLimit[7]), .C(clk16MHz), .D(n30394), 
            .S(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFS PWMLimit_i0_i8 (.Q(PWMLimit[8]), .C(clk16MHz), .D(n30393), 
            .S(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i126 (.Q(\data_in_frame[15] [5]), .C(clk16MHz), 
           .D(n29396));   // verilog/coms.v(130[12] 305[6])
    SB_DFF control_mode_i0_i5 (.Q(control_mode[5]), .C(clk16MHz), .D(n30391));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i9 (.Q(PWMLimit[9]), .C(clk16MHz), .D(n30390), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i10 (.Q(PWMLimit[10]), .C(clk16MHz), .D(n30389), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i11 (.Q(PWMLimit[11]), .C(clk16MHz), .D(n30388), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i127 (.Q(\data_in_frame[15] [6]), .C(clk16MHz), 
           .D(n29399));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i12 (.Q(PWMLimit[12]), .C(clk16MHz), .D(n30373), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i13 (.Q(PWMLimit[13]), .C(clk16MHz), .D(n30349), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i14 (.Q(PWMLimit[14]), .C(clk16MHz), .D(n30322), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i15 (.Q(PWMLimit[15]), .C(clk16MHz), .D(n30321), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i16 (.Q(PWMLimit[16]), .C(clk16MHz), .D(n30320), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i17 (.Q(PWMLimit[17]), .C(clk16MHz), .D(n30314), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i2 (.Q(\data_in[0] [1]), .C(clk16MHz), .D(n30307));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i3 (.Q(\data_in[0] [2]), .C(clk16MHz), .D(n30306));   // verilog/coms.v(130[12] 305[6])
    SB_DFF control_mode_i0_i6 (.Q(control_mode[6]), .C(clk16MHz), .D(n30305));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i4 (.Q(\data_in[0] [3]), .C(clk16MHz), .D(n30304));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i5 (.Q(\data_in[0] [4]), .C(clk16MHz), .D(n30303));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i6 (.Q(\data_in[0] [5]), .C(clk16MHz), .D(n30302));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i7 (.Q(\data_in[0] [6]), .C(clk16MHz), .D(n30301));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i8 (.Q(\data_in[0] [7]), .C(clk16MHz), .D(n30300));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i9 (.Q(\data_in[1] [0]), .C(clk16MHz), .D(n30299));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i10 (.Q(\data_in[1] [1]), .C(clk16MHz), .D(n30298));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i11 (.Q(\data_in[1] [2]), .C(clk16MHz), .D(n30297));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i12 (.Q(\data_in[1] [3]), .C(clk16MHz), .D(n30296));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i13 (.Q(\data_in[1] [4]), .C(clk16MHz), .D(n30295));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i14 (.Q(\data_in[1] [5]), .C(clk16MHz), .D(n30294));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i15 (.Q(\data_in[1] [6]), .C(clk16MHz), .D(n30293));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i16 (.Q(\data_in[1] [7]), .C(clk16MHz), .D(n30292));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i17 (.Q(\data_in[2] [0]), .C(clk16MHz), .D(n30291));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i18 (.Q(\data_in[2] [1]), .C(clk16MHz), .D(n30290));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i19 (.Q(\data_in[2] [2]), .C(clk16MHz), .D(n30289));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i20 (.Q(\data_in[2] [3]), .C(clk16MHz), .D(n30288));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i21 (.Q(\data_in[2] [4]), .C(clk16MHz), .D(n30287));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i22 (.Q(\data_in[2] [5]), .C(clk16MHz), .D(n30286));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i23 (.Q(\data_in[2] [6]), .C(clk16MHz), .D(n30285));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i24 (.Q(\data_in[2] [7]), .C(clk16MHz), .D(n30284));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i25 (.Q(\data_in[3] [0]), .C(clk16MHz), .D(n30283));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i26 (.Q(\data_in[3] [1]), .C(clk16MHz), .D(n30282));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i27 (.Q(\data_in[3] [2]), .C(clk16MHz), .D(n30281));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i28 (.Q(\data_in[3] [3]), .C(clk16MHz), .D(n30280));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i29 (.Q(\data_in[3] [4]), .C(clk16MHz), .D(n30279));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i30 (.Q(\data_in[3] [5]), .C(clk16MHz), .D(n30278));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i31 (.Q(\data_in[3] [6]), .C(clk16MHz), .D(n30277));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i32 (.Q(\data_in[3] [7]), .C(clk16MHz), .D(n30276));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i18 (.Q(PWMLimit[18]), .C(clk16MHz), .D(n30275), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i19 (.Q(PWMLimit[19]), .C(clk16MHz), .D(n30274), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFF control_mode_i0_i7 (.Q(control_mode[7]), .C(clk16MHz), .D(n30273));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i128 (.Q(\data_in_frame[15] [7]), .C(clk16MHz), 
           .D(n29407));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i20 (.Q(PWMLimit[20]), .C(clk16MHz), .D(n30271), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i47 (.Q(\data_in_frame[5] [6]), .C(clk16MHz), 
           .D(n29898));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i48 (.Q(\data_in_frame[5] [7]), .C(clk16MHz), 
           .D(n29901));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i21 (.Q(PWMLimit[21]), .C(clk16MHz), .D(n30268), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i115 (.Q(\data_in_frame[14] [2]), .C(clk16MHz), 
            .E(VCC_net), .D(n30265));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i22 (.Q(PWMLimit[22]), .C(clk16MHz), .D(n30264), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i129 (.Q(\data_in_frame[16] [0]), .C(clk16MHz), 
           .D(n57890));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i49 (.Q(\data_in_frame[6] [0]), .C(clk16MHz), 
           .D(n29904));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i50 (.Q(\data_in_frame[6] [1]), .C(clk16MHz), 
           .D(n29908));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i23 (.Q(PWMLimit[23]), .C(clk16MHz), .D(n30260), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i114 (.Q(\data_in_frame[14] [1]), .C(clk16MHz), 
            .E(VCC_net), .D(n30257));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i130 (.Q(\data_in_frame[16] [1]), .C(clk16MHz), 
           .D(n57886));   // verilog/coms.v(130[12] 305[6])
    SB_DFF current_limit_i0_i1 (.Q(current_limit[1]), .C(clk16MHz), .D(n30255));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i131 (.Q(\data_in_frame[16] [2]), .C(clk16MHz), 
           .D(n29417));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i132 (.Q(\data_in_frame[16] [3]), .C(clk16MHz), 
           .D(n29420));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i133 (.Q(\data_in_frame[16] [4]), .C(clk16MHz), 
           .D(n29423));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i134 (.Q(\data_in_frame[16] [5]), .C(clk16MHz), 
           .D(n29426));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i135 (.Q(\data_in_frame[16] [6]), .C(clk16MHz), 
           .D(n57882));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i136 (.Q(\data_in_frame[16] [7]), .C(clk16MHz), 
           .D(n29432));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i137 (.Q(\data_in_frame[17] [0]), .C(clk16MHz), 
           .D(n57878));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i138 (.Q(\data_in_frame[17] [1]), .C(clk16MHz), 
           .D(n57876));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i139 (.Q(\data_in_frame[17] [2]), .C(clk16MHz), 
           .D(n57874));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i140 (.Q(\data_in_frame[17] [3]), .C(clk16MHz), 
           .D(n57872));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i141 (.Q(\data_in_frame[17] [4]), .C(clk16MHz), 
           .D(n57868));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i142 (.Q(\data_in_frame[17] [5]), .C(clk16MHz), 
           .D(n57864));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i143 (.Q(\data_in_frame[17] [6]), .C(clk16MHz), 
           .D(n57860));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i51 (.Q(\data_in_frame[6] [2]), .C(clk16MHz), 
           .D(n29911));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i52 (.Q(\data_in_frame[6] [3]), .C(clk16MHz), 
           .D(n29914));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i53 (.Q(\data_in_frame[6] [4]), .C(clk16MHz), 
           .D(n29918));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i113 (.Q(\data_in_frame[14] [0]), .C(clk16MHz), 
            .E(VCC_net), .D(n30227));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i144 (.Q(\data_in_frame[17] [7]), .C(clk16MHz), 
           .D(n57856));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i145 (.Q(\data_in_frame[18] [0]), .C(clk16MHz), 
           .D(n57852));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i146 (.Q(\data_in_frame[18] [1]), .C(clk16MHz), 
           .D(n57850));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i54 (.Q(\data_in_frame[6] [5]), .C(clk16MHz), 
           .D(n29921));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i55 (.Q(\data_in_frame[6] [6]), .C(clk16MHz), 
           .D(n29924));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i56 (.Q(\data_in_frame[6] [7]), .C(clk16MHz), 
           .D(n29927));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i57 (.Q(\data_in_frame[7] [0]), .C(clk16MHz), 
           .D(n29930));   // verilog/coms.v(130[12] 305[6])
    SB_DFF current_limit_i0_i2 (.Q(current_limit[2]), .C(clk16MHz), .D(n30218));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i58 (.Q(\data_in_frame[7] [1]), .C(clk16MHz), 
           .D(n29934));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i59 (.Q(\data_in_frame[7] [2]), .C(clk16MHz), 
           .D(n29937));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i60 (.Q(\data_in_frame[7] [3]), .C(clk16MHz), 
           .D(n29940));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i10 (.Q(\data_out_frame[1][1] ), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5014), .S(n58666));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i61 (.Q(\data_in_frame[7] [4]), .C(clk16MHz), 
           .D(n29943));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i62 (.Q(\data_in_frame[7] [5]), .C(clk16MHz), 
           .D(n29946));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i63 (.Q(\data_in_frame[7]_c [6]), .C(clk16MHz), 
           .D(n58092));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i147 (.Q(\data_in_frame[18] [2]), .C(clk16MHz), 
           .D(n57846));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i64 (.Q(\data_in_frame[7]_c [7]), .C(clk16MHz), 
           .D(n58086));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i65 (.Q(\data_in_frame[8] [0]), .C(clk16MHz), 
           .D(n29955));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i66 (.Q(\data_in_frame[8] [1]), .C(clk16MHz), 
           .D(n29958));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i67 (.Q(\data_in_frame[8] [2]), .C(clk16MHz), 
           .D(n29961));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i68 (.Q(\data_in_frame[8] [3]), .C(clk16MHz), 
           .D(n29964));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i69 (.Q(\data_in_frame[8] [4]), .C(clk16MHz), 
           .D(n30205));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i70 (.Q(\data_in_frame[8] [5]), .C(clk16MHz), 
           .D(n29970));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i71 (.Q(\data_in_frame[8] [6]), .C(clk16MHz), 
           .D(n29973));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i72 (.Q(\data_in_frame[8] [7]), .C(clk16MHz), 
           .D(n29976));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i73 (.Q(\data_in_frame[9] [0]), .C(clk16MHz), 
           .D(n29979));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i74 (.Q(\data_in_frame[9] [1]), .C(clk16MHz), 
           .D(n29982));   // verilog/coms.v(130[12] 305[6])
    SB_DFF current_limit_i0_i3 (.Q(current_limit[3]), .C(clk16MHz), .D(n30199));   // verilog/coms.v(130[12] 305[6])
    SB_DFF current_limit_i0_i4 (.Q(current_limit[4]), .C(clk16MHz), .D(n30198));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i75 (.Q(\data_in_frame[9] [2]), .C(clk16MHz), 
           .D(n29985));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i76 (.Q(\data_in_frame[9] [3]), .C(clk16MHz), 
           .D(n29989));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i77 (.Q(\data_in_frame[9] [4]), .C(clk16MHz), 
           .D(n29992));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i78 (.Q(\data_in_frame[9] [5]), .C(clk16MHz), 
           .D(n29995));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i79 (.Q(\data_in_frame[9] [6]), .C(clk16MHz), 
           .D(n29998));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i80 (.Q(\data_in_frame[9] [7]), .C(clk16MHz), 
           .D(n30001));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i81 (.Q(\data_in_frame[10] [0]), .C(clk16MHz), 
           .D(n30004));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_775_Select_107_i2_4_lut (.I0(\data_out_frame[13] [3]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[11]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4841));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_107_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFF data_in_frame_0___i82 (.Q(\data_in_frame[10] [1]), .C(clk16MHz), 
           .D(n30007));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i83 (.Q(\data_in_frame[10] [2]), .C(clk16MHz), 
           .D(n30010));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i84 (.Q(\data_in_frame[10] [3]), .C(clk16MHz), 
           .D(n30013));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i85 (.Q(\data_in_frame[10] [4]), .C(clk16MHz), 
           .D(n30017));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i86 (.Q(\data_in_frame[10] [5]), .C(clk16MHz), 
           .D(n30020));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i87 (.Q(\data_in_frame[10] [6]), .C(clk16MHz), 
           .D(n30023));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i88 (.Q(\data_in_frame[10] [7]), .C(clk16MHz), 
           .D(n30027));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i89 (.Q(\data_in_frame[11] [0]), .C(clk16MHz), 
           .D(n30030));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i12 (.Q(\data_out_frame[1][3] ), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5015), .S(n58665));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i90 (.Q(\data_in_frame[11] [1]), .C(clk16MHz), 
           .D(n58106));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i91 (.Q(\data_in_frame[11] [2]), .C(clk16MHz), 
           .D(n58108));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i92 (.Q(\data_in_frame[11] [3]), .C(clk16MHz), 
           .D(n58060));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i93 (.Q(\data_in_frame[11] [4]), .C(clk16MHz), 
           .D(n30043));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i94 (.Q(\data_in_frame[11] [5]), .C(clk16MHz), 
           .D(n30046));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i95 (.Q(\data_in_frame[11] [6]), .C(clk16MHz), 
           .D(n30049));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i96 (.Q(\data_in_frame[11] [7]), .C(clk16MHz), 
           .D(n30053));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i97 (.Q(\data_in_frame[12] [0]), .C(clk16MHz), 
           .D(n30056));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i98 (.Q(\data_in_frame[12] [1]), .C(clk16MHz), 
           .D(n30059));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i99 (.Q(\data_in_frame[12] [2]), .C(clk16MHz), 
           .D(n30062));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i100 (.Q(\data_in_frame[12] [3]), .C(clk16MHz), 
           .D(n57932));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i101 (.Q(\data_in_frame[12] [4]), .C(clk16MHz), 
           .D(n57936));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i102 (.Q(\data_in_frame[12] [5]), .C(clk16MHz), 
           .D(n30072));   // verilog/coms.v(130[12] 305[6])
    SB_DFF current_limit_i0_i5 (.Q(current_limit[5]), .C(clk16MHz), .D(n30169));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i103 (.Q(\data_in_frame[12] [6]), .C(clk16MHz), 
           .D(n30075));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i104 (.Q(\data_in_frame[12] [7]), .C(clk16MHz), 
           .D(n30079));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i105 (.Q(\data_in_frame[13] [0]), .C(clk16MHz), 
           .D(n30082));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i106 (.Q(\data_in_frame[13] [1]), .C(clk16MHz), 
           .D(n30085));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i107 (.Q(\data_in_frame[13] [2]), .C(clk16MHz), 
           .D(n30089));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i108 (.Q(\data_in_frame[13] [3]), .C(clk16MHz), 
           .D(n30092));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i109 (.Q(\data_in_frame[13] [4]), .C(clk16MHz), 
           .D(n30095));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i110 (.Q(\data_in_frame[13] [5]), .C(clk16MHz), 
           .D(n30099));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i111 (.Q(\data_in_frame[13] [6]), .C(clk16MHz), 
           .D(n30102));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i191 (.Q(\data_in_frame[23] [6]), .C(clk16MHz), 
           .D(n57996));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i192 (.Q(\data_in_frame[23] [7]), .C(clk16MHz), 
           .D(n30110));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i112 (.Q(\data_in_frame[13] [7]), .C(clk16MHz), 
           .D(n30145));   // verilog/coms.v(130[12] 305[6])
    SB_DFF current_limit_i0_i6 (.Q(current_limit[6]), .C(clk16MHz), .D(n30154));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i148 (.Q(\data_in_frame[18] [3]), .C(clk16MHz), 
           .D(n29468));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i14 (.Q(\data_out_frame[1][5] ), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5016), .S(n58664));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i149 (.Q(\data_in_frame[18] [4]), .C(clk16MHz), 
           .D(n57842));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i150 (.Q(\data_in_frame[18] [5]), .C(clk16MHz), 
           .D(n29474));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i151 (.Q(\data_in_frame[18] [6]), .C(clk16MHz), 
           .D(n57838));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i152 (.Q(\data_in_frame[18] [7]), .C(clk16MHz), 
           .D(n57834));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i153 (.Q(\data_in_frame[19] [0]), .C(clk16MHz), 
           .D(n29483));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i154 (.Q(\data_in_frame[19] [1]), .C(clk16MHz), 
           .D(n29486));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i155 (.Q(\data_in_frame[19] [2]), .C(clk16MHz), 
           .D(n29489));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i15 (.Q(\data_out_frame[1][6] ), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5017), .S(n58663));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i156 (.Q(\data_in_frame[19] [3]), .C(clk16MHz), 
           .D(n29492));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i157 (.Q(\data_in_frame[19] [4]), .C(clk16MHz), 
           .D(n29495));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i158 (.Q(\data_in_frame[19] [5]), .C(clk16MHz), 
           .D(n29498));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i159 (.Q(\data_in_frame[19] [6]), .C(clk16MHz), 
           .D(n29501));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i160 (.Q(\data_in_frame[19] [7]), .C(clk16MHz), 
           .D(n29504));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i161 (.Q(\data_in_frame[20] [0]), .C(clk16MHz), 
           .D(n57986));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i162 (.Q(\data_in_frame[20] [1]), .C(clk16MHz), 
           .D(n30106));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i163 (.Q(\data_in_frame[20] [2]), .C(clk16MHz), 
           .D(n57980));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i164 (.Q(\data_in_frame[20] [3]), .C(clk16MHz), 
           .D(n30098));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_55402 (.I0(byte_transmit_counter[3]), 
            .I1(n71039), .I2(n67165), .I3(byte_transmit_counter[4]), .O(n71042));
    defparam byte_transmit_counter_3__bdd_4_lut_55402.LUT_INIT = 16'he4aa;
    SB_DFF data_in_frame_0___i165 (.Q(\data_in_frame[20] [4]), .C(clk16MHz), 
           .D(n29520));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_adj_1291 (.I0(byte_transmit_counter[6]), .I1(byte_transmit_counter[5]), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_5018));   // verilog/coms.v(217[11:56])
    defparam i1_2_lut_adj_1291.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_1292 (.I0(byte_transmit_counter[4]), .I1(\byte_transmit_counter[0] ), 
            .I2(\byte_transmit_counter[2] ), .I3(\byte_transmit_counter[1] ), 
            .O(n4_adj_5019));
    defparam i1_4_lut_adj_1292.LUT_INIT = 16'ha8a0;
    SB_DFF data_in_frame_0___i166 (.Q(\data_in_frame[20] [5]), .C(clk16MHz), 
           .D(n29523));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1293 (.I0(reset), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[26] [5]), 
            .O(n58468));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1293.LUT_INIT = 16'h5100;
    SB_DFF data_in_frame_0___i167 (.Q(\data_in_frame[20] [6]), .C(clk16MHz), 
           .D(n57974));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i2_3_lut_4_lut (.I0(\data_out_frame[20] [3]), .I1(n23652), .I2(n54525), 
            .I3(\data_out_frame[20] [1]), .O(n61136));
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1294 (.I0(reset), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[26] [6]), 
            .O(n58475));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1294.LUT_INIT = 16'h5100;
    SB_DFF data_in_frame_0___i168 (.Q(\data_in_frame[20] [7]), .C(clk16MHz), 
           .D(n58000));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i29667_4_lut (.I0(byte_transmit_counter[3]), .I1(byte_transmit_counter[7]), 
            .I2(n4_adj_5019), .I3(n4_adj_5018), .O(n43563));
    defparam i29667_4_lut.LUT_INIT = 16'hffec;
    SB_LUT4 i28951_2_lut (.I0(tx_active), .I1(r_SM_Main_2__N_3545[0]), .I2(GND_net), 
            .I3(GND_net), .O(n42843));
    defparam i28951_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1295 (.I0(reset), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[26] [7]), 
            .O(n58476));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1295.LUT_INIT = 16'h5100;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1296 (.I0(reset), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[27] [0]), 
            .O(n58477));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1296.LUT_INIT = 16'h5100;
    SB_DFF data_in_frame_0___i169 (.Q(\data_in_frame[21] [0]), .C(clk16MHz), 
           .D(n29535));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i170 (.Q(\data_in_frame[21] [1]), .C(clk16MHz), 
           .D(n29539));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1297 (.I0(reset), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[27] [1]), 
            .O(n58478));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1297.LUT_INIT = 16'h5100;
    SB_DFF data_in_frame_0___i171 (.Q(\data_in_frame[21] [2]), .C(clk16MHz), 
           .D(n29542));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i172 (.Q(\data_in_frame[21] [3]), .C(clk16MHz), 
           .D(n29551));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1298 (.I0(reset), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[27][2] ), 
            .O(n58479));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1298.LUT_INIT = 16'h5100;
    SB_DFF data_in_frame_0___i173 (.Q(\data_in_frame[21] [4]), .C(clk16MHz), 
           .D(n29570));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_4_lut_adj_1299 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[4] [0]), 
            .I2(ID[0]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), .O(n2_adj_5020));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1299.LUT_INIT = 16'ha088;
    SB_LUT4 select_775_Select_106_i2_4_lut (.I0(\data_out_frame[13] [2]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[10]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4840));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_106_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i51768_2_lut (.I0(n70913), .I1(\byte_transmit_counter[2] ), 
            .I2(GND_net), .I3(GND_net), .O(n67141));
    defparam i51768_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1300 (.I0(reset), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[27] [3]), 
            .O(n58471));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1300.LUT_INIT = 16'h5100;
    SB_LUT4 select_775_Select_105_i2_4_lut (.I0(\data_out_frame[13] [1]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[9]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4839));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_105_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i53421_3_lut (.I0(n71189), .I1(n70931), .I2(\byte_transmit_counter[2] ), 
            .I3(GND_net), .O(n69115));
    defparam i53421_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFESS data_out_frame_0___i16 (.Q(\data_out_frame[1][7] ), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5021), .S(n58662));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i48772_3_lut (.I0(\data_out_frame[16] [2]), .I1(\data_out_frame[17] [2]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n64466));
    defparam i48772_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1301 (.I0(reset), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[27] [4]), 
            .O(n58480));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1301.LUT_INIT = 16'h5100;
    SB_LUT4 i48773_3_lut (.I0(\data_out_frame[18] [2]), .I1(\data_out_frame[19] [2]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n64467));
    defparam i48773_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1302 (.I0(reset), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[27] [5]), 
            .O(n58469));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1302.LUT_INIT = 16'h5100;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1303 (.I0(reset), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[27] [6]), 
            .O(n58481));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1303.LUT_INIT = 16'h5100;
    SB_LUT4 i48800_3_lut (.I0(\data_out_frame[22] [2]), .I1(\data_out_frame[23] [2]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n64494));
    defparam i48800_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48799_3_lut (.I0(\data_out_frame[20] [2]), .I1(\data_out_frame[21] [2]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n64493));
    defparam i48799_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51548_2_lut (.I0(\byte_transmit_counter[0] ), .I1(\data_out_frame[0][2] ), 
            .I2(GND_net), .I3(GND_net), .O(n67049));
    defparam i51548_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i48719_3_lut (.I0(\data_out_frame[6] [2]), .I1(\data_out_frame[7] [2]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n64413));
    defparam i48719_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1304 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[13] [0]), 
            .I2(setpoint[8]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4838));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1304.LUT_INIT = 16'ha088;
    SB_DFFESS data_out_frame_0___i26 (.Q(\data_out_frame[3][1] ), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5022), .S(n58661));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i28 (.Q(\data_out_frame[3][3] ), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5023), .S(n58660));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i29 (.Q(\data_out_frame[3][4] ), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5024), .S(n58659));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i48720_4_lut (.I0(n64413), .I1(n67049), .I2(\byte_transmit_counter[2] ), 
            .I3(\byte_transmit_counter[1] ), .O(n64414));
    defparam i48720_4_lut.LUT_INIT = 16'ha0ac;
    SB_DFFESS data_out_frame_0___i31 (.Q(\data_out_frame[3][6] ), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5025), .S(n58658));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i48718_3_lut (.I0(\data_out_frame[4] [2]), .I1(\data_out_frame[5] [2]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n64412));
    defparam i48718_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1305 (.I0(reset), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[27] [7]), 
            .O(n58482));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1305.LUT_INIT = 16'h5100;
    SB_DFF data_in_frame_0___i174 (.Q(\data_in_frame[21] [5]), .C(clk16MHz), 
           .D(n29575));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i32 (.Q(\data_out_frame[3][7] ), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5026), .S(n58657));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i30065112_i1_3_lut (.I0(n70871), .I1(n70859), .I2(\byte_transmit_counter[2] ), 
            .I3(GND_net), .O(n14_adj_5027));
    defparam i30065112_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n71042_bdd_4_lut (.I0(n71042), .I1(n14_adj_5027), .I2(n7_adj_5028), 
            .I3(byte_transmit_counter[4]), .O(tx_data[2]));
    defparam n71042_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 select_775_Select_31_i2_3_lut (.I0(\data_out_frame[3][7] ), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\FRAME_MATCHER.state_31__N_2612 [3]), .I3(GND_net), .O(n2_adj_5026));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_31_i2_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_55342 (.I0(\byte_transmit_counter[1] ), 
            .I1(n64493), .I2(n64494), .I3(\byte_transmit_counter[2] ), 
            .O(n71036));
    defparam byte_transmit_counter_1__bdd_4_lut_55342.LUT_INIT = 16'he4aa;
    SB_LUT4 n71036_bdd_4_lut (.I0(n71036), .I1(n64467), .I2(n64466), .I3(\byte_transmit_counter[2] ), 
            .O(n71039));
    defparam n71036_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_55313 (.I0(byte_transmit_counter[3]), 
            .I1(n69115), .I2(n67141), .I3(byte_transmit_counter[4]), .O(n71030));
    defparam byte_transmit_counter_3__bdd_4_lut_55313.LUT_INIT = 16'he4aa;
    SB_DFFESS data_out_frame_0___i33 (.Q(\data_out_frame[4] [0]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5020), .S(n58506));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i23 (.Q(setpoint[23]), .C(clk16MHz), .E(n27674), 
            .D(n4760[23]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i22 (.Q(setpoint[22]), .C(clk16MHz), .E(n27674), 
            .D(n4760[22]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i21 (.Q(setpoint[21]), .C(clk16MHz), .E(n27674), 
            .D(n4760[21]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i20 (.Q(setpoint[20]), .C(clk16MHz), .E(n27674), 
            .D(n4760[20]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i19 (.Q(setpoint[19]), .C(clk16MHz), .E(n27674), 
            .D(n4760[19]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i18 (.Q(setpoint[18]), .C(clk16MHz), .E(n27674), 
            .D(n4760[18]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i17 (.Q(setpoint[17]), .C(clk16MHz), .E(n27674), 
            .D(n4760[17]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i16 (.Q(setpoint[16]), .C(clk16MHz), .E(n27674), 
            .D(n4760[16]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i15 (.Q(setpoint[15]), .C(clk16MHz), .E(n27674), 
            .D(n4760[15]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i14 (.Q(setpoint[14]), .C(clk16MHz), .E(n27674), 
            .D(n4760[14]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i13 (.Q(setpoint[13]), .C(clk16MHz), .E(n27674), 
            .D(n4760[13]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i12 (.Q(setpoint[12]), .C(clk16MHz), .E(n27674), 
            .D(n4760[12]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i11 (.Q(setpoint[11]), .C(clk16MHz), .E(n27674), 
            .D(n4760[11]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i10 (.Q(setpoint[10]), .C(clk16MHz), .E(n27674), 
            .D(n4760[10]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i9 (.Q(setpoint[9]), .C(clk16MHz), .E(n27674), 
            .D(n4760[9]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i8 (.Q(setpoint[8]), .C(clk16MHz), .E(n27674), 
            .D(n4760[8]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i7 (.Q(setpoint[7]), .C(clk16MHz), .E(n27674), 
            .D(n4760[7]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i6 (.Q(setpoint[6]), .C(clk16MHz), .E(n27674), 
            .D(n4760[6]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i5 (.Q(setpoint[5]), .C(clk16MHz), .E(n27674), 
            .D(n4760[5]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i4 (.Q(setpoint[4]), .C(clk16MHz), .E(n27674), 
            .D(n4760[4]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i3 (.Q(setpoint[3]), .C(clk16MHz), .E(n27674), 
            .D(n4760[3]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i2 (.Q(setpoint[2]), .C(clk16MHz), .E(n27674), 
            .D(n4760[2]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i1 (.Q(setpoint[1]), .C(clk16MHz), .E(n27674), 
            .D(n4760[1]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i34 (.Q(\data_out_frame[4] [1]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5007), .S(n58656));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i35 (.Q(\data_out_frame[4] [2]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5006), .S(n58655));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i36 (.Q(\data_out_frame[4] [3]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5005), .S(n58654));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i37 (.Q(\data_out_frame[4] [4]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5004), .S(n58653));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i38 (.Q(\data_out_frame[4] [5]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5003), .S(n58652));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i39 (.Q(\data_out_frame[4] [6]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5002), .S(n58651));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i40 (.Q(\data_out_frame[4] [7]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5001), .S(n58650));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i41 (.Q(\data_out_frame[5] [0]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5000), .S(n58649));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i42 (.Q(\data_out_frame[5] [1]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4999), .S(n58648));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i43 (.Q(\data_out_frame[5] [2]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4998), .S(n58647));   // verilog/coms.v(130[12] 305[6])
    SB_DFFS \FRAME_MATCHER.state_FSM_i9  (.Q(\FRAME_MATCHER.i_31__N_2507 ), 
            .C(clk16MHz), .D(n71283), .S(reset));   // verilog/coms.v(148[4] 304[11])
    SB_DFFR \FRAME_MATCHER.state_FSM_i8  (.Q(\FRAME_MATCHER.i_31__N_2508 ), 
            .C(clk16MHz), .D(n26964), .R(reset));   // verilog/coms.v(148[4] 304[11])
    SB_DFFR \FRAME_MATCHER.state_FSM_i7  (.Q(\FRAME_MATCHER.i_31__N_2509 ), 
            .C(clk16MHz), .D(n2048), .R(reset));   // verilog/coms.v(148[4] 304[11])
    SB_DFFR \FRAME_MATCHER.state_FSM_i6  (.Q(\FRAME_MATCHER.state[3] ), .C(clk16MHz), 
            .D(n2049), .R(reset));   // verilog/coms.v(148[4] 304[11])
    SB_DFFR \FRAME_MATCHER.state_FSM_i5  (.Q(\FRAME_MATCHER.i_31__N_2511 ), 
            .C(clk16MHz), .D(n20350), .R(reset));   // verilog/coms.v(148[4] 304[11])
    SB_DFFR \FRAME_MATCHER.state_FSM_i4  (.Q(\FRAME_MATCHER.i_31__N_2512 ), 
            .C(clk16MHz), .D(n57728), .R(reset));   // verilog/coms.v(148[4] 304[11])
    SB_DFFR \FRAME_MATCHER.state_FSM_i3  (.Q(\FRAME_MATCHER.i_31__N_2513 ), 
            .C(clk16MHz), .D(n2060), .R(reset));   // verilog/coms.v(148[4] 304[11])
    SB_DFFR \FRAME_MATCHER.state_FSM_i2  (.Q(\FRAME_MATCHER.i_31__N_2514 ), 
            .C(clk16MHz), .D(n26967), .R(reset));   // verilog/coms.v(148[4] 304[11])
    SB_DFF data_in_frame_0___i175 (.Q(\data_in_frame[21] [6]), .C(clk16MHz), 
           .D(n29578));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i44 (.Q(\data_out_frame[5] [3]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4946), .S(n58646));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i45 (.Q(\data_out_frame[5] [4]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4945), .S(n58645));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i46 (.Q(\data_out_frame[5] [5]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4944), .S(n58644));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i47 (.Q(\data_out_frame[5] [6]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4943), .S(n58643));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i48 (.Q(\data_out_frame[5] [7]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4942), .S(n58642));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i49 (.Q(\data_out_frame[6] [0]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4941), .S(n58641));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i50 (.Q(\data_out_frame[6] [1]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4939), .S(n58640));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_775_Select_30_i2_3_lut (.I0(\data_out_frame[3][6] ), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\FRAME_MATCHER.state_31__N_2612 [3]), .I3(GND_net), .O(n2_adj_5025));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_30_i2_3_lut.LUT_INIT = 16'hc8c8;
    SB_DFFESS data_out_frame_0___i51 (.Q(\data_out_frame[6] [2]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4938), .S(n58639));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_775_Select_28_i2_3_lut (.I0(\data_out_frame[3][4] ), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\FRAME_MATCHER.state_31__N_2612 [3]), .I3(GND_net), .O(n2_adj_5024));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_28_i2_3_lut.LUT_INIT = 16'hc8c8;
    SB_DFFESS data_out_frame_0___i52 (.Q(\data_out_frame[6] [3]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4937), .S(n58638));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i53 (.Q(\data_out_frame[6] [4]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4936), .S(n58637));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i54 (.Q(\data_out_frame[6] [5]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4935), .S(n58636));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_775_Select_103_i2_4_lut (.I0(\data_out_frame[12] [7]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[23]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4837));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_103_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_775_Select_102_i2_4_lut (.I0(\data_out_frame[12] [6]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[22]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4836));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_102_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFFESS data_out_frame_0___i55 (.Q(\data_out_frame[6] [6]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4934), .S(n58635));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i56 (.Q(\data_out_frame[6] [7]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4933), .S(n58634));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i57 (.Q(\data_out_frame[7] [0]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4932), .S(n58633));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i58 (.Q(\data_out_frame[7] [1]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4931), .S(n58632));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i11 (.Q(neopxl_color[11]), .C(clk16MHz), .D(n29410));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_775_Select_27_i2_3_lut (.I0(\data_out_frame[3][3] ), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\FRAME_MATCHER.state_31__N_2612 [3]), .I3(GND_net), .O(n2_adj_5023));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_27_i2_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 select_775_Select_101_i2_4_lut (.I0(\data_out_frame[12] [5]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[21]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4835));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_101_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_775_Select_100_i2_4_lut (.I0(\data_out_frame[12] [4]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[20]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4834));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_100_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_775_Select_99_i2_4_lut (.I0(\data_out_frame[12] [3]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(setpoint[19]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4833));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_99_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i2_3_lut_4_lut_adj_1306 (.I0(\data_out_frame[20] [4]), .I1(n60844), 
            .I2(\data_out_frame[20] [5]), .I3(n61261), .O(n59332));
    defparam i2_3_lut_4_lut_adj_1306.LUT_INIT = 16'h9669;
    SB_LUT4 select_775_Select_25_i2_3_lut (.I0(\data_out_frame[3][1] ), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\FRAME_MATCHER.state_31__N_2612 [3]), .I3(GND_net), .O(n2_adj_5022));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_25_i2_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 select_775_Select_98_i2_4_lut (.I0(\data_out_frame[12] [2]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(setpoint[18]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4832));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_98_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_775_Select_15_i2_3_lut (.I0(\data_out_frame[1][7] ), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\FRAME_MATCHER.state_31__N_2612 [3]), .I3(GND_net), .O(n2_adj_5021));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_15_i2_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 select_775_Select_97_i2_4_lut (.I0(\data_out_frame[12] [1]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(setpoint[17]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4831));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_97_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_775_Select_96_i2_4_lut (.I0(\data_out_frame[12] [0]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(setpoint[16]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4830));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_96_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_775_Select_95_i2_4_lut (.I0(\data_out_frame[11] [7]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[7]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4829));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_95_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1307 (.I0(\FRAME_MATCHER.i[3] ), .I1(n9_adj_5029), 
            .I2(n43501), .I3(n8_adj_4950), .O(n28337));
    defparam i1_2_lut_3_lut_4_lut_adj_1307.LUT_INIT = 16'hffef;
    SB_LUT4 i1_4_lut_adj_1308 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[11] [6]), 
            .I2(encoder1_position_scaled[6]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4828));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1308.LUT_INIT = 16'ha088;
    SB_LUT4 select_775_Select_93_i2_4_lut (.I0(\data_out_frame[11] [5]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[5]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4827));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_93_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_775_Select_92_i2_4_lut (.I0(\data_out_frame[11] [4]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[4]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4826));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_92_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_775_Select_91_i2_4_lut (.I0(\data_out_frame[11] [3]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[3]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4825));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_91_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_775_Select_90_i2_4_lut (.I0(\data_out_frame[11] [2]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[2]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4824));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_90_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_775_Select_89_i2_4_lut (.I0(\data_out_frame[11] [1]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[1]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4823));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_89_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i13_4_lut_adj_1309 (.I0(n40663), .I1(\data_in_frame[20] [7]), 
            .I2(n160), .I3(rx_data[7]), .O(n58000));   // verilog/coms.v(94[13:20])
    defparam i13_4_lut_adj_1309.LUT_INIT = 16'hc5c0;
    SB_DFFR deadband_i0_i0 (.Q(deadband[0]), .C(clk16MHz), .D(n29406), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i188 (.Q(\data_out_frame[23] [3]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4928), .S(n58547));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i12 (.Q(neopxl_color[12]), .C(clk16MHz), .D(n29405));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i13 (.Q(neopxl_color[13]), .C(clk16MHz), .D(n29403));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i52424_2_lut (.I0(n70997), .I1(\byte_transmit_counter[2] ), 
            .I2(GND_net), .I3(GND_net), .O(n67165));
    defparam i52424_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i26765_4_lut (.I0(n159), .I1(n92), .I2(rx_data[3]), .I3(\data_in_frame[20] [3]), 
            .O(n40696));   // verilog/coms.v(94[13:20])
    defparam i26765_4_lut.LUT_INIT = 16'hfac0;
    SB_DFFESS data_out_frame_0___i189 (.Q(\data_out_frame[23] [4]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4920), .S(n58548));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i26766_3_lut (.I0(n40696), .I1(\data_in_frame[20] [3]), .I2(reset), 
            .I3(GND_net), .O(n30098));   // verilog/TinyFPGA_B.v(47[5:10])
    defparam i26766_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 select_775_Select_88_i2_4_lut (.I0(\data_out_frame[11] [0]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[0]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4819));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_88_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_775_Select_87_i2_4_lut (.I0(\data_out_frame[10] [7]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[15]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4818));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_87_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_775_Select_86_i2_4_lut (.I0(\data_out_frame[10] [6]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[14]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4817));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_86_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_775_Select_85_i2_4_lut (.I0(\data_out_frame[10] [5]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[13]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4816));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_85_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFFESS data_out_frame_0___i190 (.Q(\data_out_frame[23] [5]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4919), .S(n58549));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i191 (.Q(\data_out_frame[23] [6]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4918), .S(n58550));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_adj_1310 (.I0(n40817), .I1(n132), .I2(GND_net), .I3(GND_net), 
            .O(n92));
    defparam i1_2_lut_adj_1310.LUT_INIT = 16'h8888;
    SB_LUT4 select_775_Select_84_i2_4_lut (.I0(\data_out_frame[10] [4]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[12]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4815));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_84_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_775_Select_83_i2_4_lut (.I0(\data_out_frame[10] [3]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[11]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4814));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_83_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i26780_4_lut (.I0(n159), .I1(n92), .I2(rx_data[1]), .I3(\data_in_frame[20] [1]), 
            .O(n40711));   // verilog/coms.v(94[13:20])
    defparam i26780_4_lut.LUT_INIT = 16'hfac0;
    SB_LUT4 i26781_3_lut (.I0(n40711), .I1(\data_in_frame[20] [1]), .I2(reset), 
            .I3(GND_net), .O(n30106));   // verilog/TinyFPGA_B.v(47[5:10])
    defparam i26781_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 select_775_Select_82_i2_4_lut (.I0(\data_out_frame[10] [2]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[10]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4813));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_82_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_775_Select_81_i2_4_lut (.I0(\data_out_frame[10] [1]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[9]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4812));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_81_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_6_i7_3_lut_4_lut (.I0(\byte_transmit_counter[2] ), 
            .I1(\byte_transmit_counter[1] ), .I2(n64405), .I3(n64403), 
            .O(n7_adj_5030));   // verilog/coms.v(109[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_6_i7_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 select_775_Select_80_i2_4_lut (.I0(\data_out_frame[10] [0]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[8]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4811));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_80_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFFESS data_out_frame_0___i192 (.Q(\data_out_frame[23] [7]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4917), .S(n58551));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_775_Select_79_i2_4_lut (.I0(\data_out_frame[9] [7]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[23]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4810));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_79_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_775_Select_78_i2_4_lut (.I0(\data_out_frame[9] [6]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[22]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4809));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_78_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFFESS data_out_frame_0___i193 (.Q(\data_out_frame[24] [0]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4916), .S(n58552));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i194 (.Q(\data_out_frame[24] [1]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4915), .S(n58553));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_775_Select_77_i2_4_lut (.I0(\data_out_frame[9] [5]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[21]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4808));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_77_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFFESS data_out_frame_0___i195 (.Q(\data_out_frame[24] [2]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4914), .S(n58504));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_775_Select_76_i2_4_lut (.I0(\data_out_frame[9] [4]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[20]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4807));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_76_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFFESS data_out_frame_0___i196 (.Q(\data_out_frame[24] [3]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4913), .S(n58498));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i197 (.Q(\data_out_frame[24] [4]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4912), .S(n58554));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_7_i7_3_lut_4_lut (.I0(\byte_transmit_counter[2] ), 
            .I1(\byte_transmit_counter[1] ), .I2(n64396), .I3(n64394), 
            .O(n7_adj_5031));   // verilog/coms.v(109[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_7_i7_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 select_775_Select_75_i2_4_lut (.I0(\data_out_frame[9] [3]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[19]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4806));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_75_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFFESS data_out_frame_0___i198 (.Q(\data_out_frame[24] [5]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4911), .S(n58555));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i199 (.Q(\data_out_frame[24] [6]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4910), .S(n58556));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_775_Select_74_i2_4_lut (.I0(\data_out_frame[9] [2]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[18]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4805));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_74_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFFESS data_out_frame_0___i200 (.Q(\data_out_frame[24] [7]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4909), .S(n58557));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i201 (.Q(\data_out_frame[25] [0]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4908), .S(n58558));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i202 (.Q(\data_out_frame[25] [1]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4907), .S(n58497));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_775_Select_73_i2_4_lut (.I0(\data_out_frame[9] [1]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[17]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4804));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_73_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFFESS data_out_frame_0___i203 (.Q(\data_out_frame[25] [2]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4905), .S(n58502));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i204 (.Q(\data_out_frame[25] [3]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4904), .S(n58559));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i59 (.Q(\data_out_frame[7] [2]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4903), .S(n58631));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 n71030_bdd_4_lut (.I0(n71030), .I1(n14_adj_4902), .I2(n7_adj_5032), 
            .I3(byte_transmit_counter[4]), .O(tx_data[1]));
    defparam n71030_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_4_lut_adj_1311 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[9] [0]), 
            .I2(encoder1_position_scaled[16]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4800));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1311.LUT_INIT = 16'ha088;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_0_i7_3_lut_4_lut (.I0(\byte_transmit_counter[2] ), 
            .I1(\byte_transmit_counter[1] ), .I2(n64420), .I3(n64418), 
            .O(n7_adj_5033));   // verilog/coms.v(109[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_0_i7_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 i14098_2_lut (.I0(\byte_transmit_counter[1] ), .I1(\byte_transmit_counter[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n28104));   // verilog/coms.v(109[34:55])
    defparam i14098_2_lut.LUT_INIT = 16'hbbbb;
    SB_DFFESS data_out_frame_0___i60 (.Q(\data_out_frame[7] [3]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4896), .S(n58630));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i61 (.Q(\data_out_frame[7] [4]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4895), .S(n58629));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i48713_3_lut (.I0(\data_out_frame[6] [5]), .I1(\data_out_frame[7] [5]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n64407));
    defparam i48713_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFESS data_out_frame_0___i62 (.Q(\data_out_frame[7] [5]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4893), .S(n58628));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i48714_4_lut (.I0(n64407), .I1(n28104), .I2(\byte_transmit_counter[2] ), 
            .I3(\data_out_frame[1][5] ), .O(n64408));
    defparam i48714_4_lut.LUT_INIT = 16'ha3a0;
    SB_DFFESS data_out_frame_0___i205 (.Q(\data_out_frame[25] [4]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4892), .S(n58560));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i206 (.Q(\data_out_frame[25] [5]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4891), .S(n58561));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i207 (.Q(\data_out_frame[25] [6]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4890), .S(n58562));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i208 (.Q(\data_out_frame[25] [7]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4889), .S(n58563));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i209 (.Q(\data_out_frame[26] [0]), .C(clk16MHz), 
            .E(n2873), .D(n3_adj_4887), .S(n58467));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i210 (.Q(\data_out_frame[26] [1]), .C(clk16MHz), 
            .E(n2873), .D(n3_adj_4821), .S(n58472));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i48712_3_lut (.I0(\data_out_frame[4] [5]), .I1(\data_out_frame[5] [5]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n64406));
    defparam i48712_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFESS data_out_frame_0___i211 (.Q(\data_out_frame[26][2] ), .C(clk16MHz), 
            .E(n2873), .D(n3_adj_4765), .S(n58473));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i212 (.Q(\data_out_frame[26] [3]), .C(clk16MHz), 
            .E(n2873), .D(n3_adj_4763), .S(n58470));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i213 (.Q(\data_out_frame[26] [4]), .C(clk16MHz), 
            .E(n2873), .D(n3_adj_5034), .S(n58474));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i214 (.Q(\data_out_frame[26] [5]), .C(clk16MHz), 
            .E(n2873), .D(n3_adj_4761), .S(n58468));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i215 (.Q(\data_out_frame[26] [6]), .C(clk16MHz), 
            .E(n2873), .D(n3_adj_4758), .S(n58475));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i216 (.Q(\data_out_frame[26] [7]), .C(clk16MHz), 
            .E(n2873), .D(n3_adj_4756), .S(n58476));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i217 (.Q(\data_out_frame[27] [0]), .C(clk16MHz), 
            .E(n2873), .D(n3_adj_4745), .S(n58477));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i218 (.Q(\data_out_frame[27] [1]), .C(clk16MHz), 
            .E(n2873), .D(n3_adj_4743), .S(n58478));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i219 (.Q(\data_out_frame[27][2] ), .C(clk16MHz), 
            .E(n2873), .D(n3_adj_4739), .S(n58479));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i220 (.Q(\data_out_frame[27] [3]), .C(clk16MHz), 
            .E(n2873), .D(n3_adj_4738), .S(n58471));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i221 (.Q(\data_out_frame[27] [4]), .C(clk16MHz), 
            .E(n2873), .D(n3_adj_4737), .S(n58480));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i222 (.Q(\data_out_frame[27] [5]), .C(clk16MHz), 
            .E(n2873), .D(n3_adj_4736), .S(n58469));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i223 (.Q(\data_out_frame[27] [6]), .C(clk16MHz), 
            .E(n2873), .D(n3_adj_4735), .S(n58481));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i224 (.Q(\data_out_frame[27] [7]), .C(clk16MHz), 
            .E(n2873), .D(n3), .S(n58482));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS byte_transmit_counter_i0_i1 (.Q(\byte_transmit_counter[1] ), 
            .C(clk16MHz), .E(n2873), .D(n1_adj_5035), .S(n58675));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS byte_transmit_counter_i0_i2 (.Q(\byte_transmit_counter[2] ), 
            .C(clk16MHz), .E(n2873), .D(n1_adj_5036), .S(n58676));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS byte_transmit_counter_i0_i3 (.Q(byte_transmit_counter[3]), .C(clk16MHz), 
            .E(n2873), .D(n1_adj_5037), .S(n58677));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS byte_transmit_counter_i0_i4 (.Q(byte_transmit_counter[4]), .C(clk16MHz), 
            .E(n2873), .D(n1_adj_5038), .S(n58678));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS byte_transmit_counter_i0_i5 (.Q(byte_transmit_counter[5]), .C(clk16MHz), 
            .E(n2873), .D(n1_adj_5039), .S(n58679));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS byte_transmit_counter_i0_i6 (.Q(byte_transmit_counter[6]), .C(clk16MHz), 
            .E(n2873), .D(n1_adj_5040), .S(n58680));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS byte_transmit_counter_i0_i7 (.Q(byte_transmit_counter[7]), .C(clk16MHz), 
            .E(n2873), .D(n1_adj_5041), .S(n58673));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS tx_transmit_4011 (.Q(r_SM_Main_2__N_3545[0]), .C(clk16MHz), 
            .E(n2873), .D(n1_adj_4992), .S(n28833));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS LED_4014 (.Q(LED_c), .C(clk16MHz), .E(n2873), .D(n5), 
            .S(n28832));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS driver_enable_4015 (.Q(DE_c), .C(clk16MHz), .E(n2873), .D(n26865), 
            .S(n28830));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i30089124_i1_3_lut (.I0(n71255), .I1(n70889), .I2(\byte_transmit_counter[2] ), 
            .I3(GND_net), .O(n14_adj_4798));
    defparam i30089124_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFESS byte_transmit_counter_i0_i0 (.Q(\byte_transmit_counter[0] ), 
            .C(clk16MHz), .E(n2873), .D(n1_adj_5042), .S(n58674));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i63 (.Q(\data_out_frame[7] [6]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5043), .S(n58627));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i64 (.Q(\data_out_frame[7] [7]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5044), .S(n58626));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i51551_2_lut (.I0(n70901), .I1(\byte_transmit_counter[2] ), 
            .I2(GND_net), .I3(GND_net), .O(n66954));
    defparam i51551_2_lut.LUT_INIT = 16'h2222;
    SB_DFFESS data_out_frame_0___i65 (.Q(\data_out_frame[8] [0]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5045), .S(n58625));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i66 (.Q(\data_out_frame[8] [1]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5046), .S(n58624));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 \FRAME_MATCHER.i_1938_add_4_33_lut  (.I0(n67044), .I1(n28304), 
            .I2(\FRAME_MATCHER.i [31]), .I3(n52300), .O(n27980)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1938_add_4_33_lut .LUT_INIT = 16'h8BB8;
    SB_LUT4 \FRAME_MATCHER.i_1938_add_4_32_lut  (.I0(n67043), .I1(n28304), 
            .I2(\FRAME_MATCHER.i [30]), .I3(n52299), .O(n27982)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1938_add_4_32_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_1938_add_4_32  (.CI(n52299), .I0(n28304), 
            .I1(\FRAME_MATCHER.i [30]), .CO(n52300));
    SB_LUT4 \FRAME_MATCHER.i_1938_add_4_31_lut  (.I0(n67042), .I1(n28304), 
            .I2(\FRAME_MATCHER.i [29]), .I3(n52298), .O(n27984)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1938_add_4_31_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_1938_add_4_31  (.CI(n52298), .I0(n28304), 
            .I1(\FRAME_MATCHER.i [29]), .CO(n52299));
    SB_LUT4 \FRAME_MATCHER.i_1938_add_4_30_lut  (.I0(n67037), .I1(n28304), 
            .I2(\FRAME_MATCHER.i [28]), .I3(n52297), .O(n27986)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1938_add_4_30_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_1938_add_4_30  (.CI(n52297), .I0(n28304), 
            .I1(\FRAME_MATCHER.i [28]), .CO(n52298));
    SB_LUT4 \FRAME_MATCHER.i_1938_add_4_29_lut  (.I0(n67036), .I1(n28304), 
            .I2(\FRAME_MATCHER.i [27]), .I3(n52296), .O(n27988)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1938_add_4_29_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_1938_add_4_29  (.CI(n52296), .I0(n28304), 
            .I1(\FRAME_MATCHER.i [27]), .CO(n52297));
    SB_LUT4 \FRAME_MATCHER.i_1938_add_4_28_lut  (.I0(n67028), .I1(n28304), 
            .I2(\FRAME_MATCHER.i [26]), .I3(n52295), .O(n27990)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1938_add_4_28_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_1938_add_4_28  (.CI(n52295), .I0(n28304), 
            .I1(\FRAME_MATCHER.i [26]), .CO(n52296));
    SB_LUT4 \FRAME_MATCHER.i_1938_add_4_27_lut  (.I0(n67003), .I1(n28304), 
            .I2(\FRAME_MATCHER.i [25]), .I3(n52294), .O(n27992)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1938_add_4_27_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_1938_add_4_27  (.CI(n52294), .I0(n28304), 
            .I1(\FRAME_MATCHER.i [25]), .CO(n52295));
    SB_LUT4 \FRAME_MATCHER.i_1938_add_4_26_lut  (.I0(n66999), .I1(n28304), 
            .I2(\FRAME_MATCHER.i [24]), .I3(n52293), .O(n27994)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1938_add_4_26_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_1938_add_4_26  (.CI(n52293), .I0(n28304), 
            .I1(\FRAME_MATCHER.i [24]), .CO(n52294));
    SB_LUT4 \FRAME_MATCHER.i_1938_add_4_25_lut  (.I0(n66998), .I1(n28304), 
            .I2(\FRAME_MATCHER.i [23]), .I3(n52292), .O(n27996)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1938_add_4_25_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_1938_add_4_25  (.CI(n52292), .I0(n28304), 
            .I1(\FRAME_MATCHER.i [23]), .CO(n52293));
    SB_LUT4 \FRAME_MATCHER.i_1938_add_4_24_lut  (.I0(n66997), .I1(n28304), 
            .I2(\FRAME_MATCHER.i [22]), .I3(n52291), .O(n27998)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1938_add_4_24_lut .LUT_INIT = 16'h8BB8;
    SB_LUT4 select_775_Select_71_i2_4_lut (.I0(\data_out_frame[8] [7]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder0_position_scaled[7]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4795));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_71_i2_4_lut.LUT_INIT = 16'hc088;
    SB_CARRY \FRAME_MATCHER.i_1938_add_4_24  (.CI(n52291), .I0(n28304), 
            .I1(\FRAME_MATCHER.i [22]), .CO(n52292));
    SB_LUT4 \FRAME_MATCHER.i_1938_add_4_23_lut  (.I0(n66993), .I1(n28304), 
            .I2(\FRAME_MATCHER.i [21]), .I3(n52290), .O(n28000)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1938_add_4_23_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_1938_add_4_23  (.CI(n52290), .I0(n28304), 
            .I1(\FRAME_MATCHER.i [21]), .CO(n52291));
    SB_LUT4 \FRAME_MATCHER.i_1938_add_4_22_lut  (.I0(n66992), .I1(n28304), 
            .I2(\FRAME_MATCHER.i [20]), .I3(n52289), .O(n28002)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1938_add_4_22_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_1938_add_4_22  (.CI(n52289), .I0(n28304), 
            .I1(\FRAME_MATCHER.i [20]), .CO(n52290));
    SB_LUT4 \FRAME_MATCHER.i_1938_add_4_21_lut  (.I0(n66973), .I1(n28304), 
            .I2(\FRAME_MATCHER.i [19]), .I3(n52288), .O(n28004)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1938_add_4_21_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_1938_add_4_21  (.CI(n52288), .I0(n28304), 
            .I1(\FRAME_MATCHER.i [19]), .CO(n52289));
    SB_LUT4 \FRAME_MATCHER.i_1938_add_4_20_lut  (.I0(n66972), .I1(n28304), 
            .I2(\FRAME_MATCHER.i [18]), .I3(n52287), .O(n28006)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1938_add_4_20_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_1938_add_4_20  (.CI(n52287), .I0(n28304), 
            .I1(\FRAME_MATCHER.i [18]), .CO(n52288));
    SB_LUT4 \FRAME_MATCHER.i_1938_add_4_19_lut  (.I0(n66967), .I1(n28304), 
            .I2(\FRAME_MATCHER.i [17]), .I3(n52286), .O(n28008)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1938_add_4_19_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_1938_add_4_19  (.CI(n52286), .I0(n28304), 
            .I1(\FRAME_MATCHER.i [17]), .CO(n52287));
    SB_LUT4 \FRAME_MATCHER.i_1938_add_4_18_lut  (.I0(n66966), .I1(n28304), 
            .I2(\FRAME_MATCHER.i [16]), .I3(n52285), .O(n28010)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1938_add_4_18_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_1938_add_4_18  (.CI(n52285), .I0(n28304), 
            .I1(\FRAME_MATCHER.i [16]), .CO(n52286));
    SB_LUT4 \FRAME_MATCHER.i_1938_add_4_17_lut  (.I0(n66962), .I1(n28304), 
            .I2(\FRAME_MATCHER.i [15]), .I3(n52284), .O(n28012)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1938_add_4_17_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_1938_add_4_17  (.CI(n52284), .I0(n28304), 
            .I1(\FRAME_MATCHER.i [15]), .CO(n52285));
    SB_LUT4 \FRAME_MATCHER.i_1938_add_4_16_lut  (.I0(n66959), .I1(n28304), 
            .I2(\FRAME_MATCHER.i [14]), .I3(n52283), .O(n28014)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1938_add_4_16_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_1938_add_4_16  (.CI(n52283), .I0(n28304), 
            .I1(\FRAME_MATCHER.i [14]), .CO(n52284));
    SB_LUT4 \FRAME_MATCHER.i_1938_add_4_15_lut  (.I0(n66955), .I1(n28304), 
            .I2(\FRAME_MATCHER.i [13]), .I3(n52282), .O(n28016)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1938_add_4_15_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_1938_add_4_15  (.CI(n52282), .I0(n28304), 
            .I1(\FRAME_MATCHER.i [13]), .CO(n52283));
    SB_LUT4 \FRAME_MATCHER.i_1938_add_4_14_lut  (.I0(n66953), .I1(n28304), 
            .I2(\FRAME_MATCHER.i [12]), .I3(n52281), .O(n28018)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1938_add_4_14_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_1938_add_4_14  (.CI(n52281), .I0(n28304), 
            .I1(\FRAME_MATCHER.i [12]), .CO(n52282));
    SB_LUT4 \FRAME_MATCHER.i_1938_add_4_13_lut  (.I0(n66952), .I1(n28304), 
            .I2(\FRAME_MATCHER.i [11]), .I3(n52280), .O(n28020)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1938_add_4_13_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_1938_add_4_13  (.CI(n52280), .I0(n28304), 
            .I1(\FRAME_MATCHER.i [11]), .CO(n52281));
    SB_LUT4 \FRAME_MATCHER.i_1938_add_4_12_lut  (.I0(n66951), .I1(n28304), 
            .I2(\FRAME_MATCHER.i [10]), .I3(n52279), .O(n28022)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1938_add_4_12_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_1938_add_4_12  (.CI(n52279), .I0(n28304), 
            .I1(\FRAME_MATCHER.i [10]), .CO(n52280));
    SB_LUT4 \FRAME_MATCHER.i_1938_add_4_11_lut  (.I0(n66944), .I1(n28304), 
            .I2(\FRAME_MATCHER.i [9]), .I3(n52278), .O(n28024)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1938_add_4_11_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_1938_add_4_11  (.CI(n52278), .I0(n28304), 
            .I1(\FRAME_MATCHER.i [9]), .CO(n52279));
    SB_LUT4 \FRAME_MATCHER.i_1938_add_4_10_lut  (.I0(n66942), .I1(n28304), 
            .I2(\FRAME_MATCHER.i [8]), .I3(n52277), .O(n28026)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1938_add_4_10_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_1938_add_4_10  (.CI(n52277), .I0(n28304), 
            .I1(\FRAME_MATCHER.i [8]), .CO(n52278));
    SB_LUT4 \FRAME_MATCHER.i_1938_add_4_9_lut  (.I0(n66941), .I1(n28304), 
            .I2(\FRAME_MATCHER.i [7]), .I3(n52276), .O(n28028)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1938_add_4_9_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_1938_add_4_9  (.CI(n52276), .I0(n28304), .I1(\FRAME_MATCHER.i [7]), 
            .CO(n52277));
    SB_LUT4 \FRAME_MATCHER.i_1938_add_4_8_lut  (.I0(n66940), .I1(n28304), 
            .I2(\FRAME_MATCHER.i [6]), .I3(n52275), .O(n28030)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1938_add_4_8_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_1938_add_4_8  (.CI(n52275), .I0(n28304), .I1(\FRAME_MATCHER.i [6]), 
            .CO(n52276));
    SB_LUT4 \FRAME_MATCHER.i_1938_add_4_7_lut  (.I0(n66939), .I1(n28304), 
            .I2(\FRAME_MATCHER.i[5] ), .I3(n52274), .O(n28032)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1938_add_4_7_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_1938_add_4_7  (.CI(n52274), .I0(n28304), .I1(\FRAME_MATCHER.i[5] ), 
            .CO(n52275));
    SB_LUT4 \FRAME_MATCHER.i_1938_add_4_6_lut  (.I0(n66938), .I1(n28304), 
            .I2(\FRAME_MATCHER.i[4] ), .I3(n52273), .O(n28034)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1938_add_4_6_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_1938_add_4_6  (.CI(n52273), .I0(n28304), .I1(\FRAME_MATCHER.i[4] ), 
            .CO(n52274));
    SB_LUT4 \FRAME_MATCHER.i_1938_add_4_5_lut  (.I0(n66937), .I1(n28304), 
            .I2(\FRAME_MATCHER.i[3] ), .I3(n52272), .O(n28036)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1938_add_4_5_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_1938_add_4_5  (.CI(n52272), .I0(n28304), .I1(\FRAME_MATCHER.i[3] ), 
            .CO(n52273));
    SB_LUT4 \FRAME_MATCHER.i_1938_add_4_4_lut  (.I0(n66936), .I1(n28304), 
            .I2(\FRAME_MATCHER.i [2]), .I3(n52271), .O(n28038)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1938_add_4_4_lut .LUT_INIT = 16'h8BB8;
    SB_LUT4 i13_2_lut_adj_1312 (.I0(pwm_setpoint[22]), .I1(\pwm_counter[22] ), 
            .I2(GND_net), .I3(GND_net), .O(n45));   // verilog/pwm.v(11[19:30])
    defparam i13_2_lut_adj_1312.LUT_INIT = 16'h6666;
    SB_CARRY \FRAME_MATCHER.i_1938_add_4_4  (.CI(n52271), .I0(n28304), .I1(\FRAME_MATCHER.i [2]), 
            .CO(n52272));
    SB_LUT4 \FRAME_MATCHER.i_1938_add_4_3_lut  (.I0(n66935), .I1(n28304), 
            .I2(\FRAME_MATCHER.i [1]), .I3(n52270), .O(n28040)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1938_add_4_3_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_1938_add_4_3  (.CI(n52270), .I0(n28304), .I1(\FRAME_MATCHER.i [1]), 
            .CO(n52271));
    SB_LUT4 \FRAME_MATCHER.i_1938_add_4_2_lut  (.I0(GND_net), .I1(n161_c), 
            .I2(\FRAME_MATCHER.i[0] ), .I3(GND_net), .O(n133[0])) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1938_add_4_2_lut .LUT_INIT = 16'hC33C;
    SB_CARRY \FRAME_MATCHER.i_1938_add_4_2  (.CI(GND_net), .I0(n161_c), 
            .I1(\FRAME_MATCHER.i[0] ), .CO(n52270));
    SB_LUT4 i15_2_lut (.I0(pwm_setpoint[21]), .I1(\pwm_counter[21] ), .I2(GND_net), 
            .I3(GND_net), .O(n43));   // verilog/pwm.v(11[19:30])
    defparam i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_55308 (.I0(\byte_transmit_counter[1] ), 
            .I1(n4_adj_5048), .I2(n5_adj_5049), .I3(\byte_transmit_counter[2] ), 
            .O(n71024));
    defparam byte_transmit_counter_1__bdd_4_lut_55308.LUT_INIT = 16'he4aa;
    SB_LUT4 select_775_Select_14_i2_3_lut (.I0(\data_out_frame[1][6] ), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\FRAME_MATCHER.state_31__N_2612 [3]), .I3(GND_net), .O(n2_adj_5017));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_14_i2_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_1_i7_3_lut_4_lut (.I0(\byte_transmit_counter[2] ), 
            .I1(\byte_transmit_counter[1] ), .I2(n64423), .I3(n64421), 
            .O(n7_adj_5032));   // verilog/coms.v(109[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_1_i7_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_5_i7_3_lut_4_lut (.I0(\byte_transmit_counter[2] ), 
            .I1(\byte_transmit_counter[1] ), .I2(n64408), .I3(n64406), 
            .O(n7_adj_4799));   // verilog/coms.v(109[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_5_i7_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_2_i7_3_lut_4_lut (.I0(\byte_transmit_counter[2] ), 
            .I1(\byte_transmit_counter[1] ), .I2(n64414), .I3(n64412), 
            .O(n7_adj_5028));   // verilog/coms.v(109[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_2_i7_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 select_775_Select_13_i2_3_lut (.I0(\data_out_frame[1][5] ), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\FRAME_MATCHER.state_31__N_2612 [3]), .I3(GND_net), .O(n2_adj_5016));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_13_i2_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1313 (.I0(\data_in_frame[2] [1]), .I1(\data_in_frame[2] [3]), 
            .I2(\data_in_frame[0]_c [2]), .I3(\data_in_frame[0] [1]), .O(n25815));   // verilog/coms.v(77[16:43])
    defparam i1_2_lut_3_lut_4_lut_adj_1313.LUT_INIT = 16'h6996;
    SB_LUT4 i2_2_lut_3_lut_4_lut (.I0(\data_out_frame[6] [6]), .I1(\data_out_frame[4] [5]), 
            .I2(\data_out_frame[4] [4]), .I3(\data_out_frame[9] [0]), .O(n10_adj_4869));   // verilog/coms.v(100[12:26])
    defparam i2_2_lut_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1314 (.I0(\data_out_frame[6] [6]), .I1(\data_out_frame[4] [5]), 
            .I2(\data_out_frame[4] [4]), .I3(n26039), .O(n6_adj_4859));   // verilog/coms.v(100[12:26])
    defparam i1_2_lut_3_lut_4_lut_adj_1314.LUT_INIT = 16'h6996;
    SB_LUT4 n71024_bdd_4_lut (.I0(n71024), .I1(n67066), .I2(n67065), .I3(\byte_transmit_counter[2] ), 
            .O(n71027));
    defparam n71024_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_4_i5_3_lut (.I0(\data_out_frame[6] [4]), 
            .I1(\data_out_frame[7] [4]), .I2(\byte_transmit_counter[0] ), 
            .I3(GND_net), .O(n5_adj_5049));   // verilog/coms.v(109[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_4_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_4_i4_3_lut (.I0(\data_out_frame[4] [4]), 
            .I1(\data_out_frame[5] [4]), .I2(\byte_transmit_counter[0] ), 
            .I3(GND_net), .O(n4_adj_5048));   // verilog/coms.v(109[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_4_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1315 (.I0(n54460), .I1(n54116), .I2(n54572), 
            .I3(n26689), .O(n59226));
    defparam i1_4_lut_adj_1315.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1316 (.I0(n54458), .I1(n58969), .I2(GND_net), 
            .I3(GND_net), .O(n63809));
    defparam i1_2_lut_adj_1316.LUT_INIT = 16'h6666;
    SB_LUT4 select_775_Select_11_i2_3_lut (.I0(\data_out_frame[1][3] ), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\FRAME_MATCHER.state_31__N_2612 [3]), .I3(GND_net), .O(n2_adj_5015));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_11_i2_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i1_4_lut_adj_1317 (.I0(n59232), .I1(n59380), .I2(n54447), 
            .I3(n63809), .O(n63815));
    defparam i1_4_lut_adj_1317.LUT_INIT = 16'h9669;
    SB_LUT4 i1_4_lut_adj_1318 (.I0(n61135), .I1(n58771), .I2(n59183), 
            .I3(n63815), .O(n61398));
    defparam i1_4_lut_adj_1318.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_3_lut (.I0(\FRAME_MATCHER.i_31__N_2514 ), .I1(\FRAME_MATCHER.i_31__N_2512 ), 
            .I2(\FRAME_MATCHER.i_31__N_2508 ), .I3(GND_net), .O(n3468));   // verilog/coms.v(148[4] 304[11])
    defparam i1_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1319 (.I0(\FRAME_MATCHER.i_31__N_2514 ), 
            .I1(\FRAME_MATCHER.i_31__N_2512 ), .I2(\FRAME_MATCHER.i_31__N_2511 ), 
            .I3(\FRAME_MATCHER.state[3] ), .O(n47954));   // verilog/coms.v(148[4] 304[11])
    defparam i1_2_lut_3_lut_4_lut_adj_1319.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1320 (.I0(n59235), .I1(n59379), .I2(n54411), 
            .I3(\data_in_frame[21] [0]), .O(n63951));
    defparam i1_4_lut_adj_1320.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1321 (.I0(n63951), .I1(n58771), .I2(n63743), 
            .I3(n59341), .O(n54116));
    defparam i1_4_lut_adj_1321.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1322 (.I0(n61410), .I1(n53713), .I2(GND_net), 
            .I3(GND_net), .O(Kp_23__N_1551));
    defparam i1_2_lut_adj_1322.LUT_INIT = 16'h9999;
    SB_LUT4 i1_2_lut_adj_1323 (.I0(\data_in_frame[20] [6]), .I1(\data_in_frame[18] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n59409));
    defparam i1_2_lut_adj_1323.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1324 (.I0(n59284), .I1(n25906), .I2(n53503), 
            .I3(n59427), .O(n10_adj_5050));
    defparam i4_4_lut_adj_1324.LUT_INIT = 16'h6996;
    SB_LUT4 i2_4_lut_adj_1325 (.I0(n26239), .I1(n25744), .I2(\data_in_frame[11] [5]), 
            .I3(n53442), .O(n8_adj_5051));
    defparam i2_4_lut_adj_1325.LUT_INIT = 16'h6996;
    SB_LUT4 i15795_3_lut_4_lut (.I0(n8_adj_13), .I1(n58760), .I2(rx_data[0]), 
            .I3(\data_in_frame[2] [0]), .O(n29801));
    defparam i15795_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i5_4_lut_adj_1326 (.I0(n25979), .I1(n7_adj_5053), .I2(n26435), 
            .I3(n8_adj_5051), .O(n59427));
    defparam i5_4_lut_adj_1326.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1327 (.I0(\data_in_frame[13] [7]), .I1(n59427), 
            .I2(n59368), .I3(n59083), .O(n25112));
    defparam i3_4_lut_adj_1327.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1328 (.I0(\data_in_frame[18] [3]), .I1(n54513), 
            .I2(GND_net), .I3(GND_net), .O(n54630));
    defparam i1_2_lut_adj_1328.LUT_INIT = 16'h6666;
    SB_LUT4 i2_2_lut_adj_1329 (.I0(n25112), .I1(\data_in_frame[20] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n7_adj_5054));
    defparam i2_2_lut_adj_1329.LUT_INIT = 16'h6666;
    SB_LUT4 i15798_3_lut_4_lut (.I0(n8_adj_13), .I1(n58760), .I2(rx_data[1]), 
            .I3(\data_in_frame[2] [1]), .O(n29804));
    defparam i15798_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i4_4_lut_adj_1330 (.I0(n7_adj_5054), .I1(\data_in_frame[20] [3]), 
            .I2(n54630), .I3(\data_in_frame[18] [1]), .O(n59046));
    defparam i4_4_lut_adj_1330.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1331 (.I0(\data_in_frame[15] [5]), .I1(\data_in_frame[17] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n59368));
    defparam i1_2_lut_adj_1331.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_4_lut_adj_1332 (.I0(n58812), .I1(n59259), .I2(\data_in_frame[3][6] ), 
            .I3(\data_in_frame[6] [0]), .O(n25843));   // verilog/coms.v(78[16:27])
    defparam i2_3_lut_4_lut_adj_1332.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1333 (.I0(\data_in_frame[19] [7]), .I1(n59371), 
            .I2(\data_in_frame[20] [1]), .I3(GND_net), .O(n59018));
    defparam i2_3_lut_adj_1333.LUT_INIT = 16'h9696;
    SB_LUT4 i6_2_lut_3_lut_4_lut (.I0(\data_in_frame[18] [2]), .I1(\data_in_frame[18] [4]), 
            .I2(\data_in_frame[20] [5]), .I3(n59018), .O(n22_adj_5055));
    defparam i6_2_lut_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i12_4_lut_adj_1334 (.I0(n54511), .I1(\data_in_frame[20] [0]), 
            .I2(n61410), .I3(n54411), .O(n28_adj_5056));
    defparam i12_4_lut_adj_1334.LUT_INIT = 16'h6996;
    SB_LUT4 i10_4_lut_adj_1335 (.I0(n59368), .I1(n59380), .I2(n59046), 
            .I3(n53511), .O(n26_adj_5057));
    defparam i10_4_lut_adj_1335.LUT_INIT = 16'h6996;
    SB_LUT4 i11_4_lut_adj_1336 (.I0(n59409), .I1(n22_adj_5055), .I2(\data_in_frame[19] [6]), 
            .I3(n54588), .O(n27_c));
    defparam i11_4_lut_adj_1336.LUT_INIT = 16'h9669;
    SB_LUT4 i9_4_lut_adj_1337 (.I0(n61135), .I1(n59092), .I2(n58981), 
            .I3(\data_in_frame[18] [6]), .O(n25_adj_5058));
    defparam i9_4_lut_adj_1337.LUT_INIT = 16'h9669;
    SB_LUT4 i15_4_lut_adj_1338 (.I0(n25_adj_5058), .I1(n27_c), .I2(n26_adj_5057), 
            .I3(n28_adj_5056), .O(n54460));
    defparam i15_4_lut_adj_1338.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1339 (.I0(n54447), .I1(\data_in_frame[19] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n59235));
    defparam i1_2_lut_adj_1339.LUT_INIT = 16'h6666;
    SB_LUT4 i15801_3_lut_4_lut (.I0(n8_adj_13), .I1(n58760), .I2(rx_data[2]), 
            .I3(\data_in_frame[2] [2]), .O(n29807));
    defparam i15801_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i3_4_lut_adj_1340 (.I0(\data_in_frame[18] [5]), .I1(n26605), 
            .I2(n25853), .I3(n26359), .O(n58969));   // verilog/coms.v(81[16:27])
    defparam i3_4_lut_adj_1340.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1341 (.I0(n54458), .I1(n59067), .I2(GND_net), 
            .I3(GND_net), .O(n54527));
    defparam i1_2_lut_adj_1341.LUT_INIT = 16'h6666;
    SB_LUT4 i6_4_lut_adj_1342 (.I0(n59459), .I1(\data_in_frame[11] [5]), 
            .I2(n59097), .I3(\data_in_frame[13] [7]), .O(n14_adj_5059));
    defparam i6_4_lut_adj_1342.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1343 (.I0(\data_in_frame[14] [1]), .I1(\data_in_frame[9] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n9_adj_5060));
    defparam i1_2_lut_adj_1343.LUT_INIT = 16'h6666;
    SB_LUT4 i7_4_lut_adj_1344 (.I0(n9_adj_5060), .I1(n14_adj_5059), .I2(n59374), 
            .I3(n59134), .O(n53503));
    defparam i7_4_lut_adj_1344.LUT_INIT = 16'h9669;
    SB_LUT4 i15804_3_lut_4_lut (.I0(n8_adj_13), .I1(n58760), .I2(rx_data[3]), 
            .I3(\data_in_frame[2] [3]), .O(n29810));
    defparam i15804_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15807_3_lut_4_lut (.I0(n8_adj_13), .I1(n58760), .I2(rx_data[4]), 
            .I3(\data_in_frame[2] [4]), .O(n29813));
    defparam i15807_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1345 (.I0(n53460), .I1(\data_in_frame[15] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n59206));
    defparam i1_2_lut_adj_1345.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1346 (.I0(\data_in_frame[16] [0]), .I1(\data_in_frame[13] [1]), 
            .I2(n53570), .I3(GND_net), .O(n59083));
    defparam i2_3_lut_adj_1346.LUT_INIT = 16'h9696;
    SB_LUT4 i1_4_lut_adj_1347 (.I0(\data_in_frame[15] [4]), .I1(\data_in_frame[16] [1]), 
            .I2(\data_in_frame[15] [2]), .I3(\data_in_frame[16] [4]), .O(n63675));
    defparam i1_4_lut_adj_1347.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1348 (.I0(\data_in_frame[12] [4]), .I1(\data_in_frame[15] [3]), 
            .I2(\data_in_frame[13] [2]), .I3(\data_in_frame[17] [1]), .O(n63677));
    defparam i1_4_lut_adj_1348.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1349 (.I0(n59174), .I1(n59060), .I2(n59146), 
            .I3(Kp_23__N_1389), .O(n63687));
    defparam i1_4_lut_adj_1349.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1350 (.I0(n63687), .I1(n63677), .I2(n59137), 
            .I3(n63675), .O(n63689));
    defparam i1_4_lut_adj_1350.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1351 (.I0(n26435), .I1(n58960), .I2(n25906), 
            .I3(n63689), .O(n63695));
    defparam i1_4_lut_adj_1351.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1352 (.I0(n61382), .I1(n54155), .I2(n59439), 
            .I3(n63695), .O(n63701));
    defparam i1_4_lut_adj_1352.LUT_INIT = 16'h9669;
    SB_LUT4 i1_4_lut_adj_1353 (.I0(n59083), .I1(n59206), .I2(n59471), 
            .I3(n63701), .O(n63707));
    defparam i1_4_lut_adj_1353.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1354 (.I0(n54447), .I1(n26755), .I2(n25724), 
            .I3(n63707), .O(n61135));
    defparam i1_4_lut_adj_1354.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1355 (.I0(\data_in_frame[17] [5]), .I1(n7_adj_4906), 
            .I2(\data_in_frame[15] [3]), .I3(n53570), .O(n10_adj_5061));
    defparam i4_4_lut_adj_1355.LUT_INIT = 16'h6996;
    SB_LUT4 i15811_3_lut_4_lut (.I0(n8_adj_13), .I1(n58760), .I2(rx_data[5]), 
            .I3(\data_in_frame[2] [5]), .O(n29817));
    defparam i15811_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i3_4_lut_adj_1356 (.I0(n58851), .I1(\data_in_frame[12] [7]), 
            .I2(\data_in_frame[13] [1]), .I3(n26639), .O(n61117));   // verilog/coms.v(74[16:27])
    defparam i3_4_lut_adj_1356.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut_adj_1357 (.I0(n61117), .I1(n59165), .I2(n10_adj_5061), 
            .I3(n60961), .O(n53713));
    defparam i5_4_lut_adj_1357.LUT_INIT = 16'h9669;
    SB_LUT4 i1_3_lut (.I0(n53713), .I1(n61135), .I2(\data_in_frame[18] [0]), 
            .I3(GND_net), .O(n54516));
    defparam i1_3_lut.LUT_INIT = 16'h6969;
    SB_LUT4 i1_2_lut_adj_1358 (.I0(\data_in_frame[18] [1]), .I1(\data_in_frame[18] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n26605));
    defparam i1_2_lut_adj_1358.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1359 (.I0(n54527), .I1(n54516), .I2(n58969), 
            .I3(\data_in_frame[16] [5]), .O(n54033));   // verilog/coms.v(81[16:27])
    defparam i1_4_lut_adj_1359.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1360 (.I0(n58981), .I1(\data_in_frame[18] [7]), 
            .I2(n54033), .I3(n59341), .O(n10_adj_5062));
    defparam i4_4_lut_adj_1360.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_1361 (.I0(n54475), .I1(n10_adj_5062), .I2(\data_in_frame[18] [4]), 
            .I3(GND_net), .O(Kp_23__N_1607));
    defparam i5_3_lut_adj_1361.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1362 (.I0(\data_in_frame[21] [2]), .I1(n58925), 
            .I2(\data_in_frame[21] [1]), .I3(GND_net), .O(n6_adj_5063));   // verilog/coms.v(99[12:25])
    defparam i2_3_lut_adj_1362.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_1363 (.I0(\data_in_frame[21] [7]), .I1(n6_adj_5063), 
            .I2(n59033), .I3(\data_in_frame[21] [6]), .O(n26689));   // verilog/coms.v(99[12:25])
    defparam i3_4_lut_adj_1363.LUT_INIT = 16'h6996;
    SB_LUT4 i15814_3_lut_4_lut (.I0(n8_adj_13), .I1(n58760), .I2(rx_data[6]), 
            .I3(\data_in_frame[2] [6]), .O(n29820));
    defparam i15814_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1364 (.I0(\data_in_frame[18] [7]), .I1(\data_in_frame[18] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n25853));   // verilog/coms.v(81[16:27])
    defparam i1_2_lut_adj_1364.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1365 (.I0(\data_in_frame[19] [0]), .I1(n26085), 
            .I2(n54475), .I3(GND_net), .O(n54572));
    defparam i2_3_lut_adj_1365.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1366 (.I0(n26085), .I1(n59106), .I2(GND_net), 
            .I3(GND_net), .O(n59092));
    defparam i1_2_lut_adj_1366.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1367 (.I0(\data_in_frame[23] [4]), .I1(n54572), 
            .I2(GND_net), .I3(GND_net), .O(n5_adj_5064));
    defparam i1_2_lut_adj_1367.LUT_INIT = 16'h9999;
    SB_LUT4 i1_4_lut_adj_1368 (.I0(\data_in_frame[19] [2]), .I1(\data_in_frame[17] [1]), 
            .I2(n54473), .I3(n26134), .O(n59106));
    defparam i1_4_lut_adj_1368.LUT_INIT = 16'h9669;
    SB_LUT4 i1_3_lut_adj_1369 (.I0(\data_in_frame[19] [4]), .I1(n54452), 
            .I2(n59143), .I3(GND_net), .O(n54588));
    defparam i1_3_lut_adj_1369.LUT_INIT = 16'h6969;
    SB_LUT4 i4_4_lut_adj_1370 (.I0(\data_in_frame[14] [4]), .I1(n54155), 
            .I2(\data_in_frame[9] [7]), .I3(n6_adj_5065), .O(n54458));
    defparam i4_4_lut_adj_1370.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1371 (.I0(\data_in_frame[16] [7]), .I1(\data_in_frame[16] [6]), 
            .I2(\data_in_frame[14] [6]), .I3(\data_in_frame[17] [0]), .O(n59137));
    defparam i3_4_lut_adj_1371.LUT_INIT = 16'h6996;
    SB_LUT4 i15817_3_lut_4_lut (.I0(n8_adj_13), .I1(n58760), .I2(rx_data[7]), 
            .I3(\data_in_frame[2] [7]), .O(n29823));
    defparam i15817_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i3_4_lut_adj_1372 (.I0(\data_in_frame[14] [5]), .I1(n26438), 
            .I2(n59199), .I3(\data_in_frame[12] [4]), .O(n61382));
    defparam i3_4_lut_adj_1372.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1373 (.I0(n61382), .I1(\data_in_frame[16] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n59194));
    defparam i1_2_lut_adj_1373.LUT_INIT = 16'h9999;
    SB_LUT4 i54311_3_lut (.I0(rx_data[7]), .I1(\data_in_frame[7]_c [7]), 
            .I2(n59638), .I3(GND_net), .O(n58086));   // verilog/coms.v(94[13:20])
    defparam i54311_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i54312_3_lut (.I0(rx_data[6]), .I1(\data_in_frame[7]_c [6]), 
            .I2(n59638), .I3(GND_net), .O(n58092));   // verilog/coms.v(94[13:20])
    defparam i54312_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2_4_lut_adj_1374 (.I0(n59137), .I1(n54458), .I2(n6_adj_5066), 
            .I3(\data_in_frame[12] [4]), .O(n26134));
    defparam i2_4_lut_adj_1374.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1375 (.I0(n54518), .I1(n54417), .I2(GND_net), 
            .I3(GND_net), .O(n5_adj_5067));
    defparam i1_2_lut_adj_1375.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1376 (.I0(\data_in_frame[14] [3]), .I1(n5_adj_5067), 
            .I2(n59080), .I3(n61279), .O(n59067));
    defparam i1_4_lut_adj_1376.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1377 (.I0(n59067), .I1(n26134), .I2(\data_in_frame[19] [1]), 
            .I3(n59194), .O(n10_adj_5068));
    defparam i4_4_lut_adj_1377.LUT_INIT = 16'h6996;
    SB_LUT4 i28193_3_lut (.I0(\duty[3] ), .I1(\duty[0] ), .I2(n260), .I3(GND_net), 
            .O(n7_adj_14));
    defparam i28193_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 select_775_Select_9_i2_3_lut (.I0(\data_out_frame[1][1] ), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\FRAME_MATCHER.state_31__N_2612 [3]), .I3(GND_net), .O(n2_adj_5014));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_9_i2_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i5_3_lut_adj_1378 (.I0(\data_in_frame[16] [5]), .I1(n10_adj_5068), 
            .I2(\data_in_frame[18] [7]), .I3(GND_net), .O(n26085));
    defparam i5_3_lut_adj_1378.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1379 (.I0(n26085), .I1(\data_in_frame[21] [3]), 
            .I2(\data_in_frame[21] [4]), .I3(GND_net), .O(n58925));
    defparam i2_3_lut_adj_1379.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_1380 (.I0(n53442), .I1(n59100), .I2(\data_in_frame[12] [1]), 
            .I3(n54520), .O(n61279));
    defparam i3_4_lut_adj_1380.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1381 (.I0(\data_in_frame[8] [6]), .I1(\data_in_frame[6] [3]), 
            .I2(\data_in_frame[8] [4]), .I3(\data_in_frame[8] [3]), .O(n63929));
    defparam i1_4_lut_adj_1381.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1382 (.I0(n63929), .I1(n59109), .I2(\data_in_frame[1] [6]), 
            .I3(\data_in_frame[8] [7]), .O(n63935));
    defparam i1_4_lut_adj_1382.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1383 (.I0(n59256), .I1(n63935), .I2(n58894), 
            .I3(n59412), .O(n63939));
    defparam i1_4_lut_adj_1383.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1384 (.I0(n70018), .I1(n26633), .I2(n59259), 
            .I3(n63939), .O(n63945));
    defparam i1_4_lut_adj_1384.LUT_INIT = 16'h9669;
    SB_LUT4 i1_4_lut_adj_1385 (.I0(n63945), .I1(\data_in_frame[11] [7]), 
            .I2(n54518), .I3(\data_in_frame[12] [0]), .O(n59374));
    defparam i1_4_lut_adj_1385.LUT_INIT = 16'h9669;
    SB_LUT4 i1_4_lut_adj_1386 (.I0(\data_in_frame[9] [5]), .I1(\data_in_frame[11] [6]), 
            .I2(\data_in_frame[11] [7]), .I3(\data_in_frame[7] [1]), .O(n63897));
    defparam i1_4_lut_adj_1386.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1387 (.I0(\data_in_frame[4] [7]), .I1(\data_in_frame[9] [3]), 
            .I2(\data_in_frame[5] [0]), .I3(\data_in_frame[6] [0]), .O(n63899));
    defparam i1_4_lut_adj_1387.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1388 (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(n140), .I3(n3468), .O(n40663));   // verilog/coms.v(156[9:50])
    defparam i1_2_lut_3_lut_4_lut_adj_1388.LUT_INIT = 16'hfbff;
    SB_LUT4 i1_3_lut_adj_1389 (.I0(n59121), .I1(n63899), .I2(n63897), 
            .I3(GND_net), .O(n63903));
    defparam i1_3_lut_adj_1389.LUT_INIT = 16'h9696;
    SB_LUT4 i1_4_lut_adj_1390 (.I0(n59064), .I1(n58792), .I2(n59100), 
            .I3(n63903), .O(n63909));
    defparam i1_4_lut_adj_1390.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1391 (.I0(n59474), .I1(n54113), .I2(n59397), 
            .I3(n63909), .O(n63915));
    defparam i1_4_lut_adj_1391.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1392 (.I0(n54518), .I1(n59374), .I2(n61279), 
            .I3(n63915), .O(n54468));
    defparam i1_4_lut_adj_1392.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1393 (.I0(\data_in_frame[18] [2]), .I1(\data_in_frame[18] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n26359));   // verilog/coms.v(81[16:27])
    defparam i1_2_lut_adj_1393.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1394 (.I0(n59316), .I1(\data_in_frame[14] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_5070));
    defparam i1_2_lut_adj_1394.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1395 (.I0(Kp_23__N_1271), .I1(n54468), .I2(n25925), 
            .I3(n6_adj_5070), .O(n59379));
    defparam i4_4_lut_adj_1395.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1396 (.I0(\data_in_frame[16] [3]), .I1(\data_in_frame[16] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n59146));
    defparam i1_2_lut_adj_1396.LUT_INIT = 16'h6666;
    SB_LUT4 i15768_3_lut_4_lut (.I0(n8_adj_15), .I1(n58760), .I2(rx_data[0]), 
            .I3(\data_in_frame[1] [0]), .O(n29774));
    defparam i15768_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i4_4_lut_adj_1397 (.I0(\data_in_frame[12] [7]), .I1(n25807), 
            .I2(n4_adj_5072), .I3(n59177), .O(n10_adj_5073));
    defparam i4_4_lut_adj_1397.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1398 (.I0(\data_in_frame[17] [2]), .I1(\data_in_frame[10] [6]), 
            .I2(n10_adj_5073), .I3(\data_in_frame[10] [5]), .O(n59471));
    defparam i1_4_lut_adj_1398.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1399 (.I0(\data_in_frame[13] [2]), .I1(\data_in_frame[13] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n25744));
    defparam i1_2_lut_adj_1399.LUT_INIT = 16'h6666;
    SB_LUT4 i15771_3_lut_4_lut (.I0(n8_adj_15), .I1(n58760), .I2(rx_data[1]), 
            .I3(\data_in_frame[1] [1]), .O(n29777));
    defparam i15771_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i51784_2_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n66935));   // verilog/coms.v(158[12:15])
    defparam i51784_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1_2_lut_adj_1400 (.I0(\data_in_frame[12] [3]), .I1(n59474), 
            .I2(GND_net), .I3(GND_net), .O(n59180));
    defparam i1_2_lut_adj_1400.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1401 (.I0(\data_in_frame[12] [2]), .I1(\data_in_frame[10] [1]), 
            .I2(\data_in_frame[11] [7]), .I3(GND_net), .O(n59080));
    defparam i2_3_lut_adj_1401.LUT_INIT = 16'h9696;
    SB_LUT4 i15774_3_lut_4_lut (.I0(n8_adj_15), .I1(n58760), .I2(rx_data[2]), 
            .I3(\data_in_frame[1] [2]), .O(n29780));
    defparam i15774_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_4_lut_adj_1402 (.I0(\data_in_frame[11] [2]), .I1(\data_in_frame[12] [0]), 
            .I2(\data_in_frame[11] [0]), .I3(\data_in_frame[12] [1]), .O(n63857));
    defparam i1_4_lut_adj_1402.LUT_INIT = 16'h6996;
    SB_LUT4 i51676_2_lut (.I0(\FRAME_MATCHER.i [2]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n66936));   // verilog/coms.v(158[12:15])
    defparam i51676_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1_4_lut_adj_1403 (.I0(\data_in_frame[9] [0]), .I1(\data_in_frame[11] [4]), 
            .I2(\data_in_frame[9] [5]), .I3(\data_in_frame[7] [3]), .O(n63859));
    defparam i1_4_lut_adj_1403.LUT_INIT = 16'h6996;
    SB_LUT4 i1_3_lut_adj_1404 (.I0(n63859), .I1(Kp_23__N_669), .I2(n63857), 
            .I3(GND_net), .O(n63863));
    defparam i1_3_lut_adj_1404.LUT_INIT = 16'h9696;
    SB_LUT4 i1_4_lut_adj_1405 (.I0(n59468), .I1(n59391), .I2(n63863), 
            .I3(n59080), .O(n63869));
    defparam i1_4_lut_adj_1405.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1406 (.I0(n58914), .I1(n58960), .I2(n25818), 
            .I3(n63869), .O(n63875));
    defparam i1_4_lut_adj_1406.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1407 (.I0(n26239), .I1(n61424), .I2(n63875), 
            .I3(n54417), .O(n63881));
    defparam i1_4_lut_adj_1407.LUT_INIT = 16'h9669;
    SB_LUT4 i15777_3_lut_4_lut (.I0(n8_adj_15), .I1(n58760), .I2(rx_data[3]), 
            .I3(\data_in_frame[1] [3]), .O(n29783));
    defparam i15777_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_4_lut_adj_1408 (.I0(n54436), .I1(n63749), .I2(n59180), 
            .I3(n63881), .O(n53460));
    defparam i1_4_lut_adj_1408.LUT_INIT = 16'h6996;
    SB_LUT4 data_in_frame_13__7__I_0_2_lut (.I0(\data_in_frame[13] [7]), .I1(\data_in_frame[13] [6]), 
            .I2(GND_net), .I3(GND_net), .O(Kp_23__N_1271));   // verilog/coms.v(88[17:28])
    defparam data_in_frame_13__7__I_0_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_3_lut_adj_1409 (.I0(\FRAME_MATCHER.state[3] ), .I1(\FRAME_MATCHER.i_31__N_2511 ), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n1_adj_5042));   // verilog/coms.v(148[4] 304[11])
    defparam i1_2_lut_3_lut_adj_1409.LUT_INIT = 16'h1010;
    SB_LUT4 i1_3_lut_adj_1410 (.I0(n59284), .I1(n58870), .I2(\data_in_frame[13] [2]), 
            .I3(GND_net), .O(n53832));   // verilog/coms.v(99[12:25])
    defparam i1_3_lut_adj_1410.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1411 (.I0(n25987), .I1(\data_in_frame[12] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n58960));
    defparam i1_2_lut_adj_1411.LUT_INIT = 16'h6666;
    SB_LUT4 i51512_2_lut (.I0(\FRAME_MATCHER.i[3] ), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n66937));   // verilog/coms.v(158[12:15])
    defparam i51512_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 data_in_frame_12__7__I_0_4035_2_lut (.I0(\data_in_frame[12] [7]), 
            .I1(\data_in_frame[12] [6]), .I2(GND_net), .I3(GND_net), .O(Kp_23__N_669));   // verilog/coms.v(74[16:27])
    defparam data_in_frame_12__7__I_0_4035_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1412 (.I0(\data_in_frame[14] [7]), .I1(n26435), 
            .I2(GND_net), .I3(GND_net), .O(n59177));
    defparam i1_2_lut_adj_1412.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1413 (.I0(\data_in_frame[15] [2]), .I1(n25987), 
            .I2(Kp_23__N_669), .I3(n6_adj_5074), .O(n59278));
    defparam i4_4_lut_adj_1413.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1414 (.I0(\data_in_frame[15] [1]), .I1(\data_in_frame[17] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n63629));
    defparam i1_2_lut_adj_1414.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1415 (.I0(n59156), .I1(n59278), .I2(n59177), 
            .I3(n63629), .O(n63635));
    defparam i1_4_lut_adj_1415.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1416 (.I0(n53832), .I1(n54511), .I2(n58870), 
            .I3(n63635), .O(n54452));
    defparam i1_4_lut_adj_1416.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1417 (.I0(n53570), .I1(\data_in_frame[15] [3]), 
            .I2(\data_in_frame[17] [4]), .I3(n59278), .O(n61410));
    defparam i3_4_lut_adj_1417.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1418 (.I0(\data_out_frame[12] [3]), .I1(n1513), 
            .I2(\data_out_frame[12] [2]), .I3(n1510), .O(n59055));   // verilog/coms.v(77[16:43])
    defparam i1_2_lut_3_lut_4_lut_adj_1418.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1419 (.I0(\data_in_frame[8] [1]), .I1(\data_in_frame[8] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n59412));   // verilog/coms.v(74[16:27])
    defparam i1_2_lut_adj_1419.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1420 (.I0(\data_in_frame[10] [2]), .I1(n58947), 
            .I2(n59271), .I3(n6_adj_5075), .O(n54155));
    defparam i4_4_lut_adj_1420.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1421 (.I0(n59412), .I1(n59000), .I2(\data_in_frame[10] [3]), 
            .I3(n59430), .O(n10_adj_5076));   // verilog/coms.v(79[16:43])
    defparam i4_4_lut_adj_1421.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_1422 (.I0(n59320), .I1(n10_adj_5076), .I2(n58799), 
            .I3(GND_net), .O(n26438));   // verilog/coms.v(79[16:43])
    defparam i5_3_lut_adj_1422.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1423 (.I0(\data_in_frame[14] [7]), .I1(\data_in_frame[15] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n59174));
    defparam i1_2_lut_adj_1423.LUT_INIT = 16'h6666;
    SB_LUT4 i51513_2_lut (.I0(\FRAME_MATCHER.i[4] ), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n66938));   // verilog/coms.v(158[12:15])
    defparam i51513_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1_2_lut_adj_1424 (.I0(\data_in_frame[10] [5]), .I1(n58836), 
            .I2(GND_net), .I3(GND_net), .O(n26639));   // verilog/coms.v(74[16:27])
    defparam i1_2_lut_adj_1424.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1425 (.I0(\data_in_frame[9] [7]), .I1(n26774), 
            .I2(n25843), .I3(n54002), .O(n54417));
    defparam i3_4_lut_adj_1425.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1426 (.I0(n54417), .I1(\data_in_frame[10] [1]), 
            .I2(\data_in_frame[12] [3]), .I3(GND_net), .O(n59199));
    defparam i2_3_lut_adj_1426.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1427 (.I0(\data_in_frame[10] [4]), .I1(n3_adj_5077), 
            .I2(n4_adj_5072), .I3(GND_net), .O(n25987));   // verilog/coms.v(77[16:43])
    defparam i2_3_lut_adj_1427.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1428 (.I0(n26438), .I1(n54155), .I2(GND_net), 
            .I3(GND_net), .O(n54436));
    defparam i1_2_lut_adj_1428.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1429 (.I0(n59199), .I1(\data_in_frame[16] [7]), 
            .I2(\data_in_frame[12] [5]), .I3(n59394), .O(n10_adj_5078));
    defparam i4_4_lut_adj_1429.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1430 (.I0(n59394), .I1(\data_in_frame[14] [7]), 
            .I2(\data_in_frame[15] [1]), .I3(\data_in_frame[14] [6]), .O(n14_adj_5079));   // verilog/coms.v(74[16:27])
    defparam i6_4_lut_adj_1430.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1431 (.I0(n59471), .I1(n14_adj_5079), .I2(n10_adj_5080), 
            .I3(\data_in_frame[15] [0]), .O(n59143));   // verilog/coms.v(74[16:27])
    defparam i7_4_lut_adj_1431.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1432 (.I0(\data_in_frame[17] [1]), .I1(n59143), 
            .I2(\data_in_frame[19] [3]), .I3(n54473), .O(n53511));
    defparam i3_4_lut_adj_1432.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1433 (.I0(\data_in_frame[21] [5]), .I1(\data_in_frame[19] [5]), 
            .I2(n61410), .I3(n54452), .O(n59033));
    defparam i3_4_lut_adj_1433.LUT_INIT = 16'h9669;
    SB_LUT4 i3_4_lut_adj_1434 (.I0(n58914), .I1(n25661), .I2(n26411), 
            .I3(\data_in_frame[14] [0]), .O(n59316));
    defparam i3_4_lut_adj_1434.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1435 (.I0(\data_in_frame[9] [3]), .I1(n59097), 
            .I2(\data_in_frame[11] [4]), .I3(GND_net), .O(n25925));   // verilog/coms.v(76[16:42])
    defparam i2_3_lut_adj_1435.LUT_INIT = 16'h9696;
    SB_LUT4 data_in_frame_17__7__I_0_4040_2_lut (.I0(\data_in_frame[17] [7]), 
            .I1(\data_in_frame[17] [6]), .I2(GND_net), .I3(GND_net), .O(Kp_23__N_1389));   // verilog/coms.v(73[16:27])
    defparam data_in_frame_17__7__I_0_4040_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1436 (.I0(\data_in_frame[13] [5]), .I1(\data_in_frame[15] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n59060));   // verilog/coms.v(78[16:43])
    defparam i1_2_lut_adj_1436.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1437 (.I0(\data_in_frame[16] [1]), .I1(\data_in_frame[13] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n59140));
    defparam i1_2_lut_adj_1437.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1438 (.I0(\data_in_frame[8] [6]), .I1(\data_in_frame[13] [4]), 
            .I2(n26633), .I3(n6_adj_5081), .O(n59362));   // verilog/coms.v(78[16:43])
    defparam i4_4_lut_adj_1438.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1439 (.I0(\data_in_frame[13] [6]), .I1(n59316), 
            .I2(GND_net), .I3(GND_net), .O(n59439));
    defparam i1_2_lut_adj_1439.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1440 (.I0(\data_in_frame[20] [2]), .I1(n25925), 
            .I2(n59362), .I3(\data_in_frame[18] [0]), .O(n59371));   // verilog/coms.v(78[16:43])
    defparam i3_4_lut_adj_1440.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1441 (.I0(\data_in_frame[16] [0]), .I1(n59439), 
            .I2(n59362), .I3(n59140), .O(n23833));   // verilog/coms.v(88[17:63])
    defparam i3_4_lut_adj_1441.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1442 (.I0(n25751), .I1(\data_in_frame[5] [1]), 
            .I2(n58901), .I3(n6_adj_5012), .O(n61424));   // verilog/coms.v(88[17:70])
    defparam i4_4_lut_adj_1442.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1443 (.I0(\data_in_frame[5] [2]), .I1(\data_in_frame[7] [4]), 
            .I2(n59003), .I3(n6_adj_5082), .O(n59397));
    defparam i4_4_lut_adj_1443.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1444 (.I0(n26608), .I1(n59397), .I2(GND_net), 
            .I3(GND_net), .O(n23922));
    defparam i1_2_lut_adj_1444.LUT_INIT = 16'h6666;
    SB_LUT4 i54320_2_lut (.I0(n61424), .I1(\data_in_frame[7] [3]), .I2(GND_net), 
            .I3(GND_net), .O(n70014));   // verilog/coms.v(99[12:25])
    defparam i54320_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i51514_2_lut (.I0(\FRAME_MATCHER.i[5] ), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n66939));   // verilog/coms.v(158[12:15])
    defparam i51514_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1_2_lut_adj_1445 (.I0(\data_in_frame[1] [5]), .I1(\data_in_frame[7]_c [7]), 
            .I2(GND_net), .I3(GND_net), .O(n58799));   // verilog/coms.v(78[16:27])
    defparam i1_2_lut_adj_1445.LUT_INIT = 16'h6666;
    SB_LUT4 i15783_3_lut_4_lut (.I0(n8_adj_15), .I1(n58760), .I2(rx_data[4]), 
            .I3(\data_in_frame[1] [4]), .O(n29789));
    defparam i15783_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_4_lut_adj_1446 (.I0(n26239), .I1(n58836), .I2(n3_adj_5077), 
            .I3(\data_in_frame[8] [7]), .O(n63647));
    defparam i1_4_lut_adj_1446.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1447 (.I0(n59487), .I1(n26680), .I2(n59271), 
            .I3(n63647), .O(n63653));
    defparam i1_4_lut_adj_1447.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1448 (.I0(n26426), .I1(n54404), .I2(n59459), 
            .I3(n63653), .O(n61299));
    defparam i1_4_lut_adj_1448.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1449 (.I0(\data_in_frame[9] [4]), .I1(\data_in_frame[9] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n25661));
    defparam i1_2_lut_adj_1449.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1450 (.I0(\data_in_frame[9] [1]), .I1(\data_in_frame[9] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n26219));   // verilog/coms.v(88[17:63])
    defparam i1_2_lut_adj_1450.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1451 (.I0(\data_in_frame[9] [7]), .I1(\data_in_frame[9] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n58894));   // verilog/coms.v(88[17:63])
    defparam i1_2_lut_adj_1451.LUT_INIT = 16'h6666;
    SB_LUT4 i1_3_lut_adj_1452 (.I0(n25807), .I1(n61299), .I2(\data_in_frame[9] [0]), 
            .I3(GND_net), .O(n54520));
    defparam i1_3_lut_adj_1452.LUT_INIT = 16'h6969;
    SB_LUT4 i3_4_lut_adj_1453 (.I0(\data_in_frame[9] [3]), .I1(n58894), 
            .I2(n26219), .I3(n25661), .O(Kp_23__N_1080));   // verilog/coms.v(88[17:63])
    defparam i3_4_lut_adj_1453.LUT_INIT = 16'h6996;
    SB_LUT4 i15786_3_lut_4_lut (.I0(n8_adj_15), .I1(n58760), .I2(rx_data[5]), 
            .I3(\data_in_frame[1] [5]), .O(n29792));
    defparam i15786_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i51515_2_lut (.I0(\FRAME_MATCHER.i [6]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n66940));   // verilog/coms.v(158[12:15])
    defparam i51515_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1_3_lut_adj_1454 (.I0(n61299), .I1(\data_in_frame[10] [7]), 
            .I2(\data_in_frame[11] [1]), .I3(GND_net), .O(n63749));
    defparam i1_3_lut_adj_1454.LUT_INIT = 16'h6969;
    SB_LUT4 i4_4_lut_adj_1455 (.I0(n59302), .I1(n59247), .I2(\data_in_frame[8] [7]), 
            .I3(n59391), .O(n10_adj_5083));   // verilog/coms.v(80[16:43])
    defparam i4_4_lut_adj_1455.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1456 (.I0(n53570), .I1(n25906), .I2(GND_net), 
            .I3(GND_net), .O(n59156));
    defparam i1_2_lut_adj_1456.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1457 (.I0(\data_in_frame[15] [4]), .I1(\data_in_frame[13] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_5084));
    defparam i1_2_lut_adj_1457.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1458 (.I0(n58848), .I1(\data_in_frame[9] [0]), 
            .I2(n59165), .I3(n6_adj_5084), .O(n60961));
    defparam i4_4_lut_adj_1458.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1459 (.I0(\data_in_frame[15] [5]), .I1(n54511), 
            .I2(n60961), .I3(GND_net), .O(n25724));
    defparam i2_3_lut_adj_1459.LUT_INIT = 16'h6969;
    SB_LUT4 i2_3_lut_adj_1460 (.I0(n25724), .I1(\data_in_frame[17] [6]), 
            .I2(\data_in_frame[20] [0]), .I3(GND_net), .O(n59103));
    defparam i2_3_lut_adj_1460.LUT_INIT = 16'h9696;
    SB_LUT4 i51517_2_lut (.I0(\FRAME_MATCHER.i [7]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n66941));   // verilog/coms.v(158[12:15])
    defparam i51517_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i15789_3_lut_4_lut (.I0(n8_adj_15), .I1(n58760), .I2(rx_data[6]), 
            .I3(\data_in_frame[1] [6]), .O(n29795));
    defparam i15789_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15792_3_lut_4_lut (.I0(n8_adj_15), .I1(n58760), .I2(rx_data[7]), 
            .I3(\data_in_frame[1] [7]), .O(n29798));
    defparam i15792_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i4_4_lut_adj_1461 (.I0(n26755), .I1(\data_in_frame[22] [1]), 
            .I2(\data_in_frame[21] [7]), .I3(n59103), .O(n10_adj_5085));
    defparam i4_4_lut_adj_1461.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1462 (.I0(\data_in_frame[21] [6]), .I1(n59033), 
            .I2(n53511), .I3(\data_in_frame[23] [7]), .O(n60903));
    defparam i3_4_lut_adj_1462.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1463 (.I0(n59086), .I1(\data_in_frame[18] [2]), 
            .I2(n23833), .I3(n59371), .O(n10_adj_5086));
    defparam i4_4_lut_adj_1463.LUT_INIT = 16'h6996;
    SB_LUT4 i48366_4_lut (.I0(\data_in_frame[22] [4]), .I1(n53031), .I2(n10_adj_5086), 
            .I3(\data_in_frame[20] [3]), .O(n64050));
    defparam i48366_4_lut.LUT_INIT = 16'hedde;
    SB_LUT4 i1_2_lut_3_lut_3_lut_adj_1464 (.I0(n40817), .I1(n43501), .I2(reset), 
            .I3(GND_net), .O(n40820));   // verilog/coms.v(156[9:50])
    defparam i1_2_lut_3_lut_3_lut_adj_1464.LUT_INIT = 16'h0808;
    SB_LUT4 i1_2_lut_3_lut_adj_1465 (.I0(\data_in_frame[2] [3]), .I1(\data_in_frame[0]_c [2]), 
            .I2(\data_in_frame[0] [1]), .I3(GND_net), .O(n26288));   // verilog/coms.v(78[16:43])
    defparam i1_2_lut_3_lut_adj_1465.LUT_INIT = 16'h9696;
    SB_LUT4 i54324_2_lut_3_lut_4_lut (.I0(n26608), .I1(n59397), .I2(n23926), 
            .I3(\data_in_frame[9] [6]), .O(n70018));   // verilog/coms.v(99[12:25])
    defparam i54324_2_lut_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i23377_3_lut (.I0(n375), .I1(n455), .I2(n11597), .I3(GND_net), 
            .O(n37330));
    defparam i23377_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_adj_1466 (.I0(\data_in_frame[0][3] ), .I1(\data_in_frame[0]_c [2]), 
            .I2(\data_in_frame[2] [4]), .I3(GND_net), .O(n25758));   // verilog/coms.v(169[9:87])
    defparam i1_2_lut_3_lut_adj_1466.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1467 (.I0(\FRAME_MATCHER.i[3] ), .I1(\FRAME_MATCHER.i[4] ), 
            .I2(\FRAME_MATCHER.i[5] ), .I3(n3468), .O(n58731));   // verilog/coms.v(157[7:23])
    defparam i1_2_lut_3_lut_4_lut_adj_1467.LUT_INIT = 16'hfdff;
    SB_LUT4 i1_4_lut_adj_1468 (.I0(\data_in_frame[23] [5]), .I1(n64050), 
            .I2(n58925), .I3(n53511), .O(n63719));
    defparam i1_4_lut_adj_1468.LUT_INIT = 16'h2112;
    SB_LUT4 i3_4_lut_adj_1469 (.I0(\data_in_frame[20] [4]), .I1(n59077), 
            .I2(n59380), .I3(\data_in_frame[22] [6]), .O(n61271));
    defparam i3_4_lut_adj_1469.LUT_INIT = 16'h9669;
    SB_LUT4 i3_3_lut_adj_1470 (.I0(\data_in_frame[21] [4]), .I1(n54588), 
            .I2(n59106), .I3(GND_net), .O(n8_adj_5087));
    defparam i3_3_lut_adj_1470.LUT_INIT = 16'h6969;
    SB_LUT4 i1_4_lut_adj_1471 (.I0(\data_in_frame[22] [5]), .I1(n61271), 
            .I2(n59046), .I3(n63719), .O(n63723));
    defparam i1_4_lut_adj_1471.LUT_INIT = 16'h8400;
    SB_LUT4 i1_4_lut_adj_1472 (.I0(\data_in_frame[23] [6]), .I1(n63723), 
            .I2(n8_adj_5087), .I3(\data_in_frame[21] [5]), .O(n63725));
    defparam i1_4_lut_adj_1472.LUT_INIT = 16'h4884;
    SB_LUT4 i2_3_lut_adj_1473 (.I0(\data_in_frame[21] [2]), .I1(\data_in_frame[23] [3]), 
            .I2(\data_in_frame[21] [1]), .I3(GND_net), .O(n6_adj_5088));
    defparam i2_3_lut_adj_1473.LUT_INIT = 16'h9696;
    SB_LUT4 i1_4_lut_adj_1474 (.I0(n5_adj_5064), .I1(n63725), .I2(\data_in_frame[21] [2]), 
            .I3(n25953), .O(n63727));
    defparam i1_4_lut_adj_1474.LUT_INIT = 16'h8448;
    SB_LUT4 i3_3_lut_adj_1475 (.I0(\data_in_frame[23] [1]), .I1(n26689), 
            .I2(Kp_23__N_1607), .I3(GND_net), .O(n8_adj_5089));
    defparam i3_3_lut_adj_1475.LUT_INIT = 16'h9696;
    SB_LUT4 i1_4_lut_adj_1476 (.I0(n54572), .I1(n63727), .I2(n6_adj_5088), 
            .I3(Kp_23__N_1607), .O(n63729));
    defparam i1_4_lut_adj_1476.LUT_INIT = 16'h4884;
    SB_LUT4 i1_4_lut_adj_1477 (.I0(n63729), .I1(n54572), .I2(n8_adj_5089), 
            .I3(n54460), .O(n63731));
    defparam i1_4_lut_adj_1477.LUT_INIT = 16'h8228;
    SB_LUT4 i1_4_lut_adj_1478 (.I0(n61410), .I1(\data_in_frame[19] [6]), 
            .I2(\data_in_frame[20] [1]), .I3(\data_in_frame[22] [2]), .O(n63837));
    defparam i1_4_lut_adj_1478.LUT_INIT = 16'h9669;
    SB_LUT4 i1_3_lut_adj_1479 (.I0(\data_in_frame[22] [0]), .I1(\data_in_frame[21] [7]), 
            .I2(\data_in_frame[21] [6]), .I3(GND_net), .O(n5_adj_5090));
    defparam i1_3_lut_adj_1479.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1480 (.I0(\data_in_frame[18] [1]), .I1(\data_in_frame[22] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n63825));
    defparam i1_2_lut_adj_1480.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_4_lut_adj_1481 (.I0(\data_in_frame[2] [3]), .I1(n58789), 
            .I2(\data_in_frame[0][3] ), .I3(n58815), .O(n58876));   // verilog/coms.v(78[16:43])
    defparam i1_2_lut_4_lut_adj_1481.LUT_INIT = 16'h6996;
    SB_LUT4 i48364_4_lut (.I0(\data_in_frame[19] [7]), .I1(n60903), .I2(n10_adj_5085), 
            .I3(\data_in_frame[19] [5]), .O(n64048));
    defparam i48364_4_lut.LUT_INIT = 16'hedde;
    SB_LUT4 i51518_2_lut (.I0(\FRAME_MATCHER.i [8]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n66942));   // verilog/coms.v(158[12:15])
    defparam i51518_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1_4_lut_adj_1482 (.I0(n54513), .I1(n59018), .I2(n59086), 
            .I3(n63825), .O(n63831));
    defparam i1_4_lut_adj_1482.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1483 (.I0(n5_adj_5090), .I1(\data_in_frame[19] [6]), 
            .I2(Kp_23__N_1551), .I3(n54588), .O(n61285));
    defparam i3_4_lut_adj_1483.LUT_INIT = 16'h9669;
    SB_LUT4 i1_4_lut_adj_1484 (.I0(\data_in_frame[21] [1]), .I1(n63731), 
            .I2(\data_in_frame[23] [2]), .I3(n54116), .O(n63733));
    defparam i1_4_lut_adj_1484.LUT_INIT = 16'h8448;
    SB_LUT4 i1_4_lut_adj_1485 (.I0(n59183), .I1(n54447), .I2(n54630), 
            .I3(n63801), .O(n63807));
    defparam i1_4_lut_adj_1485.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1486 (.I0(n54513), .I1(n25112), .I2(n59103), 
            .I3(n63837), .O(n63843));
    defparam i1_4_lut_adj_1486.LUT_INIT = 16'h9669;
    SB_LUT4 i1_4_lut_adj_1487 (.I0(n61285), .I1(n63831), .I2(n64048), 
            .I3(n61398), .O(n61908));
    defparam i1_4_lut_adj_1487.LUT_INIT = 16'h0802;
    SB_LUT4 i1_4_lut_adj_1488 (.I0(\data_in_frame[23] [0]), .I1(n63807), 
            .I2(n63733), .I3(n59226), .O(n63739));
    defparam i1_4_lut_adj_1488.LUT_INIT = 16'h8010;
    SB_LUT4 i1_4_lut_adj_1489 (.I0(n63739), .I1(n61908), .I2(n63843), 
            .I3(n61398), .O(n37));
    defparam i1_4_lut_adj_1489.LUT_INIT = 16'h0880;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1490 (.I0(\data_in_frame[9] [2]), .I1(n58792), 
            .I2(n59247), .I3(n26411), .O(n59097));   // verilog/coms.v(76[16:42])
    defparam i1_2_lut_3_lut_4_lut_adj_1490.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1491 (.I0(\data_in_frame[5] [0]), .I1(n26288), 
            .I2(n25758), .I3(GND_net), .O(n26282));   // verilog/coms.v(78[16:43])
    defparam i1_2_lut_3_lut_adj_1491.LUT_INIT = 16'h9696;
    SB_LUT4 equal_300_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i[0] ), .I3(GND_net), .O(n8_adj_15));   // verilog/coms.v(158[12:15])
    defparam equal_300_i8_2_lut_3_lut.LUT_INIT = 16'hefef;
    SB_LUT4 equal_293_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i[0] ), .I3(GND_net), .O(n8_adj_12));   // verilog/coms.v(158[12:15])
    defparam equal_293_i8_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_2_lut_3_lut_adj_1492 (.I0(\data_in_frame[1] [6]), .I1(\data_in_frame[1] [5]), 
            .I2(\data_in_frame[1] [7]), .I3(GND_net), .O(n25786));   // verilog/coms.v(81[16:27])
    defparam i1_2_lut_3_lut_adj_1492.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1493 (.I0(\data_in_frame[1] [3]), .I1(\data_in_frame[1] [2]), 
            .I2(\data_in_frame[3] [4]), .I3(n58947), .O(n23926));
    defparam i1_2_lut_3_lut_4_lut_adj_1493.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1494 (.I0(\data_in_frame[2] [1]), .I1(\data_in_frame[4] [2]), 
            .I2(\data_in_frame[4] [1]), .I3(\data_in_frame[3] [7]), .O(n59256));   // verilog/coms.v(73[16:69])
    defparam i1_2_lut_4_lut_adj_1494.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1495 (.I0(n26288), .I1(\data_in_frame[6] [6]), 
            .I2(\data_in_frame[4] [6]), .I3(\data_in_frame[7] [0]), .O(n58792));   // verilog/coms.v(74[16:27])
    defparam i3_4_lut_adj_1495.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1496 (.I0(n58792), .I1(n59247), .I2(GND_net), 
            .I3(GND_net), .O(n26251));   // verilog/coms.v(74[16:27])
    defparam i1_2_lut_adj_1496.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1497 (.I0(\data_in_frame[5] [0]), .I1(n59007), 
            .I2(\data_in_frame[7] [2]), .I3(GND_net), .O(n26411));
    defparam i2_3_lut_adj_1497.LUT_INIT = 16'h9696;
    SB_LUT4 i51564_2_lut (.I0(\FRAME_MATCHER.i [9]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n66944));   // verilog/coms.v(158[12:15])
    defparam i51564_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1_3_lut_adj_1498 (.I0(n59290), .I1(n54113), .I2(\data_in_frame[6] [0]), 
            .I3(GND_net), .O(n59134));   // verilog/coms.v(78[16:43])
    defparam i1_3_lut_adj_1498.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1499 (.I0(\data_in_frame[1] [6]), .I1(\data_in_frame[4] [0]), 
            .I2(\data_in_frame[3] [7]), .I3(\data_in_frame[6] [1]), .O(n59320));   // verilog/coms.v(81[16:27])
    defparam i2_3_lut_4_lut_adj_1499.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1500 (.I0(\data_in_frame[6] [4]), .I1(n59215), 
            .I2(\data_in_frame[4] [2]), .I3(\data_in_frame[1] [7]), .O(n10_adj_5091));   // verilog/coms.v(81[16:27])
    defparam i4_4_lut_adj_1500.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_1501 (.I0(\data_in_frame[1] [6]), .I1(n10_adj_5091), 
            .I2(n26316), .I3(GND_net), .O(n58818));   // verilog/coms.v(81[16:27])
    defparam i5_3_lut_adj_1501.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1502 (.I0(n58818), .I1(n58824), .I2(\data_in_frame[8] [5]), 
            .I3(GND_net), .O(n25807));   // verilog/coms.v(78[16:43])
    defparam i2_3_lut_adj_1502.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1503 (.I0(\data_in_frame[1] [3]), .I1(\data_in_frame[1] [2]), 
            .I2(\data_in_frame[3] [4]), .I3(GND_net), .O(n25860));   // verilog/coms.v(79[16:43])
    defparam i1_2_lut_3_lut_adj_1503.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1504 (.I0(n771), .I1(\FRAME_MATCHER.i_31__N_2508 ), 
            .I2(n25463), .I3(\FRAME_MATCHER.i_31__N_2507 ), .O(n63955));   // verilog/coms.v(148[4] 304[11])
    defparam i1_2_lut_3_lut_4_lut_adj_1504.LUT_INIT = 16'hfff4;
    SB_LUT4 i51570_2_lut (.I0(\FRAME_MATCHER.i [10]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n66951));   // verilog/coms.v(158[12:15])
    defparam i51570_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1_2_lut_adj_1505 (.I0(\data_in_frame[3][6] ), .I1(\data_in_frame[6] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n26343));   // verilog/coms.v(78[16:27])
    defparam i1_2_lut_adj_1505.LUT_INIT = 16'h6666;
    SB_LUT4 i1_3_lut_4_lut (.I0(\data_in_frame[20] [6]), .I1(\data_in_frame[18] [5]), 
            .I2(\data_in_frame[20] [5]), .I3(\data_in_frame[22] [7]), .O(n63801));
    defparam i1_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1506 (.I0(n61410), .I1(n53713), .I2(n54452), 
            .I3(GND_net), .O(n26755));
    defparam i1_2_lut_3_lut_adj_1506.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1507 (.I0(\data_in_frame[1] [7]), .I1(\data_in_frame[0][0] ), 
            .I2(GND_net), .I3(GND_net), .O(n59109));   // verilog/coms.v(73[16:69])
    defparam i1_2_lut_adj_1507.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_4_lut_adj_1508 (.I0(\data_in_frame[11] [2]), .I1(n58792), 
            .I2(n59247), .I3(\data_in_frame[9] [1]), .O(n58848));   // verilog/coms.v(74[16:27])
    defparam i2_3_lut_4_lut_adj_1508.LUT_INIT = 16'h6996;
    SB_LUT4 i51549_2_lut (.I0(\FRAME_MATCHER.i [11]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n66952));   // verilog/coms.v(158[12:15])
    defparam i51549_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i3_4_lut_adj_1509 (.I0(\data_in_frame[4] [3]), .I1(n59109), 
            .I2(n25815), .I3(\data_in_frame[4] [4]), .O(Kp_23__N_878));   // verilog/coms.v(73[16:69])
    defparam i3_4_lut_adj_1509.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1510 (.I0(\data_in_frame[4] [5]), .I1(Kp_23__N_878), 
            .I2(GND_net), .I3(GND_net), .O(n59064));   // verilog/coms.v(80[16:43])
    defparam i1_2_lut_adj_1510.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_3_lut_adj_1511 (.I0(n25807), .I1(Kp_23__N_974), .I2(\data_in_frame[8] [6]), 
            .I3(GND_net), .O(n59487));
    defparam i1_2_lut_3_lut_adj_1511.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1512 (.I0(n58792), .I1(n59247), .I2(n26411), 
            .I3(GND_net), .O(n26680));   // verilog/coms.v(76[16:42])
    defparam i1_2_lut_3_lut_adj_1512.LUT_INIT = 16'h9696;
    SB_LUT4 i1_3_lut_4_lut_adj_1513 (.I0(n771), .I1(\FRAME_MATCHER.i_31__N_2508 ), 
            .I2(n1951), .I3(n1954), .O(n25468));   // verilog/coms.v(148[4] 304[11])
    defparam i1_3_lut_4_lut_adj_1513.LUT_INIT = 16'h4000;
    SB_LUT4 i1_2_lut_adj_1514 (.I0(\data_in_frame[1] [6]), .I1(\data_in_frame[4] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n25869));   // verilog/coms.v(81[16:27])
    defparam i1_2_lut_adj_1514.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_4_lut_adj_1515 (.I0(n1951), .I1(n4452), .I2(n1954), 
            .I3(n1957), .O(n60750));   // verilog/coms.v(145[4] 147[7])
    defparam i2_3_lut_4_lut_adj_1515.LUT_INIT = 16'h2000;
    SB_LUT4 i3_4_lut_adj_1516 (.I0(\data_in_frame[6] [3]), .I1(\data_in_frame[0][0] ), 
            .I2(n59256), .I3(n25786), .O(n58824));   // verilog/coms.v(73[16:69])
    defparam i3_4_lut_adj_1516.LUT_INIT = 16'h6996;
    SB_LUT4 i51550_2_lut (.I0(\FRAME_MATCHER.i [12]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n66953));   // verilog/coms.v(158[12:15])
    defparam i51550_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i5_4_lut_adj_1517 (.I0(\data_in_frame[4] [1]), .I1(n58827), 
            .I2(\data_in_frame[1] [4]), .I3(\data_in_frame[3][6] ), .O(n12_adj_5092));   // verilog/coms.v(81[16:27])
    defparam i5_4_lut_adj_1517.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1518 (.I0(n25869), .I1(n12_adj_5092), .I2(\data_in_frame[6] [2]), 
            .I3(\data_in_frame[2] [0]), .O(n58922));   // verilog/coms.v(81[16:27])
    defparam i6_4_lut_adj_1518.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1519 (.I0(\data_in_frame[8] [1]), .I1(n58812), 
            .I2(n59259), .I3(n26343), .O(n59271));
    defparam i1_2_lut_4_lut_adj_1519.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1520 (.I0(n25860), .I1(n26343), .I2(\data_in_frame[1] [4]), 
            .I3(n6_adj_5093), .O(n26774));   // verilog/coms.v(79[16:43])
    defparam i4_4_lut_adj_1520.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1521 (.I0(\data_in_frame[8] [2]), .I1(n26774), 
            .I2(n25878), .I3(GND_net), .O(n3_adj_5077));   // verilog/coms.v(79[16:43])
    defparam i2_3_lut_adj_1521.LUT_INIT = 16'h9696;
    SB_LUT4 i2_2_lut_adj_1522 (.I0(\data_in_frame[8] [7]), .I1(Kp_23__N_993), 
            .I2(GND_net), .I3(GND_net), .O(n7_adj_5094));
    defparam i2_2_lut_adj_1522.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_3_lut_adj_1523 (.I0(n26608), .I1(n59397), .I2(n23926), 
            .I3(GND_net), .O(n26426));
    defparam i1_2_lut_3_lut_adj_1523.LUT_INIT = 16'h9696;
    SB_LUT4 i2_4_lut_4_lut (.I0(n1951), .I1(n4452), .I2(n63955), .I3(\FRAME_MATCHER.i_31__N_2514 ), 
            .O(n61412));   // verilog/coms.v(145[4] 147[7])
    defparam i2_4_lut_4_lut.LUT_INIT = 16'ha2a0;
    SB_LUT4 i1_2_lut_3_lut_adj_1524 (.I0(n61424), .I1(\data_in_frame[7] [3]), 
            .I2(Kp_23__N_993), .I3(GND_net), .O(n59459));
    defparam i1_2_lut_3_lut_adj_1524.LUT_INIT = 16'h9696;
    SB_LUT4 i4_4_lut_adj_1525 (.I0(\data_in_frame[7] [5]), .I1(\data_in_frame[5] [4]), 
            .I2(n59003), .I3(n6_adj_5095), .O(n54002));
    defparam i4_4_lut_adj_1525.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1526 (.I0(\data_in_frame[2] [0]), .I1(\data_in_frame[4] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n59215));   // verilog/coms.v(81[16:27])
    defparam i1_2_lut_adj_1526.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1527 (.I0(\data_in_frame[4] [2]), .I1(\data_in_frame[4] [1]), 
            .I2(\data_in_frame[3] [7]), .I3(GND_net), .O(n58805));   // verilog/coms.v(73[16:69])
    defparam i2_3_lut_adj_1527.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1528 (.I0(\data_in_frame[4] [7]), .I1(n26608), 
            .I2(GND_net), .I3(GND_net), .O(n58901));   // verilog/coms.v(80[16:43])
    defparam i1_2_lut_adj_1528.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_4_lut_adj_1529 (.I0(\data_in_frame[5] [4]), .I1(n59202), 
            .I2(\data_in_frame[5] [5]), .I3(\data_in_frame[7]_c [6]), .O(n58947));
    defparam i1_2_lut_4_lut_adj_1529.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1530 (.I0(\data_in_frame[0][6] ), .I1(n35423), 
            .I2(\data_in_frame[3] [0]), .I3(n59202), .O(n6_adj_5082));
    defparam i1_2_lut_4_lut_adj_1530.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1531 (.I0(n26282), .I1(n58901), .I2(\data_in_frame[7] [1]), 
            .I3(GND_net), .O(n59302));   // verilog/coms.v(73[16:27])
    defparam i2_3_lut_adj_1531.LUT_INIT = 16'h9696;
    SB_LUT4 i51954_2_lut (.I0(\FRAME_MATCHER.i [13]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n66955));   // verilog/coms.v(158[12:15])
    defparam i51954_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1_2_lut_3_lut_adj_1532 (.I0(\data_in_frame[9] [1]), .I1(\data_in_frame[9] [2]), 
            .I2(\data_in_frame[11] [3]), .I3(GND_net), .O(n59391));
    defparam i1_2_lut_3_lut_adj_1532.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_4_lut_adj_1533 (.I0(\data_in_frame[8] [4]), .I1(n58824), 
            .I2(n58922), .I3(\data_in_frame[10] [6]), .O(n59468));
    defparam i1_2_lut_4_lut_adj_1533.LUT_INIT = 16'h6996;
    SB_LUT4 i1_3_lut_adj_1534 (.I0(\data_in_frame[0][6] ), .I1(n35423), 
            .I2(\data_in_frame[3] [0]), .I3(GND_net), .O(n26544));
    defparam i1_3_lut_adj_1534.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1535 (.I0(\data_in_frame[2] [7]), .I1(n35423), 
            .I2(GND_net), .I3(GND_net), .O(n58997));
    defparam i1_2_lut_adj_1535.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1536 (.I0(\data_in_frame[1] [5]), .I1(\data_in_frame[1] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n58827));   // verilog/coms.v(81[16:27])
    defparam i1_2_lut_adj_1536.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_3_lut_adj_1537 (.I0(\data_in_frame[17] [7]), .I1(\data_in_frame[17] [6]), 
            .I2(n60961), .I3(GND_net), .O(n59086));
    defparam i1_2_lut_3_lut_adj_1537.LUT_INIT = 16'h6969;
    SB_LUT4 i1_2_lut_4_lut_adj_1538 (.I0(\data_in_frame[11] [2]), .I1(n26251), 
            .I2(\data_in_frame[9] [1]), .I3(n59060), .O(n6_adj_5081));   // verilog/coms.v(78[16:43])
    defparam i1_2_lut_4_lut_adj_1538.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1539 (.I0(\data_in_frame[9] [0]), .I1(\data_in_frame[6] [5]), 
            .I2(Kp_23__N_878), .I3(n58818), .O(n26633));
    defparam i1_2_lut_4_lut_adj_1539.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1540 (.I0(\FRAME_MATCHER.i[4] ), .I1(\FRAME_MATCHER.i[3] ), 
            .I2(\FRAME_MATCHER.i[5] ), .I3(GND_net), .O(n40817));   // verilog/coms.v(158[12:15])
    defparam i1_2_lut_3_lut_adj_1540.LUT_INIT = 16'h0202;
    SB_LUT4 i1_4_lut_adj_1541 (.I0(\data_in_frame[4] [6]), .I1(\data_in_frame[2] [5]), 
            .I2(\data_in_frame[5] [1]), .I3(\data_in_frame[2] [6]), .O(n63755));   // verilog/coms.v(169[9:87])
    defparam i1_4_lut_adj_1541.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1542 (.I0(n58997), .I1(n26544), .I2(n58815), 
            .I3(n63755), .O(n59007));   // verilog/coms.v(169[9:87])
    defparam i1_4_lut_adj_1542.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1543 (.I0(\data_in_frame[3] [2]), .I1(\data_in_frame[1] [0]), 
            .I2(\data_in_frame[0][6] ), .I3(\data_in_frame[1] [1]), .O(n59202));   // verilog/coms.v(73[16:27])
    defparam i3_4_lut_adj_1543.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1544 (.I0(\data_in_frame[11] [6]), .I1(n26608), 
            .I2(n59397), .I3(GND_net), .O(n58914));
    defparam i1_2_lut_3_lut_adj_1544.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1545 (.I0(\data_in_frame[4] [4]), .I1(n26316), 
            .I2(GND_net), .I3(GND_net), .O(n59153));   // verilog/coms.v(78[16:43])
    defparam i1_2_lut_adj_1545.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1546 (.I0(\data_in_frame[5] [4]), .I1(n59202), 
            .I2(\data_in_frame[5] [5]), .I3(GND_net), .O(n25700));
    defparam i2_3_lut_adj_1546.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1547 (.I0(\data_in_frame[1] [2]), .I1(\data_in_frame[3] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n58928));   // verilog/coms.v(79[16:43])
    defparam i1_2_lut_adj_1547.LUT_INIT = 16'h6666;
    SB_LUT4 i2_2_lut_3_lut (.I0(n26438), .I1(n54155), .I2(n25987), .I3(GND_net), 
            .O(n10_adj_5080));   // verilog/coms.v(74[16:27])
    defparam i2_2_lut_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i16221_3_lut_4_lut (.I0(n8_adj_5096), .I1(n58755), .I2(rx_data[0]), 
            .I3(\data_in_frame[14] [0]), .O(n30227));
    defparam i16221_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16251_3_lut_4_lut (.I0(n8_adj_5096), .I1(n58755), .I2(rx_data[1]), 
            .I3(\data_in_frame[14] [1]), .O(n30257));
    defparam i16251_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i5_3_lut_4_lut (.I0(\data_in_frame[14] [7]), .I1(\data_in_frame[15] [0]), 
            .I2(n10_adj_5078), .I3(\data_in_frame[14] [5]), .O(n54473));
    defparam i5_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1548 (.I0(\data_in_frame[12] [4]), .I1(\data_in_frame[10] [5]), 
            .I2(n58836), .I3(\data_in_frame[12] [6]), .O(n59394));
    defparam i1_2_lut_4_lut_adj_1548.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1549 (.I0(\data_in_frame[6] [6]), .I1(\data_in_frame[6] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n59365));   // verilog/coms.v(80[16:43])
    defparam i1_2_lut_adj_1549.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_3_lut_adj_1550 (.I0(\data_in_frame[12] [4]), .I1(\data_in_frame[10] [5]), 
            .I2(n58836), .I3(GND_net), .O(n25818));   // verilog/coms.v(74[16:27])
    defparam i1_2_lut_3_lut_adj_1550.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1551 (.I0(\data_in_frame[6] [7]), .I1(\data_in_frame[6] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_5097));   // verilog/coms.v(80[16:43])
    defparam i1_2_lut_adj_1551.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1552 (.I0(\data_in_frame[6] [3]), .I1(\data_in_frame[6] [4]), 
            .I2(\data_in_frame[6] [1]), .I3(n6_adj_5097), .O(n59121));   // verilog/coms.v(80[16:43])
    defparam i4_4_lut_adj_1552.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1553 (.I0(n58876), .I1(n59121), .I2(\data_in_frame[4] [5]), 
            .I3(n59365), .O(n59290));   // verilog/coms.v(80[16:43])
    defparam i3_4_lut_adj_1553.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1554 (.I0(\data_in_frame[5] [7]), .I1(\data_in_frame[3][5] ), 
            .I2(\data_in_frame[1] [3]), .I3(GND_net), .O(n58812));   // verilog/coms.v(78[16:27])
    defparam i2_3_lut_adj_1554.LUT_INIT = 16'h9696;
    SB_LUT4 i4_4_lut_adj_1555 (.I0(n58812), .I1(\data_in_frame[3][6] ), 
            .I2(\data_in_frame[1] [5]), .I3(n59290), .O(n10_adj_5098));
    defparam i4_4_lut_adj_1555.LUT_INIT = 16'h6996;
    SB_LUT4 i16259_3_lut_4_lut (.I0(n8_adj_5096), .I1(n58755), .I2(rx_data[2]), 
            .I3(\data_in_frame[14] [2]), .O(n30265));
    defparam i16259_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16390_3_lut_4_lut (.I0(n8_adj_5096), .I1(n58755), .I2(rx_data[3]), 
            .I3(\data_in_frame[14] [3]), .O(n30396));
    defparam i16390_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_4_lut_adj_1556 (.I0(\FRAME_MATCHER.i[4] ), .I1(\FRAME_MATCHER.i[3] ), 
            .I2(n43501), .I3(n87), .O(n75));   // verilog/coms.v(158[12:15])
    defparam i2_3_lut_4_lut_adj_1556.LUT_INIT = 16'h0020;
    SB_LUT4 i15372_3_lut_4_lut (.I0(n8_adj_5096), .I1(n58755), .I2(rx_data[7]), 
            .I3(\data_in_frame[14] [7]), .O(n29378));
    defparam i15372_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i48358_4_lut (.I0(\data_in_frame[8] [1]), .I1(n26239), .I2(n10_adj_5098), 
            .I3(n54113), .O(n64040));
    defparam i48358_4_lut.LUT_INIT = 16'hedde;
    SB_LUT4 i48497_4_lut (.I0(n54002), .I1(n25892), .I2(n7_adj_5094), 
            .I3(n3_adj_5077), .O(n64182));
    defparam i48497_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i10_4_lut_adj_1557 (.I0(n64040), .I1(n54404), .I2(n25807), 
            .I3(\data_in_frame[8] [0]), .O(n26_adj_5099));
    defparam i10_4_lut_adj_1557.LUT_INIT = 16'h0104;
    SB_LUT4 i48499_4_lut (.I0(n7_adj_4906), .I1(n26411), .I2(n4_adj_5072), 
            .I3(n26251), .O(n64184));
    defparam i48499_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i15369_3_lut_4_lut (.I0(n8_adj_5096), .I1(n58755), .I2(rx_data[6]), 
            .I3(\data_in_frame[14] [6]), .O(n29375));
    defparam i15369_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i9_4_lut_adj_1558 (.I0(n23926), .I1(n54308), .I2(n70014), 
            .I3(n23922), .O(n25_adj_5100));
    defparam i9_4_lut_adj_1558.LUT_INIT = 16'h0800;
    SB_LUT4 i51745_2_lut (.I0(\FRAME_MATCHER.i [14]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n66959));   // verilog/coms.v(158[12:15])
    defparam i51745_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i15366_3_lut_4_lut (.I0(n8_adj_5096), .I1(n58755), .I2(rx_data[5]), 
            .I3(\data_in_frame[14] [5]), .O(n29372));
    defparam i15366_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15363_3_lut_4_lut (.I0(n8_adj_5096), .I1(n58755), .I2(rx_data[4]), 
            .I3(\data_in_frame[14] [4]), .O(n29369));
    defparam i15363_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15_4_lut_adj_1559 (.I0(n25_adj_5100), .I1(n64184), .I2(n26_adj_5099), 
            .I3(n64182), .O(n25455));
    defparam i15_4_lut_adj_1559.LUT_INIT = 16'h0020;
    SB_LUT4 i51895_2_lut (.I0(\FRAME_MATCHER.i_31__N_2513 ), .I1(n25455), 
            .I2(GND_net), .I3(GND_net), .O(n67106));   // verilog/coms.v(18[27:29])
    defparam i51895_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 i19703_4_lut (.I0(n33697), .I1(n67106), .I2(Kp_23__N_1748), 
            .I3(n37), .O(n27674));   // verilog/coms.v(18[27:29])
    defparam i19703_4_lut.LUT_INIT = 16'hca0a;
    SB_LUT4 i1_2_lut_3_lut_adj_1560 (.I0(\data_in_frame[13] [2]), .I1(\data_in_frame[13] [0]), 
            .I2(n58851), .I3(GND_net), .O(n6_adj_5074));
    defparam i1_2_lut_3_lut_adj_1560.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_4_lut_adj_1561 (.I0(\data_in_frame[13] [0]), .I1(n26438), 
            .I2(n25987), .I3(\data_in_frame[12] [5]), .O(n26435));
    defparam i1_2_lut_4_lut_adj_1561.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1562 (.I0(\FRAME_MATCHER.i[3] ), .I1(n9_adj_5029), 
            .I2(n43501), .I3(reset), .O(n58755));   // verilog/coms.v(157[7:23])
    defparam i1_2_lut_3_lut_4_lut_adj_1562.LUT_INIT = 16'hffdf;
    SB_LUT4 i1_2_lut_3_lut_adj_1563 (.I0(n26438), .I1(n25987), .I2(\data_in_frame[12] [5]), 
            .I3(GND_net), .O(n25979));
    defparam i1_2_lut_3_lut_adj_1563.LUT_INIT = 16'h9696;
    SB_LUT4 i1_3_lut_4_lut_adj_1564 (.I0(\data_in_frame[13] [7]), .I1(\data_in_frame[13] [6]), 
            .I2(n53460), .I3(\data_in_frame[13] [5]), .O(n58870));   // verilog/coms.v(99[12:25])
    defparam i1_3_lut_4_lut_adj_1564.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1565 (.I0(n23922), .I1(n23926), .I2(\data_in_frame[9] [6]), 
            .I3(\data_in_frame[10] [0]), .O(n59474));
    defparam i1_2_lut_4_lut_adj_1565.LUT_INIT = 16'h9669;
    SB_LUT4 i4_4_lut_adj_1566 (.I0(ID[4]), .I1(\data_in_frame[0][6] ), .I2(\data_in_frame[0]_c [4]), 
            .I3(ID[6]), .O(n12_adj_5101));   // verilog/coms.v(241[12:32])
    defparam i4_4_lut_adj_1566.LUT_INIT = 16'h7bde;
    SB_LUT4 i2_4_lut_adj_1567 (.I0(\data_in_frame[0] [1]), .I1(\data_in_frame[0]_c [2]), 
            .I2(ID[1]), .I3(ID[2]), .O(n10_adj_5102));   // verilog/coms.v(241[12:32])
    defparam i2_4_lut_adj_1567.LUT_INIT = 16'h7bde;
    SB_LUT4 i3_4_lut_adj_1568 (.I0(\data_in_frame[0] [7]), .I1(\data_in_frame[0]_c [5]), 
            .I2(ID[7]), .I3(ID[5]), .O(n11));   // verilog/coms.v(241[12:32])
    defparam i3_4_lut_adj_1568.LUT_INIT = 16'h7bde;
    SB_LUT4 i1_4_lut_adj_1569 (.I0(\data_in_frame[0][0] ), .I1(\data_in_frame[0][3] ), 
            .I2(ID[0]), .I3(ID[3]), .O(n9_adj_5103));   // verilog/coms.v(241[12:32])
    defparam i1_4_lut_adj_1569.LUT_INIT = 16'h7bde;
    SB_LUT4 i7_4_lut_adj_1570 (.I0(n9_adj_5103), .I1(n11), .I2(n10_adj_5102), 
            .I3(n12_adj_5101), .O(n53031));   // verilog/coms.v(241[12:32])
    defparam i7_4_lut_adj_1570.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_3_lut_adj_1571 (.I0(\data_in_frame[2] [5]), .I1(\data_in_frame[0]_c [4]), 
            .I2(\data_in_frame[0][3] ), .I3(GND_net), .O(n25751));   // verilog/coms.v(169[9:87])
    defparam i2_3_lut_adj_1571.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1572 (.I0(\data_in_frame[0]_c [2]), .I1(\data_in_frame[2] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n58815));   // verilog/coms.v(169[9:87])
    defparam i1_2_lut_adj_1572.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1573 (.I0(\data_in_frame[2] [2]), .I1(\data_in_frame[0][0] ), 
            .I2(\data_in_frame[0] [1]), .I3(GND_net), .O(n26316));   // verilog/coms.v(99[12:25])
    defparam i2_3_lut_adj_1573.LUT_INIT = 16'h9696;
    SB_LUT4 i51580_2_lut (.I0(\FRAME_MATCHER.i [15]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n66962));   // verilog/coms.v(158[12:15])
    defparam i51580_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1_2_lut_adj_1574 (.I0(\data_in_frame[0]_c [2]), .I1(\data_in_frame[0] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n58789));   // verilog/coms.v(99[12:25])
    defparam i1_2_lut_adj_1574.LUT_INIT = 16'h6666;
    SB_LUT4 i15401_3_lut_4_lut (.I0(n98), .I1(n58755), .I2(rx_data[7]), 
            .I3(\data_in_frame[15] [7]), .O(n29407));
    defparam i15401_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i15393_3_lut_4_lut (.I0(n98), .I1(n58755), .I2(rx_data[6]), 
            .I3(\data_in_frame[15] [6]), .O(n29399));
    defparam i15393_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_3_lut_adj_1575 (.I0(\data_in_frame[18] [2]), .I1(\data_in_frame[18] [4]), 
            .I2(\data_in_frame[20] [5]), .I3(GND_net), .O(n59077));
    defparam i1_2_lut_3_lut_adj_1575.LUT_INIT = 16'h9696;
    SB_LUT4 i15390_3_lut_4_lut (.I0(n98), .I1(n58755), .I2(rx_data[5]), 
            .I3(\data_in_frame[15] [5]), .O(n29396));
    defparam i15390_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2_3_lut_4_lut_adj_1576 (.I0(\data_in_frame[16] [3]), .I1(\data_in_frame[16] [2]), 
            .I2(n59379), .I3(n23833), .O(n59380));
    defparam i2_3_lut_4_lut_adj_1576.LUT_INIT = 16'h6996;
    SB_LUT4 i16270_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(rx_data[7]), 
            .I3(\data_in[3] [7]), .O(n30276));   // verilog/coms.v(130[12] 305[6])
    defparam i16270_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_3_lut_adj_1577 (.I0(\data_in_frame[9] [1]), .I1(\data_in_frame[9] [2]), 
            .I2(\data_in_frame[9] [7]), .I3(GND_net), .O(n59100));
    defparam i1_2_lut_3_lut_adj_1577.LUT_INIT = 16'h9696;
    SB_LUT4 i15387_3_lut_4_lut (.I0(n98), .I1(n58755), .I2(rx_data[4]), 
            .I3(\data_in_frame[15] [4]), .O(n29393));
    defparam i15387_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i15384_3_lut_4_lut (.I0(n98), .I1(n58755), .I2(rx_data[3]), 
            .I3(\data_in_frame[15] [3]), .O(n29390));
    defparam i15384_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3_4_lut_adj_1578 (.I0(\data_in_frame[0] [7]), .I1(n6_adj_5104), 
            .I2(n58789), .I3(\data_in_frame[0][6] ), .O(Kp_23__N_748));   // verilog/coms.v(99[12:25])
    defparam i3_4_lut_adj_1578.LUT_INIT = 16'h6996;
    SB_LUT4 i15563_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[1] [0]), 
            .I3(\data_in[0] [0]), .O(n29569));   // verilog/coms.v(130[12] 305[6])
    defparam i15563_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i6_3_lut_adj_1579 (.I0(n26608), .I1(Kp_23__N_748), .I2(\data_in_frame[2] [1]), 
            .I3(GND_net), .O(n22_adj_5105));
    defparam i6_3_lut_adj_1579.LUT_INIT = 16'h1414;
    SB_LUT4 i54332_3_lut (.I0(\data_in_frame[0][6] ), .I1(\data_in_frame[0]_c [5]), 
            .I2(\data_in_frame[2] [7]), .I3(GND_net), .O(n70026));   // verilog/coms.v(99[12:25])
    defparam i54332_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i1_3_lut_adj_1580 (.I0(\data_in_frame[0] [7]), .I1(n1_adj_5106), 
            .I2(\data_in_frame[0][6] ), .I3(GND_net), .O(n27_adj_5107));
    defparam i1_3_lut_adj_1580.LUT_INIT = 16'hdede;
    SB_LUT4 i51829_3_lut (.I0(n1_adj_5106), .I1(\data_in_frame[0] [7]), 
            .I2(\data_in_frame[0][6] ), .I3(GND_net), .O(n67093));   // verilog/coms.v(99[12:25])
    defparam i51829_3_lut.LUT_INIT = 16'h1414;
    SB_LUT4 i10_4_lut_adj_1581 (.I0(\data_in_frame[1] [3]), .I1(\data_in_frame[1] [4]), 
            .I2(\data_in_frame[1] [6]), .I3(n26288), .O(n26_adj_5108));
    defparam i10_4_lut_adj_1581.LUT_INIT = 16'h0080;
    SB_LUT4 i16301_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[1] [1]), 
            .I3(\data_in[0] [1]), .O(n30307));   // verilog/coms.v(130[12] 305[6])
    defparam i16301_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_4_lut_adj_1582 (.I0(n67093), .I1(\data_in_frame[1] [5]), 
            .I2(n27_adj_5107), .I3(\data_in_frame[1] [0]), .O(n17_adj_5109));
    defparam i1_4_lut_adj_1582.LUT_INIT = 16'h0c88;
    SB_LUT4 i48301_2_lut (.I0(n26316), .I1(n25758), .I2(GND_net), .I3(GND_net), 
            .O(n63981));
    defparam i48301_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i16300_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[1] [2]), 
            .I3(\data_in[0] [2]), .O(n30306));   // verilog/coms.v(130[12] 305[6])
    defparam i16300_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i11_4_lut_adj_1583 (.I0(n70026), .I1(n22_adj_5105), .I2(\data_in_frame[0] [7]), 
            .I3(\data_in_frame[1] [1]), .O(n27_adj_5110));
    defparam i11_4_lut_adj_1583.LUT_INIT = 16'h4004;
    SB_LUT4 i16298_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[1] [3]), 
            .I3(\data_in[0] [3]), .O(n30304));   // verilog/coms.v(130[12] 305[6])
    defparam i16298_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i18_4_lut_adj_1584 (.I0(\FRAME_MATCHER.i [30]), .I1(\FRAME_MATCHER.i [21]), 
            .I2(\FRAME_MATCHER.i [24]), .I3(\FRAME_MATCHER.i [17]), .O(n44_adj_5111));   // verilog/coms.v(157[7:23])
    defparam i18_4_lut_adj_1584.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut_adj_1585 (.I0(\FRAME_MATCHER.i [29]), .I1(\FRAME_MATCHER.i [6]), 
            .I2(\FRAME_MATCHER.i [18]), .I3(\FRAME_MATCHER.i [23]), .O(n42_adj_5112));   // verilog/coms.v(157[7:23])
    defparam i16_4_lut_adj_1585.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_4_lut_adj_1586 (.I0(n17_adj_5109), .I1(n26_adj_5108), .I2(n53031), 
            .I3(\data_in_frame[1] [2]), .O(n29_adj_5113));
    defparam i13_4_lut_adj_1586.LUT_INIT = 16'h0800;
    SB_LUT4 i17_4_lut_adj_1587 (.I0(\FRAME_MATCHER.i [7]), .I1(\FRAME_MATCHER.i [20]), 
            .I2(\FRAME_MATCHER.i [12]), .I3(\FRAME_MATCHER.i [14]), .O(n43_adj_5114));   // verilog/coms.v(157[7:23])
    defparam i17_4_lut_adj_1587.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut_adj_1588 (.I0(\FRAME_MATCHER.i [22]), .I1(\FRAME_MATCHER.i [11]), 
            .I2(\FRAME_MATCHER.i [26]), .I3(\FRAME_MATCHER.i [16]), .O(n41_adj_5115));   // verilog/coms.v(157[7:23])
    defparam i15_4_lut_adj_1588.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut_adj_1589 (.I0(n29_adj_5113), .I1(n27_adj_5110), .I2(n23_c), 
            .I3(n63981), .O(\FRAME_MATCHER.state_31__N_2612 [3]));
    defparam i15_4_lut_adj_1589.LUT_INIT = 16'h0080;
    SB_LUT4 i1_2_lut_3_lut_adj_1590 (.I0(n40817), .I1(n43501), .I2(n8_adj_13), 
            .I3(GND_net), .O(n28309));   // verilog/coms.v(156[9:50])
    defparam i1_2_lut_3_lut_adj_1590.LUT_INIT = 16'hf7f7;
    SB_LUT4 i15381_3_lut_4_lut (.I0(n98), .I1(n58755), .I2(rx_data[2]), 
            .I3(\data_in_frame[15] [2]), .O(n29387));
    defparam i15381_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i16297_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[1] [4]), 
            .I3(\data_in[0] [4]), .O(n30303));   // verilog/coms.v(130[12] 305[6])
    defparam i16297_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i16296_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[1] [5]), 
            .I3(\data_in[0] [5]), .O(n30302));   // verilog/coms.v(130[12] 305[6])
    defparam i16296_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i14_4_lut_adj_1591 (.I0(\FRAME_MATCHER.i [13]), .I1(\FRAME_MATCHER.i [15]), 
            .I2(\FRAME_MATCHER.i [10]), .I3(\FRAME_MATCHER.i [28]), .O(n40_adj_5116));   // verilog/coms.v(157[7:23])
    defparam i14_4_lut_adj_1591.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_2_lut_adj_1592 (.I0(\FRAME_MATCHER.i [9]), .I1(\FRAME_MATCHER.i [27]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_5117));   // verilog/coms.v(157[7:23])
    defparam i13_2_lut_adj_1592.LUT_INIT = 16'heeee;
    SB_LUT4 i24_4_lut (.I0(n41_adj_5115), .I1(n43_adj_5114), .I2(n42_adj_5112), 
            .I3(n44_adj_5111), .O(n50));   // verilog/coms.v(157[7:23])
    defparam i24_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i19_4_lut_adj_1593 (.I0(\FRAME_MATCHER.i [8]), .I1(\FRAME_MATCHER.i [25]), 
            .I2(\FRAME_MATCHER.i[5] ), .I3(\FRAME_MATCHER.i [19]), .O(n45_adj_5118));   // verilog/coms.v(157[7:23])
    defparam i19_4_lut_adj_1593.LUT_INIT = 16'hfffe;
    SB_LUT4 i15378_3_lut_4_lut (.I0(n98), .I1(n58755), .I2(rx_data[1]), 
            .I3(\data_in_frame[15] [1]), .O(n29384));
    defparam i15378_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i16295_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[1] [6]), 
            .I3(\data_in[0] [6]), .O(n30301));   // verilog/coms.v(130[12] 305[6])
    defparam i16295_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2_3_lut_4_lut_adj_1594 (.I0(\data_in_frame[9] [3]), .I1(\data_in_frame[9] [4]), 
            .I2(n61424), .I3(\data_in_frame[7] [3]), .O(n53442));
    defparam i2_3_lut_4_lut_adj_1594.LUT_INIT = 16'h6996;
    SB_LUT4 select_775_Select_66_i2_4_lut (.I0(\data_out_frame[8] [2]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder0_position_scaled[2]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_66_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_3_lut_adj_1595 (.I0(n40817), .I1(n43501), .I2(n8_adj_15), 
            .I3(GND_net), .O(n28311));   // verilog/coms.v(156[9:50])
    defparam i1_2_lut_3_lut_adj_1595.LUT_INIT = 16'hf7f7;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1596 (.I0(reset), .I1(n43501), .I2(\FRAME_MATCHER.i[3] ), 
            .I3(n9_adj_5029), .O(n58760));
    defparam i1_2_lut_3_lut_4_lut_adj_1596.LUT_INIT = 16'hfffb;
    SB_LUT4 i25_4_lut (.I0(n45_adj_5118), .I1(n50), .I2(n39_adj_5117), 
            .I3(n40_adj_5116), .O(n25474));   // verilog/coms.v(157[7:23])
    defparam i25_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i29153_4_lut (.I0(\FRAME_MATCHER.i[3] ), .I1(\FRAME_MATCHER.i [31]), 
            .I2(n25474), .I3(\FRAME_MATCHER.i[4] ), .O(n4452));   // verilog/coms.v(262[9:58])
    defparam i29153_4_lut.LUT_INIT = 16'h3230;
    SB_LUT4 i30_3_lut_4_lut (.I0(n98), .I1(n58755), .I2(\data_in_frame[15] [0]), 
            .I3(rx_data[0]), .O(n22_adj_5013));
    defparam i30_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 i464_2_lut (.I0(n4452), .I1(\FRAME_MATCHER.i_31__N_2514 ), .I2(GND_net), 
            .I3(GND_net), .O(n2068));   // verilog/coms.v(148[4] 304[11])
    defparam i464_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i16294_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[1] [7]), 
            .I3(\data_in[0] [7]), .O(n30300));   // verilog/coms.v(130[12] 305[6])
    defparam i16294_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i16293_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[2] [0]), 
            .I3(\data_in[1] [0]), .O(n30299));   // verilog/coms.v(130[12] 305[6])
    defparam i16293_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i16291_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[2] [2]), 
            .I3(\data_in[1] [2]), .O(n30297));   // verilog/coms.v(130[12] 305[6])
    defparam i16291_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i16290_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[2] [3]), 
            .I3(\data_in[1] [3]), .O(n30296));   // verilog/coms.v(130[12] 305[6])
    defparam i16290_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i16289_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[2] [4]), 
            .I3(\data_in[1] [4]), .O(n30295));   // verilog/coms.v(130[12] 305[6])
    defparam i16289_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i16288_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[2] [5]), 
            .I3(\data_in[1] [5]), .O(n30294));   // verilog/coms.v(130[12] 305[6])
    defparam i16288_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i14_2_lut (.I0(deadband[9]), .I1(n367), .I2(GND_net), .I3(GND_net), 
            .O(n19_adj_16));
    defparam i14_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i16287_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[2] [6]), 
            .I3(\data_in[1] [6]), .O(n30293));   // verilog/coms.v(130[12] 305[6])
    defparam i16287_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i16286_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[2] [7]), 
            .I3(\data_in[1] [7]), .O(n30292));   // verilog/coms.v(130[12] 305[6])
    defparam i16286_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i16285_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[3] [0]), 
            .I3(\data_in[2] [0]), .O(n30291));   // verilog/coms.v(130[12] 305[6])
    defparam i16285_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i15_2_lut_adj_1597 (.I0(PWMLimit[15]), .I1(n361), .I2(GND_net), 
            .I3(GND_net), .O(n31));
    defparam i15_2_lut_adj_1597.LUT_INIT = 16'h6666;
    SB_LUT4 i2_2_lut_3_lut_adj_1598 (.I0(n25987), .I1(\data_in_frame[12] [5]), 
            .I2(n54155), .I3(GND_net), .O(n6_adj_5066));
    defparam i2_2_lut_3_lut_adj_1598.LUT_INIT = 16'h9696;
    SB_LUT4 i51899_2_lut (.I0(\FRAME_MATCHER.i [16]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n66966));   // verilog/coms.v(158[12:15])
    defparam i51899_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i16284_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[3] [1]), 
            .I3(\data_in[2] [1]), .O(n30290));   // verilog/coms.v(130[12] 305[6])
    defparam i16284_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_3_lut_adj_1599 (.I0(n40817), .I1(n43501), .I2(n8_adj_12), 
            .I3(GND_net), .O(n28313));   // verilog/coms.v(156[9:50])
    defparam i1_2_lut_3_lut_adj_1599.LUT_INIT = 16'hf7f7;
    SB_LUT4 i29610_2_lut_3_lut (.I0(n40817), .I1(n43501), .I2(n98), .I3(GND_net), 
            .O(n43503));   // verilog/coms.v(156[9:50])
    defparam i29610_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[10] [3]), .I2(\data_out_frame[11] [3]), 
            .I3(\byte_transmit_counter[1] ), .O(n71258));
    defparam byte_transmit_counter_0__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 i23677_3_lut (.I0(n18), .I1(PWMLimit[9]), .I2(n367), .I3(GND_net), 
            .O(n20));
    defparam i23677_3_lut.LUT_INIT = 16'hb2b2;
    SB_LUT4 i51666_2_lut (.I0(\FRAME_MATCHER.i [17]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n66967));   // verilog/coms.v(158[12:15])
    defparam i51666_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i15650_3_lut_4_lut (.I0(n8_adj_5096), .I1(n58720), .I2(rx_data[7]), 
            .I3(\data_in_frame[22] [7]), .O(n29656));
    defparam i15650_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 n71258_bdd_4_lut (.I0(n71258), .I1(\data_out_frame[9] [3]), 
            .I2(\data_out_frame[8] [3]), .I3(\byte_transmit_counter[1] ), 
            .O(n64471));
    defparam n71258_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i15647_3_lut_4_lut (.I0(n8_adj_5096), .I1(n58720), .I2(rx_data[6]), 
            .I3(\data_in_frame[22] [6]), .O(n29653));
    defparam i15647_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15603_3_lut_4_lut (.I0(n8_adj_5096), .I1(n58720), .I2(rx_data[5]), 
            .I3(\data_in_frame[22] [5]), .O(n29609));
    defparam i15603_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15593_3_lut_4_lut (.I0(n8_adj_5096), .I1(n58720), .I2(rx_data[4]), 
            .I3(\data_in_frame[22] [4]), .O(n29599));
    defparam i15593_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15590_3_lut_4_lut (.I0(n8_adj_5096), .I1(n58720), .I2(rx_data[3]), 
            .I3(\data_in_frame[22] [3]), .O(n29596));
    defparam i15590_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15586_3_lut_4_lut (.I0(n8_adj_5096), .I1(n58720), .I2(rx_data[2]), 
            .I3(\data_in_frame[22] [2]), .O(n29592));
    defparam i15586_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16283_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[3] [2]), 
            .I3(\data_in[2] [2]), .O(n30289));   // verilog/coms.v(130[12] 305[6])
    defparam i16283_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_3_lut_adj_1600 (.I0(\data_in_frame[12] [2]), .I1(\data_in_frame[12] [3]), 
            .I2(n59474), .I3(GND_net), .O(n6_adj_5065));
    defparam i1_2_lut_3_lut_adj_1600.LUT_INIT = 16'h9696;
    SB_LUT4 i15583_3_lut_4_lut (.I0(n8_adj_5096), .I1(n58720), .I2(rx_data[1]), 
            .I3(\data_in_frame[22] [1]), .O(n29589));
    defparam i15583_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15580_3_lut_4_lut (.I0(n8_adj_5096), .I1(n58720), .I2(rx_data[0]), 
            .I3(\data_in_frame[22] [0]), .O(n29586));
    defparam i15580_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1601 (.I0(\data_in_frame[21] [3]), .I1(n26085), 
            .I2(n59106), .I3(GND_net), .O(n25953));
    defparam i1_2_lut_3_lut_adj_1601.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1602 (.I0(\FRAME_MATCHER.i [2]), .I1(\FRAME_MATCHER.i [1]), 
            .I2(\FRAME_MATCHER.i[0] ), .I3(GND_net), .O(n98));
    defparam i1_2_lut_3_lut_adj_1602.LUT_INIT = 16'h8080;
    SB_LUT4 i16282_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[3] [3]), 
            .I3(\data_in[2] [3]), .O(n30288));   // verilog/coms.v(130[12] 305[6])
    defparam i16282_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i52423_2_lut (.I0(\FRAME_MATCHER.i [18]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n66972));   // verilog/coms.v(158[12:15])
    defparam i52423_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1_2_lut_3_lut_adj_1603 (.I0(\FRAME_MATCHER.i [2]), .I1(\FRAME_MATCHER.i [1]), 
            .I2(\FRAME_MATCHER.i[0] ), .I3(GND_net), .O(n8_adj_5096));
    defparam i1_2_lut_3_lut_adj_1603.LUT_INIT = 16'hf7f7;
    SB_LUT4 i22317_3_lut (.I0(n230), .I1(IntegralLimit[1]), .I2(n155), 
            .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3715[1] ));
    defparam i22317_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2_3_lut_4_lut_adj_1604 (.I0(n3468), .I1(n140), .I2(n40660), 
            .I3(n40817), .O(n159));
    defparam i2_3_lut_4_lut_adj_1604.LUT_INIT = 16'hfdff;
    SB_LUT4 i1_2_lut_3_lut_adj_1605 (.I0(n3468), .I1(n140), .I2(n161), 
            .I3(GND_net), .O(n163));
    defparam i1_2_lut_3_lut_adj_1605.LUT_INIT = 16'hfdfd;
    SB_LUT4 i1_2_lut_3_lut_adj_1606 (.I0(\data_out_frame[12] [3]), .I1(n1513), 
            .I2(n59329), .I3(GND_net), .O(n26849));   // verilog/coms.v(77[16:43])
    defparam i1_2_lut_3_lut_adj_1606.LUT_INIT = 16'h9696;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_55392 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[6] [3]), .I2(\data_out_frame[7] [3]), .I3(\byte_transmit_counter[1] ), 
            .O(n71018));
    defparam byte_transmit_counter_0__bdd_4_lut_55392.LUT_INIT = 16'he4aa;
    SB_LUT4 i51846_2_lut (.I0(\FRAME_MATCHER.i [19]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n66973));   // verilog/coms.v(158[12:15])
    defparam i51846_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_55492 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[10] [5]), .I2(\data_out_frame[11] [5]), 
            .I3(\byte_transmit_counter[1] ), .O(n71252));
    defparam byte_transmit_counter_0__bdd_4_lut_55492.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_2_lut_3_lut_adj_1607 (.I0(n54458), .I1(n61382), .I2(\data_in_frame[16] [6]), 
            .I3(GND_net), .O(n54411));
    defparam i1_2_lut_3_lut_adj_1607.LUT_INIT = 16'h9696;
    SB_LUT4 i51637_2_lut (.I0(\FRAME_MATCHER.i [20]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n66992));   // verilog/coms.v(158[12:15])
    defparam i51637_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i16281_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[3] [4]), 
            .I3(\data_in[2] [4]), .O(n30287));   // verilog/coms.v(130[12] 305[6])
    defparam i16281_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2_3_lut_4_lut_adj_1608 (.I0(\data_in_frame[20] [7]), .I1(n54447), 
            .I2(\data_in_frame[19] [0]), .I3(\data_in_frame[16] [3]), .O(n58981));
    defparam i2_3_lut_4_lut_adj_1608.LUT_INIT = 16'h6996;
    SB_LUT4 n71252_bdd_4_lut (.I0(n71252), .I1(\data_out_frame[9] [5]), 
            .I2(\data_out_frame[8] [5]), .I3(\byte_transmit_counter[1] ), 
            .O(n71255));
    defparam n71252_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_3_lut_4_lut_adj_1609 (.I0(\data_in_frame[18] [1]), .I1(\data_in_frame[18] [3]), 
            .I2(n54516), .I3(\data_in_frame[18] [2]), .O(n59341));
    defparam i1_3_lut_4_lut_adj_1609.LUT_INIT = 16'h6996;
    SB_LUT4 i16280_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[3] [5]), 
            .I3(\data_in[2] [5]), .O(n30286));   // verilog/coms.v(130[12] 305[6])
    defparam i16280_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i51648_2_lut (.I0(\FRAME_MATCHER.i [21]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n66993));   // verilog/coms.v(158[12:15])
    defparam i51648_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i16279_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[3] [6]), 
            .I3(\data_in[2] [6]), .O(n30285));   // verilog/coms.v(130[12] 305[6])
    defparam i16279_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i16278_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[3] [7]), 
            .I3(\data_in[2] [7]), .O(n30284));   // verilog/coms.v(130[12] 305[6])
    defparam i16278_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_55487 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[14] [3]), .I2(\data_out_frame[15] [3]), 
            .I3(\byte_transmit_counter[1] ), .O(n71246));
    defparam byte_transmit_counter_0__bdd_4_lut_55487.LUT_INIT = 16'he4aa;
    SB_LUT4 i16277_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(rx_data[0]), 
            .I3(\data_in[3] [0]), .O(n30283));   // verilog/coms.v(130[12] 305[6])
    defparam i16277_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i52352_2_lut (.I0(\FRAME_MATCHER.i [22]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n66997));   // verilog/coms.v(158[12:15])
    defparam i52352_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i2_3_lut_4_lut_adj_1610 (.I0(n40660), .I1(n140), .I2(n10_adj_4991), 
            .I3(n3468), .O(n58418));   // verilog/coms.v(156[9:50])
    defparam i2_3_lut_4_lut_adj_1610.LUT_INIT = 16'h0100;
    SB_LUT4 i16276_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(rx_data[1]), 
            .I3(\data_in[3] [1]), .O(n30282));   // verilog/coms.v(130[12] 305[6])
    defparam i16276_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i51660_2_lut (.I0(\FRAME_MATCHER.i [23]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n66998));   // verilog/coms.v(158[12:15])
    defparam i51660_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i16275_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(rx_data[2]), 
            .I3(\data_in[3] [2]), .O(n30281));   // verilog/coms.v(130[12] 305[6])
    defparam i16275_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i16274_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(rx_data[3]), 
            .I3(\data_in[3] [3]), .O(n30280));   // verilog/coms.v(130[12] 305[6])
    defparam i16274_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i14371_3_lut_4_lut (.I0(n40660), .I1(n140), .I2(n58731), .I3(reset), 
            .O(n59644));   // verilog/coms.v(156[9:50])
    defparam i14371_3_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 n71018_bdd_4_lut (.I0(n71018), .I1(\data_out_frame[5] [3]), 
            .I2(\data_out_frame[4] [3]), .I3(\byte_transmit_counter[1] ), 
            .O(n64383));
    defparam n71018_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i16273_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(rx_data[4]), 
            .I3(\data_in[3] [4]), .O(n30279));   // verilog/coms.v(130[12] 305[6])
    defparam i16273_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i51670_2_lut (.I0(\FRAME_MATCHER.i [24]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n66999));   // verilog/coms.v(158[12:15])
    defparam i51670_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 n71246_bdd_4_lut (.I0(n71246), .I1(\data_out_frame[13] [3]), 
            .I2(\data_out_frame[12] [3]), .I3(\byte_transmit_counter[1] ), 
            .O(n64480));
    defparam n71246_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut (.I0(byte_transmit_counter[3]), 
            .I1(n69205), .I2(n67162), .I3(byte_transmit_counter[4]), .O(n71240));
    defparam byte_transmit_counter_3__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n71240_bdd_4_lut (.I0(n71240), .I1(n70943), .I2(n7_adj_5033), 
            .I3(byte_transmit_counter[4]), .O(tx_data[0]));
    defparam n71240_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i16272_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(rx_data[5]), 
            .I3(\data_in[3] [5]), .O(n30278));   // verilog/coms.v(130[12] 305[6])
    defparam i16272_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2_3_lut_4_lut_adj_1611 (.I0(\data_out_frame[16] [1]), .I1(\data_out_frame[16] [2]), 
            .I2(n59481), .I3(n58785), .O(n59244));
    defparam i2_3_lut_4_lut_adj_1611.LUT_INIT = 16'h6996;
    SB_LUT4 i16271_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(rx_data[6]), 
            .I3(\data_in[3] [6]), .O(n30277));   // verilog/coms.v(130[12] 305[6])
    defparam i16271_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i23369_3_lut (.I0(n33), .I1(n375), .I2(n401), .I3(GND_net), 
            .O(n4_adj_17));
    defparam i23369_3_lut.LUT_INIT = 16'hb2b2;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_55299 (.I0(\byte_transmit_counter[1] ), 
            .I1(n64436), .I2(n64437), .I3(\byte_transmit_counter[2] ), 
            .O(n71012));
    defparam byte_transmit_counter_1__bdd_4_lut_55299.LUT_INIT = 16'he4aa;
    SB_LUT4 n71012_bdd_4_lut (.I0(n71012), .I1(n64530), .I2(n64529), .I3(\byte_transmit_counter[2] ), 
            .O(n71015));
    defparam n71012_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i16292_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[2] [1]), 
            .I3(\data_in[1] [1]), .O(n30298));   // verilog/coms.v(130[12] 305[6])
    defparam i16292_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2_3_lut_4_lut_adj_1612 (.I0(\data_out_frame[16] [1]), .I1(\data_out_frame[16] [2]), 
            .I2(n54490), .I3(n54434), .O(n59074));
    defparam i2_3_lut_4_lut_adj_1612.LUT_INIT = 16'h6996;
    SB_LUT4 i51622_2_lut (.I0(\FRAME_MATCHER.i [25]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n67003));   // verilog/coms.v(158[12:15])
    defparam i51622_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i51534_2_lut (.I0(\FRAME_MATCHER.i [26]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n67028));   // verilog/coms.v(158[12:15])
    defparam i51534_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i52336_2_lut (.I0(\FRAME_MATCHER.i [27]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n67036));   // verilog/coms.v(158[12:15])
    defparam i52336_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1_2_lut_4_lut_adj_1613 (.I0(n59284), .I1(n58870), .I2(\data_in_frame[13] [2]), 
            .I3(n59206), .O(n7_adj_5053));
    defparam i1_2_lut_4_lut_adj_1613.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_55477 (.I0(byte_transmit_counter[3]), 
            .I1(n71015), .I2(n66934), .I3(byte_transmit_counter[4]), .O(n71234));
    defparam byte_transmit_counter_3__bdd_4_lut_55477.LUT_INIT = 16'he4aa;
    SB_LUT4 i5_3_lut_4_lut_adj_1614 (.I0(\data_in_frame[16] [1]), .I1(\data_in_frame[13] [7]), 
            .I2(n10_adj_5050), .I3(\data_in_frame[16] [2]), .O(n54513));
    defparam i5_3_lut_4_lut_adj_1614.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1615 (.I0(\data_out_frame[16] [1]), .I1(\data_out_frame[16] [2]), 
            .I2(\data_out_frame[16] [7]), .I3(GND_net), .O(n58953));
    defparam i1_2_lut_3_lut_adj_1615.LUT_INIT = 16'h9696;
    SB_LUT4 i1_3_lut_4_lut_adj_1616 (.I0(n54458), .I1(n59067), .I2(\data_in_frame[16] [2]), 
            .I3(\data_in_frame[20] [6]), .O(n63743));
    defparam i1_3_lut_4_lut_adj_1616.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_55289 (.I0(\byte_transmit_counter[1] ), 
            .I1(n64553), .I2(n64554), .I3(\byte_transmit_counter[2] ), 
            .O(n71006));
    defparam byte_transmit_counter_1__bdd_4_lut_55289.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_2_lut_4_lut_adj_1617 (.I0(n59281), .I1(\data_out_frame[11] [0]), 
            .I2(n58861), .I3(\data_out_frame[8] [3]), .O(n59384));
    defparam i1_2_lut_4_lut_adj_1617.LUT_INIT = 16'h6996;
    SB_LUT4 n71006_bdd_4_lut (.I0(n71006), .I1(n64548), .I2(n64547), .I3(\byte_transmit_counter[2] ), 
            .O(n71009));
    defparam n71006_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4_2_lut_4_lut (.I0(n59281), .I1(\data_out_frame[11] [0]), .I2(n58861), 
            .I3(n59415), .O(n26_adj_4871));
    defparam i4_2_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1618 (.I0(\data_out_frame[4] [6]), .I1(\data_out_frame[5] [0]), 
            .I2(\data_out_frame[7] [2]), .I3(\data_out_frame[5] [1]), .O(n26039));   // verilog/coms.v(88[17:28])
    defparam i2_3_lut_4_lut_adj_1618.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1619 (.I0(\data_out_frame[4] [6]), .I1(\data_out_frame[5] [0]), 
            .I2(\data_out_frame[7] [0]), .I3(n58897), .O(n26298));   // verilog/coms.v(88[17:28])
    defparam i2_3_lut_4_lut_adj_1619.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1620 (.I0(\data_out_frame[6] [2]), .I1(\data_out_frame[4] [0]), 
            .I2(\data_out_frame[4] [1]), .I3(GND_net), .O(n58873));   // verilog/coms.v(77[16:43])
    defparam i1_2_lut_3_lut_adj_1620.LUT_INIT = 16'h9696;
    SB_LUT4 select_775_Select_8_i2_3_lut (.I0(\data_out_frame[1][0] ), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\FRAME_MATCHER.state_31__N_2612 [3]), .I3(GND_net), .O(n2_adj_5011));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_8_i2_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i1_2_lut_3_lut_adj_1621 (.I0(\data_out_frame[15] [5]), .I1(n54220), 
            .I2(n26210), .I3(GND_net), .O(n59308));
    defparam i1_2_lut_3_lut_adj_1621.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1622 (.I0(\data_out_frame[15] [5]), .I1(n54220), 
            .I2(\data_out_frame[15] [4]), .I3(GND_net), .O(n59305));
    defparam i1_2_lut_3_lut_adj_1622.LUT_INIT = 16'h9696;
    SB_LUT4 n71234_bdd_4_lut (.I0(n71234), .I1(n71009), .I2(n7_adj_5031), 
            .I3(byte_transmit_counter[4]), .O(tx_data[7]));
    defparam n71234_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 select_775_Select_4_i2_3_lut (.I0(\data_out_frame[0][4] ), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\FRAME_MATCHER.state_31__N_2612 [3]), .I3(GND_net), .O(n2_adj_5010));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_4_i2_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 select_775_Select_3_i2_3_lut (.I0(\data_out_frame[0][3] ), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\FRAME_MATCHER.state_31__N_2612 [3]), .I3(GND_net), .O(n2_adj_5009));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_3_i2_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i51714_2_lut (.I0(\FRAME_MATCHER.i [28]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n67037));   // verilog/coms.v(158[12:15])
    defparam i51714_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 select_775_Select_2_i2_3_lut (.I0(\data_out_frame[0][2] ), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\FRAME_MATCHER.state_31__N_2612 [3]), .I3(GND_net), .O(n2_adj_5008));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_2_i2_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_55472 (.I0(byte_transmit_counter[3]), 
            .I1(n69199), .I2(n67143), .I3(byte_transmit_counter[4]), .O(n71228));
    defparam byte_transmit_counter_3__bdd_4_lut_55472.LUT_INIT = 16'he4aa;
    SB_LUT4 i2_3_lut_4_lut_adj_1623 (.I0(n54620), .I1(n25872), .I2(n59027), 
            .I3(n59353), .O(n54479));
    defparam i2_3_lut_4_lut_adj_1623.LUT_INIT = 16'h9669;
    SB_LUT4 n71228_bdd_4_lut (.I0(n71228), .I1(n70949), .I2(n7_adj_5030), 
            .I3(byte_transmit_counter[4]), .O(tx_data[6]));
    defparam n71228_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i2_3_lut_4_lut_adj_1624 (.I0(n54620), .I1(n25872), .I2(n26849), 
            .I3(n26372), .O(n59010));
    defparam i2_3_lut_4_lut_adj_1624.LUT_INIT = 16'h9669;
    SB_LUT4 i15820_3_lut_4_lut (.I0(n28337), .I1(reset), .I2(rx_data[0]), 
            .I3(\data_in_frame[3] [0]), .O(n29826));
    defparam i15820_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15823_3_lut_4_lut (.I0(n28337), .I1(reset), .I2(rx_data[1]), 
            .I3(\data_in_frame[3] [1]), .O(n29829));
    defparam i15823_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15826_3_lut_4_lut (.I0(n28337), .I1(reset), .I2(rx_data[2]), 
            .I3(\data_in_frame[3] [2]), .O(n29832));
    defparam i15826_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15829_3_lut_4_lut (.I0(n28337), .I1(reset), .I2(rx_data[3]), 
            .I3(\data_in_frame[3] [3]), .O(n29835));
    defparam i15829_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15832_3_lut_4_lut (.I0(n28337), .I1(reset), .I2(rx_data[4]), 
            .I3(\data_in_frame[3] [4]), .O(n29838));
    defparam i15832_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15835_3_lut_4_lut (.I0(n28337), .I1(reset), .I2(rx_data[5]), 
            .I3(\data_in_frame[3][5] ), .O(n29841));
    defparam i15835_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15839_3_lut_4_lut (.I0(n28337), .I1(reset), .I2(rx_data[6]), 
            .I3(\data_in_frame[3][6] ), .O(n29845));
    defparam i15839_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11_4_lut_4_lut (.I0(n28337), .I1(reset), .I2(rx_data[7]), 
            .I3(\data_in_frame[3] [7]), .O(n58126));
    defparam i11_4_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 select_777_Select_7_i1_2_lut_3_lut (.I0(\FRAME_MATCHER.state[3] ), 
            .I1(\FRAME_MATCHER.i_31__N_2511 ), .I2(byte_transmit_counter[7]), 
            .I3(GND_net), .O(n1_adj_5041));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_7_i1_2_lut_3_lut.LUT_INIT = 16'h1010;
    SB_LUT4 i14381_3_lut_4_lut (.I0(n10_adj_4991), .I1(n43501), .I2(reset), 
            .I3(n98), .O(n59638));
    defparam i14381_3_lut_4_lut.LUT_INIT = 16'hfbff;
    SB_LUT4 i51721_2_lut (.I0(\FRAME_MATCHER.i [29]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n67042));   // verilog/coms.v(158[12:15])
    defparam i51721_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1_2_lut_4_lut_adj_1625 (.I0(n40817), .I1(n40660), .I2(n140), 
            .I3(n3468), .O(n28307));   // verilog/coms.v(148[4] 304[11])
    defparam i1_2_lut_4_lut_adj_1625.LUT_INIT = 16'hfdff;
    SB_LUT4 i14347_3_lut_4_lut (.I0(n10_adj_4991), .I1(n43501), .I2(reset), 
            .I3(n8_adj_12), .O(n7));
    defparam i14347_3_lut_4_lut.LUT_INIT = 16'hfffb;
    SB_LUT4 equal_298_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [2]), .I1(\FRAME_MATCHER.i [1]), 
            .I2(\FRAME_MATCHER.i[0] ), .I3(GND_net), .O(n8_adj_4950));   // verilog/coms.v(158[12:15])
    defparam equal_298_i8_2_lut_3_lut.LUT_INIT = 16'hbfbf;
    SB_LUT4 select_775_Select_186_i2_4_lut (.I0(\data_out_frame[23] [2]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[18]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4997));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_186_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_775_Select_185_i2_4_lut (.I0(\data_out_frame[23] [1]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[17]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4996));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_185_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i54947_2_lut_3_lut (.I0(tx_active), .I1(r_SM_Main_2__N_3545[0]), 
            .I2(n43563), .I3(GND_net), .O(tx_transmit_N_3416));
    defparam i54947_2_lut_3_lut.LUT_INIT = 16'h0101;
    SB_LUT4 select_775_Select_184_i2_4_lut (.I0(\data_out_frame[23] [0]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[16]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4995));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_184_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_775_Select_183_i2_4_lut (.I0(\data_out_frame[22] [7]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(\current[7] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4994));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_183_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i13972_4_lut (.I0(\FRAME_MATCHER.i[0] ), .I1(n133[0]), .I2(n3468), 
            .I3(\FRAME_MATCHER.i_31__N_2507 ), .O(n27978));   // verilog/coms.v(158[12:15])
    defparam i13972_4_lut.LUT_INIT = 16'hc0ca;
    SB_LUT4 equal_307_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [2]), .I1(\FRAME_MATCHER.i [1]), 
            .I2(\FRAME_MATCHER.i[0] ), .I3(GND_net), .O(n8_adj_13));   // verilog/coms.v(158[12:15])
    defparam equal_307_i8_2_lut_3_lut.LUT_INIT = 16'hfbfb;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_55462 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[22] [0]), .I2(\data_out_frame[23] [0]), 
            .I3(\byte_transmit_counter[1] ), .O(n71216));
    defparam byte_transmit_counter_0__bdd_4_lut_55462.LUT_INIT = 16'he4aa;
    SB_LUT4 i2_2_lut_3_lut_adj_1626 (.I0(\data_in_frame[0]_c [5]), .I1(\data_in_frame[0]_c [4]), 
            .I2(\data_in_frame[0][3] ), .I3(GND_net), .O(n6_adj_5104));   // verilog/coms.v(88[17:70])
    defparam i2_2_lut_3_lut_adj_1626.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1627 (.I0(\data_in_frame[0]_c [5]), .I1(\data_in_frame[0]_c [4]), 
            .I2(\data_in_frame[2] [6]), .I3(GND_net), .O(n26608));   // verilog/coms.v(88[17:70])
    defparam i1_2_lut_3_lut_adj_1627.LUT_INIT = 16'h9696;
    SB_LUT4 n71216_bdd_4_lut (.I0(n71216), .I1(\data_out_frame[21] [0]), 
            .I2(\data_out_frame[20] [0]), .I3(\byte_transmit_counter[1] ), 
            .O(n71219));
    defparam n71216_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_3_lut_adj_1628 (.I0(\data_in_frame[0][0] ), .I1(Kp_23__N_748), 
            .I2(\data_in_frame[2] [0]), .I3(GND_net), .O(n1_adj_5106));   // verilog/coms.v(73[16:69])
    defparam i1_2_lut_3_lut_adj_1628.LUT_INIT = 16'h9696;
    SB_LUT4 select_777_Select_6_i1_2_lut_3_lut (.I0(\FRAME_MATCHER.state[3] ), 
            .I1(\FRAME_MATCHER.i_31__N_2511 ), .I2(byte_transmit_counter[6]), 
            .I3(GND_net), .O(n1_adj_5040));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_6_i1_2_lut_3_lut.LUT_INIT = 16'h1010;
    SB_LUT4 i7_3_lut_4_lut (.I0(\data_in_frame[0][0] ), .I1(Kp_23__N_748), 
            .I2(n25751), .I3(\data_in_frame[1] [7]), .O(n23_c));   // verilog/coms.v(73[16:69])
    defparam i7_3_lut_4_lut.LUT_INIT = 16'h0906;
    SB_LUT4 select_775_Select_182_i2_4_lut (.I0(\data_out_frame[22] [6]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(\current[6] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4980));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_182_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_775_Select_181_i2_4_lut (.I0(\data_out_frame[22] [5]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(\current[5] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4979));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_181_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_4_lut_adj_1629 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[22] [4]), 
            .I2(\current[4] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4978));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1629.LUT_INIT = 16'ha088;
    SB_LUT4 select_775_Select_179_i2_4_lut (.I0(\data_out_frame[22] [3]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(\current[3] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4977));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_179_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i2_3_lut_4_lut_adj_1630 (.I0(n1954), .I1(n1951), .I2(\FRAME_MATCHER.i_31__N_2507 ), 
            .I3(n1957), .O(n61225));   // verilog/coms.v(148[4] 304[11])
    defparam i2_3_lut_4_lut_adj_1630.LUT_INIT = 16'h8000;
    SB_LUT4 select_775_Select_178_i2_4_lut (.I0(\data_out_frame[22] [2]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(\current[2] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4976));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_178_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_775_Select_177_i2_4_lut (.I0(\data_out_frame[22] [1]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(\current[1] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4975));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_177_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_4_lut_adj_1631 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[22] [0]), 
            .I2(\current[0] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4974));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1631.LUT_INIT = 16'ha088;
    SB_LUT4 select_775_Select_175_i2_4_lut (.I0(\data_out_frame[21] [7]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(\current[15] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4973));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_175_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i23372_3_lut (.I0(n376), .I1(n456), .I2(n11597), .I3(GND_net), 
            .O(n27629));
    defparam i23372_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 select_775_Select_174_i2_4_lut (.I0(\data_out_frame[21] [6]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(\current[15] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4972));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_174_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i51723_2_lut (.I0(\FRAME_MATCHER.i [30]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n67043));   // verilog/coms.v(158[12:15])
    defparam i51723_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 select_775_Select_173_i2_4_lut (.I0(\data_out_frame[21] [5]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(\current[15] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4971));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_173_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_4_lut_adj_1632 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[21] [4]), 
            .I2(\current[15] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4970));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1632.LUT_INIT = 16'ha088;
    SB_LUT4 i1_3_lut_4_lut_adj_1633 (.I0(\FRAME_MATCHER.i_31__N_2511 ), .I1(tx_active), 
            .I2(r_SM_Main_2__N_3545[0]), .I3(n43563), .O(n25463));   // verilog/coms.v(148[4] 304[11])
    defparam i1_3_lut_4_lut_adj_1633.LUT_INIT = 16'ha8aa;
    SB_LUT4 select_775_Select_171_i2_4_lut (.I0(\data_out_frame[21] [3]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(\current[11] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4969));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_171_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_775_Select_170_i2_4_lut (.I0(\data_out_frame[21] [2]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(\current[10] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4968));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_170_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i51724_2_lut (.I0(\FRAME_MATCHER.i [31]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n67044));   // verilog/coms.v(158[12:15])
    defparam i51724_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 select_775_Select_169_i2_4_lut (.I0(\data_out_frame[21] [1]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(\current[9] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4967));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_169_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1634 (.I0(\data_out_frame[20] [3]), .I1(n23652), 
            .I2(\data_out_frame[20] [2]), .I3(n54415), .O(n58893));
    defparam i1_2_lut_3_lut_4_lut_adj_1634.LUT_INIT = 16'h6996;
    SB_LUT4 select_775_Select_168_i2_4_lut (.I0(\data_out_frame[21] [0]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(\current[8] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4966));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_168_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_775_Select_167_i2_4_lut (.I0(\data_out_frame[20] [7]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[7]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4965));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_167_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_4_lut_adj_1635 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[20] [6]), 
            .I2(displacement[6]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4964));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1635.LUT_INIT = 16'ha088;
    SB_LUT4 i14298_1_lut (.I0(n3468), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n28304));   // verilog/coms.v(148[4] 304[11])
    defparam i14298_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_4_lut_adj_1636 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[20] [5]), 
            .I2(displacement[5]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4963));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1636.LUT_INIT = 16'ha088;
    SB_LUT4 i1_4_lut_adj_1637 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[20] [4]), 
            .I2(displacement[4]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4962));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1637.LUT_INIT = 16'ha088;
    SB_LUT4 select_777_Select_5_i1_2_lut_3_lut (.I0(\FRAME_MATCHER.state[3] ), 
            .I1(\FRAME_MATCHER.i_31__N_2511 ), .I2(byte_transmit_counter[5]), 
            .I3(GND_net), .O(n1_adj_5039));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_5_i1_2_lut_3_lut.LUT_INIT = 16'h1010;
    SB_LUT4 select_775_Select_163_i2_4_lut (.I0(\data_out_frame[20] [3]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[3]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4961));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_163_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_775_Select_162_i2_4_lut (.I0(\data_out_frame[20] [2]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[2]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4960));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_162_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_775_Select_161_i2_4_lut (.I0(\data_out_frame[20] [1]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[1]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4959));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_161_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_775_Select_160_i2_4_lut (.I0(\data_out_frame[20] [0]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[0]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4958));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_160_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_775_Select_159_i2_4_lut (.I0(\data_out_frame[19] [7]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[15]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4957));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_159_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_775_Select_158_i2_4_lut (.I0(\data_out_frame[19] [6]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[14]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4955));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_158_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_4_lut_3_lut (.I0(\data_in_frame[3] [3]), .I1(\data_in_frame[3] [1]), 
            .I2(n59250), .I3(GND_net), .O(n6_adj_5095));
    defparam i1_2_lut_4_lut_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1638 (.I0(\data_in_frame[3] [3]), .I1(n58842), 
            .I2(\data_in_frame[5] [5]), .I3(GND_net), .O(n59000));
    defparam i1_2_lut_3_lut_adj_1638.LUT_INIT = 16'h9696;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_55457 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[18] [6]), .I2(\data_out_frame[19] [6]), 
            .I3(\byte_transmit_counter[1] ), .O(n71204));
    defparam byte_transmit_counter_0__bdd_4_lut_55457.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_3_lut_4_lut_adj_1639 (.I0(\data_in_frame[3] [3]), .I1(n58842), 
            .I2(n63789), .I3(n25815), .O(n63793));
    defparam i1_3_lut_4_lut_adj_1639.LUT_INIT = 16'h6996;
    SB_LUT4 n71204_bdd_4_lut (.I0(n71204), .I1(\data_out_frame[17] [6]), 
            .I2(\data_out_frame[16] [6]), .I3(\byte_transmit_counter[1] ), 
            .O(n71207));
    defparam n71204_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_3_lut_4_lut_adj_1640 (.I0(\data_in_frame[1] [2]), .I1(\data_in_frame[1] [1]), 
            .I2(\data_in_frame[1] [0]), .I3(n59250), .O(n35423));   // verilog/coms.v(76[16:34])
    defparam i1_3_lut_4_lut_adj_1640.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1641 (.I0(\data_in_frame[1] [2]), .I1(\data_in_frame[1] [1]), 
            .I2(\data_in_frame[0] [7]), .I3(GND_net), .O(n58842));   // verilog/coms.v(76[16:34])
    defparam i1_2_lut_3_lut_adj_1641.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_4_lut_adj_1642 (.I0(\data_out_frame[23] [6]), .I1(n59253), 
            .I2(n10_adj_4883), .I3(n26716), .O(n59162));
    defparam i1_2_lut_4_lut_adj_1642.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1643 (.I0(\FRAME_MATCHER.i[0] ), .I1(rx_data_ready), 
            .I2(\FRAME_MATCHER.rx_data_ready_prev ), .I3(GND_net), .O(n140));   // verilog/coms.v(156[9:50])
    defparam i1_2_lut_3_lut_adj_1643.LUT_INIT = 16'hfbfb;
    SB_LUT4 i1_2_lut_4_lut_adj_1644 (.I0(n59250), .I1(\data_in_frame[3] [1]), 
            .I2(n58842), .I3(\data_in_frame[5] [2]), .O(n59299));   // verilog/coms.v(88[17:63])
    defparam i1_2_lut_4_lut_adj_1644.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1645 (.I0(\data_out_frame[10] [1]), .I1(\data_out_frame[5] [3]), 
            .I2(\data_out_frame[7] [5]), .I3(\data_out_frame[9] [7]), .O(n6_adj_4880));   // verilog/coms.v(78[16:27])
    defparam i1_2_lut_4_lut_adj_1645.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_55269 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[26] [0]), .I2(\data_out_frame[27] [0]), 
            .I3(\byte_transmit_counter[1] ), .O(n70970));
    defparam byte_transmit_counter_0__bdd_4_lut_55269.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_2_lut_3_lut_adj_1646 (.I0(\data_in_frame[1] [3]), .I1(\data_in_frame[1] [4]), 
            .I2(\data_in_frame[3][5] ), .I3(GND_net), .O(n26368));   // verilog/coms.v(81[16:27])
    defparam i1_2_lut_3_lut_adj_1646.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1647 (.I0(\data_in_frame[1] [3]), .I1(\data_in_frame[1] [4]), 
            .I2(n25786), .I3(GND_net), .O(n59250));   // verilog/coms.v(81[16:27])
    defparam i1_2_lut_3_lut_adj_1647.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1648 (.I0(\data_in_frame[6] [7]), .I1(n25751), 
            .I2(n59302), .I3(\data_in_frame[4] [5]), .O(n26239));   // verilog/coms.v(77[16:43])
    defparam i2_3_lut_4_lut_adj_1648.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1649 (.I0(\data_in_frame[6] [7]), .I1(n25751), 
            .I2(n59153), .I3(n25758), .O(n59247));   // verilog/coms.v(77[16:43])
    defparam i1_2_lut_3_lut_4_lut_adj_1649.LUT_INIT = 16'h6996;
    SB_LUT4 i2_2_lut_3_lut_adj_1650 (.I0(\data_out_frame[15] [0]), .I1(\data_out_frame[15] [1]), 
            .I2(n4_c), .I3(GND_net), .O(n59253));
    defparam i2_2_lut_3_lut_adj_1650.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1651 (.I0(\data_out_frame[8] [5]), .I1(\data_out_frame[8] [3]), 
            .I2(\data_out_frame[8] [2]), .I3(GND_net), .O(n58864));   // verilog/coms.v(88[17:28])
    defparam i1_2_lut_3_lut_adj_1651.LUT_INIT = 16'h9696;
    SB_LUT4 n70970_bdd_4_lut (.I0(n70970), .I1(\data_out_frame[25] [0]), 
            .I2(\data_out_frame[24] [0]), .I3(\byte_transmit_counter[1] ), 
            .O(n70973));
    defparam n70970_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_55256 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[26] [7]), .I2(\data_out_frame[27] [7]), 
            .I3(\byte_transmit_counter[1] ), .O(n70964));
    defparam byte_transmit_counter_0__bdd_4_lut_55256.LUT_INIT = 16'he4aa;
    SB_LUT4 n70964_bdd_4_lut (.I0(n70964), .I1(\data_out_frame[25] [7]), 
            .I2(\data_out_frame[24] [7]), .I3(\byte_transmit_counter[1] ), 
            .O(n70967));
    defparam n70964_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_55251 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[26] [6]), .I2(\data_out_frame[27] [6]), 
            .I3(\byte_transmit_counter[1] ), .O(n70958));
    defparam byte_transmit_counter_0__bdd_4_lut_55251.LUT_INIT = 16'he4aa;
    SB_LUT4 n70958_bdd_4_lut (.I0(n70958), .I1(\data_out_frame[25] [6]), 
            .I2(\data_out_frame[24] [6]), .I3(\byte_transmit_counter[1] ), 
            .O(n70961));
    defparam n70958_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_3_lut_adj_1652 (.I0(\data_out_frame[6] [0]), .I1(\data_out_frame[5] [7]), 
            .I2(\data_out_frame[5] [6]), .I3(GND_net), .O(n59335));   // verilog/coms.v(88[17:28])
    defparam i1_2_lut_3_lut_adj_1652.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1653 (.I0(\data_out_frame[12] [4]), .I1(\data_out_frame[12] [5]), 
            .I2(\data_out_frame[14] [6]), .I3(n26049), .O(n26716));   // verilog/coms.v(88[17:63])
    defparam i2_3_lut_4_lut_adj_1653.LUT_INIT = 16'h6996;
    SB_LUT4 i2_2_lut_3_lut_adj_1654 (.I0(\data_in_frame[8] [4]), .I1(n58824), 
            .I2(n58922), .I3(GND_net), .O(n25892));   // verilog/coms.v(88[17:28])
    defparam i2_2_lut_3_lut_adj_1654.LUT_INIT = 16'h9696;
    SB_LUT4 select_775_Select_65_i2_4_lut (.I0(\data_out_frame[8] [1]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder0_position_scaled[1]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5046));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_65_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_55467 (.I0(byte_transmit_counter[3]), 
            .I1(n69187), .I2(n67140), .I3(byte_transmit_counter[4]), .O(n71198));
    defparam byte_transmit_counter_3__bdd_4_lut_55467.LUT_INIT = 16'he4aa;
    SB_LUT4 select_775_Select_64_i2_4_lut (.I0(\data_out_frame[8] [0]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder0_position_scaled[0]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5045));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_64_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1655 (.I0(\data_in_frame[8] [4]), .I1(n58824), 
            .I2(\data_in_frame[8] [3]), .I3(n25878), .O(n58836));   // verilog/coms.v(88[17:28])
    defparam i1_2_lut_3_lut_4_lut_adj_1655.LUT_INIT = 16'h6996;
    SB_LUT4 n71198_bdd_4_lut (.I0(n71198), .I1(n70937), .I2(n71027), .I3(byte_transmit_counter[4]), 
            .O(tx_data[4]));
    defparam n71198_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i2_3_lut_4_lut_adj_1656 (.I0(\data_in_frame[1] [5]), .I1(\data_in_frame[5] [7]), 
            .I2(n26368), .I3(n59320), .O(n25878));   // verilog/coms.v(81[16:27])
    defparam i2_3_lut_4_lut_adj_1656.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1657 (.I0(\data_in_frame[1] [5]), .I1(\data_in_frame[5] [7]), 
            .I2(\data_in_frame[5] [6]), .I3(GND_net), .O(n6_adj_5093));   // verilog/coms.v(81[16:27])
    defparam i1_2_lut_3_lut_adj_1657.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1658 (.I0(\FRAME_MATCHER.state[3] ), .I1(\FRAME_MATCHER.i_31__N_2511 ), 
            .I2(byte_transmit_counter[4]), .I3(GND_net), .O(n1_adj_5038));   // verilog/coms.v(148[4] 304[11])
    defparam i1_2_lut_3_lut_adj_1658.LUT_INIT = 16'h1010;
    SB_LUT4 i1_2_lut_3_lut_adj_1659 (.I0(\FRAME_MATCHER.state[3] ), .I1(\FRAME_MATCHER.i_31__N_2511 ), 
            .I2(\byte_transmit_counter[2] ), .I3(GND_net), .O(n1_adj_5036));   // verilog/coms.v(148[4] 304[11])
    defparam i1_2_lut_3_lut_adj_1659.LUT_INIT = 16'h1010;
    SB_LUT4 i2_3_lut_4_lut_adj_1660 (.I0(n25758), .I1(n59153), .I2(n59365), 
            .I3(n59064), .O(Kp_23__N_993));   // verilog/coms.v(78[16:43])
    defparam i2_3_lut_4_lut_adj_1660.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1661 (.I0(\data_out_frame[4] [3]), .I1(\data_out_frame[6] [4]), 
            .I2(\data_out_frame[8] [6]), .I3(\data_out_frame[4] [2]), .O(n36));   // verilog/coms.v(77[16:27])
    defparam i1_2_lut_4_lut_adj_1661.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1662 (.I0(n26368), .I1(n59134), .I2(\data_in_frame[5] [6]), 
            .I3(n54308), .O(n6_adj_5075));
    defparam i1_2_lut_4_lut_adj_1662.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_4_lut_adj_1663 (.I0(n26368), .I1(n59134), .I2(\data_in_frame[5] [6]), 
            .I3(n25860), .O(n54404));
    defparam i1_2_lut_4_lut_adj_1663.LUT_INIT = 16'h9669;
    SB_LUT4 i2_2_lut_3_lut_adj_1664 (.I0(n25878), .I1(\data_in_frame[8] [3]), 
            .I2(n58922), .I3(GND_net), .O(n4_adj_5072));   // verilog/coms.v(239[9:81])
    defparam i2_2_lut_3_lut_adj_1664.LUT_INIT = 16'h9696;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_55246 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[22] [6]), .I2(\data_out_frame[23] [6]), 
            .I3(\byte_transmit_counter[1] ), .O(n70952));
    defparam byte_transmit_counter_0__bdd_4_lut_55246.LUT_INIT = 16'he4aa;
    SB_LUT4 i5_3_lut_4_lut_adj_1665 (.I0(\data_in_frame[6] [5]), .I1(Kp_23__N_878), 
            .I2(\data_in_frame[6] [6]), .I3(n10_adj_5083), .O(n25906));   // verilog/coms.v(78[16:43])
    defparam i5_3_lut_4_lut_adj_1665.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1666 (.I0(\data_in_frame[6] [5]), .I1(Kp_23__N_878), 
            .I2(n58818), .I3(GND_net), .O(Kp_23__N_974));   // verilog/coms.v(78[16:43])
    defparam i1_2_lut_3_lut_adj_1666.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1667 (.I0(n53933), .I1(n58987), .I2(n25142), 
            .I3(GND_net), .O(n59338));
    defparam i1_2_lut_3_lut_adj_1667.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1668 (.I0(\FRAME_MATCHER.state[3] ), .I1(\FRAME_MATCHER.i_31__N_2511 ), 
            .I2(byte_transmit_counter[3]), .I3(GND_net), .O(n1_adj_5037));   // verilog/coms.v(148[4] 304[11])
    defparam i1_2_lut_3_lut_adj_1668.LUT_INIT = 16'h1010;
    SB_LUT4 i2_2_lut_3_lut_adj_1669 (.I0(n53933), .I1(n58987), .I2(n54570), 
            .I3(GND_net), .O(n6_adj_4760));
    defparam i2_2_lut_3_lut_adj_1669.LUT_INIT = 16'h9696;
    SB_LUT4 n70952_bdd_4_lut (.I0(n70952), .I1(\data_out_frame[21] [6]), 
            .I2(\data_out_frame[20] [6]), .I3(\byte_transmit_counter[1] ), 
            .O(n70955));
    defparam n70952_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_3_lut_adj_1670 (.I0(\data_in_frame[13] [3]), .I1(\data_in_frame[13] [4]), 
            .I2(\data_in_frame[13] [1]), .I3(GND_net), .O(n59284));   // verilog/coms.v(88[17:63])
    defparam i1_2_lut_3_lut_adj_1670.LUT_INIT = 16'h9696;
    SB_LUT4 i1_4_lut_3_lut (.I0(n54520), .I1(n63749), .I2(n7_adj_5094), 
            .I3(GND_net), .O(n53570));
    defparam i1_4_lut_3_lut.LUT_INIT = 16'h6969;
    SB_LUT4 i1_2_lut_3_lut_adj_1671 (.I0(Kp_23__N_1080), .I1(n54520), .I2(n54002), 
            .I3(GND_net), .O(n54518));
    defparam i1_2_lut_3_lut_adj_1671.LUT_INIT = 16'h6969;
    SB_LUT4 i2_3_lut_4_lut_adj_1672 (.I0(n25860), .I1(n59000), .I2(\data_in_frame[8] [0]), 
            .I3(n58799), .O(n59259));
    defparam i2_3_lut_4_lut_adj_1672.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1673 (.I0(n25860), .I1(n59000), .I2(\data_in_frame[7]_c [7]), 
            .I3(n59134), .O(n54308));
    defparam i2_3_lut_4_lut_adj_1673.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1674 (.I0(\data_in_frame[11] [0]), .I1(\data_in_frame[10] [7]), 
            .I2(\data_in_frame[13] [2]), .I3(n59468), .O(n59165));   // verilog/coms.v(74[16:27])
    defparam i2_3_lut_4_lut_adj_1674.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1675 (.I0(\data_in_frame[11] [0]), .I1(\data_in_frame[10] [7]), 
            .I2(n59487), .I3(GND_net), .O(n58851));   // verilog/coms.v(74[16:27])
    defparam i1_2_lut_3_lut_adj_1675.LUT_INIT = 16'h9696;
    SB_LUT4 i15921_3_lut_4_lut (.I0(n8_adj_5096), .I1(n58760), .I2(rx_data[7]), 
            .I3(\data_in_frame[6] [7]), .O(n29927));
    defparam i15921_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15918_3_lut_4_lut (.I0(n8_adj_5096), .I1(n58760), .I2(rx_data[6]), 
            .I3(\data_in_frame[6] [6]), .O(n29924));
    defparam i15918_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15915_3_lut_4_lut (.I0(n8_adj_5096), .I1(n58760), .I2(rx_data[5]), 
            .I3(\data_in_frame[6] [5]), .O(n29921));
    defparam i15915_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15912_3_lut_4_lut (.I0(n8_adj_5096), .I1(n58760), .I2(rx_data[4]), 
            .I3(\data_in_frame[6] [4]), .O(n29918));
    defparam i15912_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_55447 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[18] [1]), .I2(\data_out_frame[19] [1]), 
            .I3(\byte_transmit_counter[1] ), .O(n71186));
    defparam byte_transmit_counter_0__bdd_4_lut_55447.LUT_INIT = 16'he4aa;
    SB_LUT4 i15908_3_lut_4_lut (.I0(n8_adj_5096), .I1(n58760), .I2(rx_data[3]), 
            .I3(\data_in_frame[6] [3]), .O(n29914));
    defparam i15908_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15905_3_lut_4_lut (.I0(n8_adj_5096), .I1(n58760), .I2(rx_data[2]), 
            .I3(\data_in_frame[6] [2]), .O(n29911));
    defparam i15905_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15902_3_lut_4_lut (.I0(n8_adj_5096), .I1(n58760), .I2(rx_data[1]), 
            .I3(\data_in_frame[6] [1]), .O(n29908));
    defparam i15902_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15898_3_lut_4_lut (.I0(n8_adj_5096), .I1(n58760), .I2(rx_data[0]), 
            .I3(\data_in_frame[6] [0]), .O(n29904));
    defparam i15898_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_4_lut_adj_1676 (.I0(\data_out_frame[11] [6]), .I1(n25614), 
            .I2(n58931), .I3(n26039), .O(n59012));
    defparam i1_2_lut_4_lut_adj_1676.LUT_INIT = 16'h6996;
    SB_LUT4 n71186_bdd_4_lut (.I0(n71186), .I1(\data_out_frame[17] [1]), 
            .I2(\data_out_frame[16] [1]), .I3(\byte_transmit_counter[1] ), 
            .O(n71189));
    defparam n71186_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_3_lut_adj_1677 (.I0(\data_out_frame[5] [3]), .I1(\data_out_frame[4] [7]), 
            .I2(\data_out_frame[7] [3]), .I3(GND_net), .O(n6_adj_4865));   // verilog/coms.v(76[16:34])
    defparam i1_2_lut_3_lut_adj_1677.LUT_INIT = 16'h9696;
    SB_LUT4 i14373_3_lut_4_lut (.I0(n161_c), .I1(n58731), .I2(reset), 
            .I3(n8_adj_4950), .O(n7_adj_18));
    defparam i14373_3_lut_4_lut.LUT_INIT = 16'hfffd;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_55284 (.I0(\byte_transmit_counter[1] ), 
            .I1(n64367), .I2(n64368), .I3(\byte_transmit_counter[2] ), 
            .O(n70946));
    defparam byte_transmit_counter_1__bdd_4_lut_55284.LUT_INIT = 16'he4aa;
    SB_LUT4 i14379_3_lut_4_lut (.I0(n161_c), .I1(n58731), .I2(reset), 
            .I3(n8_adj_12), .O(n28385));
    defparam i14379_3_lut_4_lut.LUT_INIT = 16'hfffd;
    SB_LUT4 n70946_bdd_4_lut (.I0(n70946), .I1(n64488), .I2(n64487), .I3(\byte_transmit_counter[2] ), 
            .O(n70949));
    defparam n70946_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i2_3_lut_4_lut_adj_1678 (.I0(n59067), .I1(n59232), .I2(n54411), 
            .I3(n25853), .O(n54475));
    defparam i2_3_lut_4_lut_adj_1678.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1679 (.I0(n59067), .I1(n59232), .I2(\data_in_frame[16] [3]), 
            .I3(GND_net), .O(n59183));
    defparam i1_2_lut_3_lut_adj_1679.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1680 (.I0(\data_in_frame[14] [2]), .I1(n54468), 
            .I2(\data_in_frame[16] [4]), .I3(GND_net), .O(n59232));
    defparam i1_2_lut_3_lut_adj_1680.LUT_INIT = 16'h6969;
    SB_LUT4 i1_2_lut_3_lut_adj_1681 (.I0(\data_in_frame[14] [2]), .I1(n54468), 
            .I2(n53503), .I3(GND_net), .O(n54447));
    defparam i1_2_lut_3_lut_adj_1681.LUT_INIT = 16'h6969;
    SB_LUT4 i15995_3_lut_4_lut (.I0(n8_adj_15), .I1(n58755), .I2(rx_data[7]), 
            .I3(\data_in_frame[9] [7]), .O(n30001));
    defparam i15995_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15992_3_lut_4_lut (.I0(n8_adj_15), .I1(n58755), .I2(rx_data[6]), 
            .I3(\data_in_frame[9] [6]), .O(n29998));
    defparam i15992_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15989_3_lut_4_lut (.I0(n8_adj_15), .I1(n58755), .I2(rx_data[5]), 
            .I3(\data_in_frame[9] [5]), .O(n29995));
    defparam i15989_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15986_3_lut_4_lut (.I0(n8_adj_15), .I1(n58755), .I2(rx_data[4]), 
            .I3(\data_in_frame[9] [4]), .O(n29992));
    defparam i15986_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15983_3_lut_4_lut (.I0(n8_adj_15), .I1(n58755), .I2(rx_data[3]), 
            .I3(\data_in_frame[9] [3]), .O(n29989));
    defparam i15983_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15979_3_lut_4_lut (.I0(n8_adj_15), .I1(n58755), .I2(rx_data[2]), 
            .I3(\data_in_frame[9] [2]), .O(n29985));
    defparam i15979_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15976_3_lut_4_lut (.I0(n8_adj_15), .I1(n58755), .I2(rx_data[1]), 
            .I3(\data_in_frame[9] [1]), .O(n29982));
    defparam i15976_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_55236 (.I0(\byte_transmit_counter[1] ), 
            .I1(n64400), .I2(n64401), .I3(\byte_transmit_counter[2] ), 
            .O(n70940));
    defparam byte_transmit_counter_1__bdd_4_lut_55236.LUT_INIT = 16'he4aa;
    SB_LUT4 i15973_3_lut_4_lut (.I0(n8_adj_15), .I1(n58755), .I2(rx_data[0]), 
            .I3(\data_in_frame[9] [0]), .O(n29979));
    defparam i15973_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16021_3_lut_4_lut (.I0(n8_adj_13), .I1(n58755), .I2(rx_data[7]), 
            .I3(\data_in_frame[10] [7]), .O(n30027));
    defparam i16021_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16017_3_lut_4_lut (.I0(n8_adj_13), .I1(n58755), .I2(rx_data[6]), 
            .I3(\data_in_frame[10] [6]), .O(n30023));
    defparam i16017_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16014_3_lut_4_lut (.I0(n8_adj_13), .I1(n58755), .I2(rx_data[5]), 
            .I3(\data_in_frame[10] [5]), .O(n30020));
    defparam i16014_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16011_3_lut_4_lut (.I0(n8_adj_13), .I1(n58755), .I2(rx_data[4]), 
            .I3(\data_in_frame[10] [4]), .O(n30017));
    defparam i16011_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 n70940_bdd_4_lut (.I0(n70940), .I1(n64485), .I2(n64484), .I3(\byte_transmit_counter[2] ), 
            .O(n70943));
    defparam n70940_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i16007_3_lut_4_lut (.I0(n8_adj_13), .I1(n58755), .I2(rx_data[3]), 
            .I3(\data_in_frame[10] [3]), .O(n30013));
    defparam i16007_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i54326_3_lut_4_lut (.I0(n53515), .I1(\data_out_frame[14] [3]), 
            .I2(n54114), .I3(n59010), .O(n70020));
    defparam i54326_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i16004_3_lut_4_lut (.I0(n8_adj_13), .I1(n58755), .I2(rx_data[2]), 
            .I3(\data_in_frame[10] [2]), .O(n30010));
    defparam i16004_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16001_3_lut_4_lut (.I0(n8_adj_13), .I1(n58755), .I2(rx_data[1]), 
            .I3(\data_in_frame[10] [1]), .O(n30007));
    defparam i16001_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15998_3_lut_4_lut (.I0(n8_adj_13), .I1(n58755), .I2(rx_data[0]), 
            .I3(\data_in_frame[10] [0]), .O(n30004));
    defparam i15998_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1682 (.I0(n53031), .I1(n25455), .I2(\FRAME_MATCHER.i_31__N_2513 ), 
            .I3(GND_net), .O(n33697));   // verilog/coms.v(241[12:32])
    defparam i1_2_lut_3_lut_adj_1682.LUT_INIT = 16'h4040;
    SB_LUT4 select_775_Select_157_i2_4_lut (.I0(\data_out_frame[19] [5]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[13]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4948));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_157_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_55231 (.I0(\byte_transmit_counter[1] ), 
            .I1(n64457), .I2(n64458), .I3(\byte_transmit_counter[2] ), 
            .O(n70934));
    defparam byte_transmit_counter_1__bdd_4_lut_55231.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_2_lut_4_lut_adj_1683 (.I0(\data_out_frame[16] [0]), .I1(\data_out_frame[15] [5]), 
            .I2(n54220), .I3(n26210), .O(n54620));
    defparam i1_2_lut_4_lut_adj_1683.LUT_INIT = 16'h6996;
    SB_LUT4 n70934_bdd_4_lut (.I0(n70934), .I1(n64473), .I2(n64472), .I3(\byte_transmit_counter[2] ), 
            .O(n70937));
    defparam n70934_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_3_lut_adj_1684 (.I0(n53031), .I1(n25455), .I2(LED_c), 
            .I3(GND_net), .O(n33_adj_5126));   // verilog/coms.v(241[12:32])
    defparam i1_2_lut_3_lut_adj_1684.LUT_INIT = 16'hf4f4;
    SB_LUT4 i1_2_lut_3_lut_adj_1685 (.I0(Kp_23__N_1748), .I1(n37), .I2(n33693), 
            .I3(GND_net), .O(n5));   // verilog/coms.v(148[4] 304[11])
    defparam i1_2_lut_3_lut_adj_1685.LUT_INIT = 16'hf8f8;
    SB_LUT4 select_775_Select_156_i2_4_lut (.I0(\data_out_frame[19] [4]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[12]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4947));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_156_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i23370_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n37), .I2(\data_in_frame[16] [0]), 
            .I3(deadband[0]), .O(n29406));   // verilog/coms.v(148[4] 304[11])
    defparam i23370_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_55241 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[22] [1]), .I2(\data_out_frame[23] [1]), 
            .I3(\byte_transmit_counter[1] ), .O(n70928));
    defparam byte_transmit_counter_0__bdd_4_lut_55241.LUT_INIT = 16'he4aa;
    SB_LUT4 mux_1052_i2_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n37), .I2(\data_in_frame[3] [1]), 
            .I3(\data_in_frame[19] [1]), .O(n4760[1]));   // verilog/coms.v(148[4] 304[11])
    defparam mux_1052_i2_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 i1_2_lut_4_lut_adj_1686 (.I0(\data_out_frame[12] [2]), .I1(n1510), 
            .I2(\data_out_frame[12] [1]), .I3(n25052), .O(n54114));
    defparam i1_2_lut_4_lut_adj_1686.LUT_INIT = 16'h6996;
    SB_LUT4 mux_1052_i3_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n37), .I2(\data_in_frame[3] [2]), 
            .I3(\data_in_frame[19] [2]), .O(n4760[2]));   // verilog/coms.v(148[4] 304[11])
    defparam mux_1052_i3_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 mux_1052_i4_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n37), .I2(\data_in_frame[3] [3]), 
            .I3(\data_in_frame[19] [3]), .O(n4760[3]));   // verilog/coms.v(148[4] 304[11])
    defparam mux_1052_i4_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 mux_1052_i5_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n37), .I2(\data_in_frame[3] [4]), 
            .I3(\data_in_frame[19] [4]), .O(n4760[4]));   // verilog/coms.v(148[4] 304[11])
    defparam mux_1052_i5_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 mux_1052_i6_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n37), .I2(\data_in_frame[3][5] ), 
            .I3(\data_in_frame[19] [5]), .O(n4760[5]));   // verilog/coms.v(148[4] 304[11])
    defparam mux_1052_i6_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 i2_3_lut_4_lut_adj_1687 (.I0(\data_out_frame[7] [6]), .I1(\data_out_frame[7] [5]), 
            .I2(n59323), .I3(\data_out_frame[11] [7]), .O(n25052));   // verilog/coms.v(78[16:27])
    defparam i2_3_lut_4_lut_adj_1687.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1688 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[19] [3]), 
            .I2(displacement[11]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4940));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1688.LUT_INIT = 16'ha088;
    SB_LUT4 mux_1052_i7_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n37), .I2(\data_in_frame[3][6] ), 
            .I3(\data_in_frame[19] [6]), .O(n4760[6]));   // verilog/coms.v(148[4] 304[11])
    defparam mux_1052_i7_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 i21811_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n37), .I2(\data_in_frame[3] [7]), 
            .I3(\data_in_frame[19] [7]), .O(n4760[7]));   // verilog/coms.v(148[4] 304[11])
    defparam i21811_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 n70928_bdd_4_lut (.I0(n70928), .I1(\data_out_frame[21] [1]), 
            .I2(\data_out_frame[20] [1]), .I3(\byte_transmit_counter[1] ), 
            .O(n70931));
    defparam n70928_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 mux_1052_i9_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n37), .I2(\data_in_frame[2] [0]), 
            .I3(\data_in_frame[18] [0]), .O(n4760[8]));   // verilog/coms.v(148[4] 304[11])
    defparam mux_1052_i9_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 mux_1052_i10_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n37), .I2(\data_in_frame[2] [1]), 
            .I3(\data_in_frame[18] [1]), .O(n4760[9]));   // verilog/coms.v(148[4] 304[11])
    defparam mux_1052_i10_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 mux_1052_i11_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n37), .I2(\data_in_frame[2] [2]), 
            .I3(\data_in_frame[18] [2]), .O(n4760[10]));   // verilog/coms.v(148[4] 304[11])
    defparam mux_1052_i11_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 mux_1052_i12_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n37), .I2(\data_in_frame[2] [3]), 
            .I3(\data_in_frame[18] [3]), .O(n4760[11]));   // verilog/coms.v(148[4] 304[11])
    defparam mux_1052_i12_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 mux_1052_i13_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n37), .I2(\data_in_frame[2] [4]), 
            .I3(\data_in_frame[18] [4]), .O(n4760[12]));   // verilog/coms.v(148[4] 304[11])
    defparam mux_1052_i13_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 byte_transmit_counter_2__bdd_4_lut (.I0(\byte_transmit_counter[2] ), 
            .I1(n64471), .I2(n64480), .I3(byte_transmit_counter[3]), .O(n70922));
    defparam byte_transmit_counter_2__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 mux_1052_i14_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n37), .I2(\data_in_frame[2] [5]), 
            .I3(\data_in_frame[18] [5]), .O(n4760[13]));   // verilog/coms.v(148[4] 304[11])
    defparam mux_1052_i14_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 n70922_bdd_4_lut (.I0(n70922), .I1(n64383), .I2(n64382), .I3(byte_transmit_counter[3]), 
            .O(n70925));
    defparam n70922_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 mux_1052_i15_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n37), .I2(\data_in_frame[2] [6]), 
            .I3(\data_in_frame[18] [6]), .O(n4760[14]));   // verilog/coms.v(148[4] 304[11])
    defparam mux_1052_i15_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 select_775_Select_63_i2_4_lut (.I0(\data_out_frame[7] [7]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder0_position_scaled[15]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5044));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_63_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 mux_1052_i16_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n37), .I2(\data_in_frame[2] [7]), 
            .I3(\data_in_frame[18] [7]), .O(n4760[15]));   // verilog/coms.v(148[4] 304[11])
    defparam mux_1052_i16_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 mux_1052_i17_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n37), .I2(\data_in_frame[1] [0]), 
            .I3(\data_in_frame[17] [0]), .O(n4760[16]));   // verilog/coms.v(148[4] 304[11])
    defparam mux_1052_i17_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 mux_1052_i18_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n37), .I2(\data_in_frame[1] [1]), 
            .I3(\data_in_frame[17] [1]), .O(n4760[17]));   // verilog/coms.v(148[4] 304[11])
    defparam mux_1052_i18_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 mux_1052_i19_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n37), .I2(\data_in_frame[1] [2]), 
            .I3(\data_in_frame[17] [2]), .O(n4760[18]));   // verilog/coms.v(148[4] 304[11])
    defparam mux_1052_i19_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 mux_1052_i20_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n37), .I2(\data_in_frame[1] [3]), 
            .I3(\data_in_frame[17] [3]), .O(n4760[19]));   // verilog/coms.v(148[4] 304[11])
    defparam mux_1052_i20_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 mux_1052_i21_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n37), .I2(\data_in_frame[1] [4]), 
            .I3(\data_in_frame[17] [4]), .O(n4760[20]));   // verilog/coms.v(148[4] 304[11])
    defparam mux_1052_i21_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 i1_2_lut_4_lut_adj_1689 (.I0(n26716), .I1(\data_out_frame[16] [6]), 
            .I2(n26817), .I3(n59244), .O(n54450));
    defparam i1_2_lut_4_lut_adj_1689.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1690 (.I0(n26716), .I1(\data_out_frame[16] [6]), 
            .I2(n26817), .I3(GND_net), .O(n25678));   // verilog/coms.v(88[17:28])
    defparam i1_2_lut_3_lut_adj_1690.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1691 (.I0(\data_out_frame[14] [4]), .I1(n59124), 
            .I2(n70022), .I3(GND_net), .O(n59353));
    defparam i1_2_lut_3_lut_adj_1691.LUT_INIT = 16'h6969;
    SB_LUT4 i54328_2_lut_3_lut (.I0(n53515), .I1(\data_out_frame[18] [7]), 
            .I2(\data_out_frame[18] [6]), .I3(GND_net), .O(n70022));
    defparam i54328_2_lut_3_lut.LUT_INIT = 16'h6969;
    SB_LUT4 i1_2_lut_4_lut_adj_1692 (.I0(n26376), .I1(n36), .I2(\data_out_frame[10] [7]), 
            .I3(n59462), .O(n6_adj_4822));   // verilog/coms.v(77[16:27])
    defparam i1_2_lut_4_lut_adj_1692.LUT_INIT = 16'h6996;
    SB_LUT4 mux_1052_i22_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n37), .I2(\data_in_frame[1] [5]), 
            .I3(\data_in_frame[17] [5]), .O(n4760[21]));   // verilog/coms.v(148[4] 304[11])
    defparam mux_1052_i22_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 select_775_Select_62_i2_4_lut (.I0(\data_out_frame[7] [6]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder0_position_scaled[14]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5043));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_62_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_55222 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[26] [4]), .I2(\data_out_frame[27] [4]), 
            .I3(\byte_transmit_counter[1] ), .O(n70916));
    defparam byte_transmit_counter_0__bdd_4_lut_55222.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_2_lut_3_lut_adj_1693 (.I0(\data_out_frame[13] [6]), .I1(n26347), 
            .I2(n53470), .I3(GND_net), .O(n54432));
    defparam i1_2_lut_3_lut_adj_1693.LUT_INIT = 16'h9696;
    SB_LUT4 n70916_bdd_4_lut (.I0(n70916), .I1(\data_out_frame[25] [4]), 
            .I2(\data_out_frame[24] [4]), .I3(\byte_transmit_counter[1] ), 
            .O(n70919));
    defparam n70916_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_4_lut_adj_1694 (.I0(\data_out_frame[16] [3]), .I1(n59455), 
            .I2(\data_out_frame[16] [4]), .I3(n59424), .O(n6_adj_4791));
    defparam i1_2_lut_4_lut_adj_1694.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_55213 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[26] [1]), .I2(\data_out_frame[27] [1]), 
            .I3(\byte_transmit_counter[1] ), .O(n70910));
    defparam byte_transmit_counter_0__bdd_4_lut_55213.LUT_INIT = 16'he4aa;
    SB_LUT4 n70910_bdd_4_lut (.I0(n70910), .I1(\data_out_frame[25] [1]), 
            .I2(\data_out_frame[24] [1]), .I3(\byte_transmit_counter[1] ), 
            .O(n70913));
    defparam n70910_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_55208 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[26] [3]), .I2(\data_out_frame[27] [3]), 
            .I3(\byte_transmit_counter[1] ), .O(n70904));
    defparam byte_transmit_counter_0__bdd_4_lut_55208.LUT_INIT = 16'he4aa;
    SB_LUT4 n70904_bdd_4_lut (.I0(n70904), .I1(\data_out_frame[25] [3]), 
            .I2(\data_out_frame[24] [3]), .I3(\byte_transmit_counter[1] ), 
            .O(n70907));
    defparam n70904_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_4_lut_adj_1695 (.I0(n25650), .I1(\data_out_frame[15] [5]), 
            .I2(n54220), .I3(\data_out_frame[15] [4]), .O(n54552));
    defparam i1_2_lut_4_lut_adj_1695.LUT_INIT = 16'h6996;
    SB_LUT4 mux_1052_i23_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n37), .I2(\data_in_frame[1] [6]), 
            .I3(\data_in_frame[17] [6]), .O(n4760[22]));   // verilog/coms.v(148[4] 304[11])
    defparam mux_1052_i23_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 mux_1052_i24_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n37), .I2(\data_in_frame[1] [7]), 
            .I3(\data_in_frame[17] [7]), .O(n4760[23]));   // verilog/coms.v(148[4] 304[11])
    defparam mux_1052_i24_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 i16254_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n37), .I2(\data_in_frame[8] [7]), 
            .I3(PWMLimit[23]), .O(n30260));   // verilog/coms.v(148[4] 304[11])
    defparam i16254_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_55203 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[26] [5]), .I2(\data_out_frame[27] [5]), 
            .I3(\byte_transmit_counter[1] ), .O(n70898));
    defparam byte_transmit_counter_0__bdd_4_lut_55203.LUT_INIT = 16'he4aa;
    SB_LUT4 n70898_bdd_4_lut (.I0(n70898), .I1(\data_out_frame[25] [5]), 
            .I2(\data_out_frame[24] [5]), .I3(\byte_transmit_counter[1] ), 
            .O(n70901));
    defparam n70898_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i16258_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n37), .I2(\data_in_frame[8] [6]), 
            .I3(PWMLimit[22]), .O(n30264));   // verilog/coms.v(148[4] 304[11])
    defparam i16258_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_55198 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[14] [1]), .I2(\data_out_frame[15] [1]), 
            .I3(\byte_transmit_counter[1] ), .O(n70892));
    defparam byte_transmit_counter_0__bdd_4_lut_55198.LUT_INIT = 16'he4aa;
    SB_LUT4 n70892_bdd_4_lut (.I0(n70892), .I1(\data_out_frame[13] [1]), 
            .I2(\data_out_frame[12] [1]), .I3(\byte_transmit_counter[1] ), 
            .O(n70895));
    defparam n70892_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i16262_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n37), .I2(\data_in_frame[8] [5]), 
            .I3(PWMLimit[21]), .O(n30268));   // verilog/coms.v(148[4] 304[11])
    defparam i16262_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i23888_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n37), .I2(\data_in_frame[8] [4]), 
            .I3(PWMLimit[20]), .O(n30271));   // verilog/coms.v(148[4] 304[11])
    defparam i23888_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2_3_lut_4_lut_adj_1696 (.I0(n26347), .I1(n26649), .I2(\data_out_frame[13] [7]), 
            .I3(\data_out_frame[13] [6]), .O(n59186));
    defparam i2_3_lut_4_lut_adj_1696.LUT_INIT = 16'h6996;
    SB_LUT4 i16268_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n37), .I2(\data_in_frame[8] [3]), 
            .I3(PWMLimit[19]), .O(n30274));   // verilog/coms.v(148[4] 304[11])
    defparam i16268_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_2_lut_3_lut_adj_1697 (.I0(\FRAME_MATCHER.state[3] ), .I1(\FRAME_MATCHER.i_31__N_2511 ), 
            .I2(\byte_transmit_counter[1] ), .I3(GND_net), .O(n1_adj_5035));   // verilog/coms.v(148[4] 304[11])
    defparam i1_2_lut_3_lut_adj_1697.LUT_INIT = 16'h1010;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_55193 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[14] [5]), .I2(\data_out_frame[15] [5]), 
            .I3(\byte_transmit_counter[1] ), .O(n70886));
    defparam byte_transmit_counter_0__bdd_4_lut_55193.LUT_INIT = 16'he4aa;
    SB_LUT4 i2_3_lut_4_lut_adj_1698 (.I0(\data_out_frame[18] [4]), .I1(n53707), 
            .I2(\data_out_frame[16] [4]), .I3(n59055), .O(n59452));
    defparam i2_3_lut_4_lut_adj_1698.LUT_INIT = 16'h6996;
    SB_LUT4 i16269_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n37), .I2(\data_in_frame[8] [2]), 
            .I3(PWMLimit[18]), .O(n30275));   // verilog/coms.v(148[4] 304[11])
    defparam i16269_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i16308_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n37), .I2(\data_in_frame[8] [1]), 
            .I3(PWMLimit[17]), .O(n30314));   // verilog/coms.v(148[4] 304[11])
    defparam i16308_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i16314_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n37), .I2(\data_in_frame[8] [0]), 
            .I3(PWMLimit[16]), .O(n30320));   // verilog/coms.v(148[4] 304[11])
    defparam i16314_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n70886_bdd_4_lut (.I0(n70886), .I1(\data_out_frame[13] [5]), 
            .I2(\data_out_frame[12] [5]), .I3(\byte_transmit_counter[1] ), 
            .O(n70889));
    defparam n70886_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i2_3_lut_4_lut_adj_1699 (.I0(n53707), .I1(n59074), .I2(\data_out_frame[18] [4]), 
            .I3(\data_out_frame[18] [3]), .O(n61261));
    defparam i2_3_lut_4_lut_adj_1699.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1700 (.I0(\data_out_frame[18] [4]), .I1(n53707), 
            .I2(\data_out_frame[20] [0]), .I3(GND_net), .O(n6_adj_4801));
    defparam i1_2_lut_3_lut_adj_1700.LUT_INIT = 16'h9696;
    SB_LUT4 i20838_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n37), .I2(\data_in_frame[9] [7]), 
            .I3(PWMLimit[15]), .O(n30321));   // verilog/coms.v(148[4] 304[11])
    defparam i20838_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i16316_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n37), .I2(\data_in_frame[9] [6]), 
            .I3(PWMLimit[14]), .O(n30322));   // verilog/coms.v(148[4] 304[11])
    defparam i16316_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_55188 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[18] [0]), .I2(\data_out_frame[19] [0]), 
            .I3(\byte_transmit_counter[1] ), .O(n70880));
    defparam byte_transmit_counter_0__bdd_4_lut_55188.LUT_INIT = 16'he4aa;
    SB_LUT4 i16343_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n37), .I2(\data_in_frame[9] [5]), 
            .I3(PWMLimit[13]), .O(n30349));   // verilog/coms.v(148[4] 304[11])
    defparam i16343_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n70880_bdd_4_lut (.I0(n70880), .I1(\data_out_frame[17] [0]), 
            .I2(\data_out_frame[16] [0]), .I3(\byte_transmit_counter[1] ), 
            .O(n70883));
    defparam n70880_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i16367_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n37), .I2(\data_in_frame[9] [4]), 
            .I3(PWMLimit[12]), .O(n30373));   // verilog/coms.v(148[4] 304[11])
    defparam i16367_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_2_lut_4_lut_adj_1701 (.I0(n60980), .I1(n26347), .I2(n26649), 
            .I3(n1699), .O(n54434));
    defparam i1_2_lut_4_lut_adj_1701.LUT_INIT = 16'h9669;
    SB_LUT4 i16382_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n37), .I2(\data_in_frame[9] [3]), 
            .I3(PWMLimit[11]), .O(n30388));   // verilog/coms.v(148[4] 304[11])
    defparam i16382_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_2_lut_3_lut_adj_1702 (.I0(\data_out_frame[19] [7]), .I1(\data_out_frame[19] [6]), 
            .I2(n53610), .I3(GND_net), .O(n6_adj_4767));
    defparam i1_2_lut_3_lut_adj_1702.LUT_INIT = 16'h9696;
    SB_LUT4 i16383_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n37), .I2(\data_in_frame[9] [2]), 
            .I3(PWMLimit[10]), .O(n30389));   // verilog/coms.v(148[4] 304[11])
    defparam i16383_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i14_2_lut_adj_1703 (.I0(rx_data_ready), .I1(\FRAME_MATCHER.rx_data_ready_prev ), 
            .I2(GND_net), .I3(GND_net), .O(n161_c));   // verilog/coms.v(156[9:50])
    defparam i14_2_lut_adj_1703.LUT_INIT = 16'h2222;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_55183 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[10] [2]), .I2(\data_out_frame[11] [2]), 
            .I3(\byte_transmit_counter[1] ), .O(n70868));
    defparam byte_transmit_counter_0__bdd_4_lut_55183.LUT_INIT = 16'he4aa;
    SB_LUT4 i23671_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n37), .I2(\data_in_frame[9] [1]), 
            .I3(PWMLimit[9]), .O(n30390));   // verilog/coms.v(148[4] 304[11])
    defparam i23671_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n70868_bdd_4_lut (.I0(n70868), .I1(\data_out_frame[9] [2]), 
            .I2(\data_out_frame[8] [2]), .I3(\byte_transmit_counter[1] ), 
            .O(n70871));
    defparam n70868_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i16387_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n37), .I2(\data_in_frame[9] [0]), 
            .I3(PWMLimit[8]), .O(n30393));   // verilog/coms.v(148[4] 304[11])
    defparam i16387_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2_3_lut_4_lut_adj_1704 (.I0(\data_out_frame[25] [7]), .I1(\data_out_frame[22] [5]), 
            .I2(n53928), .I3(\data_out_frame[24] [0]), .O(n59448));
    defparam i2_3_lut_4_lut_adj_1704.LUT_INIT = 16'h9669;
    SB_LUT4 i16388_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n37), .I2(\data_in_frame[10] [7]), 
            .I3(PWMLimit[7]), .O(n30394));   // verilog/coms.v(148[4] 304[11])
    defparam i16388_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i16421_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n37), .I2(\data_in_frame[10] [6]), 
            .I3(PWMLimit[6]), .O(n30427));   // verilog/coms.v(148[4] 304[11])
    defparam i16421_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i16422_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n37), .I2(\data_in_frame[10] [5]), 
            .I3(PWMLimit[5]), .O(n30428));   // verilog/coms.v(148[4] 304[11])
    defparam i16422_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2_2_lut_4_lut (.I0(n53735), .I1(n59218), .I2(\data_out_frame[23] [7]), 
            .I3(\data_out_frame[24] [2]), .O(n6_adj_4762));
    defparam i2_2_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 select_775_Select_212_i3_3_lut_4_lut (.I0(\data_out_frame[24] [2]), 
            .I1(\data_out_frame[24] [3]), .I2(\FRAME_MATCHER.state[3] ), 
            .I3(n59338), .O(n3_adj_5034));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_212_i3_3_lut_4_lut.LUT_INIT = 16'h9060;
    SB_LUT4 i1_2_lut_adj_1705 (.I0(\FRAME_MATCHER.i[4] ), .I1(\FRAME_MATCHER.i[5] ), 
            .I2(GND_net), .I3(GND_net), .O(n9_adj_5029));   // verilog/coms.v(158[12:15])
    defparam i1_2_lut_adj_1705.LUT_INIT = 16'heeee;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_55173 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[14] [2]), .I2(\data_out_frame[15] [2]), 
            .I3(\byte_transmit_counter[1] ), .O(n70856));
    defparam byte_transmit_counter_0__bdd_4_lut_55173.LUT_INIT = 16'he4aa;
    SB_LUT4 i16426_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n37), .I2(\data_in_frame[10] [4]), 
            .I3(PWMLimit[4]), .O(n30432));   // verilog/coms.v(148[4] 304[11])
    defparam i16426_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i3_3_lut_4_lut (.I0(\data_out_frame[24] [5]), .I1(n61136), .I2(n59448), 
            .I3(n59356), .O(n8_adj_4755));
    defparam i3_3_lut_4_lut.LUT_INIT = 16'h9669;
    SB_LUT4 i16428_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n37), .I2(\data_in_frame[10] [3]), 
            .I3(PWMLimit[3]), .O(n30434));   // verilog/coms.v(148[4] 304[11])
    defparam i16428_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 select_775_Select_154_i2_4_lut (.I0(\data_out_frame[19] [2]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[10]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4930));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_154_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_775_Select_153_i2_4_lut (.I0(\data_out_frame[19] [1]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[9]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4929));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_153_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i16429_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n37), .I2(\data_in_frame[10] [2]), 
            .I3(PWMLimit[2]), .O(n30435));   // verilog/coms.v(148[4] 304[11])
    defparam i16429_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i20843_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n37), .I2(\data_in_frame[10] [1]), 
            .I3(PWMLimit[1]), .O(n30436));   // verilog/coms.v(148[4] 304[11])
    defparam i20843_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2_2_lut_4_lut_adj_1706 (.I0(n1835), .I1(n59168), .I2(n54220), 
            .I3(\data_out_frame[16] [1]), .O(n7_c));
    defparam i2_2_lut_4_lut_adj_1706.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1707 (.I0(n70020), .I1(n54620), .I2(\data_out_frame[20] [7]), 
            .I3(GND_net), .O(n8_adj_4747));
    defparam i1_2_lut_3_lut_adj_1707.LUT_INIT = 16'h9696;
    SB_LUT4 select_775_Select_152_i2_4_lut (.I0(\data_out_frame[19] [0]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[8]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4927));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_152_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i15528_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n37), .I2(\data_in_frame[13] [0]), 
            .I3(IntegralLimit[0]), .O(n29534));   // verilog/coms.v(148[4] 304[11])
    defparam i15528_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i15548_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n37), .I2(\data_in_frame[3] [0]), 
            .I3(\Kp[0] ), .O(n29554));   // verilog/coms.v(148[4] 304[11])
    defparam i15548_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_2_lut_4_lut_adj_1708 (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i[3] ), .I3(n9_adj_5029), .O(n161));
    defparam i1_2_lut_4_lut_adj_1708.LUT_INIT = 16'hfffb;
    SB_LUT4 i1_2_lut_4_lut_adj_1709 (.I0(n1835), .I1(n59168), .I2(n54220), 
            .I3(\data_out_frame[18] [3]), .O(n6_adj_4802));
    defparam i1_2_lut_4_lut_adj_1709.LUT_INIT = 16'h6996;
    SB_LUT4 i15549_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n37), .I2(\data_in_frame[5] [0]), 
            .I3(\Ki[0] ), .O(n29555));   // verilog/coms.v(148[4] 304[11])
    defparam i15549_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_4_lut_adj_1710 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[18] [7]), 
            .I2(displacement[23]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4926));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1710.LUT_INIT = 16'ha088;
    SB_LUT4 i29608_2_lut_3_lut (.I0(n3468), .I1(rx_data_ready), .I2(\FRAME_MATCHER.rx_data_ready_prev ), 
            .I3(GND_net), .O(n43501));
    defparam i29608_2_lut_3_lut.LUT_INIT = 16'h0808;
    SB_LUT4 i23376_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n37), .I2(\data_in_frame[10] [0]), 
            .I3(PWMLimit[0]), .O(n29559));   // verilog/coms.v(148[4] 304[11])
    defparam i23376_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_4_lut_adj_1711 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[18] [6]), 
            .I2(displacement[22]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4925));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1711.LUT_INIT = 16'ha088;
    SB_LUT4 select_775_Select_149_i2_4_lut (.I0(\data_out_frame[18] [5]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[21]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4924));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_149_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i2_2_lut_4_lut_adj_1712 (.I0(\data_out_frame[22] [7]), .I1(\data_out_frame[20] [6]), 
            .I2(\data_out_frame[22] [6]), .I3(n26350), .O(n10_adj_4740));
    defparam i2_2_lut_4_lut_adj_1712.LUT_INIT = 16'h6996;
    SB_LUT4 select_775_Select_148_i2_4_lut (.I0(\data_out_frame[18] [4]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[20]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4923));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_148_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i15674_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n37), .I2(\data_in_frame[4] [7]), 
            .I3(\Ki[15] ), .O(n29680));   // verilog/coms.v(148[4] 304[11])
    defparam i15674_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i15675_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n37), .I2(\data_in_frame[4] [6]), 
            .I3(\Ki[14] ), .O(n29681));   // verilog/coms.v(148[4] 304[11])
    defparam i15675_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i15676_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n37), .I2(\data_in_frame[4] [5]), 
            .I3(\Ki[13] ), .O(n29682));   // verilog/coms.v(148[4] 304[11])
    defparam i15676_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_4_lut_adj_1713 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(DE_c), 
            .I2(n47954), .I3(n33690), .O(n26865));
    defparam i1_4_lut_adj_1713.LUT_INIT = 16'hccc8;
    SB_LUT4 i1_4_lut_adj_1714 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[18] [3]), 
            .I2(displacement[19]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4922));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1714.LUT_INIT = 16'ha088;
    SB_LUT4 i1_2_lut_4_lut_adj_1715 (.I0(\data_out_frame[25] [4]), .I1(\data_out_frame[23] [3]), 
            .I2(n59241), .I3(n53546), .O(n58994));
    defparam i1_2_lut_4_lut_adj_1715.LUT_INIT = 16'h6996;
    SB_LUT4 select_775_Select_146_i2_4_lut (.I0(\data_out_frame[18] [2]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[18]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4921));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_146_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i15677_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n37), .I2(\data_in_frame[4] [4]), 
            .I3(\Ki[12] ), .O(n29683));   // verilog/coms.v(148[4] 304[11])
    defparam i15677_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_3_lut_adj_1716 (.I0(LED_c), .I1(\FRAME_MATCHER.i_31__N_2508 ), 
            .I2(n47954), .I3(GND_net), .O(n27233));   // verilog/coms.v(148[4] 304[11])
    defparam i1_3_lut_adj_1716.LUT_INIT = 16'ha8a8;
    SB_LUT4 i15678_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n37), .I2(\data_in_frame[4] [3]), 
            .I3(\Ki[11] ), .O(n29684));   // verilog/coms.v(148[4] 304[11])
    defparam i15678_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i15679_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n37), .I2(\data_in_frame[4] [2]), 
            .I3(\Ki[10] ), .O(n29685));   // verilog/coms.v(148[4] 304[11])
    defparam i15679_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i15680_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n37), .I2(\data_in_frame[4] [1]), 
            .I3(\Ki[9] ), .O(n29686));   // verilog/coms.v(148[4] 304[11])
    defparam i15680_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i14826_4_lut (.I0(n2873), .I1(n33_adj_5126), .I2(n27233), 
            .I3(\FRAME_MATCHER.i_31__N_2513 ), .O(n28832));   // verilog/coms.v(130[12] 305[6])
    defparam i14826_4_lut.LUT_INIT = 16'ha8a0;
    SB_LUT4 n70856_bdd_4_lut (.I0(n70856), .I1(\data_out_frame[13] [2]), 
            .I2(\data_out_frame[12] [2]), .I3(\byte_transmit_counter[1] ), 
            .O(n70859));
    defparam n70856_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i15681_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n37), .I2(\data_in_frame[4] [0]), 
            .I3(\Ki[8] ), .O(n29687));   // verilog/coms.v(148[4] 304[11])
    defparam i15681_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i19687_4_lut (.I0(Kp_23__N_1748), .I1(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(LED_c), .O(n33693));   // verilog/coms.v(118[11:12])
    defparam i19687_4_lut.LUT_INIT = 16'hfac0;
    SB_LUT4 i14827_2_lut_2_lut (.I0(reset), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(GND_net), .I3(GND_net), .O(n28833));   // verilog/coms.v(130[12] 305[6])
    defparam i14827_2_lut_2_lut.LUT_INIT = 16'h4444;
    uart_tx tx (.r_SM_Main({r_SM_Main}), .GND_net(GND_net), .tx_o(tx_o), 
            .clk16MHz(clk16MHz), .tx_data({tx_data}), .r_Clock_Count({r_Clock_Count}), 
            .VCC_net(VCC_net), .n4938(n4938), .n29(n29), .n23(n23), 
            .\o_Rx_DV_N_3488[12] (\o_Rx_DV_N_3488[12] ), .\o_Rx_DV_N_3488[24] (\o_Rx_DV_N_3488[24] ), 
            .n27(n27), .n29581(n29581), .tx_active(tx_active), .\r_SM_Main_2__N_3536[1] (\r_SM_Main_2__N_3536[1] ), 
            .\r_SM_Main_2__N_3545[0] (r_SM_Main_2__N_3545[0]), .n59648(n59648), 
            .n60274(n60274), .n6(n6), .tx_enable(tx_enable)) /* synthesis syn_module_defined=1 */ ;   // verilog/coms.v(110[25:94])
    uart_rx rx (.GND_net(GND_net), .baudrate({baudrate}), .r_Clock_Count({r_Clock_Count_adj_29}), 
            .\o_Rx_DV_N_3488[2] (\o_Rx_DV_N_3488[2] ), .\o_Rx_DV_N_3488[1] (\o_Rx_DV_N_3488[1] ), 
            .\o_Rx_DV_N_3488[3] (\o_Rx_DV_N_3488[3] ), .\o_Rx_DV_N_3488[4] (\o_Rx_DV_N_3488[4] ), 
            .\o_Rx_DV_N_3488[5] (\o_Rx_DV_N_3488[5] ), .\o_Rx_DV_N_3488[6] (\o_Rx_DV_N_3488[6] ), 
            .\o_Rx_DV_N_3488[8] (\o_Rx_DV_N_3488[8] ), .\o_Rx_DV_N_3488[7] (\o_Rx_DV_N_3488[7] ), 
            .\r_Bit_Index[0] (\r_Bit_Index[0] ), .n61449(n61449), .\o_Rx_DV_N_3488[12] (\o_Rx_DV_N_3488[12] ), 
            .\o_Rx_DV_N_3488[24] (\o_Rx_DV_N_3488[24] ), .n29(n29), .n23(n23), 
            .n62163(n62163), .\r_SM_Main_2__N_3446[1] (\r_SM_Main_2__N_3446[1] ), 
            .n27(n27), .r_Rx_Data(r_Rx_Data), .\r_SM_Main[1] (\r_SM_Main[1]_adj_27 ), 
            .clk16MHz(clk16MHz), .\r_SM_Main[2] (\r_SM_Main[2]_adj_28 ), 
            .RX_N_2(RX_N_2), .VCC_net(VCC_net), .n25515(n25515), .n62091(n62091), 
            .n60815(n60815), .n62089(n62089), .\o_Rx_DV_N_3488[0] (\o_Rx_DV_N_3488[0] ), 
            .n4935(n4935), .n27901(n27901), .n59702(n59702), .n62513(n62513), 
            .n62417(n62417), .n62465(n62465), .n62401(n62401), .n30420(n30420), 
            .rx_data({rx_data}), .n54640(n54640), .rx_data_ready(rx_data_ready), 
            .n30416(n30416), .n62433(n62433), .n30126(n30126), .n30125(n30125), 
            .n30124(n30124), .n30123(n30123), .n30122(n30122), .n30121(n30121), 
            .n30120(n30120), .n62481(n62481), .n58684(n58684), .n62497(n62497), 
            .n62449(n62449), .n27661(n27661)) /* synthesis syn_module_defined=1 */ ;   // verilog/coms.v(96[25:68])
    
endmodule
//
// Verilog Description of module uart_tx
//

module uart_tx (r_SM_Main, GND_net, tx_o, clk16MHz, tx_data, r_Clock_Count, 
            VCC_net, n4938, n29, n23, \o_Rx_DV_N_3488[12] , \o_Rx_DV_N_3488[24] , 
            n27, n29581, tx_active, \r_SM_Main_2__N_3536[1] , \r_SM_Main_2__N_3545[0] , 
            n59648, n60274, n6, tx_enable) /* synthesis syn_module_defined=1 */ ;
    output [2:0]r_SM_Main;
    input GND_net;
    output tx_o;
    input clk16MHz;
    input [7:0]tx_data;
    output [8:0]r_Clock_Count;
    input VCC_net;
    input n4938;
    input n29;
    input n23;
    input \o_Rx_DV_N_3488[12] ;
    input \o_Rx_DV_N_3488[24] ;
    input n27;
    input n29581;
    output tx_active;
    input \r_SM_Main_2__N_3536[1] ;
    input \r_SM_Main_2__N_3545[0] ;
    input n59648;
    input n60274;
    output n6;
    output tx_enable;
    
    wire clk16MHz /* synthesis SET_AS_NETWORK=clk16MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    
    wire n40445, n70979, n3, n25019;
    wire [7:0]r_Tx_Data;   // verilog/uart_tx.v(35[16:25])
    
    wire n54672;
    wire [8:0]n41;
    
    wire n52390, n52389, n52388, n52387, n52386, n52385, n52384, 
        n52383;
    wire [2:0]r_Bit_Index;   // verilog/uart_tx.v(34[16:27])
    
    wire n64526, n64527, n64533, n64532, n62239, n62245, n3_adj_4732;
    wire [2:0]n460;
    
    wire n59740, n29120, n40417, n54670, n71281, n14, n15, n66996, 
        n58489, n66980, n66977, n9, n60245, n70976;
    
    SB_LUT4 i1_1_lut (.I0(r_SM_Main[2]), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n40445));
    defparam i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 r_SM_Main_2__I_0_62_i3_3_lut (.I0(r_SM_Main[0]), .I1(n70979), 
            .I2(r_SM_Main[1]), .I3(GND_net), .O(n3));   // verilog/uart_tx.v(44[7] 143[14])
    defparam r_SM_Main_2__I_0_62_i3_3_lut.LUT_INIT = 16'he5e5;
    SB_DFFE o_Tx_Serial_51 (.Q(tx_o), .C(clk16MHz), .E(n40445), .D(n3));   // verilog/uart_tx.v(41[10] 144[8])
    SB_DFFE r_Tx_Data_i0 (.Q(r_Tx_Data[0]), .C(clk16MHz), .E(n25019), 
            .D(tx_data[0]));   // verilog/uart_tx.v(41[10] 144[8])
    SB_DFFSR r_SM_Main_i0 (.Q(r_SM_Main[0]), .C(clk16MHz), .D(n54672), 
            .R(r_SM_Main[2]));   // verilog/uart_tx.v(41[10] 144[8])
    SB_LUT4 r_Clock_Count_1949_add_4_10_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[8]), .I3(n52390), .O(n41[8])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1949_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 r_Clock_Count_1949_add_4_9_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[7]), .I3(n52389), .O(n41[7])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1949_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1949_add_4_9 (.CI(n52389), .I0(GND_net), .I1(r_Clock_Count[7]), 
            .CO(n52390));
    SB_LUT4 r_Clock_Count_1949_add_4_8_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[6]), .I3(n52388), .O(n41[6])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1949_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1949_add_4_8 (.CI(n52388), .I0(GND_net), .I1(r_Clock_Count[6]), 
            .CO(n52389));
    SB_LUT4 r_Clock_Count_1949_add_4_7_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[5]), .I3(n52387), .O(n41[5])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1949_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1949_add_4_7 (.CI(n52387), .I0(GND_net), .I1(r_Clock_Count[5]), 
            .CO(n52388));
    SB_LUT4 r_Clock_Count_1949_add_4_6_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[4]), .I3(n52386), .O(n41[4])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1949_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1949_add_4_6 (.CI(n52386), .I0(GND_net), .I1(r_Clock_Count[4]), 
            .CO(n52387));
    SB_LUT4 r_Clock_Count_1949_add_4_5_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[3]), .I3(n52385), .O(n41[3])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1949_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1949_add_4_5 (.CI(n52385), .I0(GND_net), .I1(r_Clock_Count[3]), 
            .CO(n52386));
    SB_LUT4 r_Clock_Count_1949_add_4_4_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[2]), .I3(n52384), .O(n41[2])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1949_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1949_add_4_4 (.CI(n52384), .I0(GND_net), .I1(r_Clock_Count[2]), 
            .CO(n52385));
    SB_LUT4 r_Clock_Count_1949_add_4_3_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[1]), .I3(n52383), .O(n41[1])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1949_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1949_add_4_3 (.CI(n52383), .I0(GND_net), .I1(r_Clock_Count[1]), 
            .CO(n52384));
    SB_LUT4 r_Clock_Count_1949_add_4_2_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[0]), .I3(VCC_net), .O(n41[0])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1949_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1949_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(r_Clock_Count[0]), 
            .CO(n52383));
    SB_LUT4 i48832_3_lut (.I0(r_Tx_Data[0]), .I1(r_Tx_Data[1]), .I2(r_Bit_Index[0]), 
            .I3(GND_net), .O(n64526));
    defparam i48832_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48833_3_lut (.I0(r_Tx_Data[4]), .I1(r_Tx_Data[5]), .I2(r_Bit_Index[0]), 
            .I3(GND_net), .O(n64527));
    defparam i48833_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48839_3_lut (.I0(r_Tx_Data[6]), .I1(r_Tx_Data[7]), .I2(r_Bit_Index[0]), 
            .I3(GND_net), .O(n64533));
    defparam i48839_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48838_3_lut (.I0(r_Tx_Data[2]), .I1(r_Tx_Data[3]), .I2(r_Bit_Index[0]), 
            .I3(GND_net), .O(n64532));
    defparam i48838_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut (.I0(n4938), .I1(r_SM_Main[0]), .I2(GND_net), .I3(GND_net), 
            .O(n62239));
    defparam i1_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i1_4_lut (.I0(n29), .I1(n23), .I2(\o_Rx_DV_N_3488[12] ), .I3(n62239), 
            .O(n62245));
    defparam i1_4_lut.LUT_INIT = 16'h0100;
    SB_LUT4 i10_4_lut (.I0(\o_Rx_DV_N_3488[24] ), .I1(r_SM_Main[1]), .I2(n27), 
            .I3(n62245), .O(n3_adj_4732));   // verilog/uart_tx.v(32[16:25])
    defparam i10_4_lut.LUT_INIT = 16'hc9cc;
    SB_DFF r_Tx_Active_53 (.Q(tx_active), .C(clk16MHz), .D(n29581));   // verilog/uart_tx.v(41[10] 144[8])
    SB_DFFESR r_Bit_Index_i1 (.Q(r_Bit_Index[1]), .C(clk16MHz), .E(n59740), 
            .D(n460[1]), .R(n29120));   // verilog/uart_tx.v(41[10] 144[8])
    SB_DFFESR r_Bit_Index_i2 (.Q(r_Bit_Index[2]), .C(clk16MHz), .E(n59740), 
            .D(n460[2]), .R(n29120));   // verilog/uart_tx.v(41[10] 144[8])
    SB_DFFESR r_Clock_Count_1949__i1 (.Q(r_Clock_Count[1]), .C(clk16MHz), 
            .E(n40445), .D(n41[1]), .R(n40417));   // verilog/uart_tx.v(119[34:51])
    SB_DFFESR r_Clock_Count_1949__i2 (.Q(r_Clock_Count[2]), .C(clk16MHz), 
            .E(n40445), .D(n41[2]), .R(n40417));   // verilog/uart_tx.v(119[34:51])
    SB_DFFESR r_Clock_Count_1949__i3 (.Q(r_Clock_Count[3]), .C(clk16MHz), 
            .E(n40445), .D(n41[3]), .R(n40417));   // verilog/uart_tx.v(119[34:51])
    SB_DFFESR r_Clock_Count_1949__i4 (.Q(r_Clock_Count[4]), .C(clk16MHz), 
            .E(n40445), .D(n41[4]), .R(n40417));   // verilog/uart_tx.v(119[34:51])
    SB_DFFESR r_Clock_Count_1949__i5 (.Q(r_Clock_Count[5]), .C(clk16MHz), 
            .E(n40445), .D(n41[5]), .R(n40417));   // verilog/uart_tx.v(119[34:51])
    SB_DFFESR r_Clock_Count_1949__i6 (.Q(r_Clock_Count[6]), .C(clk16MHz), 
            .E(n40445), .D(n41[6]), .R(n40417));   // verilog/uart_tx.v(119[34:51])
    SB_DFFESR r_Clock_Count_1949__i7 (.Q(r_Clock_Count[7]), .C(clk16MHz), 
            .E(n40445), .D(n41[7]), .R(n40417));   // verilog/uart_tx.v(119[34:51])
    SB_DFFESR r_Clock_Count_1949__i8 (.Q(r_Clock_Count[8]), .C(clk16MHz), 
            .E(n40445), .D(n41[8]), .R(n40417));   // verilog/uart_tx.v(119[34:51])
    SB_DFFESR r_Clock_Count_1949__i0 (.Q(r_Clock_Count[0]), .C(clk16MHz), 
            .E(n40445), .D(n41[0]), .R(n40417));   // verilog/uart_tx.v(119[34:51])
    SB_DFFE r_Bit_Index_i0 (.Q(r_Bit_Index[0]), .C(clk16MHz), .E(VCC_net), 
            .D(n54670));   // verilog/uart_tx.v(41[10] 144[8])
    SB_DFF r_SM_Main_i2 (.Q(r_SM_Main[2]), .C(clk16MHz), .D(n71281));   // verilog/uart_tx.v(41[10] 144[8])
    SB_DFFSR r_SM_Main_i1 (.Q(r_SM_Main[1]), .C(clk16MHz), .D(n3_adj_4732), 
            .R(r_SM_Main[2]));   // verilog/uart_tx.v(41[10] 144[8])
    SB_DFFE r_Tx_Data_i7 (.Q(r_Tx_Data[7]), .C(clk16MHz), .E(n25019), 
            .D(tx_data[7]));   // verilog/uart_tx.v(41[10] 144[8])
    SB_DFFE r_Tx_Data_i6 (.Q(r_Tx_Data[6]), .C(clk16MHz), .E(n25019), 
            .D(tx_data[6]));   // verilog/uart_tx.v(41[10] 144[8])
    SB_DFFE r_Tx_Data_i5 (.Q(r_Tx_Data[5]), .C(clk16MHz), .E(n25019), 
            .D(tx_data[5]));   // verilog/uart_tx.v(41[10] 144[8])
    SB_DFFE r_Tx_Data_i4 (.Q(r_Tx_Data[4]), .C(clk16MHz), .E(n25019), 
            .D(tx_data[4]));   // verilog/uart_tx.v(41[10] 144[8])
    SB_DFFE r_Tx_Data_i3 (.Q(r_Tx_Data[3]), .C(clk16MHz), .E(n25019), 
            .D(tx_data[3]));   // verilog/uart_tx.v(41[10] 144[8])
    SB_DFFE r_Tx_Data_i2 (.Q(r_Tx_Data[2]), .C(clk16MHz), .E(n25019), 
            .D(tx_data[2]));   // verilog/uart_tx.v(41[10] 144[8])
    SB_DFFE r_Tx_Data_i1 (.Q(r_Tx_Data[1]), .C(clk16MHz), .E(n25019), 
            .D(tx_data[1]));   // verilog/uart_tx.v(41[10] 144[8])
    SB_LUT4 i55146_2_lut_4_lut (.I0(\r_SM_Main_2__N_3536[1] ), .I1(r_SM_Main[1]), 
            .I2(r_SM_Main[2]), .I3(r_SM_Main[0]), .O(n59740));
    defparam i55146_2_lut_4_lut.LUT_INIT = 16'h0007;
    SB_LUT4 i5_3_lut (.I0(r_SM_Main[0]), .I1(\o_Rx_DV_N_3488[24] ), .I2(n27), 
            .I3(GND_net), .O(n14));
    defparam i5_3_lut.LUT_INIT = 16'h0202;
    SB_LUT4 i6_4_lut (.I0(n29), .I1(\o_Rx_DV_N_3488[12] ), .I2(n23), .I3(n4938), 
            .O(n15));
    defparam i6_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i8_4_lut (.I0(n15), .I1(n40445), .I2(n14), .I3(r_SM_Main[1]), 
            .O(n71281));
    defparam i8_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i52351_2_lut_3_lut (.I0(r_SM_Main[2]), .I1(r_SM_Main[0]), .I2(r_SM_Main[1]), 
            .I3(GND_net), .O(n66996));   // verilog/uart_tx.v(32[16:25])
    defparam i52351_2_lut_3_lut.LUT_INIT = 16'h1010;
    SB_LUT4 i2_3_lut_4_lut (.I0(r_SM_Main[1]), .I1(r_SM_Main[2]), .I2(r_SM_Main[0]), 
            .I3(\r_SM_Main_2__N_3545[0] ), .O(n25019));
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h0100;
    SB_LUT4 i2_3_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[0]), .I2(r_Bit_Index[2]), 
            .I3(GND_net), .O(n58489));   // verilog/uart_tx.v(41[10] 144[8])
    defparam i2_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i52340_3_lut (.I0(n58489), .I1(\o_Rx_DV_N_3488[12] ), .I2(n4938), 
            .I3(GND_net), .O(n66980));   // verilog/uart_tx.v(32[16:25])
    defparam i52340_3_lut.LUT_INIT = 16'h0202;
    SB_LUT4 i52337_4_lut (.I0(n66980), .I1(\o_Rx_DV_N_3488[24] ), .I2(n29), 
            .I3(n23), .O(n66977));   // verilog/uart_tx.v(32[16:25])
    defparam i52337_4_lut.LUT_INIT = 16'h0002;
    SB_LUT4 i23_4_lut (.I0(\r_SM_Main_2__N_3545[0] ), .I1(n66977), .I2(r_SM_Main[1]), 
            .I3(n27), .O(n9));   // verilog/uart_tx.v(32[16:25])
    defparam i23_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i22_3_lut (.I0(n9), .I1(\r_SM_Main_2__N_3536[1] ), .I2(r_SM_Main[0]), 
            .I3(GND_net), .O(n54672));   // verilog/uart_tx.v(32[16:25])
    defparam i22_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12_4_lut (.I0(n66996), .I1(n59740), .I2(r_Bit_Index[0]), 
            .I3(n60245), .O(n54670));   // verilog/uart_tx.v(32[16:25])
    defparam i12_4_lut.LUT_INIT = 16'h303a;
    SB_LUT4 i55085_4_lut (.I0(\r_SM_Main_2__N_3536[1] ), .I1(r_SM_Main[2]), 
            .I2(r_SM_Main[1]), .I3(r_SM_Main[0]), .O(n40417));
    defparam i55085_4_lut.LUT_INIT = 16'h1113;
    SB_LUT4 i26503_3_lut (.I0(r_Bit_Index[2]), .I1(r_Bit_Index[1]), .I2(r_Bit_Index[0]), 
            .I3(GND_net), .O(n460[2]));   // verilog/uart_tx.v(34[16:27])
    defparam i26503_3_lut.LUT_INIT = 16'h6a6a;
    SB_LUT4 i43866_rep_29_2_lut (.I0(\r_SM_Main_2__N_3536[1] ), .I1(r_SM_Main[1]), 
            .I2(GND_net), .I3(GND_net), .O(n60245));
    defparam i43866_rep_29_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut_adj_1056 (.I0(n59648), .I1(n60245), .I2(r_SM_Main[1]), 
            .I3(n58489), .O(n29120));
    defparam i1_4_lut_adj_1056.LUT_INIT = 16'h1101;
    SB_LUT4 i16_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[0]), .I2(GND_net), 
            .I3(GND_net), .O(n460[1]));   // verilog/uart_tx.v(34[16:27])
    defparam i16_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 r_Bit_Index_2__bdd_4_lut (.I0(r_Bit_Index[2]), .I1(n64532), 
            .I2(n64533), .I3(r_Bit_Index[1]), .O(n70976));
    defparam r_Bit_Index_2__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n70976_bdd_4_lut (.I0(n70976), .I1(n64527), .I2(n64526), .I3(r_Bit_Index[1]), 
            .O(n70979));
    defparam n70976_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i17_4_lut (.I0(r_SM_Main[0]), .I1(n60274), .I2(r_SM_Main[1]), 
            .I3(\r_SM_Main_2__N_3545[0] ), .O(n6));
    defparam i17_4_lut.LUT_INIT = 16'h3530;
    SB_LUT4 o_Tx_Serial_I_0_1_lut (.I0(tx_o), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(tx_enable));   // verilog/uart_tx.v(39[24:36])
    defparam o_Tx_Serial_I_0_1_lut.LUT_INIT = 16'h5555;
    
endmodule
//
// Verilog Description of module uart_rx
//

module uart_rx (GND_net, baudrate, r_Clock_Count, \o_Rx_DV_N_3488[2] , 
            \o_Rx_DV_N_3488[1] , \o_Rx_DV_N_3488[3] , \o_Rx_DV_N_3488[4] , 
            \o_Rx_DV_N_3488[5] , \o_Rx_DV_N_3488[6] , \o_Rx_DV_N_3488[8] , 
            \o_Rx_DV_N_3488[7] , \r_Bit_Index[0] , n61449, \o_Rx_DV_N_3488[12] , 
            \o_Rx_DV_N_3488[24] , n29, n23, n62163, \r_SM_Main_2__N_3446[1] , 
            n27, r_Rx_Data, \r_SM_Main[1] , clk16MHz, \r_SM_Main[2] , 
            RX_N_2, VCC_net, n25515, n62091, n60815, n62089, \o_Rx_DV_N_3488[0] , 
            n4935, n27901, n59702, n62513, n62417, n62465, n62401, 
            n30420, rx_data, n54640, rx_data_ready, n30416, n62433, 
            n30126, n30125, n30124, n30123, n30122, n30121, n30120, 
            n62481, n58684, n62497, n62449, n27661) /* synthesis syn_module_defined=1 */ ;
    input GND_net;
    input [31:0]baudrate;
    output [7:0]r_Clock_Count;
    output \o_Rx_DV_N_3488[2] ;
    output \o_Rx_DV_N_3488[1] ;
    output \o_Rx_DV_N_3488[3] ;
    output \o_Rx_DV_N_3488[4] ;
    output \o_Rx_DV_N_3488[5] ;
    output \o_Rx_DV_N_3488[6] ;
    output \o_Rx_DV_N_3488[8] ;
    output \o_Rx_DV_N_3488[7] ;
    output \r_Bit_Index[0] ;
    output n61449;
    output \o_Rx_DV_N_3488[12] ;
    output \o_Rx_DV_N_3488[24] ;
    output n29;
    output n23;
    input n62163;
    input \r_SM_Main_2__N_3446[1] ;
    output n27;
    output r_Rx_Data;
    output \r_SM_Main[1] ;
    input clk16MHz;
    output \r_SM_Main[2] ;
    input RX_N_2;
    input VCC_net;
    output n25515;
    input n62091;
    output n60815;
    output n62089;
    output \o_Rx_DV_N_3488[0] ;
    input n4935;
    output n27901;
    output n59702;
    output n62513;
    output n62417;
    output n62465;
    output n62401;
    input n30420;
    output [7:0]rx_data;
    input n54640;
    output rx_data_ready;
    input n30416;
    output n62433;
    input n30126;
    input n30125;
    input n30124;
    input n30123;
    input n30122;
    input n30121;
    input n30120;
    output n62481;
    input n58684;
    output n62497;
    output n62449;
    output n27661;
    
    wire clk16MHz /* synthesis SET_AS_NETWORK=clk16MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    
    wire n52189, n3056, n2144, n52190;
    wire [23:0]n8391;
    
    wire n3057, n2013, n52188;
    wire [23:0]n8079;
    
    wire n1557, n1011, n52010, n3058, n1879, n52187, n52011, n538, 
        n858, n1558, n856, n52009, n63061, n25574, n59806, n3, 
        n63065, n5, n63069, n8, n58444;
    wire [2:0]r_Bit_Index;   // verilog/uart_rx.v(34[17:28])
    
    wire n3059, n1742, n52186, n1559, n698, n52008, n64168, n64268;
    wire [2:0]r_SM_Main;   // verilog/uart_rx.v(37[17:26])
    
    wire n2, n11632, n3_adj_4458, n3060, n1602, n52185, n2957;
    wire [23:0]n8365;
    wire [23:0]n294;
    
    wire n3065, n3061, n1459, n52184, n3062, n1460, n52183, n3063, 
        n52182, n3064, n52181, n52180, n3066, n52179, n1560, n52007, 
        r_Rx_Data_R, n62057, n59790;
    wire [23:0]n8053;
    
    wire n1408, n52006, n1409, n52005, n2938, n3188, n52178, n1410, 
        n52004, n2939, n3084, n52177, n2940, n2977, n52176, n2956, 
        n1411, n52003, n2941, n2867, n52175, n2942, n2754, n52174, 
        n2955, n2943, n2638, n52173, n2954, n2953, n3154;
    wire [23:0]n8417;
    
    wire n41, n3155, n39, n3158, n33, n3157, n35, n3156, n37, 
        n3163, n23_adj_4459, n3162, n25, n2952, n3160, n29_adj_4460, 
        n3159, n31, n3171, n7, n3152, n45, n3153, n43, n3169, 
        n11, n3168, n13, n3167, n15, n3161, n27_adj_4461, n1412, 
        n52002, n3170, n9, n3166, n17, n2944, n2519, n52172, 
        n1413, n52001, n2951, n2945, n2397, n52171, n1414, n52000, 
        n3165, n19, n2946, n2272, n52170, n3164, n21, n67236, 
        n67246, n16, n67204, n8_adj_4462, n24, n3172, n3274, n67270, 
        n2947, n52169, n2948, n52168, n2949, n52167, n2950, n52166, 
        n52165, n68175, n68170, n1415, n51999, n69549, n68894, 
        n69780, n12, n52164, n62039, n59836, n62059, n48, n4;
    wire [23:0]n8027;
    
    wire n1261, n51998, n1262, n51997, n69482, n69483, n52163, 
        n67225, n10, n30, n67230, n69843, n69421, n69974, n51141, 
        n1263, n51996, n69975, n6, n69484, n69485, n67214, n52162, 
        n52161, n69424, n69419, n69911, n1264, n51995, n67216, 
        n51140, n61999, n69670, n40, n61987, n1265, n51994, n52160, 
        n64284, n51139, n62093, n52159, n62055, n59794, n3151, 
        n3253, n69672, n63609, n63463, n63461, n61995, n60953, 
        n1266, n51993, n1267, n51992, n62037, n59840;
    wire [23:0]n8339;
    
    wire n2827, n52158, n2828, n52157;
    wire [23:0]n8001;
    
    wire n1111, n51991, n2829, n52156, n2830, n52155, n2831, n52154, 
        n1112, n51990, n2832, n52153, n2833, n52152, n2834, n52151, 
        n2835, n52150;
    wire [7:0]n1;
    
    wire n52382, n52381, n52380, n1113, n51989, n52379, n3046, 
        n3047, n3049, n3048, n3050, n3053, n52378, n2836, n52149, 
        n1114, n51988, n33_adj_4466, n3054, n2837, n52148, n52377, 
        n52376, n31_adj_4468, n3051, n37_adj_4469, n3052, n35_adj_4470, 
        n2838, n52147, n25_adj_4471, n27_adj_4472, n51138;
    wire [24:0]o_Rx_DV_N_3488;
    
    wire n9_adj_4473, n21_adj_4474, n51137, n23_adj_4475, n3055, n1115, 
        n51987, n13_adj_4476, n15_adj_4477, n1116, n51986, n2839, 
        n52146, n62035, n59844, n17_adj_4479, n29_adj_4480, n11_adj_4481, 
        n19_adj_4482, n63613, n63615, n63611, n25589, n67294, n2840, 
        n52145, n68221, n68924, n68922, n67296, n6_adj_4483, n69490, 
        n2841, n52144, n2842, n52143, n2843, n52142, n14, n32, 
        n2844, n52141, n69491, n2845, n52140, n62053, n59798, 
        n67290, n12_adj_4484, n67283, n69841, n69411;
    wire [23:0]n8313;
    
    wire n2713, n52139, n51136, n62253, n8_adj_4485, n69492, n69493, 
        n67307, n68211, n10_adj_4486, n69408, n51135, n69407, n2714, 
        n52138, n69237, n69972, n69486, n2715, n52137, n69994, 
        n69995, n69987, n69764, n51134, n69765, n51133, n62251, 
        n2716, n52136, n35_adj_4487, n51132, n61997, n39_adj_4488, 
        n2717, n52135, n51131, n2718, n52134, n51130, n33_adj_4489, 
        n37_adj_4490, n23_adj_4491, n25_adj_4492, n51129, n2719, n52133, 
        n51128, n2720, n52132, n27_adj_4493, n29_adj_4494, n11_adj_4495, 
        n13_adj_4496, n21_adj_4497, n15_adj_4498, n2721, n52131, n17_adj_4499, 
        n19_adj_4500, n31_adj_4501, n67338, n68310, n68944, n68938, 
        n67340, n8_adj_4502, n69496, n51127, n69497, n51126, n2722, 
        n52130, n16_adj_4503, n34, n67332, n14_adj_4504, n67329, 
        n69839, n69399, n10_adj_4505, n69498, n69499, n51125, n67365, 
        n68239, n12_adj_4506, n20, n69397, n69243, n69970, n69402, 
        n69996, n69997, n69985, n69404, n2106, n31_adj_4507, n2107, 
        n29_adj_4508, n2105, n33_adj_4509, n51124, n2104, n35_adj_4510, 
        n2723, n52129, n2102, n39_adj_4511, n2487, n25_adj_4512, 
        n1556, n39_adj_4513, n51123, n2724, n52128, n1555, n41_adj_4514, 
        n2725, n52127, n37_adj_4515, n2726, n52126, n51122, n2727, 
        n52125, n1838, n33_adj_4516, n1839, n31_adj_4517, n1837, 
        n35_adj_4518, n1836, n37_adj_4519, n1834, n41_adj_4520, n2728, 
        n52124, n2729, n52123, n2730, n52122, n1835, n39_adj_4521, 
        n2236, n29_adj_4522, n2235, n31_adj_4523, n2237, n27_adj_4524, 
        n2233, n35_adj_4525, n2238, n25_adj_4526, n25577, n59802, 
        n2232, n37_adj_4527, n2231, n39_adj_4528, n51121, n62051, 
        n2230, n41_adj_4529, n2234, n33_adj_4530;
    wire [23:0]n8287;
    
    wire n2596, n52121, n51120, n2597, n52120, n2229, n43_adj_4531, 
        n2598, n52119, n2599, n52118, n64170, n43066, n804, n20902, 
        n20904, n2600, n52117, n961, n962, n20912, n2601, n52116, 
        n41_adj_4532, n2363, n27_adj_4533, n51119, n2362, n29_adj_4534, 
        n2602, n52115, n2603, n52114, n2604, n52113, n2605, n52112, 
        n2606, n52111, n51118, n2607, n52110, n2608, n52109, n25598, 
        n2609, n52108, n2610, n52107, n2611, n52106, n2612, n52105, 
        n62049;
    wire [23:0]n8261;
    
    wire n2476, n52104, n2477, n52103, n2478, n52102, n2479, n52101, 
        n2480, n52100, n2481, n52099, n2482, n52098, n2483, n52097, 
        n67076, n67082, n67073, n67079, n3_adj_4535, n37_adj_4536, 
        n41_adj_4537, n35_adj_4538, n39_adj_4539, n23_adj_4540, n25_adj_4541, 
        n27_adj_4542, n25580, n29_adj_4543, n31_adj_4544, n69731, 
        n64246, n13_adj_4545, n15_adj_4546, n33_adj_4547, n17_adj_4548, 
        n19_adj_4549, n21_adj_4550, n64192, n63505, n64190, n63459, 
        n64248, n2484, n52096, n67401, n68350, n68960, n68958, 
        n67404, n10_adj_4551, n69502, n69503, n18, n36, n67397, 
        n16_adj_4552, n67394, n69837, n69391, n14_adj_4553, n22, 
        n12_adj_4554, n67420, n69835, n69836, n69715, n69281, n69968, 
        n69661, n69992, n69993, n69989;
    wire [2:0]n479;
    
    wire n27701, n29076, n39_adj_4555, n62551, n48_adj_4556, n37_adj_4557, 
        n43_adj_4558, n4_adj_4559, n41_adj_4560, n31_adj_4561, n33_adj_4562, 
        n25_adj_4563, n27_adj_4564, n29_adj_4565, n59818, n48_adj_4566, 
        n15_adj_4567, n17_adj_4568, n2485, n52095, n41_adj_4569, n45_adj_4570, 
        n43_adj_4571, n27_adj_4572, n29_adj_4573, n31_adj_4574, n59814, 
        n39_adj_4575, n62549, n62541, n62545, n62547, n63959, n63961, 
        n62543, n64214, n64124, n59613, n64280, n17_adj_4576, n19_adj_4577, 
        n33_adj_4578, n35_adj_4579, n2364;
    wire [23:0]n8235;
    
    wire n37_adj_4580, n43_adj_4581, n2356, n41_adj_4582, n39_adj_4583, 
        n31_adj_4584, n33_adj_4585, n35_adj_4586, n11253, n1975;
    wire [23:0]n8157;
    wire [23:0]n8183;
    
    wire n2486, n52094;
    wire [23:0]n8209;
    
    wire n27_adj_4587, n29_adj_4588, n2367, n2490, n52093, n2489, 
        n19_adj_4589, n2488, n52092, n21_adj_4590, n62045, n2491, 
        n2355, n2353, n52091, n2357, n39_adj_4591, n2358, n37_adj_4592, 
        n2359, n35_adj_4593, n2103, n37_adj_4594, n2101, n41_adj_4595, 
        n2108, n27_adj_4596, n71282, n67709, n30_adj_4597, n38_adj_4598, 
        n59821, n2109, n26, n69267, n69268, n67703, n28, n67701, 
        n69748, n68483, n69934, n2100, n69935, n2099, n69866, 
        n2098, n48_adj_4599, n52090, n63515, n63465, n63513, n62569, 
        n63523, n63519, n63521, n25562, n2240, n2366, n21_adj_4600, 
        n2360, n33_adj_4601, n2354, n45_adj_4602, n52089, n23_adj_4603, 
        n2361, n64194, n59827, n31_adj_4604, n1976, n27_adj_4605, 
        n29_adj_4606, n62047, n59810, n41_adj_4607, n43_adj_4608, 
        n19_adj_4609, n67615, n67600, n69428, n18_adj_4610, n69649, 
        n69650, n67613, n68504, n24_adj_4611, n26_adj_4612, n42_adj_4613, 
        n48_adj_4614, n22_adj_4615, n30_adj_4616, n20_adj_4617, n67598, 
        n69758, n69759, n69568, n68506, n69028, n68503, n69030, 
        n52088, n52087, n2227, n1695, n43_adj_4618, n1698, n37_adj_4619, 
        n1696, n41_adj_4620, n1697, n39_adj_4621, n59830, n1701, 
        n32_adj_4622, n69279, n69280, n67757, n68642, n34_adj_4623, 
        n69349, n68466, n69599, n1694, n69600, n3082, n1693, n48_adj_4624, 
        n63491, n63493, n63481, n63369, n25553, n1841, n1971, 
        n37_adj_4625, n1972, n35_adj_4626, n1970, n39_adj_4627, n1974, 
        n31_adj_4628, n1973, n33_adj_4629, n1554, n43_adj_4630, n32_adj_4631, 
        n69283, n69284, n3186, n52086, n67767, n68650, n34_adj_4632, 
        n69347, n68459, n69603, n1553, n69604, n1552, n48_adj_4633, 
        n64228, n1702;
    wire [23:0]n8105;
    
    wire n1840;
    wire [23:0]n8131;
    
    wire n29_adj_4634, n1969, n41_adj_4635, n27_adj_4636, n67729, 
        n30_adj_4637, n38_adj_4638, n26_adj_4639, n69275, n69276, 
        n67723, n28_adj_4640, n67719, n69746, n68475, n69930, n1968, 
        n69931, n1967, n69870, n1966, n48_adj_4641, n2110, n2239, 
        n45_adj_4642, n39_adj_4643, n43_adj_4644, n41_adj_4645, n52085, 
        n34_adj_4646, n69285, n69286, n67776, n68656, n36_adj_4647, 
        n38_adj_4648, n68455, n69345, n2228, n1833, n40_adj_4649, 
        n41_adj_4650, n63509, n63511, n63507, n63401, n63391, n25586, 
        n805, n59847, n42_adj_4651, n960, n69293, n959, n69294, 
        n59530, n48_adj_4652, n63383, n63381, n25605, n37_adj_4653, 
        n63375, n63373, n62683, n43068, n67096, n70030, n48_adj_4654, 
        n46, n59526, n48_adj_4655, n63371, n62695, n52084, n62687, 
        n25608, n52083, n14_adj_4656, n15_adj_4657, n52082, n52081, 
        n52080, n52079, n52078, n52077, n2365, n52076, n52075, 
        n52074, n64242, n52073, n52072, n52071, n52070, n52069, 
        n52068, n52067, n52066, n52065, n52064, n52063, n52062, 
        n52061, n52060, n62043, n52059, n52058, n52057, n52056, 
        n52055, n52054, n52053, n52052, n52051, n52050, n52049, 
        n52048, n52047, n52046, n52045, n52044, n52043, n52042, 
        n52041, n52040, n52039, n52038, n52037, n42_adj_4658, n69295, 
        n803, n69296, n1977, n52036, n59528, n1831, n52035, n1832, 
        n52034, n52033, n52032, n39_adj_4659, n52222, n52031, n52030, 
        n23_adj_4660, n43_adj_4661, n52029, n52221, n52028, n52220, 
        n52219, n38_adj_4662, n40_adj_4663, n42_adj_4664, n67796, 
        n69730, n52218, n52027, n52217, n52216, n1699, n35_adj_4665, 
        n52215, n52214, n52026, n52025, n52213, n62041, n52212, 
        n52024, n52023, n67382, n52211, n52210, n11417, n42_adj_4666, 
        n42_adj_4667, n52022, n52021, n52209, n52020, n52208, n43_adj_4668, 
        n29_adj_4669, n67745, n1700, n52019, n52207, n52018, n52206, 
        n52205, n52204, n52203, n52017, n52202, n52201, n52200, 
        n59786, n52199, n52198, n52016, n52197, n52196, n52195, 
        n32_adj_4670, n40_adj_4671, n28_adj_4672, n69277, n52194, 
        n52015, n69278, n67741, n52014, n52013, n52193, n52192, 
        n30_adj_4673, n67739, n69726, n52012, n52191, n68471, n69918, 
        n69919, n63979, n25_adj_4674, n62363, n64202, n62391, n64128, 
        n64274, n64262, n67378, n44_adj_4675, n44_adj_4676, n44_adj_4677, 
        n23_adj_4678, n67683, n67677, n22_adj_4679, n28_adj_4680, 
        n30_adj_4681, n26_adj_4682, n34_adj_4683, n24_adj_4684, n67675, 
        n69754, n69755, n69574, n69448, n67681, n69526, n68493, 
        n69722, n69723, n48_adj_4685, n64142, n61975, n61167, n62307, 
        n62325, n64208, n64276, n60333, n62563, n62565, n62629, 
        n67007, n67008, n46_adj_4686, n11424, n20914, n46_adj_4687, 
        n36_adj_4688, n38_adj_4689, n40_adj_4690, n67786, n69742, 
        n69743, n69608, n48_adj_4691, n6_adj_4692, n33_adj_4693, n31_adj_4694, 
        n21_adj_4695, n67651, n67645, n26_adj_4696, n28_adj_4697, 
        n24_adj_4698, n32_adj_4699, n22_adj_4700, n67642, n69756, 
        n69757, n69570, n69432, n20_adj_4701, n67649, n69829, n68499, 
        n69922, n69923, n69888, n23_adj_4702, n25_adj_4703, n62017, 
        n62015, n17_adj_4704, n67571, n67566, n69341, n16_adj_4705, 
        n69520, n69521, n67569, n68439, n22_adj_4706, n69031, n69374, 
        n20_adj_4707, n28_adj_4708, n18_adj_4709, n67564, n69877, 
        n69878, n69811, n68442, n69518, n69652, n69849, n69850, 
        n14_adj_4710, n67483, n16_adj_4711, n18_adj_4712, n67452, 
        n21_adj_4713, n23_adj_4714, n25_adj_4715, n20_adj_4716, n16_adj_4717, 
        n67536, n18_adj_4718, n37_adj_4719, n20_adj_4720, n67512, 
        n22_adj_4721, n62589, n67521, n68432, n69012, n69010, n67526, 
        n14_adj_4722, n69514, n69515, n40_adj_4723, n67515, n69033, 
        n69381, n26_adj_4724, n69831, n69832, n69719, n69311, n69655, 
        n69654, n69657, n19_adj_4725, n21_adj_4726, n23_adj_4727, 
        n35_adj_4728, n62711, n67464, n68398, n68994, n68984, n67469, 
        n12_adj_4729, n69510, n38_adj_4730, n69511, n67456, n69508, 
        n69385, n24_adj_4731, n69833, n69834, n69717, n69303, n69821, 
        n69659, n69976, n69977, n67033, n67030, n67056, n67053, 
        n67050, n62117, n62123;
    
    SB_CARRY add_2793_13 (.CI(n52189), .I0(n3056), .I1(n2144), .CO(n52190));
    SB_LUT4 add_2793_12_lut (.I0(GND_net), .I1(n3057), .I2(n2013), .I3(n52188), 
            .O(n8391[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2793_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2793_12 (.CI(n52188), .I0(n3057), .I1(n2013), .CO(n52189));
    SB_LUT4 add_2781_6_lut (.I0(GND_net), .I1(n1557), .I2(n1011), .I3(n52010), 
            .O(n8079[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2781_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2793_11_lut (.I0(GND_net), .I1(n3058), .I2(n1879), .I3(n52187), 
            .O(n8391[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2793_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2781_6 (.CI(n52010), .I0(n1557), .I1(n1011), .CO(n52011));
    SB_LUT4 div_37_i2175_1_lut (.I0(baudrate[0]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n538));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2175_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i2174_1_lut (.I0(baudrate[1]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n858));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2174_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_2781_5_lut (.I0(GND_net), .I1(n1558), .I2(n856), .I3(n52009), 
            .O(n8079[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2781_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut (.I0(r_Clock_Count[1]), .I1(r_Clock_Count[0]), .I2(\o_Rx_DV_N_3488[2] ), 
            .I3(\o_Rx_DV_N_3488[1] ), .O(n63061));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 i44160_1_lut (.I0(n25574), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n59806));
    defparam i44160_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 equal_267_i3_2_lut (.I0(r_Clock_Count[2]), .I1(\o_Rx_DV_N_3488[3] ), 
            .I2(GND_net), .I3(GND_net), .O(n3));   // verilog/uart_rx.v(69[17:62])
    defparam equal_267_i3_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_963 (.I0(r_Clock_Count[3]), .I1(n3), .I2(\o_Rx_DV_N_3488[4] ), 
            .I3(n63061), .O(n63065));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_963.LUT_INIT = 16'hffde;
    SB_CARRY add_2793_11 (.CI(n52187), .I0(n3058), .I1(n1879), .CO(n52188));
    SB_LUT4 equal_267_i5_2_lut (.I0(r_Clock_Count[4]), .I1(\o_Rx_DV_N_3488[5] ), 
            .I2(GND_net), .I3(GND_net), .O(n5));   // verilog/uart_rx.v(69[17:62])
    defparam equal_267_i5_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_2781_5 (.CI(n52009), .I0(n1558), .I1(n856), .CO(n52010));
    SB_LUT4 i1_4_lut_adj_964 (.I0(r_Clock_Count[5]), .I1(n5), .I2(\o_Rx_DV_N_3488[6] ), 
            .I3(n63065), .O(n63069));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_964.LUT_INIT = 16'hffde;
    SB_LUT4 equal_267_i8_2_lut (.I0(r_Clock_Count[7]), .I1(\o_Rx_DV_N_3488[8] ), 
            .I2(GND_net), .I3(GND_net), .O(n8));   // verilog/uart_rx.v(69[17:62])
    defparam equal_267_i8_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_965 (.I0(r_Clock_Count[6]), .I1(n8), .I2(n63069), 
            .I3(\o_Rx_DV_N_3488[7] ), .O(n58444));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_965.LUT_INIT = 16'hfdfe;
    SB_LUT4 i2_3_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), .I2(\r_Bit_Index[0] ), 
            .I3(GND_net), .O(n61449));
    defparam i2_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 add_2793_10_lut (.I0(GND_net), .I1(n3059), .I2(n1742), .I3(n52186), 
            .O(n8391[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2793_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2781_4_lut (.I0(GND_net), .I1(n1559), .I2(n698), .I3(n52008), 
            .O(n8079[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2781_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i48483_2_lut (.I0(\o_Rx_DV_N_3488[12] ), .I1(n58444), .I2(GND_net), 
            .I3(GND_net), .O(n64168));
    defparam i48483_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i48583_4_lut (.I0(\o_Rx_DV_N_3488[24] ), .I1(n29), .I2(n23), 
            .I3(n64168), .O(n64268));
    defparam i48583_4_lut.LUT_INIT = 16'hfffe;
    SB_CARRY add_2793_10 (.CI(n52186), .I0(n3059), .I1(n1742), .CO(n52187));
    SB_LUT4 r_SM_Main_2__I_0_62_Mux_0_i2_4_lut (.I0(n62163), .I1(\r_SM_Main_2__N_3446[1] ), 
            .I2(r_SM_Main[0]), .I3(n27), .O(n2));   // verilog/uart_rx.v(53[7] 144[14])
    defparam r_SM_Main_2__I_0_62_Mux_0_i2_4_lut.LUT_INIT = 16'hc0c5;
    SB_LUT4 r_SM_Main_2__I_0_62_Mux_0_i1_4_lut (.I0(r_Rx_Data), .I1(n64268), 
            .I2(r_SM_Main[0]), .I3(n27), .O(n11632));   // verilog/uart_rx.v(53[7] 144[14])
    defparam r_SM_Main_2__I_0_62_Mux_0_i1_4_lut.LUT_INIT = 16'h0a3a;
    SB_LUT4 r_SM_Main_2__I_0_62_Mux_0_i3_3_lut (.I0(n11632), .I1(n2), .I2(\r_SM_Main[1] ), 
            .I3(GND_net), .O(n3_adj_4458));   // verilog/uart_rx.v(53[7] 144[14])
    defparam r_SM_Main_2__I_0_62_Mux_0_i3_3_lut.LUT_INIT = 16'hc5c5;
    SB_LUT4 add_2793_9_lut (.I0(GND_net), .I1(n3060), .I2(n1602), .I3(n52185), 
            .O(n8391[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2793_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2793_9 (.CI(n52185), .I0(n3060), .I1(n1602), .CO(n52186));
    SB_LUT4 div_37_i2066_3_lut (.I0(n2957), .I1(n8365[4]), .I2(n294[3]), 
            .I3(GND_net), .O(n3065));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2066_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2793_8_lut (.I0(GND_net), .I1(n3061), .I2(n1459), .I3(n52184), 
            .O(n8391[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2793_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2793_8 (.CI(n52184), .I0(n3061), .I1(n1459), .CO(n52185));
    SB_LUT4 add_2793_7_lut (.I0(GND_net), .I1(n3062), .I2(n1460), .I3(n52183), 
            .O(n8391[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2793_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2793_7 (.CI(n52183), .I0(n3062), .I1(n1460), .CO(n52184));
    SB_LUT4 add_2793_6_lut (.I0(GND_net), .I1(n3063), .I2(n1011), .I3(n52182), 
            .O(n8391[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2793_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2793_6 (.CI(n52182), .I0(n3063), .I1(n1011), .CO(n52183));
    SB_LUT4 add_2793_5_lut (.I0(GND_net), .I1(n3064), .I2(n856), .I3(n52181), 
            .O(n8391[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2793_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2793_5 (.CI(n52181), .I0(n3064), .I1(n856), .CO(n52182));
    SB_LUT4 add_2793_4_lut (.I0(GND_net), .I1(n3065), .I2(n698), .I3(n52180), 
            .O(n8391[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2793_4_lut.LUT_INIT = 16'hC33C;
    SB_DFFSR r_SM_Main_i0 (.Q(r_SM_Main[0]), .C(clk16MHz), .D(n3_adj_4458), 
            .R(\r_SM_Main[2] ));   // verilog/uart_rx.v(50[10] 145[8])
    SB_CARRY add_2781_4 (.CI(n52008), .I0(n1559), .I1(n698), .CO(n52009));
    SB_CARRY add_2793_4 (.CI(n52180), .I0(n3065), .I1(n698), .CO(n52181));
    SB_LUT4 add_2793_3_lut (.I0(GND_net), .I1(n3066), .I2(n858), .I3(n52179), 
            .O(n8391[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2793_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2781_3_lut (.I0(GND_net), .I1(n1560), .I2(n858), .I3(n52007), 
            .O(n8079[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2781_3_lut.LUT_INIT = 16'hC33C;
    SB_DFF r_Rx_Data_56 (.Q(r_Rx_Data), .C(clk16MHz), .D(r_Rx_Data_R));   // verilog/uart_rx.v(42[10] 46[8])
    SB_CARRY add_2793_3 (.CI(n52179), .I0(n3066), .I1(n858), .CO(n52180));
    SB_DFF r_Rx_Data_R_55 (.Q(r_Rx_Data_R), .C(clk16MHz), .D(RX_N_2));   // verilog/uart_rx.v(42[10] 46[8])
    SB_CARRY add_2781_3 (.CI(n52007), .I0(n1560), .I1(n858), .CO(n52008));
    SB_LUT4 add_2781_2_lut (.I0(GND_net), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n8079[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2781_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2781_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n52007));
    SB_LUT4 add_2793_2_lut (.I0(n59790), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n62057)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2793_2_lut.LUT_INIT = 16'h8228;
    SB_LUT4 add_2780_10_lut (.I0(GND_net), .I1(n1408), .I2(n1742), .I3(n52006), 
            .O(n8053[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2780_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2780_9_lut (.I0(GND_net), .I1(n1409), .I2(n1602), .I3(n52005), 
            .O(n8053[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2780_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2793_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n52179));
    SB_CARRY add_2780_9 (.CI(n52005), .I0(n1409), .I1(n1602), .CO(n52006));
    SB_LUT4 add_2792_22_lut (.I0(GND_net), .I1(n2938), .I2(n3188), .I3(n52178), 
            .O(n8365[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2792_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2780_8_lut (.I0(GND_net), .I1(n1410), .I2(n1459), .I3(n52004), 
            .O(n8053[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2780_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2780_8 (.CI(n52004), .I0(n1410), .I1(n1459), .CO(n52005));
    SB_LUT4 add_2792_21_lut (.I0(GND_net), .I1(n2939), .I2(n3084), .I3(n52177), 
            .O(n8365[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2792_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2792_21 (.CI(n52177), .I0(n2939), .I1(n3084), .CO(n52178));
    SB_LUT4 add_2792_20_lut (.I0(GND_net), .I1(n2940), .I2(n2977), .I3(n52176), 
            .O(n8365[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2792_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2792_20 (.CI(n52176), .I0(n2940), .I1(n2977), .CO(n52177));
    SB_LUT4 div_37_i2065_3_lut (.I0(n2956), .I1(n8365[5]), .I2(n294[3]), 
            .I3(GND_net), .O(n3064));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2065_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2780_7_lut (.I0(GND_net), .I1(n1411), .I2(n1460), .I3(n52003), 
            .O(n8053[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2780_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2792_19_lut (.I0(GND_net), .I1(n2941), .I2(n2867), .I3(n52175), 
            .O(n8365[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2792_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2792_19 (.CI(n52175), .I0(n2941), .I1(n2867), .CO(n52176));
    SB_LUT4 add_2792_18_lut (.I0(GND_net), .I1(n2942), .I2(n2754), .I3(n52174), 
            .O(n8365[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2792_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2792_18 (.CI(n52174), .I0(n2942), .I1(n2754), .CO(n52175));
    SB_LUT4 div_37_i2064_3_lut (.I0(n2955), .I1(n8365[6]), .I2(n294[3]), 
            .I3(GND_net), .O(n3063));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2064_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2170_1_lut (.I0(baudrate[5]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1460));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2170_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_2792_17_lut (.I0(GND_net), .I1(n2943), .I2(n2638), .I3(n52173), 
            .O(n8365[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2792_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_i2063_3_lut (.I0(n2954), .I1(n8365[7]), .I2(n294[3]), 
            .I3(GND_net), .O(n3062));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2063_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2169_1_lut (.I0(baudrate[6]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1459));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2169_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i2062_3_lut (.I0(n2953), .I1(n8365[8]), .I2(n294[3]), 
            .I3(GND_net), .O(n3061));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2062_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2210_i41_4_lut (.I0(n3154), .I1(baudrate[20]), 
            .I2(n8417[20]), .I3(n294[1]), .O(n41));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i41_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_LessThan_2210_i39_4_lut (.I0(n3155), .I1(baudrate[19]), 
            .I2(n8417[19]), .I3(n294[1]), .O(n39));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i39_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_LessThan_2210_i33_4_lut (.I0(n3158), .I1(baudrate[16]), 
            .I2(n8417[16]), .I3(n294[1]), .O(n33));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i33_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_LessThan_2210_i35_4_lut (.I0(n3157), .I1(baudrate[17]), 
            .I2(n8417[17]), .I3(n294[1]), .O(n35));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i35_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_LessThan_2210_i37_4_lut (.I0(n3156), .I1(baudrate[18]), 
            .I2(n8417[18]), .I3(n294[1]), .O(n37));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i37_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_LessThan_2210_i23_4_lut (.I0(n3163), .I1(baudrate[11]), 
            .I2(n8417[11]), .I3(n294[1]), .O(n23_adj_4459));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i23_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_LessThan_2210_i25_4_lut (.I0(n3162), .I1(baudrate[12]), 
            .I2(n8417[12]), .I3(n294[1]), .O(n25));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i25_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_i2168_1_lut (.I0(baudrate[7]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1602));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2168_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i2061_3_lut (.I0(n2952), .I1(n8365[9]), .I2(n294[3]), 
            .I3(GND_net), .O(n3060));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2061_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2210_i29_4_lut (.I0(n3160), .I1(baudrate[14]), 
            .I2(n8417[14]), .I3(n294[1]), .O(n29_adj_4460));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i29_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_LessThan_2210_i31_4_lut (.I0(n3159), .I1(baudrate[15]), 
            .I2(n8417[15]), .I3(n294[1]), .O(n31));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i31_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_LessThan_2210_i7_4_lut (.I0(n3171), .I1(baudrate[3]), 
            .I2(n8417[3]), .I3(n294[1]), .O(n7));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i7_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_LessThan_2210_i45_4_lut (.I0(n3152), .I1(baudrate[22]), 
            .I2(n8417[22]), .I3(n294[1]), .O(n45));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i45_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_LessThan_2210_i43_4_lut (.I0(n3153), .I1(baudrate[21]), 
            .I2(n8417[21]), .I3(n294[1]), .O(n43));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i43_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_LessThan_2210_i11_4_lut (.I0(n3169), .I1(baudrate[5]), 
            .I2(n8417[5]), .I3(n294[1]), .O(n11));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i11_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_LessThan_2210_i13_4_lut (.I0(n3168), .I1(baudrate[6]), 
            .I2(n8417[6]), .I3(n294[1]), .O(n13));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i13_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_LessThan_2210_i15_4_lut (.I0(n3167), .I1(baudrate[7]), 
            .I2(n8417[7]), .I3(n294[1]), .O(n15));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i15_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_LessThan_2210_i27_4_lut (.I0(n3161), .I1(baudrate[13]), 
            .I2(n8417[13]), .I3(n294[1]), .O(n27_adj_4461));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i27_4_lut.LUT_INIT = 16'h3c66;
    SB_CARRY add_2792_17 (.CI(n52173), .I0(n2943), .I1(n2638), .CO(n52174));
    SB_CARRY add_2780_7 (.CI(n52003), .I0(n1411), .I1(n1460), .CO(n52004));
    SB_LUT4 add_2780_6_lut (.I0(GND_net), .I1(n1412), .I2(n1011), .I3(n52002), 
            .O(n8053[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2780_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_2210_i9_4_lut (.I0(n3170), .I1(baudrate[4]), 
            .I2(n8417[4]), .I3(n294[1]), .O(n9));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i9_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_LessThan_2210_i17_4_lut (.I0(n3166), .I1(baudrate[8]), 
            .I2(n8417[8]), .I3(n294[1]), .O(n17));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i17_4_lut.LUT_INIT = 16'h3c66;
    SB_CARRY add_2780_6 (.CI(n52002), .I0(n1412), .I1(n1011), .CO(n52003));
    SB_LUT4 add_2792_16_lut (.I0(GND_net), .I1(n2944), .I2(n2519), .I3(n52172), 
            .O(n8365[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2792_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2780_5_lut (.I0(GND_net), .I1(n1413), .I2(n856), .I3(n52001), 
            .O(n8053[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2780_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2780_5 (.CI(n52001), .I0(n1413), .I1(n856), .CO(n52002));
    SB_CARRY add_2792_16 (.CI(n52172), .I0(n2944), .I1(n2519), .CO(n52173));
    SB_LUT4 div_37_i2173_1_lut (.I0(baudrate[2]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n698));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2173_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i2167_1_lut (.I0(baudrate[8]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1742));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2167_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i2060_3_lut (.I0(n2951), .I1(n8365[10]), .I2(n294[3]), 
            .I3(GND_net), .O(n3059));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2060_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2792_15_lut (.I0(GND_net), .I1(n2945), .I2(n2397), .I3(n52171), 
            .O(n8365[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2792_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2792_15 (.CI(n52171), .I0(n2945), .I1(n2397), .CO(n52172));
    SB_LUT4 add_2780_4_lut (.I0(GND_net), .I1(n1414), .I2(n698), .I3(n52000), 
            .O(n8053[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2780_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_2210_i19_4_lut (.I0(n3165), .I1(baudrate[9]), 
            .I2(n8417[9]), .I3(n294[1]), .O(n19));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i19_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 add_2792_14_lut (.I0(GND_net), .I1(n2946), .I2(n2272), .I3(n52170), 
            .O(n8365[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2792_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_2210_i21_4_lut (.I0(n3164), .I1(baudrate[10]), 
            .I2(n8417[10]), .I3(n294[1]), .O(n21));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i21_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 i51542_4_lut (.I0(n27_adj_4461), .I1(n15), .I2(n13), .I3(n11), 
            .O(n67236));
    defparam i51542_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i51552_4_lut (.I0(n21), .I1(n19), .I2(n17), .I3(n9), .O(n67246));
    defparam i51552_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_37_LessThan_2210_i16_3_lut (.I0(baudrate[9]), .I1(baudrate[21]), 
            .I2(n43), .I3(GND_net), .O(n16));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51510_2_lut (.I0(n43), .I1(n19), .I2(GND_net), .I3(GND_net), 
            .O(n67204));
    defparam i51510_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 div_37_LessThan_2210_i8_3_lut (.I0(baudrate[4]), .I1(baudrate[8]), 
            .I2(n17), .I3(GND_net), .O(n8_adj_4462));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2210_i24_3_lut (.I0(n16), .I1(baudrate[22]), 
            .I2(n45), .I3(GND_net), .O(n24));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2208_3_lut (.I0(n3172), .I1(n8417[2]), .I2(n294[1]), 
            .I3(GND_net), .O(n3274));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2208_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51576_3_lut (.I0(n7), .I1(n3274), .I2(baudrate[2]), .I3(GND_net), 
            .O(n67270));
    defparam i51576_3_lut.LUT_INIT = 16'hbebe;
    SB_CARRY add_2792_14 (.CI(n52170), .I0(n2946), .I1(n2272), .CO(n52171));
    SB_LUT4 add_2792_13_lut (.I0(GND_net), .I1(n2947), .I2(n2144), .I3(n52169), 
            .O(n8365[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2792_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2792_13 (.CI(n52169), .I0(n2947), .I1(n2144), .CO(n52170));
    SB_LUT4 add_2792_12_lut (.I0(GND_net), .I1(n2948), .I2(n2013), .I3(n52168), 
            .O(n8365[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2792_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2780_4 (.CI(n52000), .I0(n1414), .I1(n698), .CO(n52001));
    SB_CARRY add_2792_12 (.CI(n52168), .I0(n2948), .I1(n2013), .CO(n52169));
    SB_LUT4 add_2792_11_lut (.I0(GND_net), .I1(n2949), .I2(n1879), .I3(n52167), 
            .O(n8365[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2792_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2792_11 (.CI(n52167), .I0(n2949), .I1(n1879), .CO(n52168));
    SB_LUT4 add_2792_10_lut (.I0(GND_net), .I1(n2950), .I2(n1742), .I3(n52166), 
            .O(n8365[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2792_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2792_10 (.CI(n52166), .I0(n2950), .I1(n1742), .CO(n52167));
    SB_LUT4 add_2792_9_lut (.I0(GND_net), .I1(n2951), .I2(n1602), .I3(n52165), 
            .O(n8365[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2792_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2792_9 (.CI(n52165), .I0(n2951), .I1(n1602), .CO(n52166));
    SB_LUT4 i52481_4_lut (.I0(n13), .I1(n11), .I2(n9), .I3(n67270), 
            .O(n68175));
    defparam i52481_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i52476_4_lut (.I0(n19), .I1(n17), .I2(n15), .I3(n68175), 
            .O(n68170));
    defparam i52476_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 add_2780_3_lut (.I0(GND_net), .I1(n1415), .I2(n858), .I3(n51999), 
            .O(n8053[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2780_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i53855_4_lut (.I0(n25), .I1(n23_adj_4459), .I2(n21), .I3(n68170), 
            .O(n69549));
    defparam i53855_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i53200_4_lut (.I0(n31), .I1(n29_adj_4460), .I2(n27_adj_4461), 
            .I3(n69549), .O(n68894));
    defparam i53200_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i54086_4_lut (.I0(n37), .I1(n35), .I2(n33), .I3(n68894), 
            .O(n69780));
    defparam i54086_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_LessThan_2210_i12_3_lut (.I0(baudrate[7]), .I1(baudrate[16]), 
            .I2(n33), .I3(GND_net), .O(n12));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2792_8_lut (.I0(GND_net), .I1(n2952), .I2(n1459), .I3(n52164), 
            .O(n8365[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2792_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2780_3 (.CI(n51999), .I0(n1415), .I1(n858), .CO(n52000));
    SB_LUT4 add_2780_2_lut (.I0(n59836), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n62039)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2780_2_lut.LUT_INIT = 16'h8228;
    SB_LUT4 div_37_LessThan_2210_i4_4_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n62059), .I3(n48), .O(n4));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i4_4_lut.LUT_INIT = 16'hee8e;
    SB_CARRY add_2792_8 (.CI(n52164), .I0(n2952), .I1(n1459), .CO(n52165));
    SB_CARRY add_2780_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n51999));
    SB_LUT4 add_2779_9_lut (.I0(GND_net), .I1(n1261), .I2(n1602), .I3(n51998), 
            .O(n8027[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2779_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2779_8_lut (.I0(GND_net), .I1(n1262), .I2(n1459), .I3(n51997), 
            .O(n8027[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2779_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2779_8 (.CI(n51997), .I0(n1262), .I1(n1459), .CO(n51998));
    SB_LUT4 i53788_3_lut (.I0(n4), .I1(baudrate[13]), .I2(n27_adj_4461), 
            .I3(GND_net), .O(n69482));   // verilog/uart_rx.v(119[33:55])
    defparam i53788_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53789_3_lut (.I0(n69482), .I1(baudrate[14]), .I2(n29_adj_4460), 
            .I3(GND_net), .O(n69483));   // verilog/uart_rx.v(119[33:55])
    defparam i53789_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2792_7_lut (.I0(GND_net), .I1(n2953), .I2(n1460), .I3(n52163), 
            .O(n8365[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2792_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i51531_2_lut (.I0(n33), .I1(n15), .I2(GND_net), .I3(GND_net), 
            .O(n67225));
    defparam i51531_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 div_37_LessThan_2210_i10_3_lut (.I0(baudrate[5]), .I1(baudrate[6]), 
            .I2(n13), .I3(GND_net), .O(n10));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2210_i30_3_lut (.I0(n12), .I1(baudrate[17]), 
            .I2(n35), .I3(GND_net), .O(n30));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51536_4_lut (.I0(n33), .I1(n31), .I2(n29_adj_4460), .I3(n67236), 
            .O(n67230));
    defparam i51536_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i54149_4_lut (.I0(n30), .I1(n10), .I2(n35), .I3(n67225), 
            .O(n69843));   // verilog/uart_rx.v(119[33:55])
    defparam i54149_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i53727_3_lut (.I0(n69483), .I1(baudrate[15]), .I2(n31), .I3(GND_net), 
            .O(n69421));   // verilog/uart_rx.v(119[33:55])
    defparam i53727_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i54280_4_lut (.I0(n69421), .I1(n69843), .I2(n35), .I3(n67230), 
            .O(n69974));   // verilog/uart_rx.v(119[33:55])
    defparam i54280_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 sub_38_add_2_26_lut (.I0(GND_net), .I1(GND_net), .I2(VCC_net), 
            .I3(n51141), .O(\o_Rx_DV_N_3488[24] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2792_7 (.CI(n52163), .I0(n2953), .I1(n1460), .CO(n52164));
    SB_LUT4 add_2779_7_lut (.I0(GND_net), .I1(n1263), .I2(n1460), .I3(n51996), 
            .O(n8027[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2779_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i54281_3_lut (.I0(n69974), .I1(baudrate[18]), .I2(n37), .I3(GND_net), 
            .O(n69975));   // verilog/uart_rx.v(119[33:55])
    defparam i54281_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2210_i6_3_lut (.I0(baudrate[2]), .I1(baudrate[3]), 
            .I2(n7), .I3(GND_net), .O(n6));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53790_3_lut (.I0(n6), .I1(baudrate[10]), .I2(n21), .I3(GND_net), 
            .O(n69484));   // verilog/uart_rx.v(119[33:55])
    defparam i53790_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53791_3_lut (.I0(n69484), .I1(baudrate[11]), .I2(n23_adj_4459), 
            .I3(GND_net), .O(n69485));   // verilog/uart_rx.v(119[33:55])
    defparam i53791_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51520_4_lut (.I0(n43), .I1(n25), .I2(n23_adj_4459), .I3(n67246), 
            .O(n67214));
    defparam i51520_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 add_2792_6_lut (.I0(GND_net), .I1(n2954), .I2(n1011), .I3(n52162), 
            .O(n8365[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2792_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2792_6 (.CI(n52162), .I0(n2954), .I1(n1011), .CO(n52163));
    SB_LUT4 add_2792_5_lut (.I0(GND_net), .I1(n2955), .I2(n856), .I3(n52161), 
            .O(n8365[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2792_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2779_7 (.CI(n51996), .I0(n1263), .I1(n1460), .CO(n51997));
    SB_CARRY add_2792_5 (.CI(n52161), .I0(n2955), .I1(n856), .CO(n52162));
    SB_LUT4 i53730_4_lut (.I0(n24), .I1(n8_adj_4462), .I2(n45), .I3(n67204), 
            .O(n69424));   // verilog/uart_rx.v(119[33:55])
    defparam i53730_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i53725_3_lut (.I0(n69485), .I1(baudrate[12]), .I2(n25), .I3(GND_net), 
            .O(n69419));   // verilog/uart_rx.v(119[33:55])
    defparam i53725_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i54217_3_lut (.I0(n69975), .I1(baudrate[19]), .I2(n39), .I3(GND_net), 
            .O(n69911));   // verilog/uart_rx.v(119[33:55])
    defparam i54217_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2779_6_lut (.I0(GND_net), .I1(n1264), .I2(n1011), .I3(n51995), 
            .O(n8027[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2779_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2779_6 (.CI(n51995), .I0(n1264), .I1(n1011), .CO(n51996));
    SB_LUT4 i51522_4_lut (.I0(n43), .I1(n41), .I2(n39), .I3(n69780), 
            .O(n67216));
    defparam i51522_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 sub_38_add_2_25_lut (.I0(n61999), .I1(n25515), .I2(VCC_net), 
            .I3(n51140), .O(n27)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_25_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_38_add_2_25 (.CI(n51140), .I0(n25515), .I1(VCC_net), 
            .CO(n51141));
    SB_LUT4 i53976_4_lut (.I0(n69419), .I1(n69424), .I2(n45), .I3(n67214), 
            .O(n69670));   // verilog/uart_rx.v(119[33:55])
    defparam i53976_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i54207_3_lut (.I0(n69911), .I1(baudrate[20]), .I2(n41), .I3(GND_net), 
            .O(n40));   // verilog/uart_rx.v(119[33:55])
    defparam i54207_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut (.I0(baudrate[25]), .I1(baudrate[31]), .I2(GND_net), 
            .I3(GND_net), .O(n61987));
    defparam i1_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 add_2779_5_lut (.I0(GND_net), .I1(n1265), .I2(n856), .I3(n51994), 
            .O(n8027[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2779_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2792_4_lut (.I0(GND_net), .I1(n2956), .I2(n698), .I3(n52160), 
            .O(n8365[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2792_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_38_add_2_24_lut (.I0(n62093), .I1(n64284), .I2(VCC_net), 
            .I3(n51139), .O(n29)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_24_lut.LUT_INIT = 16'hebbe;
    SB_CARRY add_2792_4 (.CI(n52160), .I0(n2956), .I1(n698), .CO(n52161));
    SB_LUT4 add_2792_3_lut (.I0(GND_net), .I1(n2957), .I2(n858), .I3(n52159), 
            .O(n8365[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2792_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_38_add_2_24 (.CI(n51139), .I0(n64284), .I1(VCC_net), 
            .CO(n51140));
    SB_CARRY add_2792_3 (.CI(n52159), .I0(n2957), .I1(n858), .CO(n52160));
    SB_LUT4 add_2792_2_lut (.I0(n59794), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n62055)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2792_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_2779_5 (.CI(n51994), .I0(n1265), .I1(n856), .CO(n51995));
    SB_LUT4 div_37_i2187_3_lut (.I0(n3151), .I1(n8417[23]), .I2(n294[1]), 
            .I3(GND_net), .O(n3253));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2187_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53978_4_lut (.I0(n40), .I1(n69670), .I2(n45), .I3(n67216), 
            .O(n69672));   // verilog/uart_rx.v(119[33:55])
    defparam i53978_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i1_4_lut_adj_966 (.I0(n63609), .I1(n63463), .I2(n61987), .I3(n63461), 
            .O(n61995));
    defparam i1_4_lut_adj_966.LUT_INIT = 16'hfffe;
    SB_LUT4 i54707_4_lut (.I0(n61995), .I1(n69672), .I2(baudrate[23]), 
            .I3(n3253), .O(n60953));   // verilog/uart_rx.v(119[33:55])
    defparam i54707_4_lut.LUT_INIT = 16'h1501;
    SB_CARRY add_2792_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n52159));
    SB_LUT4 add_2779_4_lut (.I0(GND_net), .I1(n1266), .I2(n698), .I3(n51993), 
            .O(n8027[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2779_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2779_4 (.CI(n51993), .I0(n1266), .I1(n698), .CO(n51994));
    SB_LUT4 add_2779_3_lut (.I0(GND_net), .I1(n1267), .I2(n858), .I3(n51992), 
            .O(n8027[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2779_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2779_3 (.CI(n51992), .I0(n1267), .I1(n858), .CO(n51993));
    SB_LUT4 add_2779_2_lut (.I0(n59840), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n62037)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2779_2_lut.LUT_INIT = 16'h8228;
    SB_LUT4 add_2791_21_lut (.I0(GND_net), .I1(n2827), .I2(n3084), .I3(n52158), 
            .O(n8339[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2791_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2779_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n51992));
    SB_LUT4 add_2791_20_lut (.I0(GND_net), .I1(n2828), .I2(n2977), .I3(n52157), 
            .O(n8339[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2791_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2791_20 (.CI(n52157), .I0(n2828), .I1(n2977), .CO(n52158));
    SB_LUT4 add_2778_8_lut (.I0(GND_net), .I1(n1111), .I2(n1459), .I3(n51991), 
            .O(n8001[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2778_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2791_19_lut (.I0(GND_net), .I1(n2829), .I2(n2867), .I3(n52156), 
            .O(n8339[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2791_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2791_19 (.CI(n52156), .I0(n2829), .I1(n2867), .CO(n52157));
    SB_LUT4 add_2791_18_lut (.I0(GND_net), .I1(n2830), .I2(n2754), .I3(n52155), 
            .O(n8339[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2791_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2791_18 (.CI(n52155), .I0(n2830), .I1(n2754), .CO(n52156));
    SB_LUT4 add_2791_17_lut (.I0(GND_net), .I1(n2831), .I2(n2638), .I3(n52154), 
            .O(n8339[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2791_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2778_7_lut (.I0(GND_net), .I1(n1112), .I2(n1460), .I3(n51990), 
            .O(n8001[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2778_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2791_17 (.CI(n52154), .I0(n2831), .I1(n2638), .CO(n52155));
    SB_LUT4 add_2791_16_lut (.I0(GND_net), .I1(n2832), .I2(n2519), .I3(n52153), 
            .O(n8339[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2791_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2791_16 (.CI(n52153), .I0(n2832), .I1(n2519), .CO(n52154));
    SB_LUT4 add_2791_15_lut (.I0(GND_net), .I1(n2833), .I2(n2397), .I3(n52152), 
            .O(n8339[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2791_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2791_15 (.CI(n52152), .I0(n2833), .I1(n2397), .CO(n52153));
    SB_LUT4 add_2791_14_lut (.I0(GND_net), .I1(n2834), .I2(n2272), .I3(n52151), 
            .O(n8339[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2791_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2791_14 (.CI(n52151), .I0(n2834), .I1(n2272), .CO(n52152));
    SB_CARRY add_2778_7 (.CI(n51990), .I0(n1112), .I1(n1460), .CO(n51991));
    SB_LUT4 add_2791_13_lut (.I0(GND_net), .I1(n2835), .I2(n2144), .I3(n52150), 
            .O(n8339[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2791_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2791_13 (.CI(n52150), .I0(n2835), .I1(n2144), .CO(n52151));
    SB_LUT4 r_Clock_Count_1947_add_4_9_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[7]), .I3(n52382), .O(n1[7])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1947_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 r_Clock_Count_1947_add_4_8_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[6]), .I3(n52381), .O(n1[6])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1947_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1947_add_4_8 (.CI(n52381), .I0(GND_net), .I1(r_Clock_Count[6]), 
            .CO(n52382));
    SB_LUT4 r_Clock_Count_1947_add_4_7_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[5]), .I3(n52380), .O(n1[5])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1947_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2778_6_lut (.I0(GND_net), .I1(n1113), .I2(n1011), .I3(n51989), 
            .O(n8001[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2778_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1947_add_4_7 (.CI(n52380), .I0(GND_net), .I1(r_Clock_Count[5]), 
            .CO(n52381));
    SB_LUT4 r_Clock_Count_1947_add_4_6_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[4]), .I3(n52379), .O(n1[4])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1947_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2778_6 (.CI(n51989), .I0(n1113), .I1(n1011), .CO(n51990));
    SB_CARRY r_Clock_Count_1947_add_4_6 (.CI(n52379), .I0(GND_net), .I1(r_Clock_Count[4]), 
            .CO(n52380));
    SB_LUT4 div_37_i2118_3_lut (.I0(n3046), .I1(n8391[23]), .I2(n294[2]), 
            .I3(GND_net), .O(n3151));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2118_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2135_3_lut (.I0(n3063), .I1(n8391[6]), .I2(n294[2]), 
            .I3(GND_net), .O(n3168));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2135_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2119_3_lut (.I0(n3047), .I1(n8391[22]), .I2(n294[2]), 
            .I3(GND_net), .O(n3152));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2119_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2121_3_lut (.I0(n3049), .I1(n8391[20]), .I2(n294[2]), 
            .I3(GND_net), .O(n3154));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2121_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2120_3_lut (.I0(n3048), .I1(n8391[21]), .I2(n294[2]), 
            .I3(GND_net), .O(n3153));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2120_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2122_3_lut (.I0(n3050), .I1(n8391[19]), .I2(n294[2]), 
            .I3(GND_net), .O(n3155));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2122_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2125_3_lut (.I0(n3053), .I1(n8391[16]), .I2(n294[2]), 
            .I3(GND_net), .O(n3158));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2125_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 r_Clock_Count_1947_add_4_5_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[3]), .I3(n52378), .O(n1[3])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1947_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2791_12_lut (.I0(GND_net), .I1(n2836), .I2(n2013), .I3(n52149), 
            .O(n8339[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2791_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2791_12 (.CI(n52149), .I0(n2836), .I1(n2013), .CO(n52150));
    SB_LUT4 add_2778_5_lut (.I0(GND_net), .I1(n1114), .I2(n856), .I3(n51988), 
            .O(n8001[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2778_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_2141_i33_2_lut (.I0(n3158), .I1(baudrate[15]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_4466));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i2126_3_lut (.I0(n3054), .I1(n8391[15]), .I2(n294[2]), 
            .I3(GND_net), .O(n3159));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2126_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2791_11_lut (.I0(GND_net), .I1(n2837), .I2(n1879), .I3(n52148), 
            .O(n8339[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2791_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1947_add_4_5 (.CI(n52378), .I0(GND_net), .I1(r_Clock_Count[3]), 
            .CO(n52379));
    SB_LUT4 r_Clock_Count_1947_add_4_4_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[2]), .I3(n52377), .O(n1[2])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1947_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2791_11 (.CI(n52148), .I0(n2837), .I1(n1879), .CO(n52149));
    SB_CARRY r_Clock_Count_1947_add_4_4 (.CI(n52377), .I0(GND_net), .I1(r_Clock_Count[2]), 
            .CO(n52378));
    SB_LUT4 r_Clock_Count_1947_add_4_3_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[1]), .I3(n52376), .O(n1[1])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1947_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_2141_i31_2_lut (.I0(n3159), .I1(baudrate[14]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_4468));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i2123_3_lut (.I0(n3051), .I1(n8391[18]), .I2(n294[2]), 
            .I3(GND_net), .O(n3156));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2123_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2141_i37_2_lut (.I0(n3156), .I1(baudrate[17]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_4469));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i2124_3_lut (.I0(n3052), .I1(n8391[17]), .I2(n294[2]), 
            .I3(GND_net), .O(n3157));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2124_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2141_i35_2_lut (.I0(n3157), .I1(baudrate[16]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_4470));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_2791_10_lut (.I0(GND_net), .I1(n2838), .I2(n1742), .I3(n52147), 
            .O(n8339[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2791_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1947_add_4_3 (.CI(n52376), .I0(GND_net), .I1(r_Clock_Count[1]), 
            .CO(n52377));
    SB_LUT4 div_37_i2128_3_lut (.I0(n3056), .I1(n8391[13]), .I2(n294[2]), 
            .I3(GND_net), .O(n3161));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2128_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2129_3_lut (.I0(n3057), .I1(n8391[12]), .I2(n294[2]), 
            .I3(GND_net), .O(n3162));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2129_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2778_5 (.CI(n51988), .I0(n1114), .I1(n856), .CO(n51989));
    SB_CARRY add_2791_10 (.CI(n52147), .I0(n2838), .I1(n1742), .CO(n52148));
    SB_LUT4 div_37_LessThan_2141_i25_2_lut (.I0(n3162), .I1(baudrate[11]), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_4471));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_2141_i27_2_lut (.I0(n3161), .I1(baudrate[12]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_4472));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 sub_38_add_2_23_lut (.I0(o_Rx_DV_N_3488[18]), .I1(n294[21]), 
            .I2(VCC_net), .I3(n51138), .O(n23)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_23_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_38_add_2_23 (.CI(n51138), .I0(n294[21]), .I1(VCC_net), 
            .CO(n51139));
    SB_LUT4 div_37_i2137_3_lut (.I0(n3065), .I1(n8391[4]), .I2(n294[2]), 
            .I3(GND_net), .O(n3170));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2137_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2138_3_lut (.I0(n3066), .I1(n8391[3]), .I2(n294[2]), 
            .I3(GND_net), .O(n3171));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2138_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2141_i9_2_lut (.I0(n3170), .I1(baudrate[3]), 
            .I2(GND_net), .I3(GND_net), .O(n9_adj_4473));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i2130_3_lut (.I0(n3058), .I1(n8391[11]), .I2(n294[2]), 
            .I3(GND_net), .O(n3163));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2130_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2131_3_lut (.I0(n3059), .I1(n8391[10]), .I2(n294[2]), 
            .I3(GND_net), .O(n3164));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2131_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2141_i21_2_lut (.I0(n3164), .I1(baudrate[9]), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_4474));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 sub_38_add_2_22_lut (.I0(n62091), .I1(n294[20]), .I2(VCC_net), 
            .I3(n51137), .O(n62093)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_22_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 div_37_LessThan_2141_i23_2_lut (.I0(n3163), .I1(baudrate[10]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_4475));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i2127_3_lut (.I0(n3055), .I1(n8391[14]), .I2(n294[2]), 
            .I3(GND_net), .O(n3160));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2127_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2134_3_lut (.I0(n3062), .I1(n8391[7]), .I2(n294[2]), 
            .I3(GND_net), .O(n3167));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2134_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2133_3_lut (.I0(n3061), .I1(n8391[8]), .I2(n294[2]), 
            .I3(GND_net), .O(n3166));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2133_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2778_4_lut (.I0(GND_net), .I1(n1115), .I2(n698), .I3(n51987), 
            .O(n8001[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2778_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_2141_i13_2_lut (.I0(n3168), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n13_adj_4476));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_2141_i15_2_lut (.I0(n3167), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_4477));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i15_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_2778_4 (.CI(n51987), .I0(n1115), .I1(n698), .CO(n51988));
    SB_LUT4 add_2778_3_lut (.I0(GND_net), .I1(n1116), .I2(n858), .I3(n51986), 
            .O(n8001[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2778_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2778_3 (.CI(n51986), .I0(n1116), .I1(n858), .CO(n51987));
    SB_LUT4 r_Clock_Count_1947_add_4_2_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[0]), .I3(VCC_net), .O(n1[0])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1947_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_38_add_2_22 (.CI(n51137), .I0(n294[20]), .I1(VCC_net), 
            .CO(n51138));
    SB_LUT4 add_2791_9_lut (.I0(GND_net), .I1(n2839), .I2(n1602), .I3(n52146), 
            .O(n8339[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2791_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2778_2_lut (.I0(n59844), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n62035)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2778_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_2791_9 (.CI(n52146), .I0(n2839), .I1(n1602), .CO(n52147));
    SB_CARRY r_Clock_Count_1947_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(r_Clock_Count[0]), 
            .CO(n52376));
    SB_LUT4 div_37_LessThan_2141_i17_2_lut (.I0(n3166), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_4479));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_2141_i29_2_lut (.I0(n3160), .I1(baudrate[13]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_4480));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i2136_3_lut (.I0(n3064), .I1(n8391[5]), .I2(n294[2]), 
            .I3(GND_net), .O(n3169));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2136_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2778_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n51986));
    SB_LUT4 div_37_i2132_3_lut (.I0(n3060), .I1(n8391[9]), .I2(n294[2]), 
            .I3(GND_net), .O(n3165));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2132_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2141_i11_2_lut (.I0(n3169), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_4481));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_2141_i19_2_lut (.I0(n3165), .I1(baudrate[8]), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_4482));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_967 (.I0(baudrate[26]), .I1(baudrate[30]), .I2(GND_net), 
            .I3(GND_net), .O(n63609));
    defparam i1_2_lut_adj_967.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_968 (.I0(n63613), .I1(n63615), .I2(n63461), .I3(n63611), 
            .O(n25589));
    defparam i1_4_lut_adj_968.LUT_INIT = 16'hfffe;
    SB_LUT4 i51600_4_lut (.I0(n29_adj_4480), .I1(n17_adj_4479), .I2(n15_adj_4477), 
            .I3(n13_adj_4476), .O(n67294));
    defparam i51600_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 add_2791_8_lut (.I0(GND_net), .I1(n2840), .I2(n1459), .I3(n52145), 
            .O(n8339[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2791_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i52527_4_lut (.I0(n11_adj_4481), .I1(n9_adj_4473), .I2(n3171), 
            .I3(baudrate[2]), .O(n68221));
    defparam i52527_4_lut.LUT_INIT = 16'heffe;
    SB_LUT4 i53230_4_lut (.I0(n17_adj_4479), .I1(n15_adj_4477), .I2(n13_adj_4476), 
            .I3(n68221), .O(n68924));
    defparam i53230_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i53228_4_lut (.I0(n23_adj_4475), .I1(n21_adj_4474), .I2(n19_adj_4482), 
            .I3(n68924), .O(n68922));
    defparam i53228_4_lut.LUT_INIT = 16'hfeff;
    SB_CARRY add_2791_8 (.CI(n52145), .I0(n2840), .I1(n1459), .CO(n52146));
    SB_LUT4 i51602_4_lut (.I0(n29_adj_4480), .I1(n27_adj_4472), .I2(n25_adj_4471), 
            .I3(n68922), .O(n67296));
    defparam i51602_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_37_LessThan_2141_i6_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n3172), .I3(GND_net), .O(n6_adj_4483));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i6_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i53796_3_lut (.I0(n6_adj_4483), .I1(baudrate[13]), .I2(n29_adj_4480), 
            .I3(GND_net), .O(n69490));   // verilog/uart_rx.v(119[33:55])
    defparam i53796_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2791_7_lut (.I0(GND_net), .I1(n2841), .I2(n1460), .I3(n52144), 
            .O(n8339[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2791_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2791_7 (.CI(n52144), .I0(n2841), .I1(n1460), .CO(n52145));
    SB_LUT4 add_2791_6_lut (.I0(GND_net), .I1(n2842), .I2(n1011), .I3(n52143), 
            .O(n8339[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2791_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2791_6 (.CI(n52143), .I0(n2842), .I1(n1011), .CO(n52144));
    SB_LUT4 add_2791_5_lut (.I0(GND_net), .I1(n2843), .I2(n856), .I3(n52142), 
            .O(n8339[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2791_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_2141_i32_3_lut (.I0(n14), .I1(baudrate[17]), 
            .I2(n37_adj_4469), .I3(GND_net), .O(n32));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i32_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2791_5 (.CI(n52142), .I0(n2843), .I1(n856), .CO(n52143));
    SB_LUT4 add_2791_4_lut (.I0(GND_net), .I1(n2844), .I2(n698), .I3(n52141), 
            .O(n8339[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2791_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2791_4 (.CI(n52141), .I0(n2844), .I1(n698), .CO(n52142));
    SB_LUT4 i53797_3_lut (.I0(n69490), .I1(baudrate[14]), .I2(n31_adj_4468), 
            .I3(GND_net), .O(n69491));   // verilog/uart_rx.v(119[33:55])
    defparam i53797_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2791_3_lut (.I0(GND_net), .I1(n2845), .I2(n858), .I3(n52140), 
            .O(n8339[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2791_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2791_3 (.CI(n52140), .I0(n2845), .I1(n858), .CO(n52141));
    SB_LUT4 add_2791_2_lut (.I0(n59798), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n62053)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2791_2_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i51596_4_lut (.I0(n35_adj_4470), .I1(n33_adj_4466), .I2(n31_adj_4468), 
            .I3(n67294), .O(n67290));
    defparam i51596_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i54147_4_lut (.I0(n32), .I1(n12_adj_4484), .I2(n37_adj_4469), 
            .I3(n67283), .O(n69841));   // verilog/uart_rx.v(119[33:55])
    defparam i54147_4_lut.LUT_INIT = 16'haaac;
    SB_CARRY add_2791_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n52140));
    SB_LUT4 i53717_3_lut (.I0(n69491), .I1(baudrate[15]), .I2(n33_adj_4466), 
            .I3(GND_net), .O(n69411));   // verilog/uart_rx.v(119[33:55])
    defparam i53717_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2790_20_lut (.I0(GND_net), .I1(n2713), .I2(n2977), .I3(n52139), 
            .O(n8313[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2790_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_38_add_2_21_lut (.I0(n62253), .I1(n294[19]), .I2(VCC_net), 
            .I3(n51136), .O(n60815)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_21_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_38_add_2_21 (.CI(n51136), .I0(n294[19]), .I1(VCC_net), 
            .CO(n51137));
    SB_LUT4 i53798_3_lut (.I0(n8_adj_4485), .I1(baudrate[10]), .I2(n23_adj_4475), 
            .I3(GND_net), .O(n69492));   // verilog/uart_rx.v(119[33:55])
    defparam i53798_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53799_3_lut (.I0(n69492), .I1(baudrate[11]), .I2(n25_adj_4471), 
            .I3(GND_net), .O(n69493));   // verilog/uart_rx.v(119[33:55])
    defparam i53799_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52517_4_lut (.I0(n25_adj_4471), .I1(n23_adj_4475), .I2(n21_adj_4474), 
            .I3(n67307), .O(n68211));
    defparam i52517_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i53714_3_lut (.I0(n10_adj_4486), .I1(baudrate[9]), .I2(n21_adj_4474), 
            .I3(GND_net), .O(n69408));   // verilog/uart_rx.v(119[33:55])
    defparam i53714_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 sub_38_add_2_20_lut (.I0(GND_net), .I1(n294[18]), .I2(VCC_net), 
            .I3(n51135), .O(o_Rx_DV_N_3488[18])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i53713_3_lut (.I0(n69493), .I1(baudrate[12]), .I2(n27_adj_4472), 
            .I3(GND_net), .O(n69407));   // verilog/uart_rx.v(119[33:55])
    defparam i53713_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2790_19_lut (.I0(GND_net), .I1(n2714), .I2(n2867), .I3(n52138), 
            .O(n8313[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2790_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_38_add_2_20 (.CI(n51135), .I0(n294[18]), .I1(VCC_net), 
            .CO(n51136));
    SB_CARRY add_2790_19 (.CI(n52138), .I0(n2714), .I1(n2867), .CO(n52139));
    SB_LUT4 i53543_4_lut (.I0(n35_adj_4470), .I1(n33_adj_4466), .I2(n31_adj_4468), 
            .I3(n67296), .O(n69237));
    defparam i53543_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i54278_4_lut (.I0(n69411), .I1(n69841), .I2(n37_adj_4469), 
            .I3(n67290), .O(n69972));   // verilog/uart_rx.v(119[33:55])
    defparam i54278_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i53792_4_lut (.I0(n69407), .I1(n69408), .I2(n27_adj_4472), 
            .I3(n68211), .O(n69486));   // verilog/uart_rx.v(119[33:55])
    defparam i53792_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 add_2790_18_lut (.I0(GND_net), .I1(n2715), .I2(n2754), .I3(n52137), 
            .O(n8313[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2790_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i54300_4_lut (.I0(n69486), .I1(n69972), .I2(n37_adj_4469), 
            .I3(n69237), .O(n69994));   // verilog/uart_rx.v(119[33:55])
    defparam i54300_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i54301_3_lut (.I0(n69994), .I1(baudrate[18]), .I2(n3155), 
            .I3(GND_net), .O(n69995));   // verilog/uart_rx.v(119[33:55])
    defparam i54301_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i54293_3_lut (.I0(n69995), .I1(baudrate[19]), .I2(n3154), 
            .I3(GND_net), .O(n69987));   // verilog/uart_rx.v(119[33:55])
    defparam i54293_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i54070_3_lut (.I0(n69987), .I1(baudrate[20]), .I2(n3153), 
            .I3(GND_net), .O(n69764));   // verilog/uart_rx.v(119[33:55])
    defparam i54070_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 sub_38_add_2_19_lut (.I0(o_Rx_DV_N_3488[10]), .I1(n294[17]), 
            .I2(VCC_net), .I3(n51134), .O(n62089)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_19_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 i54071_3_lut (.I0(n69764), .I1(baudrate[21]), .I2(n3152), 
            .I3(GND_net), .O(n69765));   // verilog/uart_rx.v(119[33:55])
    defparam i54071_3_lut.LUT_INIT = 16'h8e8e;
    SB_CARRY sub_38_add_2_19 (.CI(n51134), .I0(n294[17]), .I1(VCC_net), 
            .CO(n51135));
    SB_LUT4 i53723_3_lut (.I0(n69765), .I1(baudrate[22]), .I2(n3151), 
            .I3(GND_net), .O(n48));   // verilog/uart_rx.v(119[33:55])
    defparam i53723_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 sub_38_add_2_18_lut (.I0(n62251), .I1(n294[16]), .I2(VCC_net), 
            .I3(n51133), .O(n62253)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_18_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_38_add_2_18 (.CI(n51133), .I0(n294[16]), .I1(VCC_net), 
            .CO(n51134));
    SB_CARRY add_2790_18 (.CI(n52137), .I0(n2715), .I1(n2754), .CO(n52138));
    SB_LUT4 div_37_i2047_3_lut (.I0(n2938), .I1(n8365[23]), .I2(n294[3]), 
            .I3(GND_net), .O(n3046));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2047_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2790_17_lut (.I0(GND_net), .I1(n2716), .I2(n2638), .I3(n52136), 
            .O(n8313[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2790_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_i2055_3_lut (.I0(n2946), .I1(n8365[15]), .I2(n294[3]), 
            .I3(GND_net), .O(n3054));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2055_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2048_3_lut (.I0(n2939), .I1(n8365[22]), .I2(n294[3]), 
            .I3(GND_net), .O(n3047));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2048_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2049_3_lut (.I0(n2940), .I1(n8365[21]), .I2(n294[3]), 
            .I3(GND_net), .O(n3048));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2049_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2050_3_lut (.I0(n2941), .I1(n8365[20]), .I2(n294[3]), 
            .I3(GND_net), .O(n3049));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2050_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2053_3_lut (.I0(n2944), .I1(n8365[17]), .I2(n294[3]), 
            .I3(GND_net), .O(n3052));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2053_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2070_i35_2_lut (.I0(n3052), .I1(baudrate[15]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_4487));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 sub_38_add_2_17_lut (.I0(n61997), .I1(n294[15]), .I2(VCC_net), 
            .I3(n51132), .O(n61999)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_17_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_38_add_2_17 (.CI(n51132), .I0(n294[15]), .I1(VCC_net), 
            .CO(n51133));
    SB_LUT4 div_37_i2051_3_lut (.I0(n2942), .I1(n8365[19]), .I2(n294[3]), 
            .I3(GND_net), .O(n3050));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2051_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2790_17 (.CI(n52136), .I0(n2716), .I1(n2638), .CO(n52137));
    SB_LUT4 div_37_LessThan_2070_i39_2_lut (.I0(n3050), .I1(baudrate[17]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_4488));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_2790_16_lut (.I0(GND_net), .I1(n2717), .I2(n2519), .I3(n52135), 
            .O(n8313[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2790_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_38_add_2_16_lut (.I0(o_Rx_DV_N_3488[13]), .I1(n294[14]), 
            .I2(VCC_net), .I3(n51131), .O(n62251)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_16_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_38_add_2_16 (.CI(n51131), .I0(n294[14]), .I1(VCC_net), 
            .CO(n51132));
    SB_LUT4 div_37_i2054_3_lut (.I0(n2945), .I1(n8365[16]), .I2(n294[3]), 
            .I3(GND_net), .O(n3053));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2054_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2790_16 (.CI(n52135), .I0(n2717), .I1(n2519), .CO(n52136));
    SB_LUT4 add_2790_15_lut (.I0(GND_net), .I1(n2718), .I2(n2397), .I3(n52134), 
            .O(n8313[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2790_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_38_add_2_15_lut (.I0(GND_net), .I1(n294[13]), .I2(VCC_net), 
            .I3(n51130), .O(o_Rx_DV_N_3488[13])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_38_add_2_15 (.CI(n51130), .I0(n294[13]), .I1(VCC_net), 
            .CO(n51131));
    SB_LUT4 div_37_LessThan_2070_i33_2_lut (.I0(n3053), .I1(baudrate[14]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_4489));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i2052_3_lut (.I0(n2943), .I1(n8365[18]), .I2(n294[3]), 
            .I3(GND_net), .O(n3051));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2052_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2070_i37_2_lut (.I0(n3051), .I1(baudrate[16]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_4490));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_2070_i23_2_lut (.I0(n3058), .I1(baudrate[9]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_4491));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_2070_i25_2_lut (.I0(n3057), .I1(baudrate[10]), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_4492));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i2056_3_lut (.I0(n2947), .I1(n8365[14]), .I2(n294[3]), 
            .I3(GND_net), .O(n3055));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2056_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2790_15 (.CI(n52134), .I0(n2718), .I1(n2397), .CO(n52135));
    SB_LUT4 sub_38_add_2_14_lut (.I0(GND_net), .I1(n294[12]), .I2(VCC_net), 
            .I3(n51129), .O(\o_Rx_DV_N_3488[12] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_38_add_2_14 (.CI(n51129), .I0(n294[12]), .I1(VCC_net), 
            .CO(n51130));
    SB_LUT4 add_2790_14_lut (.I0(GND_net), .I1(n2719), .I2(n2272), .I3(n52133), 
            .O(n8313[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2790_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2790_14 (.CI(n52133), .I0(n2719), .I1(n2272), .CO(n52134));
    SB_LUT4 sub_38_add_2_13_lut (.I0(o_Rx_DV_N_3488[9]), .I1(n294[11]), 
            .I2(VCC_net), .I3(n51128), .O(n61997)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_13_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 add_2790_13_lut (.I0(GND_net), .I1(n2720), .I2(n2144), .I3(n52132), 
            .O(n8313[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2790_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_2070_i27_2_lut (.I0(n3056), .I1(baudrate[11]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_4493));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_2070_i29_2_lut (.I0(n3055), .I1(baudrate[12]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_4494));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i29_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_2790_13 (.CI(n52132), .I0(n2720), .I1(n2144), .CO(n52133));
    SB_LUT4 div_37_LessThan_2070_i11_2_lut (.I0(n3064), .I1(baudrate[3]), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_4495));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_2070_i13_2_lut (.I0(n3063), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n13_adj_4496));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_2070_i21_2_lut (.I0(n3059), .I1(baudrate[8]), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_4497));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_2070_i15_2_lut (.I0(n3062), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_4498));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_2790_12_lut (.I0(GND_net), .I1(n2721), .I2(n2013), .I3(n52131), 
            .O(n8313[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2790_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_2070_i17_2_lut (.I0(n3061), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_4499));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_2070_i19_2_lut (.I0(n3060), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_4500));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_2070_i31_2_lut (.I0(n3054), .I1(baudrate[13]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_4501));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i51644_4_lut (.I0(n31_adj_4501), .I1(n19_adj_4500), .I2(n17_adj_4499), 
            .I3(n15_adj_4498), .O(n67338));
    defparam i51644_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i52616_4_lut (.I0(n13_adj_4496), .I1(n11_adj_4495), .I2(n3065), 
            .I3(baudrate[2]), .O(n68310));
    defparam i52616_4_lut.LUT_INIT = 16'heffe;
    SB_LUT4 i53250_4_lut (.I0(n19_adj_4500), .I1(n17_adj_4499), .I2(n15_adj_4498), 
            .I3(n68310), .O(n68944));
    defparam i53250_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i53244_4_lut (.I0(n25_adj_4492), .I1(n23_adj_4491), .I2(n21_adj_4497), 
            .I3(n68944), .O(n68938));
    defparam i53244_4_lut.LUT_INIT = 16'hfeff;
    SB_CARRY sub_38_add_2_13 (.CI(n51128), .I0(n294[11]), .I1(VCC_net), 
            .CO(n51129));
    SB_LUT4 i51646_4_lut (.I0(n31_adj_4501), .I1(n29_adj_4494), .I2(n27_adj_4493), 
            .I3(n68938), .O(n67340));
    defparam i51646_4_lut.LUT_INIT = 16'haaab;
    SB_CARRY add_2790_12 (.CI(n52131), .I0(n2721), .I1(n2013), .CO(n52132));
    SB_LUT4 div_37_LessThan_2070_i8_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n3066), .I3(GND_net), .O(n8_adj_4502));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i8_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i53802_3_lut (.I0(n8_adj_4502), .I1(baudrate[13]), .I2(n31_adj_4501), 
            .I3(GND_net), .O(n69496));   // verilog/uart_rx.v(119[33:55])
    defparam i53802_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 sub_38_add_2_12_lut (.I0(GND_net), .I1(n294[10]), .I2(VCC_net), 
            .I3(n51127), .O(o_Rx_DV_N_3488[10])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_38_add_2_12 (.CI(n51127), .I0(n294[10]), .I1(VCC_net), 
            .CO(n51128));
    SB_LUT4 i53803_3_lut (.I0(n69496), .I1(baudrate[14]), .I2(n33_adj_4489), 
            .I3(GND_net), .O(n69497));   // verilog/uart_rx.v(119[33:55])
    defparam i53803_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 sub_38_add_2_11_lut (.I0(GND_net), .I1(n294[9]), .I2(VCC_net), 
            .I3(n51126), .O(o_Rx_DV_N_3488[9])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2790_11_lut (.I0(GND_net), .I1(n2722), .I2(n1879), .I3(n52130), 
            .O(n8313[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2790_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_2070_i34_3_lut (.I0(n16_adj_4503), .I1(baudrate[17]), 
            .I2(n39_adj_4488), .I3(GND_net), .O(n34));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i34_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51638_4_lut (.I0(n37_adj_4490), .I1(n35_adj_4487), .I2(n33_adj_4489), 
            .I3(n67338), .O(n67332));
    defparam i51638_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i54145_4_lut (.I0(n34), .I1(n14_adj_4504), .I2(n39_adj_4488), 
            .I3(n67329), .O(n69839));   // verilog/uart_rx.v(119[33:55])
    defparam i54145_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i53705_3_lut (.I0(n69497), .I1(baudrate[15]), .I2(n35_adj_4487), 
            .I3(GND_net), .O(n69399));   // verilog/uart_rx.v(119[33:55])
    defparam i53705_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53804_3_lut (.I0(n10_adj_4505), .I1(baudrate[10]), .I2(n25_adj_4492), 
            .I3(GND_net), .O(n69498));   // verilog/uart_rx.v(119[33:55])
    defparam i53804_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY sub_38_add_2_11 (.CI(n51126), .I0(n294[9]), .I1(VCC_net), 
            .CO(n51127));
    SB_LUT4 i53805_3_lut (.I0(n69498), .I1(baudrate[11]), .I2(n27_adj_4493), 
            .I3(GND_net), .O(n69499));   // verilog/uart_rx.v(119[33:55])
    defparam i53805_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 sub_38_add_2_10_lut (.I0(GND_net), .I1(n294[8]), .I2(VCC_net), 
            .I3(n51125), .O(\o_Rx_DV_N_3488[8] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i52545_4_lut (.I0(n27_adj_4493), .I1(n25_adj_4492), .I2(n23_adj_4491), 
            .I3(n67365), .O(n68239));
    defparam i52545_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 div_37_LessThan_2070_i20_3_lut (.I0(n12_adj_4506), .I1(baudrate[9]), 
            .I2(n23_adj_4491), .I3(GND_net), .O(n20));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i20_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53703_3_lut (.I0(n69499), .I1(baudrate[12]), .I2(n29_adj_4494), 
            .I3(GND_net), .O(n69397));   // verilog/uart_rx.v(119[33:55])
    defparam i53703_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53549_4_lut (.I0(n37_adj_4490), .I1(n35_adj_4487), .I2(n33_adj_4489), 
            .I3(n67340), .O(n69243));
    defparam i53549_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i54276_4_lut (.I0(n69399), .I1(n69839), .I2(n39_adj_4488), 
            .I3(n67332), .O(n69970));   // verilog/uart_rx.v(119[33:55])
    defparam i54276_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i53708_4_lut (.I0(n69397), .I1(n20), .I2(n29_adj_4494), .I3(n68239), 
            .O(n69402));   // verilog/uart_rx.v(119[33:55])
    defparam i53708_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i54302_4_lut (.I0(n69402), .I1(n69970), .I2(n39_adj_4488), 
            .I3(n69243), .O(n69996));   // verilog/uart_rx.v(119[33:55])
    defparam i54302_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i54303_3_lut (.I0(n69996), .I1(baudrate[18]), .I2(n3049), 
            .I3(GND_net), .O(n69997));   // verilog/uart_rx.v(119[33:55])
    defparam i54303_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i54291_3_lut (.I0(n69997), .I1(baudrate[19]), .I2(n3048), 
            .I3(GND_net), .O(n69985));   // verilog/uart_rx.v(119[33:55])
    defparam i54291_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i53710_3_lut (.I0(n69985), .I1(baudrate[20]), .I2(n3047), 
            .I3(GND_net), .O(n69404));   // verilog/uart_rx.v(119[33:55])
    defparam i53710_3_lut.LUT_INIT = 16'h8e8e;
    SB_CARRY sub_38_add_2_10 (.CI(n51125), .I0(n294[8]), .I1(VCC_net), 
            .CO(n51126));
    SB_LUT4 div_37_LessThan_1430_i31_2_lut (.I0(n2106), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_4507));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1430_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1430_i29_2_lut (.I0(n2107), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_4508));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1430_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1430_i33_2_lut (.I0(n2105), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_4509));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1430_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 sub_38_add_2_9_lut (.I0(GND_net), .I1(n294[7]), .I2(VCC_net), 
            .I3(n51124), .O(\o_Rx_DV_N_3488[7] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_1430_i35_2_lut (.I0(n2104), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_4510));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1430_i35_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_2790_11 (.CI(n52130), .I0(n2722), .I1(n1879), .CO(n52131));
    SB_LUT4 add_2790_10_lut (.I0(GND_net), .I1(n2723), .I2(n1742), .I3(n52129), 
            .O(n8313[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2790_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_1430_i39_2_lut (.I0(n2102), .I1(baudrate[9]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_4511));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1430_i39_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_2790_10 (.CI(n52129), .I0(n2723), .I1(n1742), .CO(n52130));
    SB_CARRY sub_38_add_2_9 (.CI(n51124), .I0(n294[7]), .I1(VCC_net), 
            .CO(n51125));
    SB_LUT4 div_37_LessThan_1685_i25_2_lut (.I0(n2487), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_4512));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1062_i39_2_lut (.I0(n1556), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_4513));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1062_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 sub_38_add_2_8_lut (.I0(GND_net), .I1(n294[6]), .I2(VCC_net), 
            .I3(n51123), .O(\o_Rx_DV_N_3488[6] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2790_9_lut (.I0(GND_net), .I1(n2724), .I2(n1602), .I3(n52128), 
            .O(n8313[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2790_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_38_add_2_8 (.CI(n51123), .I0(n294[6]), .I1(VCC_net), 
            .CO(n51124));
    SB_LUT4 div_37_LessThan_1062_i41_2_lut (.I0(n1555), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_4514));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1062_i41_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_2790_9 (.CI(n52128), .I0(n2724), .I1(n1602), .CO(n52129));
    SB_LUT4 add_2790_8_lut (.I0(GND_net), .I1(n2725), .I2(n1459), .I3(n52127), 
            .O(n8313[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2790_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2790_8 (.CI(n52127), .I0(n2725), .I1(n1459), .CO(n52128));
    SB_LUT4 div_37_LessThan_1062_i37_2_lut (.I0(n1557), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_4515));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1062_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_2790_7_lut (.I0(GND_net), .I1(n2726), .I2(n1460), .I3(n52126), 
            .O(n8313[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2790_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2790_7 (.CI(n52126), .I0(n2726), .I1(n1460), .CO(n52127));
    SB_LUT4 sub_38_add_2_7_lut (.I0(GND_net), .I1(n294[5]), .I2(VCC_net), 
            .I3(n51122), .O(\o_Rx_DV_N_3488[5] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2790_6_lut (.I0(GND_net), .I1(n2727), .I2(n1011), .I3(n52125), 
            .O(n8313[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2790_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2790_6 (.CI(n52125), .I0(n2727), .I1(n1011), .CO(n52126));
    SB_LUT4 div_37_LessThan_1250_i33_2_lut (.I0(n1838), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_4516));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1250_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1250_i31_2_lut (.I0(n1839), .I1(baudrate[3]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_4517));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1250_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1250_i35_2_lut (.I0(n1837), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_4518));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1250_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1250_i37_2_lut (.I0(n1836), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_4519));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1250_i37_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY sub_38_add_2_7 (.CI(n51122), .I0(n294[5]), .I1(VCC_net), 
            .CO(n51123));
    SB_LUT4 div_37_LessThan_1250_i41_2_lut (.I0(n1834), .I1(baudrate[8]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_4520));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1250_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_2790_5_lut (.I0(GND_net), .I1(n2728), .I2(n856), .I3(n52124), 
            .O(n8313[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2790_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2790_5 (.CI(n52124), .I0(n2728), .I1(n856), .CO(n52125));
    SB_LUT4 add_2790_4_lut (.I0(GND_net), .I1(n2729), .I2(n698), .I3(n52123), 
            .O(n8313[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2790_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2790_4 (.CI(n52123), .I0(n2729), .I1(n698), .CO(n52124));
    SB_LUT4 add_2790_3_lut (.I0(GND_net), .I1(n2730), .I2(n858), .I3(n52122), 
            .O(n8313[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2790_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_1250_i39_2_lut (.I0(n1835), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_4521));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1250_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1517_i29_2_lut (.I0(n2236), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_4522));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1517_i31_2_lut (.I0(n2235), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_4523));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1517_i27_2_lut (.I0(n2237), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_4524));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1517_i35_2_lut (.I0(n2233), .I1(baudrate[8]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_4525));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1517_i25_2_lut (.I0(n2238), .I1(baudrate[3]), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_4526));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i44156_1_lut (.I0(n25577), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n59802));
    defparam i44156_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_LessThan_1517_i37_2_lut (.I0(n2232), .I1(baudrate[9]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_4527));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1517_i39_2_lut (.I0(n2231), .I1(baudrate[10]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_4528));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i39_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_2790_3 (.CI(n52122), .I0(n2730), .I1(n858), .CO(n52123));
    SB_LUT4 sub_38_add_2_6_lut (.I0(GND_net), .I1(n294[4]), .I2(VCC_net), 
            .I3(n51121), .O(\o_Rx_DV_N_3488[4] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2790_2_lut (.I0(n59802), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n62051)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2790_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY sub_38_add_2_6 (.CI(n51121), .I0(n294[4]), .I1(VCC_net), 
            .CO(n51122));
    SB_CARRY add_2790_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n52122));
    SB_LUT4 div_37_LessThan_1517_i41_2_lut (.I0(n2230), .I1(baudrate[11]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_4529));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1517_i33_2_lut (.I0(n2234), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_4530));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_2789_19_lut (.I0(GND_net), .I1(n2596), .I2(n2867), .I3(n52121), 
            .O(n8287[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2789_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_38_add_2_5_lut (.I0(GND_net), .I1(n294[3]), .I2(VCC_net), 
            .I3(n51120), .O(\o_Rx_DV_N_3488[3] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_38_add_2_5 (.CI(n51120), .I0(n294[3]), .I1(VCC_net), 
            .CO(n51121));
    SB_LUT4 add_2789_18_lut (.I0(GND_net), .I1(n2597), .I2(n2754), .I3(n52120), 
            .O(n8287[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2789_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2789_18 (.CI(n52120), .I0(n2597), .I1(n2754), .CO(n52121));
    SB_LUT4 div_37_LessThan_1517_i43_2_lut (.I0(n2229), .I1(baudrate[12]), 
            .I2(GND_net), .I3(GND_net), .O(n43_adj_4531));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_2789_17_lut (.I0(GND_net), .I1(n2598), .I2(n2638), .I3(n52119), 
            .O(n8287[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2789_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2789_17 (.CI(n52119), .I0(n2598), .I1(n2638), .CO(n52120));
    SB_LUT4 add_2789_16_lut (.I0(GND_net), .I1(n2599), .I2(n2519), .I3(n52118), 
            .O(n8287[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2789_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2789_16 (.CI(n52118), .I0(n2599), .I1(n2519), .CO(n52119));
    SB_LUT4 i48485_2_lut (.I0(baudrate[3]), .I1(baudrate[4]), .I2(GND_net), 
            .I3(GND_net), .O(n64170));
    defparam i48485_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i29173_2_lut (.I0(baudrate[1]), .I1(baudrate[0]), .I2(GND_net), 
            .I3(GND_net), .O(n43066));
    defparam i29173_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i7218_4_lut (.I0(n804), .I1(n43066), .I2(n20902), .I3(baudrate[2]), 
            .O(n20904));   // verilog/uart_rx.v(119[33:55])
    defparam i7218_4_lut.LUT_INIT = 16'ha2aa;
    SB_LUT4 add_2789_15_lut (.I0(GND_net), .I1(n2600), .I2(n2397), .I3(n52117), 
            .O(n8287[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2789_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i7224_4_lut (.I0(n961), .I1(baudrate[2]), .I2(n962), .I3(baudrate[1]), 
            .O(n20912));   // verilog/uart_rx.v(119[33:55])
    defparam i7224_4_lut.LUT_INIT = 16'ha2aa;
    SB_CARRY add_2789_15 (.CI(n52117), .I0(n2600), .I1(n2397), .CO(n52118));
    SB_LUT4 add_2789_14_lut (.I0(GND_net), .I1(n2601), .I2(n2272), .I3(n52116), 
            .O(n8287[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2789_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2789_14 (.CI(n52116), .I0(n2601), .I1(n2272), .CO(n52117));
    SB_LUT4 div_37_i2172_1_lut (.I0(baudrate[3]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n856));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2172_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_LessThan_866_i41_2_lut (.I0(n1264), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_4532));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_866_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1602_i27_2_lut (.I0(n2363), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_4533));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 sub_38_add_2_4_lut (.I0(GND_net), .I1(n294[2]), .I2(VCC_net), 
            .I3(n51119), .O(\o_Rx_DV_N_3488[2] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_1602_i29_2_lut (.I0(n2362), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_4534));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_2789_13_lut (.I0(GND_net), .I1(n2602), .I2(n2144), .I3(n52115), 
            .O(n8287[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2789_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2789_13 (.CI(n52115), .I0(n2602), .I1(n2144), .CO(n52116));
    SB_LUT4 add_2789_12_lut (.I0(GND_net), .I1(n2603), .I2(n2013), .I3(n52114), 
            .O(n8287[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2789_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_38_add_2_4 (.CI(n51119), .I0(n294[2]), .I1(VCC_net), 
            .CO(n51120));
    SB_CARRY add_2789_12 (.CI(n52114), .I0(n2603), .I1(n2013), .CO(n52115));
    SB_LUT4 add_2789_11_lut (.I0(GND_net), .I1(n2604), .I2(n1879), .I3(n52113), 
            .O(n8287[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2789_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2789_11 (.CI(n52113), .I0(n2604), .I1(n1879), .CO(n52114));
    SB_LUT4 add_2789_10_lut (.I0(GND_net), .I1(n2605), .I2(n1742), .I3(n52112), 
            .O(n8287[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2789_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2789_10 (.CI(n52112), .I0(n2605), .I1(n1742), .CO(n52113));
    SB_LUT4 add_2789_9_lut (.I0(GND_net), .I1(n2606), .I2(n1602), .I3(n52111), 
            .O(n8287[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2789_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_38_add_2_3_lut (.I0(GND_net), .I1(n294[1]), .I2(VCC_net), 
            .I3(n51118), .O(\o_Rx_DV_N_3488[1] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2789_9 (.CI(n52111), .I0(n2606), .I1(n1602), .CO(n52112));
    SB_LUT4 add_2789_8_lut (.I0(GND_net), .I1(n2607), .I2(n1459), .I3(n52110), 
            .O(n8287[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2789_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2789_8 (.CI(n52110), .I0(n2607), .I1(n1459), .CO(n52111));
    SB_LUT4 add_2789_7_lut (.I0(GND_net), .I1(n2608), .I2(n1460), .I3(n52109), 
            .O(n8287[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2789_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_38_add_2_3 (.CI(n51118), .I0(n294[1]), .I1(VCC_net), 
            .CO(n51119));
    SB_CARRY add_2789_7 (.CI(n52109), .I0(n2608), .I1(n1460), .CO(n52110));
    SB_LUT4 sub_38_add_2_2_lut (.I0(GND_net), .I1(n60953), .I2(GND_net), 
            .I3(VCC_net), .O(\o_Rx_DV_N_3488[0] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_38_add_2_2 (.CI(VCC_net), .I0(n60953), .I1(GND_net), 
            .CO(n51118));
    SB_LUT4 i54477_3_lut (.I0(n25598), .I1(baudrate[1]), .I2(baudrate[2]), 
            .I3(GND_net), .O(n25515));   // verilog/uart_rx.v(119[33:55])
    defparam i54477_3_lut.LUT_INIT = 16'h0101;
    SB_LUT4 add_2789_6_lut (.I0(GND_net), .I1(n2609), .I2(n1011), .I3(n52108), 
            .O(n8287[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2789_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2789_6 (.CI(n52108), .I0(n2609), .I1(n1011), .CO(n52109));
    SB_LUT4 add_2789_5_lut (.I0(GND_net), .I1(n2610), .I2(n856), .I3(n52107), 
            .O(n8287[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2789_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2789_5 (.CI(n52107), .I0(n2610), .I1(n856), .CO(n52108));
    SB_LUT4 add_2789_4_lut (.I0(GND_net), .I1(n2611), .I2(n698), .I3(n52106), 
            .O(n8287[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2789_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2789_4 (.CI(n52106), .I0(n2611), .I1(n698), .CO(n52107));
    SB_LUT4 add_2789_3_lut (.I0(GND_net), .I1(n2612), .I2(n858), .I3(n52105), 
            .O(n8287[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2789_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2789_3 (.CI(n52105), .I0(n2612), .I1(n858), .CO(n52106));
    SB_LUT4 add_2789_2_lut (.I0(n59806), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n62049)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2789_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_2789_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n52105));
    SB_LUT4 add_2788_18_lut (.I0(GND_net), .I1(n2476), .I2(n2754), .I3(n52104), 
            .O(n8261[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2788_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_i2166_1_lut (.I0(baudrate[9]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1879));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2166_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_2788_17_lut (.I0(GND_net), .I1(n2477), .I2(n2638), .I3(n52103), 
            .O(n8261[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2788_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2788_17 (.CI(n52103), .I0(n2477), .I1(n2638), .CO(n52104));
    SB_LUT4 div_37_i2059_3_lut (.I0(n2950), .I1(n8365[11]), .I2(n294[3]), 
            .I3(GND_net), .O(n3058));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2059_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2788_16_lut (.I0(GND_net), .I1(n2478), .I2(n2519), .I3(n52102), 
            .O(n8261[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2788_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_i2171_1_lut (.I0(baudrate[4]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1011));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2171_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_2788_16 (.CI(n52102), .I0(n2478), .I1(n2519), .CO(n52103));
    SB_LUT4 add_2788_15_lut (.I0(GND_net), .I1(n2479), .I2(n2397), .I3(n52101), 
            .O(n8261[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2788_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2788_15 (.CI(n52101), .I0(n2479), .I1(n2397), .CO(n52102));
    SB_LUT4 add_2788_14_lut (.I0(GND_net), .I1(n2480), .I2(n2272), .I3(n52100), 
            .O(n8261[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2788_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2788_14 (.CI(n52100), .I0(n2480), .I1(n2272), .CO(n52101));
    SB_LUT4 add_2788_13_lut (.I0(GND_net), .I1(n2481), .I2(n2144), .I3(n52099), 
            .O(n8261[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2788_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2788_13 (.CI(n52099), .I0(n2481), .I1(n2144), .CO(n52100));
    SB_LUT4 add_2788_12_lut (.I0(GND_net), .I1(n2482), .I2(n2013), .I3(n52098), 
            .O(n8261[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2788_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2788_12 (.CI(n52098), .I0(n2482), .I1(n2013), .CO(n52099));
    SB_LUT4 add_2788_11_lut (.I0(GND_net), .I1(n2483), .I2(n1879), .I3(n52097), 
            .O(n8261[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2788_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i52238_4_lut (.I0(r_SM_Main[0]), .I1(\o_Rx_DV_N_3488[12] ), 
            .I2(n4935), .I3(\o_Rx_DV_N_3488[8] ), .O(n67076));   // verilog/uart_rx.v(53[7] 144[14])
    defparam i52238_4_lut.LUT_INIT = 16'hfffd;
    SB_LUT4 i52278_4_lut (.I0(r_Rx_Data), .I1(\o_Rx_DV_N_3488[12] ), .I2(n58444), 
            .I3(r_SM_Main[0]), .O(n67082));   // verilog/uart_rx.v(53[7] 144[14])
    defparam i52278_4_lut.LUT_INIT = 16'h0100;
    SB_LUT4 div_37_i2165_1_lut (.I0(baudrate[10]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2013));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2165_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i2058_3_lut (.I0(n2949), .I1(n8365[12]), .I2(n294[3]), 
            .I3(GND_net), .O(n3057));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2058_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2788_11 (.CI(n52097), .I0(n2483), .I1(n1879), .CO(n52098));
    SB_LUT4 i52235_4_lut (.I0(n67076), .I1(\o_Rx_DV_N_3488[24] ), .I2(n29), 
            .I3(n23), .O(n67073));   // verilog/uart_rx.v(53[7] 144[14])
    defparam i52235_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_i1974_3_lut (.I0(n2827), .I1(n8339[23]), .I2(n294[4]), 
            .I3(GND_net), .O(n2938));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1974_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52243_4_lut (.I0(n67082), .I1(\o_Rx_DV_N_3488[24] ), .I2(n29), 
            .I3(n23), .O(n67079));   // verilog/uart_rx.v(53[7] 144[14])
    defparam i52243_4_lut.LUT_INIT = 16'h0002;
    SB_LUT4 r_SM_Main_2__I_0_62_Mux_1_i3_4_lut (.I0(n67079), .I1(n67073), 
            .I2(\r_SM_Main[1] ), .I3(n27), .O(n3_adj_4535));   // verilog/uart_rx.v(53[7] 144[14])
    defparam r_SM_Main_2__I_0_62_Mux_1_i3_4_lut.LUT_INIT = 16'hf0ca;
    SB_LUT4 div_37_i1976_3_lut (.I0(n2829), .I1(n8339[21]), .I2(n294[4]), 
            .I3(GND_net), .O(n2940));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1976_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1975_3_lut (.I0(n2828), .I1(n8339[22]), .I2(n294[4]), 
            .I3(GND_net), .O(n2939));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1975_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1979_3_lut (.I0(n2832), .I1(n8339[18]), .I2(n294[4]), 
            .I3(GND_net), .O(n2943));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1979_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1997_i37_2_lut (.I0(n2943), .I1(baudrate[15]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_4536));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1977_3_lut (.I0(n2830), .I1(n8339[20]), .I2(n294[4]), 
            .I3(GND_net), .O(n2941));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1977_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1997_i41_2_lut (.I0(n2941), .I1(baudrate[17]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_4537));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1980_3_lut (.I0(n2833), .I1(n8339[17]), .I2(n294[4]), 
            .I3(GND_net), .O(n2944));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1980_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1997_i35_2_lut (.I0(n2944), .I1(baudrate[14]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_4538));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1978_3_lut (.I0(n2831), .I1(n8339[19]), .I2(n294[4]), 
            .I3(GND_net), .O(n2942));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1978_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1997_i39_2_lut (.I0(n2942), .I1(baudrate[16]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_4539));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1986_3_lut (.I0(n2839), .I1(n8339[11]), .I2(n294[4]), 
            .I3(GND_net), .O(n2950));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1986_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1985_3_lut (.I0(n2838), .I1(n8339[12]), .I2(n294[4]), 
            .I3(GND_net), .O(n2949));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1985_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1997_i23_2_lut (.I0(n2950), .I1(baudrate[8]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_4540));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1997_i25_2_lut (.I0(n2949), .I1(baudrate[9]), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_4541));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1997_i27_2_lut (.I0(n2948), .I1(baudrate[10]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_4542));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i44152_1_lut (.I0(n25580), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n59798));
    defparam i44152_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i1983_3_lut (.I0(n2836), .I1(n8339[14]), .I2(n294[4]), 
            .I3(GND_net), .O(n2947));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1983_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1982_3_lut (.I0(n2835), .I1(n8339[15]), .I2(n294[4]), 
            .I3(GND_net), .O(n2946));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1982_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1997_i29_2_lut (.I0(n2947), .I1(baudrate[11]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_4543));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1997_i31_2_lut (.I0(n2946), .I1(baudrate[12]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_4544));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_4_lut (.I0(n69731), .I1(baudrate[6]), .I2(n1111), 
            .I3(n62035), .O(n1267));   // verilog/uart_rx.v(119[33:55])
    defparam i1_2_lut_4_lut.LUT_INIT = 16'h7100;
    SB_LUT4 i55097_2_lut_4_lut (.I0(n69731), .I1(baudrate[6]), .I2(n1111), 
            .I3(n64246), .O(n294[17]));   // verilog/uart_rx.v(119[33:55])
    defparam i55097_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_LUT4 i48562_1_lut (.I0(n64246), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n59844));
    defparam i48562_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i1990_3_lut (.I0(n2843), .I1(n8339[7]), .I2(n294[4]), 
            .I3(GND_net), .O(n2954));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1990_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1991_3_lut (.I0(n2844), .I1(n8339[6]), .I2(n294[4]), 
            .I3(GND_net), .O(n2955));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1991_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1992_3_lut (.I0(n2845), .I1(n8339[5]), .I2(n294[4]), 
            .I3(GND_net), .O(n2956));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1992_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1997_i13_2_lut (.I0(n2955), .I1(baudrate[3]), 
            .I2(GND_net), .I3(GND_net), .O(n13_adj_4545));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1997_i15_2_lut (.I0(n2954), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_4546));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1981_3_lut (.I0(n2834), .I1(n8339[16]), .I2(n294[4]), 
            .I3(GND_net), .O(n2945));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1981_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1997_i33_2_lut (.I0(n2945), .I1(baudrate[13]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_4547));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1987_3_lut (.I0(n2840), .I1(n8339[10]), .I2(n294[4]), 
            .I3(GND_net), .O(n2951));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1987_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1988_3_lut (.I0(n2841), .I1(n8339[9]), .I2(n294[4]), 
            .I3(GND_net), .O(n2952));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1988_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1989_3_lut (.I0(n2842), .I1(n8339[8]), .I2(n294[4]), 
            .I3(GND_net), .O(n2953));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1989_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1997_i17_2_lut (.I0(n2953), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_4548));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1997_i19_2_lut (.I0(n2952), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_4549));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1997_i21_2_lut (.I0(n2951), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_4550));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i48507_3_lut (.I0(baudrate[31]), .I1(baudrate[21]), .I2(baudrate[27]), 
            .I3(GND_net), .O(n64192));
    defparam i48507_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i48563_4_lut (.I0(n64192), .I1(n63505), .I2(n64190), .I3(n63459), 
            .O(n64248));
    defparam i48563_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 add_2788_10_lut (.I0(GND_net), .I1(n2484), .I2(n1742), .I3(n52096), 
            .O(n8261[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2788_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i51707_4_lut (.I0(n33_adj_4547), .I1(n21_adj_4550), .I2(n19_adj_4549), 
            .I3(n17_adj_4548), .O(n67401));
    defparam i51707_4_lut.LUT_INIT = 16'haaab;
    SB_CARRY add_2788_10 (.CI(n52096), .I0(n2484), .I1(n1742), .CO(n52097));
    SB_LUT4 i52656_4_lut (.I0(n15_adj_4546), .I1(n13_adj_4545), .I2(n2956), 
            .I3(baudrate[2]), .O(n68350));
    defparam i52656_4_lut.LUT_INIT = 16'heffe;
    SB_LUT4 i53266_4_lut (.I0(n21_adj_4550), .I1(n19_adj_4549), .I2(n17_adj_4548), 
            .I3(n68350), .O(n68960));
    defparam i53266_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i53264_4_lut (.I0(n27_adj_4542), .I1(n25_adj_4541), .I2(n23_adj_4540), 
            .I3(n68960), .O(n68958));
    defparam i53264_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i51710_4_lut (.I0(n33_adj_4547), .I1(n31_adj_4544), .I2(n29_adj_4543), 
            .I3(n68958), .O(n67404));
    defparam i51710_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_37_LessThan_1997_i10_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n2957), .I3(GND_net), .O(n10_adj_4551));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i10_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i53808_3_lut (.I0(n10_adj_4551), .I1(baudrate[13]), .I2(n33_adj_4547), 
            .I3(GND_net), .O(n69502));   // verilog/uart_rx.v(119[33:55])
    defparam i53808_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53809_3_lut (.I0(n69502), .I1(baudrate[14]), .I2(n35_adj_4538), 
            .I3(GND_net), .O(n69503));   // verilog/uart_rx.v(119[33:55])
    defparam i53809_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1997_i36_3_lut (.I0(n18), .I1(baudrate[17]), 
            .I2(n41_adj_4537), .I3(GND_net), .O(n36));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i36_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51703_4_lut (.I0(n39_adj_4539), .I1(n37_adj_4536), .I2(n35_adj_4538), 
            .I3(n67401), .O(n67397));
    defparam i51703_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i54143_4_lut (.I0(n36), .I1(n16_adj_4552), .I2(n41_adj_4537), 
            .I3(n67394), .O(n69837));   // verilog/uart_rx.v(119[33:55])
    defparam i54143_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i53697_3_lut (.I0(n69503), .I1(baudrate[15]), .I2(n37_adj_4536), 
            .I3(GND_net), .O(n69391));   // verilog/uart_rx.v(119[33:55])
    defparam i53697_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1997_i22_3_lut (.I0(n14_adj_4553), .I1(baudrate[9]), 
            .I2(n25_adj_4541), .I3(GND_net), .O(n22));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i22_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i54141_4_lut (.I0(n22), .I1(n12_adj_4554), .I2(n25_adj_4541), 
            .I3(n67420), .O(n69835));   // verilog/uart_rx.v(119[33:55])
    defparam i54141_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i54142_3_lut (.I0(n69835), .I1(baudrate[10]), .I2(n27_adj_4542), 
            .I3(GND_net), .O(n69836));   // verilog/uart_rx.v(119[33:55])
    defparam i54142_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i54021_3_lut (.I0(n69836), .I1(baudrate[11]), .I2(n29_adj_4543), 
            .I3(GND_net), .O(n69715));   // verilog/uart_rx.v(119[33:55])
    defparam i54021_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53587_4_lut (.I0(n39_adj_4539), .I1(n37_adj_4536), .I2(n35_adj_4538), 
            .I3(n67404), .O(n69281));
    defparam i53587_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i54274_4_lut (.I0(n69391), .I1(n69837), .I2(n41_adj_4537), 
            .I3(n67397), .O(n69968));   // verilog/uart_rx.v(119[33:55])
    defparam i54274_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i53967_3_lut (.I0(n69715), .I1(baudrate[12]), .I2(n31_adj_4544), 
            .I3(GND_net), .O(n69661));   // verilog/uart_rx.v(119[33:55])
    defparam i53967_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i54298_4_lut (.I0(n69661), .I1(n69968), .I2(n41_adj_4537), 
            .I3(n69281), .O(n69992));   // verilog/uart_rx.v(119[33:55])
    defparam i54298_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i54299_3_lut (.I0(n69992), .I1(baudrate[18]), .I2(n2940), 
            .I3(GND_net), .O(n69993));   // verilog/uart_rx.v(119[33:55])
    defparam i54299_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i54295_3_lut (.I0(n69993), .I1(baudrate[19]), .I2(n2939), 
            .I3(GND_net), .O(n69989));   // verilog/uart_rx.v(119[33:55])
    defparam i54295_3_lut.LUT_INIT = 16'h8e8e;
    SB_DFFESR r_Bit_Index_i1 (.Q(r_Bit_Index[1]), .C(clk16MHz), .E(n27901), 
            .D(n479[1]), .R(n59702));   // verilog/uart_rx.v(50[10] 145[8])
    SB_DFFESR r_Bit_Index_i2 (.Q(r_Bit_Index[2]), .C(clk16MHz), .E(n27901), 
            .D(n479[2]), .R(n59702));   // verilog/uart_rx.v(50[10] 145[8])
    SB_DFFESR r_Clock_Count_1947__i1 (.Q(r_Clock_Count[1]), .C(clk16MHz), 
            .E(n27701), .D(n1[1]), .R(n29076));   // verilog/uart_rx.v(121[34:51])
    SB_DFFESR r_Clock_Count_1947__i2 (.Q(r_Clock_Count[2]), .C(clk16MHz), 
            .E(n27701), .D(n1[2]), .R(n29076));   // verilog/uart_rx.v(121[34:51])
    SB_DFFESR r_Clock_Count_1947__i3 (.Q(r_Clock_Count[3]), .C(clk16MHz), 
            .E(n27701), .D(n1[3]), .R(n29076));   // verilog/uart_rx.v(121[34:51])
    SB_DFFESR r_Clock_Count_1947__i4 (.Q(r_Clock_Count[4]), .C(clk16MHz), 
            .E(n27701), .D(n1[4]), .R(n29076));   // verilog/uart_rx.v(121[34:51])
    SB_DFFESR r_Clock_Count_1947__i5 (.Q(r_Clock_Count[5]), .C(clk16MHz), 
            .E(n27701), .D(n1[5]), .R(n29076));   // verilog/uart_rx.v(121[34:51])
    SB_DFFESR r_Clock_Count_1947__i6 (.Q(r_Clock_Count[6]), .C(clk16MHz), 
            .E(n27701), .D(n1[6]), .R(n29076));   // verilog/uart_rx.v(121[34:51])
    SB_DFFESR r_Clock_Count_1947__i7 (.Q(r_Clock_Count[7]), .C(clk16MHz), 
            .E(n27701), .D(n1[7]), .R(n29076));   // verilog/uart_rx.v(121[34:51])
    SB_LUT4 div_37_i1899_3_lut (.I0(n2713), .I1(n8313[23]), .I2(n294[5]), 
            .I3(GND_net), .O(n2827));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1899_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1900_3_lut (.I0(n2714), .I1(n8313[22]), .I2(n294[5]), 
            .I3(GND_net), .O(n2828));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1900_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1903_3_lut (.I0(n2717), .I1(n8313[19]), .I2(n294[5]), 
            .I3(GND_net), .O(n2831));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1903_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1922_i39_2_lut (.I0(n2831), .I1(baudrate[15]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_4555));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1904_3_lut (.I0(n2718), .I1(n8313[18]), .I2(n294[5]), 
            .I3(GND_net), .O(n2832));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1904_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut_4_lut (.I0(n62551), .I1(n64246), .I2(baudrate[0]), 
            .I3(n48_adj_4556), .O(n962));
    defparam i1_3_lut_4_lut.LUT_INIT = 16'h0010;
    SB_LUT4 div_37_LessThan_1922_i37_2_lut (.I0(n2832), .I1(baudrate[14]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_4557));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1901_3_lut (.I0(n2715), .I1(n8313[21]), .I2(n294[5]), 
            .I3(GND_net), .O(n2829));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1901_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1922_i43_2_lut (.I0(n2829), .I1(baudrate[17]), 
            .I2(GND_net), .I3(GND_net), .O(n43_adj_4558));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1902_3_lut (.I0(n2716), .I1(n8313[20]), .I2(n294[5]), 
            .I3(GND_net), .O(n2830));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1902_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut_4_lut_adj_969 (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(\r_Bit_Index[0] ), .I3(n4_adj_4559), .O(n62513));
    defparam i1_3_lut_4_lut_adj_969.LUT_INIT = 16'hfff7;
    SB_LUT4 div_37_LessThan_1922_i41_2_lut (.I0(n2830), .I1(baudrate[16]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_4560));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1906_3_lut (.I0(n2720), .I1(n8313[16]), .I2(n294[5]), 
            .I3(GND_net), .O(n2834));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1906_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1907_3_lut (.I0(n2721), .I1(n8313[15]), .I2(n294[5]), 
            .I3(GND_net), .O(n2835));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1907_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut_4_lut_adj_970 (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(\r_Bit_Index[0] ), .I3(n4_adj_4559), .O(n62417));
    defparam i1_3_lut_4_lut_adj_970.LUT_INIT = 16'hff7f;
    SB_LUT4 div_37_LessThan_1922_i31_2_lut (.I0(n2835), .I1(baudrate[11]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_4561));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1922_i33_2_lut (.I0(n2834), .I1(baudrate[12]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_4562));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1908_3_lut (.I0(n2722), .I1(n8313[14]), .I2(n294[5]), 
            .I3(GND_net), .O(n2836));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1908_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1910_3_lut (.I0(n2724), .I1(n8313[12]), .I2(n294[5]), 
            .I3(GND_net), .O(n2838));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1910_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut_4_lut_adj_971 (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(\r_Bit_Index[0] ), .I3(n4_adj_4559), .O(n62465));   // verilog/uart_rx.v(98[17:39])
    defparam i1_3_lut_4_lut_adj_971.LUT_INIT = 16'hffbf;
    SB_LUT4 div_37_LessThan_1922_i25_2_lut (.I0(n2838), .I1(baudrate[8]), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_4563));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1922_i27_2_lut (.I0(n2837), .I1(baudrate[9]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_4564));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1922_i29_2_lut (.I0(n2836), .I1(baudrate[10]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_4565));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1914_3_lut (.I0(n2728), .I1(n8313[8]), .I2(n294[5]), 
            .I3(GND_net), .O(n2842));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1914_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1915_3_lut (.I0(n2729), .I1(n8313[7]), .I2(n294[5]), 
            .I3(GND_net), .O(n2843));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1915_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1916_3_lut (.I0(n2730), .I1(n8313[6]), .I2(n294[5]), 
            .I3(GND_net), .O(n2844));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1916_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48564_1_lut (.I0(n64248), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n59794));
    defparam i48564_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i48348_1_lut_2_lut_3_lut_4_lut (.I0(baudrate[16]), .I1(baudrate[17]), 
            .I2(n25574), .I3(baudrate[15]), .O(n59818));
    defparam i48348_1_lut_2_lut_3_lut_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i55121_2_lut_3_lut_4_lut (.I0(baudrate[16]), .I1(baudrate[17]), 
            .I2(n25574), .I3(n48_adj_4566), .O(n294[8]));
    defparam i55121_2_lut_3_lut_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 div_37_LessThan_1922_i15_2_lut (.I0(n2843), .I1(baudrate[3]), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_4567));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_3_lut_4_lut_adj_972 (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(\r_Bit_Index[0] ), .I3(n4_adj_4559), .O(n62401));   // verilog/uart_rx.v(98[17:39])
    defparam i1_3_lut_4_lut_adj_972.LUT_INIT = 16'hfffb;
    SB_LUT4 div_37_LessThan_1922_i17_2_lut (.I0(n2842), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_4568));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1905_3_lut (.I0(n2719), .I1(n8313[17]), .I2(n294[5]), 
            .I3(GND_net), .O(n2833));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1905_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFESR r_Clock_Count_1947__i0 (.Q(r_Clock_Count[0]), .C(clk16MHz), 
            .E(n27701), .D(n1[0]), .R(n29076));   // verilog/uart_rx.v(121[34:51])
    SB_LUT4 div_37_i1912_3_lut (.I0(n2726), .I1(n8313[10]), .I2(n294[5]), 
            .I3(GND_net), .O(n2840));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1912_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1822_3_lut (.I0(n2596), .I1(n8287[23]), .I2(n294[6]), 
            .I3(GND_net), .O(n2713));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1822_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1825_3_lut (.I0(n2599), .I1(n8287[20]), .I2(n294[6]), 
            .I3(GND_net), .O(n2716));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1825_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2788_9_lut (.I0(GND_net), .I1(n2485), .I2(n1602), .I3(n52095), 
            .O(n8261[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2788_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_1845_i41_2_lut (.I0(n2716), .I1(baudrate[15]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_4569));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1823_3_lut (.I0(n2597), .I1(n8287[22]), .I2(n294[6]), 
            .I3(GND_net), .O(n2714));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1823_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1845_i45_2_lut (.I0(n2714), .I1(baudrate[17]), 
            .I2(GND_net), .I3(GND_net), .O(n45_adj_4570));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i45_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1824_3_lut (.I0(n2598), .I1(n8287[21]), .I2(n294[6]), 
            .I3(GND_net), .O(n2715));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1824_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1845_i43_2_lut (.I0(n2715), .I1(baudrate[16]), 
            .I2(GND_net), .I3(GND_net), .O(n43_adj_4571));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1830_3_lut (.I0(n2604), .I1(n8287[15]), .I2(n294[6]), 
            .I3(GND_net), .O(n2721));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1830_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1832_3_lut (.I0(n2606), .I1(n8287[13]), .I2(n294[6]), 
            .I3(GND_net), .O(n2723));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1832_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1831_3_lut (.I0(n2605), .I1(n8287[14]), .I2(n294[6]), 
            .I3(GND_net), .O(n2722));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1831_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1845_i27_2_lut (.I0(n2723), .I1(baudrate[8]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_4572));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1845_i29_2_lut (.I0(n2722), .I1(baudrate[9]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_4573));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1845_i31_2_lut (.I0(n2721), .I1(baudrate[10]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_4574));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i48324_1_lut_2_lut_3_lut (.I0(baudrate[16]), .I1(baudrate[17]), 
            .I2(n25574), .I3(GND_net), .O(n59814));
    defparam i48324_1_lut_2_lut_3_lut.LUT_INIT = 16'h0101;
    SB_LUT4 div_37_i1826_3_lut (.I0(n2600), .I1(n8287[19]), .I2(n294[6]), 
            .I3(GND_net), .O(n2717));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1826_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1845_i39_2_lut (.I0(n2717), .I1(baudrate[14]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_4575));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_973 (.I0(baudrate[7]), .I1(baudrate[8]), .I2(GND_net), 
            .I3(GND_net), .O(n62549));
    defparam i1_2_lut_adj_973.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_974 (.I0(baudrate[15]), .I1(baudrate[16]), .I2(GND_net), 
            .I3(GND_net), .O(n62541));
    defparam i1_2_lut_adj_974.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_975 (.I0(baudrate[11]), .I1(baudrate[12]), .I2(GND_net), 
            .I3(GND_net), .O(n62545));
    defparam i1_2_lut_adj_975.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_976 (.I0(baudrate[9]), .I1(baudrate[10]), .I2(GND_net), 
            .I3(GND_net), .O(n62547));
    defparam i1_2_lut_adj_976.LUT_INIT = 16'heeee;
    SB_LUT4 i48281_2_lut (.I0(baudrate[19]), .I1(baudrate[20]), .I2(GND_net), 
            .I3(GND_net), .O(n63959));
    defparam i48281_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 div_37_i1836_3_lut (.I0(n2610), .I1(n8287[9]), .I2(n294[6]), 
            .I3(GND_net), .O(n2727));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1836_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1837_3_lut (.I0(n2611), .I1(n8287[8]), .I2(n294[6]), 
            .I3(GND_net), .O(n2728));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1837_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_977 (.I0(baudrate[17]), .I1(baudrate[18]), .I2(GND_net), 
            .I3(GND_net), .O(n63961));
    defparam i1_2_lut_adj_977.LUT_INIT = 16'heeee;
    SB_LUT4 i48529_4_lut (.I0(n62547), .I1(n62543), .I2(n62545), .I3(n62541), 
            .O(n64214));
    defparam i48529_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_i1838_3_lut (.I0(n2612), .I1(n8287[7]), .I2(n294[6]), 
            .I3(GND_net), .O(n2729));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1838_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48595_4_lut (.I0(n64248), .I1(n64124), .I2(n59613), .I3(baudrate[4]), 
            .O(n64280));
    defparam i48595_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_LessThan_1845_i17_2_lut (.I0(n2728), .I1(baudrate[3]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_4576));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i54352_4_lut (.I0(n64214), .I1(n63961), .I2(n64280), .I3(n63959), 
            .O(n64284));
    defparam i54352_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 div_37_LessThan_1845_i19_2_lut (.I0(n2727), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_4577));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1828_3_lut (.I0(n2602), .I1(n8287[17]), .I2(n294[6]), 
            .I3(GND_net), .O(n2719));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1828_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1829_3_lut (.I0(n2603), .I1(n8287[16]), .I2(n294[6]), 
            .I3(GND_net), .O(n2720));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1829_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1845_i33_2_lut (.I0(n2720), .I1(baudrate[11]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_4578));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1845_i35_2_lut (.I0(n2719), .I1(baudrate[12]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_4579));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1744_3_lut (.I0(n2477), .I1(n8261[22]), .I2(n294[7]), 
            .I3(GND_net), .O(n2597));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1744_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1827_3_lut (.I0(n2601), .I1(n8287[18]), .I2(n294[6]), 
            .I3(GND_net), .O(n2718));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1827_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1673_3_lut (.I0(n2364), .I1(n8235[12]), .I2(n294[8]), 
            .I3(GND_net), .O(n2487));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1673_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1743_3_lut (.I0(n2476), .I1(n8261[23]), .I2(n294[7]), 
            .I3(GND_net), .O(n2596));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1743_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1748_3_lut (.I0(n2481), .I1(n8261[18]), .I2(n294[7]), 
            .I3(GND_net), .O(n2601));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1748_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1766_i37_2_lut (.I0(n2601), .I1(baudrate[12]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_4580));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1745_3_lut (.I0(n2478), .I1(n8261[21]), .I2(n294[7]), 
            .I3(GND_net), .O(n2598));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1745_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1766_i43_2_lut (.I0(n2598), .I1(baudrate[15]), 
            .I2(GND_net), .I3(GND_net), .O(n43_adj_4581));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1665_3_lut (.I0(n2356), .I1(n8235[20]), .I2(n294[8]), 
            .I3(GND_net), .O(n2479));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1665_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2788_9 (.CI(n52095), .I0(n2485), .I1(n1602), .CO(n52096));
    SB_LUT4 div_37_i1746_3_lut (.I0(n2479), .I1(n8261[20]), .I2(n294[7]), 
            .I3(GND_net), .O(n2599));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1746_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1766_i41_2_lut (.I0(n2599), .I1(baudrate[14]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_4582));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1747_3_lut (.I0(n2480), .I1(n8261[19]), .I2(n294[7]), 
            .I3(GND_net), .O(n2600));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1747_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1766_i39_2_lut (.I0(n2600), .I1(baudrate[13]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_4583));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1749_3_lut (.I0(n2482), .I1(n8261[17]), .I2(n294[7]), 
            .I3(GND_net), .O(n2602));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1749_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1751_3_lut (.I0(n2484), .I1(n8261[15]), .I2(n294[7]), 
            .I3(GND_net), .O(n2604));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1751_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1750_3_lut (.I0(n2483), .I1(n8261[16]), .I2(n294[7]), 
            .I3(GND_net), .O(n2603));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1750_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1766_i31_2_lut (.I0(n2604), .I1(baudrate[9]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_4584));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1766_i33_2_lut (.I0(n2603), .I1(baudrate[10]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_4585));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1766_i35_2_lut (.I0(n2602), .I1(baudrate[11]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_4586));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i35_2_lut.LUT_INIT = 16'h6666;
    SB_DFF r_Rx_Byte_i0 (.Q(rx_data[0]), .C(clk16MHz), .D(n30420));   // verilog/uart_rx.v(50[10] 145[8])
    SB_LUT4 i5572_2_lut_3_lut_4_lut (.I0(baudrate[2]), .I1(n20902), .I2(baudrate[1]), 
            .I3(baudrate[0]), .O(n11253));   // verilog/uart_rx.v(119[33:55])
    defparam i5572_2_lut_3_lut_4_lut.LUT_INIT = 16'h4445;
    SB_DFFE r_Rx_DV_58 (.Q(rx_data_ready), .C(clk16MHz), .E(VCC_net), 
            .D(n54640));   // verilog/uart_rx.v(50[10] 145[8])
    SB_DFFE r_Bit_Index_i0 (.Q(\r_Bit_Index[0] ), .C(clk16MHz), .E(VCC_net), 
            .D(n30416));   // verilog/uart_rx.v(50[10] 145[8])
    SB_LUT4 div_37_i1416_3_lut (.I0(n1975), .I1(n8157[14]), .I2(n294[11]), 
            .I3(GND_net), .O(n2107));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1416_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1503_3_lut (.I0(n2107), .I1(n8183[14]), .I2(n294[10]), 
            .I3(GND_net), .O(n2236));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1503_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2788_8_lut (.I0(GND_net), .I1(n2486), .I2(n1459), .I3(n52094), 
            .O(n8261[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2788_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_i1588_3_lut (.I0(n2236), .I1(n8209[14]), .I2(n294[9]), 
            .I3(GND_net), .O(n2362));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1588_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1671_3_lut (.I0(n2362), .I1(n8235[14]), .I2(n294[8]), 
            .I3(GND_net), .O(n2485));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1671_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1753_3_lut (.I0(n2486), .I1(n8261[13]), .I2(n294[7]), 
            .I3(GND_net), .O(n2606));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1753_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1752_3_lut (.I0(n2485), .I1(n8261[14]), .I2(n294[7]), 
            .I3(GND_net), .O(n2605));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1752_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1766_i27_2_lut (.I0(n2606), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_4587));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1766_i29_2_lut (.I0(n2605), .I1(baudrate[8]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_4588));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1676_3_lut (.I0(n2367), .I1(n8235[9]), .I2(n294[8]), 
            .I3(GND_net), .O(n2490));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1676_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2788_8 (.CI(n52094), .I0(n2486), .I1(n1459), .CO(n52095));
    SB_LUT4 add_2788_7_lut (.I0(GND_net), .I1(n2487), .I2(n1460), .I3(n52093), 
            .O(n8261[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2788_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2788_7 (.CI(n52093), .I0(n2487), .I1(n1460), .CO(n52094));
    SB_LUT4 div_37_i1756_3_lut (.I0(n2489), .I1(n8261[10]), .I2(n294[7]), 
            .I3(GND_net), .O(n2609));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1756_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1757_3_lut (.I0(n2490), .I1(n8261[9]), .I2(n294[7]), 
            .I3(GND_net), .O(n2610));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1757_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1766_i19_2_lut (.I0(n2610), .I1(baudrate[3]), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_4589));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_2788_6_lut (.I0(GND_net), .I1(n2488), .I2(n1011), .I3(n52092), 
            .O(n8261[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2788_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2788_6 (.CI(n52092), .I0(n2488), .I1(n1011), .CO(n52093));
    SB_LUT4 div_37_LessThan_1766_i21_2_lut (.I0(n2609), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_4590));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_978 (.I0(n62045), .I1(n48_adj_4566), .I2(GND_net), 
            .I3(GND_net), .O(n2491));
    defparam i1_2_lut_adj_978.LUT_INIT = 16'h2222;
    SB_LUT4 div_37_i1758_3_lut (.I0(n2491), .I1(n8261[8]), .I2(n294[7]), 
            .I3(GND_net), .O(n2611));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1758_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1664_3_lut (.I0(n2355), .I1(n8235[21]), .I2(n294[8]), 
            .I3(GND_net), .O(n2478));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1664_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1662_3_lut (.I0(n2353), .I1(n8235[23]), .I2(n294[8]), 
            .I3(GND_net), .O(n2476));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1662_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2788_5_lut (.I0(GND_net), .I1(n2489), .I2(n856), .I3(n52091), 
            .O(n8261[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2788_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_3_lut_4_lut_adj_979 (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(\r_Bit_Index[0] ), .I3(n4_adj_4559), .O(n62433));   // verilog/uart_rx.v(98[17:39])
    defparam i1_3_lut_4_lut_adj_979.LUT_INIT = 16'hfffd;
    SB_LUT4 div_37_i1666_3_lut (.I0(n2357), .I1(n8235[19]), .I2(n294[8]), 
            .I3(GND_net), .O(n2480));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1666_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1685_i39_2_lut (.I0(n2480), .I1(baudrate[12]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_4591));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1667_3_lut (.I0(n2358), .I1(n8235[18]), .I2(n294[8]), 
            .I3(GND_net), .O(n2481));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1667_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1685_i37_2_lut (.I0(n2481), .I1(baudrate[11]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_4592));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1668_3_lut (.I0(n2359), .I1(n8235[17]), .I2(n294[8]), 
            .I3(GND_net), .O(n2482));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1668_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1685_i35_2_lut (.I0(n2482), .I1(baudrate[10]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_4593));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i35_2_lut.LUT_INIT = 16'h6666;
    SB_DFF r_Rx_Byte_i7 (.Q(rx_data[7]), .C(clk16MHz), .D(n30126));   // verilog/uart_rx.v(50[10] 145[8])
    SB_LUT4 div_37_LessThan_1430_i37_2_lut (.I0(n2103), .I1(baudrate[8]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_4594));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1430_i37_2_lut.LUT_INIT = 16'h6666;
    SB_DFF r_Rx_Byte_i6 (.Q(rx_data[6]), .C(clk16MHz), .D(n30125));   // verilog/uart_rx.v(50[10] 145[8])
    SB_DFF r_Rx_Byte_i5 (.Q(rx_data[5]), .C(clk16MHz), .D(n30124));   // verilog/uart_rx.v(50[10] 145[8])
    SB_LUT4 div_37_LessThan_1430_i41_2_lut (.I0(n2101), .I1(baudrate[10]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_4595));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1430_i41_2_lut.LUT_INIT = 16'h6666;
    SB_DFF r_Rx_Byte_i4 (.Q(rx_data[4]), .C(clk16MHz), .D(n30123));   // verilog/uart_rx.v(50[10] 145[8])
    SB_LUT4 div_37_LessThan_1430_i27_2_lut (.I0(n2108), .I1(baudrate[3]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_4596));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1430_i27_2_lut.LUT_INIT = 16'h6666;
    SB_DFF r_Rx_Byte_i3 (.Q(rx_data[3]), .C(clk16MHz), .D(n30122));   // verilog/uart_rx.v(50[10] 145[8])
    SB_DFF r_Rx_Byte_i2 (.Q(rx_data[2]), .C(clk16MHz), .D(n30121));   // verilog/uart_rx.v(50[10] 145[8])
    SB_DFF r_Rx_Byte_i1 (.Q(rx_data[1]), .C(clk16MHz), .D(n30120));   // verilog/uart_rx.v(50[10] 145[8])
    SB_DFF r_SM_Main_i2 (.Q(\r_SM_Main[2] ), .C(clk16MHz), .D(n71282));   // verilog/uart_rx.v(50[10] 145[8])
    SB_LUT4 i52015_4_lut (.I0(n33_adj_4509), .I1(n31_adj_4507), .I2(n29_adj_4508), 
            .I3(n27_adj_4596), .O(n67709));
    defparam i52015_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_37_LessThan_1430_i38_3_lut (.I0(n30_adj_4597), .I1(baudrate[10]), 
            .I2(n41_adj_4595), .I3(GND_net), .O(n38_adj_4598));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1430_i38_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29200_rep_4_2_lut (.I0(n8157[11]), .I1(n294[11]), .I2(GND_net), 
            .I3(GND_net), .O(n59821));   // verilog/uart_rx.v(119[33:55])
    defparam i29200_rep_4_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 div_37_LessThan_1430_i26_4_lut (.I0(n59821), .I1(baudrate[2]), 
            .I2(n2109), .I3(baudrate[1]), .O(n26));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1430_i26_4_lut.LUT_INIT = 16'h4d0c;
    SB_CARRY add_2788_5 (.CI(n52091), .I0(n2489), .I1(n856), .CO(n52092));
    SB_LUT4 i53573_3_lut (.I0(n26), .I1(baudrate[6]), .I2(n33_adj_4509), 
            .I3(GND_net), .O(n69267));   // verilog/uart_rx.v(119[33:55])
    defparam i53573_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53574_3_lut (.I0(n69267), .I1(baudrate[7]), .I2(n35_adj_4510), 
            .I3(GND_net), .O(n69268));   // verilog/uart_rx.v(119[33:55])
    defparam i53574_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52009_4_lut (.I0(n39_adj_4511), .I1(n37_adj_4594), .I2(n35_adj_4510), 
            .I3(n67709), .O(n67703));
    defparam i52009_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i54054_4_lut (.I0(n38_adj_4598), .I1(n28), .I2(n41_adj_4595), 
            .I3(n67701), .O(n69748));   // verilog/uart_rx.v(119[33:55])
    defparam i54054_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i52789_3_lut (.I0(n69268), .I1(baudrate[8]), .I2(n37_adj_4594), 
            .I3(GND_net), .O(n68483));   // verilog/uart_rx.v(119[33:55])
    defparam i52789_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i54240_4_lut (.I0(n68483), .I1(n69748), .I2(n41_adj_4595), 
            .I3(n67703), .O(n69934));   // verilog/uart_rx.v(119[33:55])
    defparam i54240_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i54241_3_lut (.I0(n69934), .I1(baudrate[11]), .I2(n2100), 
            .I3(GND_net), .O(n69935));   // verilog/uart_rx.v(119[33:55])
    defparam i54241_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i54172_3_lut (.I0(n69935), .I1(baudrate[12]), .I2(n2099), 
            .I3(GND_net), .O(n69866));   // verilog/uart_rx.v(119[33:55])
    defparam i54172_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i52795_3_lut (.I0(n69866), .I1(baudrate[13]), .I2(n2098), 
            .I3(GND_net), .O(n48_adj_4599));   // verilog/uart_rx.v(119[33:55])
    defparam i52795_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 add_2788_4_lut (.I0(GND_net), .I1(n2490), .I2(n698), .I3(n52090), 
            .O(n8261[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2788_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_980 (.I0(baudrate[27]), .I1(baudrate[24]), .I2(baudrate[29]), 
            .I3(baudrate[30]), .O(n63515));
    defparam i1_4_lut_adj_980.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_3_lut (.I0(n63465), .I1(n63513), .I2(n62569), .I3(GND_net), 
            .O(n63523));
    defparam i1_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_4_lut_adj_981 (.I0(n63523), .I1(n63519), .I2(n63521), .I3(n63515), 
            .O(n25562));
    defparam i1_4_lut_adj_981.LUT_INIT = 16'hfffe;
    SB_CARRY add_2788_4 (.CI(n52090), .I0(n2490), .I1(n698), .CO(n52091));
    SB_LUT4 i1_3_lut_adj_982 (.I0(n25562), .I1(n48_adj_4599), .I2(baudrate[0]), 
            .I3(GND_net), .O(n2240));
    defparam i1_3_lut_adj_982.LUT_INIT = 16'hefef;
    SB_LUT4 div_37_i1592_3_lut (.I0(n2240), .I1(n8209[10]), .I2(n294[9]), 
            .I3(GND_net), .O(n2366));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1592_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1675_3_lut (.I0(n2366), .I1(n8235[10]), .I2(n294[8]), 
            .I3(GND_net), .O(n2489));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1675_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1685_i21_2_lut (.I0(n2489), .I1(baudrate[3]), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_4600));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1669_3_lut (.I0(n2360), .I1(n8235[16]), .I2(n294[8]), 
            .I3(GND_net), .O(n2483));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1669_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1685_i33_2_lut (.I0(n2483), .I1(baudrate[9]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_4601));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1663_3_lut (.I0(n2354), .I1(n8235[22]), .I2(n294[8]), 
            .I3(GND_net), .O(n2477));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1663_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1685_i45_2_lut (.I0(n2477), .I1(baudrate[15]), 
            .I2(GND_net), .I3(GND_net), .O(n45_adj_4602));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i45_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_2788_3_lut (.I0(GND_net), .I1(n2491), .I2(n858), .I3(n52089), 
            .O(n8261[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2788_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_3_lut_4_lut_adj_983 (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(\r_Bit_Index[0] ), .I3(n4_adj_4559), .O(n62481));   // verilog/uart_rx.v(98[17:39])
    defparam i1_3_lut_4_lut_adj_983.LUT_INIT = 16'hffdf;
    SB_LUT4 div_37_LessThan_1685_i23_2_lut (.I0(n2488), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_4603));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1670_3_lut (.I0(n2361), .I1(n8235[15]), .I2(n294[8]), 
            .I3(GND_net), .O(n2484));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1670_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2788_3 (.CI(n52089), .I0(n2491), .I1(n858), .CO(n52090));
    SB_LUT4 i48536_1_lut_2_lut (.I0(baudrate[12]), .I1(n64194), .I2(GND_net), 
            .I3(GND_net), .O(n59827));
    defparam i48536_1_lut_2_lut.LUT_INIT = 16'h1111;
    SB_LUT4 div_37_LessThan_1685_i31_2_lut (.I0(n2484), .I1(baudrate[8]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_4604));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1417_3_lut (.I0(n1976), .I1(n8157[13]), .I2(n294[11]), 
            .I3(GND_net), .O(n2108));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1417_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1504_3_lut (.I0(n2108), .I1(n8183[13]), .I2(n294[10]), 
            .I3(GND_net), .O(n2237));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1504_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1589_3_lut (.I0(n2237), .I1(n8209[13]), .I2(n294[9]), 
            .I3(GND_net), .O(n2363));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1589_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1672_3_lut (.I0(n2363), .I1(n8235[13]), .I2(n294[8]), 
            .I3(GND_net), .O(n2486));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1672_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1685_i27_2_lut (.I0(n2486), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_4605));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1685_i29_2_lut (.I0(n2485), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_4606));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_2788_2_lut (.I0(n59810), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n62047)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2788_2_lut.LUT_INIT = 16'h8228;
    SB_LUT4 div_37_LessThan_1685_i41_2_lut (.I0(n2479), .I1(baudrate[13]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_4607));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1685_i43_2_lut (.I0(n2478), .I1(baudrate[14]), 
            .I2(GND_net), .I3(GND_net), .O(n43_adj_4608));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1685_i19_2_lut (.I0(n2490), .I1(baudrate[2]), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_4609));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i51921_4_lut (.I0(n25_adj_4512), .I1(n23_adj_4603), .I2(n21_adj_4600), 
            .I3(n19_adj_4609), .O(n67615));
    defparam i51921_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i51906_4_lut (.I0(n31_adj_4604), .I1(n29_adj_4606), .I2(n27_adj_4605), 
            .I3(n67615), .O(n67600));
    defparam i51906_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i53734_4_lut (.I0(n37_adj_4592), .I1(n35_adj_4593), .I2(n33_adj_4601), 
            .I3(n67600), .O(n69428));
    defparam i53734_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i53955_3_lut (.I0(n18_adj_4610), .I1(baudrate[13]), .I2(n41_adj_4607), 
            .I3(GND_net), .O(n69649));   // verilog/uart_rx.v(119[33:55])
    defparam i53955_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53956_3_lut (.I0(n69649), .I1(baudrate[14]), .I2(n43_adj_4608), 
            .I3(GND_net), .O(n69650));   // verilog/uart_rx.v(119[33:55])
    defparam i53956_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52810_4_lut (.I0(n43_adj_4608), .I1(n41_adj_4607), .I2(n29_adj_4606), 
            .I3(n67613), .O(n68504));
    defparam i52810_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 div_37_LessThan_1685_i26_3_lut (.I0(n24_adj_4611), .I1(baudrate[7]), 
            .I2(n29_adj_4606), .I3(GND_net), .O(n26_adj_4612));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i26_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2788_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n52089));
    SB_LUT4 i53674_3_lut (.I0(n69650), .I1(baudrate[15]), .I2(n45_adj_4602), 
            .I3(GND_net), .O(n42_adj_4613));   // verilog/uart_rx.v(119[33:55])
    defparam i53674_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i55112_2_lut_3_lut (.I0(baudrate[12]), .I1(n64194), .I2(n48_adj_4614), 
            .I3(GND_net), .O(n294[12]));
    defparam i55112_2_lut_3_lut.LUT_INIT = 16'h0101;
    SB_LUT4 div_37_LessThan_1685_i30_3_lut (.I0(n22_adj_4615), .I1(baudrate[9]), 
            .I2(n33_adj_4601), .I3(GND_net), .O(n30_adj_4616));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i54064_4_lut (.I0(n30_adj_4616), .I1(n20_adj_4617), .I2(n33_adj_4601), 
            .I3(n67598), .O(n69758));   // verilog/uart_rx.v(119[33:55])
    defparam i54064_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i54065_3_lut (.I0(n69758), .I1(baudrate[10]), .I2(n35_adj_4593), 
            .I3(GND_net), .O(n69759));   // verilog/uart_rx.v(119[33:55])
    defparam i54065_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53874_3_lut (.I0(n69759), .I1(baudrate[11]), .I2(n37_adj_4592), 
            .I3(GND_net), .O(n69568));   // verilog/uart_rx.v(119[33:55])
    defparam i53874_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52812_4_lut (.I0(n43_adj_4608), .I1(n41_adj_4607), .I2(n39_adj_4591), 
            .I3(n69428), .O(n68506));
    defparam i52812_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i53334_4_lut (.I0(n42_adj_4613), .I1(n26_adj_4612), .I2(n45_adj_4602), 
            .I3(n68504), .O(n69028));   // verilog/uart_rx.v(119[33:55])
    defparam i53334_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i52809_3_lut (.I0(n69568), .I1(baudrate[12]), .I2(n39_adj_4591), 
            .I3(GND_net), .O(n68503));   // verilog/uart_rx.v(119[33:55])
    defparam i52809_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53336_4_lut (.I0(n68503), .I1(n69028), .I2(n45_adj_4602), 
            .I3(n68506), .O(n69030));   // verilog/uart_rx.v(119[33:55])
    defparam i53336_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 add_2787_17_lut (.I0(GND_net), .I1(n2353), .I2(n2638), .I3(n52088), 
            .O(n8235[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2787_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2787_16_lut (.I0(GND_net), .I1(n2354), .I2(n2519), .I3(n52087), 
            .O(n8235[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2787_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_i1579_3_lut (.I0(n2227), .I1(n8209[23]), .I2(n294[9]), 
            .I3(GND_net), .O(n2353));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1579_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_984 (.I0(baudrate[27]), .I1(baudrate[28]), .I2(GND_net), 
            .I3(GND_net), .O(n63461));
    defparam i1_2_lut_adj_984.LUT_INIT = 16'heeee;
    SB_LUT4 div_37_LessThan_1157_i43_2_lut (.I0(n1695), .I1(baudrate[8]), 
            .I2(GND_net), .I3(GND_net), .O(n43_adj_4618));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1157_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1157_i37_2_lut (.I0(n1698), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_4619));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1157_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1157_i41_2_lut (.I0(n1696), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_4620));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1157_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1157_i39_2_lut (.I0(n1697), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_4621));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1157_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i29197_rep_5_2_lut (.I0(n8079[14]), .I1(n294[14]), .I2(GND_net), 
            .I3(GND_net), .O(n59830));   // verilog/uart_rx.v(119[33:55])
    defparam i29197_rep_5_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 div_37_LessThan_1157_i32_4_lut (.I0(n59830), .I1(baudrate[2]), 
            .I2(n1701), .I3(baudrate[1]), .O(n32_adj_4622));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1157_i32_4_lut.LUT_INIT = 16'h4d0c;
    SB_DFFSR r_SM_Main_i1 (.Q(\r_SM_Main[1] ), .C(clk16MHz), .D(n3_adj_4535), 
            .R(\r_SM_Main[2] ));   // verilog/uart_rx.v(50[10] 145[8])
    SB_LUT4 i53585_3_lut (.I0(n32_adj_4622), .I1(baudrate[6]), .I2(n39_adj_4621), 
            .I3(GND_net), .O(n69279));   // verilog/uart_rx.v(119[33:55])
    defparam i53585_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53586_3_lut (.I0(n69279), .I1(baudrate[7]), .I2(n41_adj_4620), 
            .I3(GND_net), .O(n69280));   // verilog/uart_rx.v(119[33:55])
    defparam i53586_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52948_4_lut (.I0(n41_adj_4620), .I1(n39_adj_4621), .I2(n37_adj_4619), 
            .I3(n67757), .O(n68642));
    defparam i52948_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i53655_3_lut (.I0(n34_adj_4623), .I1(baudrate[5]), .I2(n37_adj_4619), 
            .I3(GND_net), .O(n69349));   // verilog/uart_rx.v(119[33:55])
    defparam i53655_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52772_3_lut (.I0(n69280), .I1(baudrate[8]), .I2(n43_adj_4618), 
            .I3(GND_net), .O(n68466));   // verilog/uart_rx.v(119[33:55])
    defparam i52772_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53905_4_lut (.I0(n68466), .I1(n69349), .I2(n43_adj_4618), 
            .I3(n68642), .O(n69599));   // verilog/uart_rx.v(119[33:55])
    defparam i53905_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i53906_3_lut (.I0(n69599), .I1(baudrate[9]), .I2(n1694), .I3(GND_net), 
            .O(n69600));   // verilog/uart_rx.v(119[33:55])
    defparam i53906_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_i2083_1_lut (.I0(baudrate[21]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n3082));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2083_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_LessThan_1157_i48_3_lut (.I0(n69600), .I1(baudrate[10]), 
            .I2(n1693), .I3(GND_net), .O(n48_adj_4624));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1157_i48_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i1_4_lut_adj_985 (.I0(n63505), .I1(n63461), .I2(n63463), .I3(baudrate[11]), 
            .O(n63491));
    defparam i1_4_lut_adj_985.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_986 (.I0(n63491), .I1(n63493), .I2(n63481), .I3(n63369), 
            .O(n25553));
    defparam i1_4_lut_adj_986.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_3_lut_adj_987 (.I0(n25553), .I1(n48_adj_4624), .I2(baudrate[0]), 
            .I3(GND_net), .O(n1841));
    defparam i1_3_lut_adj_987.LUT_INIT = 16'hefef;
    SB_CARRY add_2787_16 (.CI(n52087), .I0(n2354), .I1(n2519), .CO(n52088));
    SB_LUT4 div_37_LessThan_1341_i37_2_lut (.I0(n1971), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_4625));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1341_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1341_i35_2_lut (.I0(n1972), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_4626));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1341_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1341_i39_2_lut (.I0(n1970), .I1(baudrate[8]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_4627));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1341_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1341_i31_2_lut (.I0(n1974), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_4628));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1341_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1341_i33_2_lut (.I0(n1973), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_4629));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1341_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1062_i43_2_lut (.I0(n1554), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n43_adj_4630));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1062_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1062_i32_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n1560), .I3(GND_net), .O(n32_adj_4631));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1062_i32_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i53589_3_lut (.I0(n32_adj_4631), .I1(baudrate[5]), .I2(n39_adj_4513), 
            .I3(GND_net), .O(n69283));   // verilog/uart_rx.v(119[33:55])
    defparam i53589_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53590_3_lut (.I0(n69283), .I1(baudrate[6]), .I2(n41_adj_4514), 
            .I3(GND_net), .O(n69284));   // verilog/uart_rx.v(119[33:55])
    defparam i53590_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2153_1_lut (.I0(baudrate[22]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n3186));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2153_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_2787_15_lut (.I0(GND_net), .I1(n2355), .I2(n2397), .I3(n52086), 
            .O(n8235[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2787_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i52956_4_lut (.I0(n41_adj_4514), .I1(n39_adj_4513), .I2(n37_adj_4515), 
            .I3(n67767), .O(n68650));
    defparam i52956_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i53653_3_lut (.I0(n34_adj_4632), .I1(baudrate[4]), .I2(n37_adj_4515), 
            .I3(GND_net), .O(n69347));   // verilog/uart_rx.v(119[33:55])
    defparam i53653_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52765_3_lut (.I0(n69284), .I1(baudrate[7]), .I2(n43_adj_4630), 
            .I3(GND_net), .O(n68459));   // verilog/uart_rx.v(119[33:55])
    defparam i52765_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53909_4_lut (.I0(n68459), .I1(n69347), .I2(n43_adj_4630), 
            .I3(n68650), .O(n69603));   // verilog/uart_rx.v(119[33:55])
    defparam i53909_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i53910_3_lut (.I0(n69603), .I1(baudrate[8]), .I2(n1553), .I3(GND_net), 
            .O(n69604));   // verilog/uart_rx.v(119[33:55])
    defparam i53910_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_1062_i48_3_lut (.I0(n69604), .I1(baudrate[9]), 
            .I2(n1552), .I3(GND_net), .O(n48_adj_4633));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1062_i48_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i1_3_lut_adj_988 (.I0(n64228), .I1(n48_adj_4633), .I2(n8079[14]), 
            .I3(GND_net), .O(n1702));
    defparam i1_3_lut_adj_988.LUT_INIT = 16'h1010;
    SB_LUT4 div_37_i1236_3_lut (.I0(n1702), .I1(n8105[14]), .I2(n294[13]), 
            .I3(GND_net), .O(n1840));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1236_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1327_3_lut (.I0(n1840), .I1(n8131[14]), .I2(n294[12]), 
            .I3(GND_net), .O(n1975));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1327_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1341_i29_2_lut (.I0(n1975), .I1(baudrate[3]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_4634));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1341_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1341_i41_2_lut (.I0(n1969), .I1(baudrate[9]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_4635));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1341_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1328_3_lut (.I0(n1841), .I1(n8131[13]), .I2(n294[12]), 
            .I3(GND_net), .O(n1976));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1328_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1341_i27_2_lut (.I0(n1976), .I1(baudrate[2]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_4636));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1341_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i2163_1_lut (.I0(baudrate[12]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2272));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2163_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i52035_4_lut (.I0(n33_adj_4629), .I1(n31_adj_4628), .I2(n29_adj_4634), 
            .I3(n27_adj_4636), .O(n67729));
    defparam i52035_4_lut.LUT_INIT = 16'haaab;
    SB_CARRY add_2787_15 (.CI(n52086), .I0(n2355), .I1(n2397), .CO(n52087));
    SB_LUT4 div_37_LessThan_1341_i38_3_lut (.I0(n30_adj_4637), .I1(baudrate[9]), 
            .I2(n41_adj_4635), .I3(GND_net), .O(n38_adj_4638));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1341_i38_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53581_3_lut (.I0(n26_adj_4639), .I1(baudrate[5]), .I2(n33_adj_4629), 
            .I3(GND_net), .O(n69275));   // verilog/uart_rx.v(119[33:55])
    defparam i53581_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53582_3_lut (.I0(n69275), .I1(baudrate[6]), .I2(n35_adj_4626), 
            .I3(GND_net), .O(n69276));   // verilog/uart_rx.v(119[33:55])
    defparam i53582_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2162_1_lut (.I0(baudrate[13]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2397));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2162_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i52029_4_lut (.I0(n39_adj_4627), .I1(n37_adj_4625), .I2(n35_adj_4626), 
            .I3(n67729), .O(n67723));
    defparam i52029_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_37_i2161_1_lut (.I0(baudrate[14]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2519));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2161_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i54052_4_lut (.I0(n38_adj_4638), .I1(n28_adj_4640), .I2(n41_adj_4635), 
            .I3(n67719), .O(n69746));   // verilog/uart_rx.v(119[33:55])
    defparam i54052_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i52781_3_lut (.I0(n69276), .I1(baudrate[7]), .I2(n37_adj_4625), 
            .I3(GND_net), .O(n68475));   // verilog/uart_rx.v(119[33:55])
    defparam i52781_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i54236_4_lut (.I0(n68475), .I1(n69746), .I2(n41_adj_4635), 
            .I3(n67723), .O(n69930));   // verilog/uart_rx.v(119[33:55])
    defparam i54236_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i54237_3_lut (.I0(n69930), .I1(baudrate[10]), .I2(n1968), 
            .I3(GND_net), .O(n69931));   // verilog/uart_rx.v(119[33:55])
    defparam i54237_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i54176_3_lut (.I0(n69931), .I1(baudrate[11]), .I2(n1967), 
            .I3(GND_net), .O(n69870));   // verilog/uart_rx.v(119[33:55])
    defparam i54176_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i52787_3_lut (.I0(n69870), .I1(baudrate[12]), .I2(n1966), 
            .I3(GND_net), .O(n48_adj_4641));   // verilog/uart_rx.v(119[33:55])
    defparam i52787_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i1_3_lut_adj_989 (.I0(n64194), .I1(n48_adj_4641), .I2(n8157[11]), 
            .I3(GND_net), .O(n2110));
    defparam i1_3_lut_adj_989.LUT_INIT = 16'h1010;
    SB_LUT4 div_37_i1506_3_lut (.I0(n2110), .I1(n8183[11]), .I2(n294[10]), 
            .I3(GND_net), .O(n2239));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1506_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_965_i45_2_lut (.I0(n1409), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n45_adj_4642));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_965_i45_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_965_i39_2_lut (.I0(n1412), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_4643));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_965_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_965_i43_2_lut (.I0(n1410), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n43_adj_4644));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_965_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_965_i41_2_lut (.I0(n1411), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_4645));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_965_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_2787_14_lut (.I0(GND_net), .I1(n2356), .I2(n2272), .I3(n52085), 
            .O(n8235[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2787_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i53591_3_lut (.I0(n34_adj_4646), .I1(baudrate[5]), .I2(n41_adj_4645), 
            .I3(GND_net), .O(n69285));   // verilog/uart_rx.v(119[33:55])
    defparam i53591_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53592_3_lut (.I0(n69285), .I1(baudrate[6]), .I2(n43_adj_4644), 
            .I3(GND_net), .O(n69286));   // verilog/uart_rx.v(119[33:55])
    defparam i53592_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52962_4_lut (.I0(n43_adj_4644), .I1(n41_adj_4645), .I2(n39_adj_4643), 
            .I3(n67776), .O(n68656));
    defparam i52962_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 div_37_LessThan_965_i38_3_lut (.I0(n36_adj_4647), .I1(baudrate[4]), 
            .I2(n39_adj_4643), .I3(GND_net), .O(n38_adj_4648));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_965_i38_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52761_3_lut (.I0(n69286), .I1(baudrate[7]), .I2(n45_adj_4642), 
            .I3(GND_net), .O(n68455));   // verilog/uart_rx.v(119[33:55])
    defparam i52761_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53651_4_lut (.I0(n68455), .I1(n38_adj_4648), .I2(n45_adj_4642), 
            .I3(n68656), .O(n69345));   // verilog/uart_rx.v(119[33:55])
    defparam i53651_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 div_37_i1142_3_lut (.I0(n1560), .I1(n8079[15]), .I2(n294[14]), 
            .I3(GND_net), .O(n1701));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1142_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1235_3_lut (.I0(n1701), .I1(n8105[15]), .I2(n294[13]), 
            .I3(GND_net), .O(n1839));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1235_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1326_3_lut (.I0(n1839), .I1(n8131[15]), .I2(n294[12]), 
            .I3(GND_net), .O(n1974));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1326_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1415_3_lut (.I0(n1974), .I1(n8157[15]), .I2(n294[11]), 
            .I3(GND_net), .O(n2106));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1415_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1502_3_lut (.I0(n2106), .I1(n8183[15]), .I2(n294[10]), 
            .I3(GND_net), .O(n2235));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1502_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1587_3_lut (.I0(n2235), .I1(n8209[15]), .I2(n294[9]), 
            .I3(GND_net), .O(n2361));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1587_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1580_3_lut (.I0(n2228), .I1(n8209[22]), .I2(n294[9]), 
            .I3(GND_net), .O(n2354));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1580_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1320_3_lut (.I0(n1833), .I1(n8131[21]), .I2(n294[12]), 
            .I3(GND_net), .O(n1968));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1320_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1409_3_lut (.I0(n1968), .I1(n8157[21]), .I2(n294[11]), 
            .I3(GND_net), .O(n2100));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1409_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1496_3_lut (.I0(n2100), .I1(n8183[21]), .I2(n294[10]), 
            .I3(GND_net), .O(n2229));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1496_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1581_3_lut (.I0(n2229), .I1(n8209[21]), .I2(n294[9]), 
            .I3(GND_net), .O(n2355));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1581_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5730_2_lut (.I0(n962), .I1(baudrate[1]), .I2(GND_net), .I3(GND_net), 
            .O(n40_adj_4649));   // verilog/uart_rx.v(119[33:55])
    defparam i5730_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 div_37_i745_4_lut (.I0(n961), .I1(n40_adj_4649), .I2(n294[18]), 
            .I3(baudrate[2]), .O(n1114));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i745_4_lut.LUT_INIT = 16'h6a9a;
    SB_LUT4 div_37_i846_3_lut (.I0(n1114), .I1(n8001[20]), .I2(n294[17]), 
            .I3(GND_net), .O(n1264));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i846_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i945_3_lut (.I0(n1264), .I1(n8027[20]), .I2(n294[16]), 
            .I3(GND_net), .O(n1411));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i945_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1042_3_lut (.I0(n1411), .I1(n8053[20]), .I2(n294[15]), 
            .I3(GND_net), .O(n1555));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1042_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1137_3_lut (.I0(n1555), .I1(n8079[20]), .I2(n294[14]), 
            .I3(GND_net), .O(n1696));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1137_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1230_3_lut (.I0(n1696), .I1(n8105[20]), .I2(n294[13]), 
            .I3(GND_net), .O(n1834));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1230_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1321_3_lut (.I0(n1834), .I1(n8131[20]), .I2(n294[12]), 
            .I3(GND_net), .O(n1969));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1321_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1410_3_lut (.I0(n1969), .I1(n8157[20]), .I2(n294[11]), 
            .I3(GND_net), .O(n2101));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1410_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1497_3_lut (.I0(n2101), .I1(n8183[20]), .I2(n294[10]), 
            .I3(GND_net), .O(n2230));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1497_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1582_3_lut (.I0(n2230), .I1(n8209[20]), .I2(n294[9]), 
            .I3(GND_net), .O(n2356));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1582_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1602_i41_2_lut (.I0(n2356), .I1(baudrate[12]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_4650));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_990 (.I0(baudrate[25]), .I1(baudrate[29]), .I2(GND_net), 
            .I3(GND_net), .O(n63611));
    defparam i1_2_lut_adj_990.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_991 (.I0(baudrate[24]), .I1(baudrate[31]), .I2(GND_net), 
            .I3(GND_net), .O(n63613));
    defparam i1_2_lut_adj_991.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_992 (.I0(n63513), .I1(n63509), .I2(n63511), .I3(n63507), 
            .O(n63493));
    defparam i1_4_lut_adj_992.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_993 (.I0(n63611), .I1(n63401), .I2(n63505), .I3(n63391), 
            .O(n25586));
    defparam i1_4_lut_adj_993.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_i642_4_lut (.I0(n805), .I1(baudrate[1]), .I2(n294[19]), 
            .I3(baudrate[0]), .O(n961));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i642_4_lut.LUT_INIT = 16'h9a6a;
    SB_LUT4 i29182_rep_6_2_lut (.I0(baudrate[0]), .I1(n294[19]), .I2(GND_net), 
            .I3(GND_net), .O(n59847));   // verilog/uart_rx.v(119[33:55])
    defparam i29182_rep_6_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 div_37_LessThan_662_i42_4_lut (.I0(n59847), .I1(baudrate[2]), 
            .I2(n961), .I3(baudrate[1]), .O(n42_adj_4651));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_662_i42_4_lut.LUT_INIT = 16'h4d0c;
    SB_LUT4 i53599_3_lut (.I0(n42_adj_4651), .I1(baudrate[3]), .I2(n960), 
            .I3(GND_net), .O(n69293));   // verilog/uart_rx.v(119[33:55])
    defparam i53599_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i53600_3_lut (.I0(n69293), .I1(baudrate[4]), .I2(n959), .I3(GND_net), 
            .O(n69294));   // verilog/uart_rx.v(119[33:55])
    defparam i53600_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_662_i48_3_lut (.I0(n69294), .I1(baudrate[5]), 
            .I2(n59530), .I3(GND_net), .O(n48_adj_4652));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_662_i48_3_lut.LUT_INIT = 16'he8e8;
    SB_LUT4 i1_4_lut_adj_994 (.I0(n63383), .I1(n25586), .I2(n63493), .I3(n63381), 
            .O(n25605));
    defparam i1_4_lut_adj_994.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_3_lut_adj_995 (.I0(n25605), .I1(n48_adj_4652), .I2(baudrate[0]), 
            .I3(GND_net), .O(n1116));
    defparam i1_3_lut_adj_995.LUT_INIT = 16'hefef;
    SB_LUT4 div_37_i848_3_lut (.I0(n1116), .I1(n8001[18]), .I2(n294[17]), 
            .I3(GND_net), .O(n1266));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i848_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i947_3_lut (.I0(n1266), .I1(n8027[18]), .I2(n294[16]), 
            .I3(GND_net), .O(n1413));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i947_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1044_3_lut (.I0(n1413), .I1(n8053[18]), .I2(n294[15]), 
            .I3(GND_net), .O(n1557));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1044_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1139_3_lut (.I0(n1557), .I1(n8079[18]), .I2(n294[14]), 
            .I3(GND_net), .O(n1698));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1139_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1232_3_lut (.I0(n1698), .I1(n8105[18]), .I2(n294[13]), 
            .I3(GND_net), .O(n1836));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1232_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1323_3_lut (.I0(n1836), .I1(n8131[18]), .I2(n294[12]), 
            .I3(GND_net), .O(n1971));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1323_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1412_3_lut (.I0(n1971), .I1(n8157[18]), .I2(n294[11]), 
            .I3(GND_net), .O(n2103));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1412_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1499_3_lut (.I0(n2103), .I1(n8183[18]), .I2(n294[10]), 
            .I3(GND_net), .O(n2232));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1499_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1584_3_lut (.I0(n2232), .I1(n8209[18]), .I2(n294[9]), 
            .I3(GND_net), .O(n2358));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1584_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1602_i37_2_lut (.I0(n2358), .I1(baudrate[10]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_4653));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_996 (.I0(baudrate[16]), .I1(baudrate[17]), .I2(GND_net), 
            .I3(GND_net), .O(n63511));
    defparam i1_2_lut_adj_996.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_997 (.I0(baudrate[6]), .I1(baudrate[7]), .I2(GND_net), 
            .I3(GND_net), .O(n63375));
    defparam i1_2_lut_adj_997.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_998 (.I0(baudrate[8]), .I1(baudrate[9]), .I2(GND_net), 
            .I3(GND_net), .O(n63373));
    defparam i1_2_lut_adj_998.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_999 (.I0(baudrate[4]), .I1(baudrate[5]), .I2(GND_net), 
            .I3(GND_net), .O(n62683));
    defparam i1_2_lut_adj_999.LUT_INIT = 16'heeee;
    SB_LUT4 i29175_2_lut (.I0(baudrate[1]), .I1(baudrate[0]), .I2(GND_net), 
            .I3(GND_net), .O(n43068));
    defparam i29175_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 div_37_LessThan_450_i46_4_lut (.I0(n67096), .I1(baudrate[2]), 
            .I2(n70030), .I3(n48_adj_4654), .O(n46));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_450_i46_4_lut.LUT_INIT = 16'hc0e8;
    SB_LUT4 div_37_LessThan_450_i48_3_lut (.I0(n46), .I1(baudrate[3]), .I2(n59526), 
            .I3(GND_net), .O(n48_adj_4655));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_450_i48_3_lut.LUT_INIT = 16'he8e8;
    SB_LUT4 i1_4_lut_adj_1000 (.I0(n62683), .I1(n63373), .I2(n63375), 
            .I3(n63371), .O(n62695));
    defparam i1_4_lut_adj_1000.LUT_INIT = 16'hfffe;
    SB_CARRY add_2787_14 (.CI(n52085), .I0(n2356), .I1(n2272), .CO(n52086));
    SB_LUT4 add_2787_13_lut (.I0(GND_net), .I1(n2357), .I2(n2144), .I3(n52084), 
            .O(n8235[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2787_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1001 (.I0(n62695), .I1(n25580), .I2(n62687), 
            .I3(n63521), .O(n25608));
    defparam i1_4_lut_adj_1001.LUT_INIT = 16'hfffe;
    SB_CARRY add_2787_13 (.CI(n52084), .I0(n2357), .I1(n2144), .CO(n52085));
    SB_LUT4 add_2787_12_lut (.I0(GND_net), .I1(n2358), .I2(n2013), .I3(n52083), 
            .O(n8235[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2787_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i5_3_lut (.I0(r_SM_Main[0]), .I1(\o_Rx_DV_N_3488[24] ), .I2(n27), 
            .I3(GND_net), .O(n14_adj_4656));
    defparam i5_3_lut.LUT_INIT = 16'h0202;
    SB_LUT4 i6_4_lut (.I0(n29), .I1(\o_Rx_DV_N_3488[12] ), .I2(n23), .I3(n4935), 
            .O(n15_adj_4657));
    defparam i6_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i8_4_lut (.I0(n15_adj_4657), .I1(\o_Rx_DV_N_3488[8] ), .I2(n14_adj_4656), 
            .I3(n58684), .O(n71282));
    defparam i8_4_lut.LUT_INIT = 16'h2000;
    SB_CARRY add_2787_12 (.CI(n52083), .I0(n2358), .I1(n2013), .CO(n52084));
    SB_LUT4 add_2787_11_lut (.I0(GND_net), .I1(n2359), .I2(n1879), .I3(n52082), 
            .O(n8235[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2787_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2787_11 (.CI(n52082), .I0(n2359), .I1(n1879), .CO(n52083));
    SB_LUT4 i1_2_lut_adj_1002 (.I0(baudrate[13]), .I1(baudrate[14]), .I2(GND_net), 
            .I3(GND_net), .O(n62543));
    defparam i1_2_lut_adj_1002.LUT_INIT = 16'heeee;
    SB_LUT4 add_2787_10_lut (.I0(GND_net), .I1(n2360), .I2(n1742), .I3(n52081), 
            .O(n8235[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2787_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2787_10 (.CI(n52081), .I0(n2360), .I1(n1742), .CO(n52082));
    SB_LUT4 add_2787_9_lut (.I0(GND_net), .I1(n2361), .I2(n1602), .I3(n52080), 
            .O(n8235[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2787_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2787_9 (.CI(n52080), .I0(n2361), .I1(n1602), .CO(n52081));
    SB_LUT4 add_2787_8_lut (.I0(GND_net), .I1(n2362), .I2(n1459), .I3(n52079), 
            .O(n8235[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2787_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2787_8 (.CI(n52079), .I0(n2362), .I1(n1459), .CO(n52080));
    SB_LUT4 add_2787_7_lut (.I0(GND_net), .I1(n2363), .I2(n1460), .I3(n52078), 
            .O(n8235[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2787_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2787_7 (.CI(n52078), .I0(n2363), .I1(n1460), .CO(n52079));
    SB_LUT4 add_2787_6_lut (.I0(GND_net), .I1(n2364), .I2(n1011), .I3(n52077), 
            .O(n8235[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2787_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2787_6 (.CI(n52077), .I0(n2364), .I1(n1011), .CO(n52078));
    SB_LUT4 add_2787_5_lut (.I0(GND_net), .I1(n2365), .I2(n856), .I3(n52076), 
            .O(n8235[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2787_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2787_5 (.CI(n52076), .I0(n2365), .I1(n856), .CO(n52077));
    SB_LUT4 add_2787_4_lut (.I0(GND_net), .I1(n2366), .I2(n698), .I3(n52075), 
            .O(n8235[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2787_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2787_4 (.CI(n52075), .I0(n2366), .I1(n698), .CO(n52076));
    SB_LUT4 add_2787_3_lut (.I0(GND_net), .I1(n2367), .I2(n858), .I3(n52074), 
            .O(n8235[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2787_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_i2160_1_lut (.I0(baudrate[15]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2638));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2160_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_2787_3 (.CI(n52074), .I0(n2367), .I1(n858), .CO(n52075));
    SB_LUT4 add_2787_2_lut (.I0(n59814), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n62045)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2787_2_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i48557_2_lut (.I0(baudrate[9]), .I1(n64228), .I2(GND_net), 
            .I3(GND_net), .O(n64242));
    defparam i48557_2_lut.LUT_INIT = 16'heeee;
    SB_CARRY add_2787_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n52074));
    SB_LUT4 add_2786_16_lut (.I0(GND_net), .I1(n2227), .I2(n2519), .I3(n52073), 
            .O(n8209[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2786_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2786_15_lut (.I0(GND_net), .I1(n2228), .I2(n2397), .I3(n52072), 
            .O(n8209[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2786_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2786_15 (.CI(n52072), .I0(n2228), .I1(n2397), .CO(n52073));
    SB_LUT4 add_2786_14_lut (.I0(GND_net), .I1(n2229), .I2(n2272), .I3(n52071), 
            .O(n8209[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2786_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2786_14 (.CI(n52071), .I0(n2229), .I1(n2272), .CO(n52072));
    SB_LUT4 add_2786_13_lut (.I0(GND_net), .I1(n2230), .I2(n2144), .I3(n52070), 
            .O(n8209[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2786_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2786_13 (.CI(n52070), .I0(n2230), .I1(n2144), .CO(n52071));
    SB_LUT4 add_2786_12_lut (.I0(GND_net), .I1(n2231), .I2(n2013), .I3(n52069), 
            .O(n8209[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2786_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2786_12 (.CI(n52069), .I0(n2231), .I1(n2013), .CO(n52070));
    SB_LUT4 add_2786_11_lut (.I0(GND_net), .I1(n2232), .I2(n1879), .I3(n52068), 
            .O(n8209[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2786_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2786_11 (.CI(n52068), .I0(n2232), .I1(n1879), .CO(n52069));
    SB_LUT4 add_2786_10_lut (.I0(GND_net), .I1(n2233), .I2(n1742), .I3(n52067), 
            .O(n8209[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2786_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2786_10 (.CI(n52067), .I0(n2233), .I1(n1742), .CO(n52068));
    SB_LUT4 add_2786_9_lut (.I0(GND_net), .I1(n2234), .I2(n1602), .I3(n52066), 
            .O(n8209[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2786_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2786_9 (.CI(n52066), .I0(n2234), .I1(n1602), .CO(n52067));
    SB_LUT4 add_2786_8_lut (.I0(GND_net), .I1(n2235), .I2(n1459), .I3(n52065), 
            .O(n8209[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2786_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_adj_1003 (.I0(baudrate[5]), .I1(baudrate[6]), .I2(GND_net), 
            .I3(GND_net), .O(n62551));
    defparam i1_2_lut_adj_1003.LUT_INIT = 16'heeee;
    SB_CARRY add_2786_8 (.CI(n52065), .I0(n2235), .I1(n1459), .CO(n52066));
    SB_LUT4 add_2786_7_lut (.I0(GND_net), .I1(n2236), .I2(n1460), .I3(n52064), 
            .O(n8209[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2786_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2786_7 (.CI(n52064), .I0(n2236), .I1(n1460), .CO(n52065));
    SB_LUT4 add_2786_6_lut (.I0(GND_net), .I1(n2237), .I2(n1011), .I3(n52063), 
            .O(n8209[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2786_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2786_6 (.CI(n52063), .I0(n2237), .I1(n1011), .CO(n52064));
    SB_LUT4 add_2786_5_lut (.I0(GND_net), .I1(n2238), .I2(n856), .I3(n52062), 
            .O(n8209[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2786_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2786_5 (.CI(n52062), .I0(n2238), .I1(n856), .CO(n52063));
    SB_LUT4 add_2786_4_lut (.I0(GND_net), .I1(n2239), .I2(n698), .I3(n52061), 
            .O(n8209[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2786_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2786_4 (.CI(n52061), .I0(n2239), .I1(n698), .CO(n52062));
    SB_LUT4 add_2786_3_lut (.I0(GND_net), .I1(n2240), .I2(n858), .I3(n52060), 
            .O(n8209[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2786_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2786_3 (.CI(n52060), .I0(n2240), .I1(n858), .CO(n52061));
    SB_LUT4 add_2786_2_lut (.I0(n59818), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n62043)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2786_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_2786_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n52060));
    SB_LUT4 add_2785_14_lut (.I0(GND_net), .I1(n2098), .I2(n2397), .I3(n52059), 
            .O(n8183[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2785_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2785_13_lut (.I0(GND_net), .I1(n2099), .I2(n2272), .I3(n52058), 
            .O(n8183[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2785_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2785_13 (.CI(n52058), .I0(n2099), .I1(n2272), .CO(n52059));
    SB_LUT4 add_2785_12_lut (.I0(GND_net), .I1(n2100), .I2(n2144), .I3(n52057), 
            .O(n8183[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2785_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2785_12 (.CI(n52057), .I0(n2100), .I1(n2144), .CO(n52058));
    SB_LUT4 add_2785_11_lut (.I0(GND_net), .I1(n2101), .I2(n2013), .I3(n52056), 
            .O(n8183[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2785_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2785_11 (.CI(n52056), .I0(n2101), .I1(n2013), .CO(n52057));
    SB_LUT4 add_2785_10_lut (.I0(GND_net), .I1(n2102), .I2(n1879), .I3(n52055), 
            .O(n8183[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2785_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2785_10 (.CI(n52055), .I0(n2102), .I1(n1879), .CO(n52056));
    SB_LUT4 add_2785_9_lut (.I0(GND_net), .I1(n2103), .I2(n1742), .I3(n52054), 
            .O(n8183[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2785_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2785_9 (.CI(n52054), .I0(n2103), .I1(n1742), .CO(n52055));
    SB_LUT4 add_2785_8_lut (.I0(GND_net), .I1(n2104), .I2(n1602), .I3(n52053), 
            .O(n8183[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2785_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2785_8 (.CI(n52053), .I0(n2104), .I1(n1602), .CO(n52054));
    SB_LUT4 add_2785_7_lut (.I0(GND_net), .I1(n2105), .I2(n1459), .I3(n52052), 
            .O(n8183[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2785_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2785_7 (.CI(n52052), .I0(n2105), .I1(n1459), .CO(n52053));
    SB_LUT4 add_2785_6_lut (.I0(GND_net), .I1(n2106), .I2(n1460), .I3(n52051), 
            .O(n8183[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2785_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2785_6 (.CI(n52051), .I0(n2106), .I1(n1460), .CO(n52052));
    SB_LUT4 add_2785_5_lut (.I0(GND_net), .I1(n2107), .I2(n1011), .I3(n52050), 
            .O(n8183[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2785_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_3_lut_adj_1004 (.I0(n25608), .I1(n48_adj_4655), .I2(baudrate[0]), 
            .I3(GND_net), .O(n805));
    defparam i1_3_lut_adj_1004.LUT_INIT = 16'hefef;
    SB_CARRY add_2785_5 (.CI(n52050), .I0(n2107), .I1(n1011), .CO(n52051));
    SB_LUT4 add_2785_4_lut (.I0(GND_net), .I1(n2108), .I2(n856), .I3(n52049), 
            .O(n8183[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2785_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2785_4 (.CI(n52049), .I0(n2108), .I1(n856), .CO(n52050));
    SB_LUT4 add_2785_3_lut (.I0(GND_net), .I1(n2109), .I2(n698), .I3(n52048), 
            .O(n8183[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2785_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2785_3 (.CI(n52048), .I0(n2109), .I1(n698), .CO(n52049));
    SB_LUT4 add_2785_2_lut (.I0(GND_net), .I1(n2110), .I2(n858), .I3(VCC_net), 
            .O(n8183[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2785_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2785_2 (.CI(VCC_net), .I0(n2110), .I1(n858), .CO(n52048));
    SB_LUT4 add_2784_14_lut (.I0(GND_net), .I1(n1966), .I2(n2272), .I3(n52047), 
            .O(n8157[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2784_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2784_13_lut (.I0(GND_net), .I1(n1967), .I2(n2144), .I3(n52046), 
            .O(n8157[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2784_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2784_13 (.CI(n52046), .I0(n1967), .I1(n2144), .CO(n52047));
    SB_LUT4 add_2784_12_lut (.I0(GND_net), .I1(n1968), .I2(n2013), .I3(n52045), 
            .O(n8157[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2784_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2784_12 (.CI(n52045), .I0(n1968), .I1(n2013), .CO(n52046));
    SB_LUT4 add_2784_11_lut (.I0(GND_net), .I1(n1969), .I2(n1879), .I3(n52044), 
            .O(n8157[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2784_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2784_11 (.CI(n52044), .I0(n1969), .I1(n1879), .CO(n52045));
    SB_LUT4 add_2784_10_lut (.I0(GND_net), .I1(n1970), .I2(n1742), .I3(n52043), 
            .O(n8157[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2784_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2784_10 (.CI(n52043), .I0(n1970), .I1(n1742), .CO(n52044));
    SB_LUT4 add_2784_9_lut (.I0(GND_net), .I1(n1971), .I2(n1602), .I3(n52042), 
            .O(n8157[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2784_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2784_9 (.CI(n52042), .I0(n1971), .I1(n1602), .CO(n52043));
    SB_LUT4 add_2784_8_lut (.I0(GND_net), .I1(n1972), .I2(n1459), .I3(n52041), 
            .O(n8157[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2784_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2784_8 (.CI(n52041), .I0(n1972), .I1(n1459), .CO(n52042));
    SB_LUT4 add_2784_7_lut (.I0(GND_net), .I1(n1973), .I2(n1460), .I3(n52040), 
            .O(n8157[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2784_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2784_7 (.CI(n52040), .I0(n1973), .I1(n1460), .CO(n52041));
    SB_LUT4 add_2784_6_lut (.I0(GND_net), .I1(n1974), .I2(n1011), .I3(n52039), 
            .O(n8157[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2784_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2784_6 (.CI(n52039), .I0(n1974), .I1(n1011), .CO(n52040));
    SB_LUT4 add_2784_5_lut (.I0(GND_net), .I1(n1975), .I2(n856), .I3(n52038), 
            .O(n8157[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2784_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2784_5 (.CI(n52038), .I0(n1975), .I1(n856), .CO(n52039));
    SB_LUT4 add_2784_4_lut (.I0(GND_net), .I1(n1976), .I2(n698), .I3(n52037), 
            .O(n8157[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2784_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_557_i42_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n805), .I3(GND_net), .O(n42_adj_4658));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_557_i42_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i53601_3_lut (.I0(n42_adj_4658), .I1(baudrate[2]), .I2(n804), 
            .I3(GND_net), .O(n69295));   // verilog/uart_rx.v(119[33:55])
    defparam i53601_3_lut.LUT_INIT = 16'h8e8e;
    SB_CARRY add_2784_4 (.CI(n52037), .I0(n1976), .I1(n698), .CO(n52038));
    SB_LUT4 i53602_3_lut (.I0(n69295), .I1(baudrate[3]), .I2(n803), .I3(GND_net), 
            .O(n69296));   // verilog/uart_rx.v(119[33:55])
    defparam i53602_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 add_2784_3_lut (.I0(GND_net), .I1(n1977), .I2(n858), .I3(n52036), 
            .O(n8157[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2784_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2784_3 (.CI(n52036), .I0(n1977), .I1(n858), .CO(n52037));
    SB_LUT4 add_2784_2_lut (.I0(GND_net), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n8157[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2784_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_557_i48_3_lut (.I0(n69296), .I1(baudrate[4]), 
            .I2(n59528), .I3(GND_net), .O(n48_adj_4556));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_557_i48_3_lut.LUT_INIT = 16'he8e8;
    SB_LUT4 div_37_i847_3_lut (.I0(n1115), .I1(n8001[19]), .I2(n294[17]), 
            .I3(GND_net), .O(n1265));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i847_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i946_3_lut (.I0(n1265), .I1(n8027[19]), .I2(n294[16]), 
            .I3(GND_net), .O(n1412));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i946_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1043_3_lut (.I0(n1412), .I1(n8053[19]), .I2(n294[15]), 
            .I3(GND_net), .O(n1556));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1043_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1138_3_lut (.I0(n1556), .I1(n8079[19]), .I2(n294[14]), 
            .I3(GND_net), .O(n1697));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1138_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1231_3_lut (.I0(n1697), .I1(n8105[19]), .I2(n294[13]), 
            .I3(GND_net), .O(n1835));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1231_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1322_3_lut (.I0(n1835), .I1(n8131[19]), .I2(n294[12]), 
            .I3(GND_net), .O(n1970));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1322_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1411_3_lut (.I0(n1970), .I1(n8157[19]), .I2(n294[11]), 
            .I3(GND_net), .O(n2102));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1411_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1498_3_lut (.I0(n2102), .I1(n8183[19]), .I2(n294[10]), 
            .I3(GND_net), .O(n2231));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1498_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2784_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n52036));
    SB_LUT4 add_2783_13_lut (.I0(GND_net), .I1(n1831), .I2(n2144), .I3(n52035), 
            .O(n8131[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2783_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2783_12_lut (.I0(GND_net), .I1(n1832), .I2(n2013), .I3(n52034), 
            .O(n8131[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2783_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2783_12 (.CI(n52034), .I0(n1832), .I1(n2013), .CO(n52035));
    SB_LUT4 div_37_i1583_3_lut (.I0(n2231), .I1(n8209[19]), .I2(n294[9]), 
            .I3(GND_net), .O(n2357));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1583_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2783_11_lut (.I0(GND_net), .I1(n1833), .I2(n1879), .I3(n52033), 
            .O(n8131[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2783_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2783_11 (.CI(n52033), .I0(n1833), .I1(n1879), .CO(n52034));
    SB_LUT4 add_2783_10_lut (.I0(GND_net), .I1(n1834), .I2(n1742), .I3(n52032), 
            .O(n8131[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2783_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2783_10 (.CI(n52032), .I0(n1834), .I1(n1742), .CO(n52033));
    SB_LUT4 div_37_LessThan_1602_i39_2_lut (.I0(n2357), .I1(baudrate[11]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_4659));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i2159_1_lut (.I0(baudrate[16]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2754));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2159_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_2794_25_lut (.I0(GND_net), .I1(n3151), .I2(n3186), .I3(n52222), 
            .O(n8417[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2794_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2783_9_lut (.I0(GND_net), .I1(n1835), .I2(n1602), .I3(n52031), 
            .O(n8131[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2783_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2783_9 (.CI(n52031), .I0(n1835), .I1(n1602), .CO(n52032));
    SB_LUT4 add_2783_8_lut (.I0(GND_net), .I1(n1836), .I2(n1459), .I3(n52030), 
            .O(n8131[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2783_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_i2158_1_lut (.I0(baudrate[17]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2867));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2158_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_LessThan_1602_i23_2_lut (.I0(n2365), .I1(baudrate[3]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_4660));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_765_i43_2_lut (.I0(n1113), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n43_adj_4661));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_765_i43_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_2783_8 (.CI(n52030), .I0(n1836), .I1(n1459), .CO(n52031));
    SB_LUT4 add_2783_7_lut (.I0(GND_net), .I1(n1837), .I2(n1460), .I3(n52029), 
            .O(n8131[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2783_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2794_24_lut (.I0(GND_net), .I1(n3152), .I2(n3082), .I3(n52221), 
            .O(n8417[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2794_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2794_24 (.CI(n52221), .I0(n3152), .I1(n3082), .CO(n52222));
    SB_CARRY add_2783_7 (.CI(n52029), .I0(n1837), .I1(n1460), .CO(n52030));
    SB_LUT4 add_2783_6_lut (.I0(GND_net), .I1(n1838), .I2(n1011), .I3(n52028), 
            .O(n8131[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2783_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2794_23_lut (.I0(GND_net), .I1(n3153), .I2(n3188), .I3(n52220), 
            .O(n8417[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2794_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2794_23 (.CI(n52220), .I0(n3153), .I1(n3188), .CO(n52221));
    SB_CARRY add_2783_6 (.CI(n52028), .I0(n1838), .I1(n1011), .CO(n52029));
    SB_LUT4 add_2794_22_lut (.I0(GND_net), .I1(n3154), .I2(n3084), .I3(n52219), 
            .O(n8417[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2794_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_i2157_1_lut (.I0(baudrate[18]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2977));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2157_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_LessThan_765_i38_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n1116), .I3(GND_net), .O(n38_adj_4662));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_765_i38_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_i2156_1_lut (.I0(baudrate[19]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n3084));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2156_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_LessThan_765_i42_3_lut (.I0(n40_adj_4663), .I1(baudrate[4]), 
            .I2(n43_adj_4661), .I3(GND_net), .O(n42_adj_4664));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_765_i42_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i54036_4_lut (.I0(n42_adj_4664), .I1(n38_adj_4662), .I2(n43_adj_4661), 
            .I3(n67796), .O(n69730));   // verilog/uart_rx.v(119[33:55])
    defparam i54036_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i54037_3_lut (.I0(n69730), .I1(baudrate[5]), .I2(n1112), .I3(GND_net), 
            .O(n69731));   // verilog/uart_rx.v(119[33:55])
    defparam i54037_3_lut.LUT_INIT = 16'h8e8e;
    SB_CARRY add_2794_22 (.CI(n52219), .I0(n3154), .I1(n3084), .CO(n52220));
    SB_LUT4 add_2794_21_lut (.I0(GND_net), .I1(n3155), .I2(n2977), .I3(n52218), 
            .O(n8417[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2794_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2794_21 (.CI(n52218), .I0(n3155), .I1(n2977), .CO(n52219));
    SB_LUT4 add_2783_5_lut (.I0(GND_net), .I1(n1839), .I2(n856), .I3(n52027), 
            .O(n8131[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2783_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2794_20_lut (.I0(GND_net), .I1(n3156), .I2(n2867), .I3(n52217), 
            .O(n8417[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2794_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2794_20 (.CI(n52217), .I0(n3156), .I1(n2867), .CO(n52218));
    SB_LUT4 add_2794_19_lut (.I0(GND_net), .I1(n3157), .I2(n2754), .I3(n52216), 
            .O(n8417[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2794_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2794_19 (.CI(n52216), .I0(n3157), .I1(n2754), .CO(n52217));
    SB_LUT4 div_37_i948_3_lut (.I0(n1267), .I1(n8027[17]), .I2(n294[16]), 
            .I3(GND_net), .O(n1414));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i948_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1045_3_lut (.I0(n1414), .I1(n8053[17]), .I2(n294[15]), 
            .I3(GND_net), .O(n1558));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1045_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1140_3_lut (.I0(n1558), .I1(n8079[17]), .I2(n294[14]), 
            .I3(GND_net), .O(n1699));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1140_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1233_3_lut (.I0(n1699), .I1(n8105[17]), .I2(n294[13]), 
            .I3(GND_net), .O(n1837));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1233_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_adj_1005 (.I0(n69345), .I1(baudrate[8]), .I2(n1408), 
            .I3(n62039), .O(n1560));   // verilog/uart_rx.v(119[33:55])
    defparam i1_2_lut_4_lut_adj_1005.LUT_INIT = 16'h7100;
    SB_LUT4 div_37_i1324_3_lut (.I0(n1837), .I1(n8131[17]), .I2(n294[12]), 
            .I3(GND_net), .O(n1972));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1324_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1413_3_lut (.I0(n1972), .I1(n8157[17]), .I2(n294[11]), 
            .I3(GND_net), .O(n2104));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1413_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1500_3_lut (.I0(n2104), .I1(n8183[17]), .I2(n294[10]), 
            .I3(GND_net), .O(n2233));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1500_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1585_3_lut (.I0(n2233), .I1(n8209[17]), .I2(n294[9]), 
            .I3(GND_net), .O(n2359));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1585_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1602_i35_2_lut (.I0(n2359), .I1(baudrate[9]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_4665));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_2794_18_lut (.I0(GND_net), .I1(n3158), .I2(n2638), .I3(n52215), 
            .O(n8417[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2794_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2783_5 (.CI(n52027), .I0(n1839), .I1(n856), .CO(n52028));
    SB_CARRY add_2794_18 (.CI(n52215), .I0(n3158), .I1(n2638), .CO(n52216));
    SB_LUT4 add_2794_17_lut (.I0(GND_net), .I1(n3159), .I2(n2519), .I3(n52214), 
            .O(n8417[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2794_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2783_4_lut (.I0(GND_net), .I1(n1840), .I2(n698), .I3(n52026), 
            .O(n8131[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2783_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2783_4 (.CI(n52026), .I0(n1840), .I1(n698), .CO(n52027));
    SB_LUT4 add_2783_3_lut (.I0(GND_net), .I1(n1841), .I2(n858), .I3(n52025), 
            .O(n8131[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2783_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2794_17 (.CI(n52214), .I0(n3159), .I1(n2519), .CO(n52215));
    SB_LUT4 add_2794_16_lut (.I0(GND_net), .I1(n3160), .I2(n2397), .I3(n52213), 
            .O(n8417[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2794_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2783_3 (.CI(n52025), .I0(n1841), .I1(n858), .CO(n52026));
    SB_CARRY add_2794_16 (.CI(n52213), .I0(n3160), .I1(n2397), .CO(n52214));
    SB_LUT4 add_2783_2_lut (.I0(n59827), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n62041)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2783_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_2783_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n52025));
    SB_LUT4 add_2794_15_lut (.I0(GND_net), .I1(n3161), .I2(n2272), .I3(n52212), 
            .O(n8417[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2794_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_i2155_1_lut (.I0(baudrate[20]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n3188));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2155_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_2782_11_lut (.I0(GND_net), .I1(n1693), .I2(n2013), .I3(n52024), 
            .O(n8105[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2782_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2794_15 (.CI(n52212), .I0(n3161), .I1(n2272), .CO(n52213));
    SB_LUT4 add_2782_10_lut (.I0(GND_net), .I1(n1694), .I2(n1879), .I3(n52023), 
            .O(n8105[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2782_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i52356_4_lut (.I0(n25598), .I1(n67382), .I2(n48_adj_4654), 
            .I3(baudrate[0]), .O(n804));
    defparam i52356_4_lut.LUT_INIT = 16'h3633;
    SB_LUT4 i55106_2_lut_4_lut (.I0(n69345), .I1(baudrate[8]), .I2(n1408), 
            .I3(n64242), .O(n294[15]));   // verilog/uart_rx.v(119[33:55])
    defparam i55106_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_LUT4 i52082_3_lut_4_lut (.I0(n1413), .I1(baudrate[3]), .I2(baudrate[2]), 
            .I3(n1414), .O(n67776));   // verilog/uart_rx.v(119[33:55])
    defparam i52082_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 add_2794_14_lut (.I0(GND_net), .I1(n3162), .I2(n2144), .I3(n52211), 
            .O(n8417[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2794_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2794_14 (.CI(n52211), .I0(n3162), .I1(n2144), .CO(n52212));
    SB_LUT4 add_2794_13_lut (.I0(GND_net), .I1(n3163), .I2(n2013), .I3(n52210), 
            .O(n8417[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2794_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2782_10 (.CI(n52023), .I0(n1694), .I1(n1879), .CO(n52024));
    SB_LUT4 i5738_2_lut (.I0(n20912), .I1(n11417), .I2(GND_net), .I3(GND_net), 
            .O(n42_adj_4666));   // verilog/uart_rx.v(119[33:55])
    defparam i5738_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 div_37_i641_4_lut (.I0(n804), .I1(n42_adj_4667), .I2(n294[19]), 
            .I3(baudrate[2]), .O(n960));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i641_4_lut.LUT_INIT = 16'h6a9a;
    SB_LUT4 add_2782_9_lut (.I0(GND_net), .I1(n1695), .I2(n1742), .I3(n52022), 
            .O(n8105[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2782_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2782_9 (.CI(n52022), .I0(n1695), .I1(n1742), .CO(n52023));
    SB_CARRY add_2794_13 (.CI(n52210), .I0(n3163), .I1(n2013), .CO(n52211));
    SB_LUT4 div_37_i744_4_lut (.I0(n960), .I1(baudrate[3]), .I2(n294[18]), 
            .I3(n42_adj_4666), .O(n1113));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i744_4_lut.LUT_INIT = 16'h6a9a;
    SB_LUT4 add_2782_8_lut (.I0(GND_net), .I1(n1696), .I2(n1602), .I3(n52021), 
            .O(n8105[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2782_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_965_i36_3_lut_3_lut (.I0(n1413), .I1(baudrate[3]), 
            .I2(baudrate[2]), .I3(GND_net), .O(n36_adj_4647));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_965_i36_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 div_37_i845_3_lut (.I0(n1113), .I1(n8001[21]), .I2(n294[17]), 
            .I3(GND_net), .O(n1263));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i845_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i944_3_lut (.I0(n1263), .I1(n8027[21]), .I2(n294[16]), 
            .I3(GND_net), .O(n1410));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i944_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1041_3_lut (.I0(n1410), .I1(n8053[21]), .I2(n294[15]), 
            .I3(GND_net), .O(n1554));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1041_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1136_3_lut (.I0(n1554), .I1(n8079[21]), .I2(n294[14]), 
            .I3(GND_net), .O(n1695));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1136_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2794_12_lut (.I0(GND_net), .I1(n3164), .I2(n1879), .I3(n52209), 
            .O(n8417[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2794_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2782_8 (.CI(n52021), .I0(n1696), .I1(n1602), .CO(n52022));
    SB_LUT4 add_2782_7_lut (.I0(GND_net), .I1(n1697), .I2(n1459), .I3(n52020), 
            .O(n8105[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2782_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2794_12 (.CI(n52209), .I0(n3164), .I1(n1879), .CO(n52210));
    SB_LUT4 add_2794_11_lut (.I0(GND_net), .I1(n3165), .I2(n1742), .I3(n52208), 
            .O(n8417[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2794_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_i1229_3_lut (.I0(n1695), .I1(n8105[21]), .I2(n294[13]), 
            .I3(GND_net), .O(n1833));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1229_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1250_i43_2_lut (.I0(n1833), .I1(baudrate[9]), 
            .I2(GND_net), .I3(GND_net), .O(n43_adj_4668));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1250_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1250_i29_2_lut (.I0(n1840), .I1(baudrate[2]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_4669));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1250_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i52051_4_lut (.I0(n35_adj_4518), .I1(n33_adj_4516), .I2(n31_adj_4517), 
            .I3(n29_adj_4669), .O(n67745));
    defparam i52051_4_lut.LUT_INIT = 16'haaab;
    SB_CARRY add_2794_11 (.CI(n52208), .I0(n3165), .I1(n1742), .CO(n52209));
    SB_LUT4 i52063_3_lut_4_lut (.I0(n1699), .I1(baudrate[4]), .I2(baudrate[3]), 
            .I3(n1700), .O(n67757));   // verilog/uart_rx.v(119[33:55])
    defparam i52063_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_CARRY add_2782_7 (.CI(n52020), .I0(n1697), .I1(n1459), .CO(n52021));
    SB_LUT4 div_37_LessThan_1157_i34_3_lut_3_lut (.I0(n1699), .I1(baudrate[4]), 
            .I2(baudrate[3]), .I3(GND_net), .O(n34_adj_4623));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1157_i34_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 i1_2_lut_4_lut_adj_1006 (.I0(n69030), .I1(baudrate[16]), .I2(n2476), 
            .I3(n62047), .O(n2612));   // verilog/uart_rx.v(119[33:55])
    defparam i1_2_lut_4_lut_adj_1006.LUT_INIT = 16'h7100;
    SB_LUT4 add_2782_6_lut (.I0(GND_net), .I1(n1698), .I2(n1460), .I3(n52019), 
            .O(n8105[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2782_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2782_6 (.CI(n52019), .I0(n1698), .I1(n1460), .CO(n52020));
    SB_LUT4 add_2794_10_lut (.I0(GND_net), .I1(n3166), .I2(n1602), .I3(n52207), 
            .O(n8417[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2794_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2782_5_lut (.I0(GND_net), .I1(n1699), .I2(n1011), .I3(n52018), 
            .O(n8105[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2782_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2794_10 (.CI(n52207), .I0(n3166), .I1(n1602), .CO(n52208));
    SB_LUT4 add_2794_9_lut (.I0(GND_net), .I1(n3167), .I2(n1459), .I3(n52206), 
            .O(n8417[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2794_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2794_9 (.CI(n52206), .I0(n3167), .I1(n1459), .CO(n52207));
    SB_LUT4 add_2794_8_lut (.I0(GND_net), .I1(n3168), .I2(n1460), .I3(n52205), 
            .O(n8417[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2794_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2794_8 (.CI(n52205), .I0(n3168), .I1(n1460), .CO(n52206));
    SB_LUT4 add_2794_7_lut (.I0(GND_net), .I1(n3169), .I2(n1011), .I3(n52204), 
            .O(n8417[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2794_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2794_7 (.CI(n52204), .I0(n3169), .I1(n1011), .CO(n52205));
    SB_LUT4 add_2794_6_lut (.I0(GND_net), .I1(n3170), .I2(n856), .I3(n52203), 
            .O(n8417[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2794_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2782_5 (.CI(n52018), .I0(n1699), .I1(n1011), .CO(n52019));
    SB_CARRY add_2794_6 (.CI(n52203), .I0(n3170), .I1(n856), .CO(n52204));
    SB_LUT4 add_2782_4_lut (.I0(GND_net), .I1(n1700), .I2(n856), .I3(n52017), 
            .O(n8105[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2782_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2794_5_lut (.I0(GND_net), .I1(n3171), .I2(n698), .I3(n52202), 
            .O(n8417[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2794_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2794_5 (.CI(n52202), .I0(n3171), .I1(n698), .CO(n52203));
    SB_LUT4 add_2794_4_lut (.I0(GND_net), .I1(n3172), .I2(n858), .I3(n52201), 
            .O(n8417[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2794_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2782_4 (.CI(n52017), .I0(n1700), .I1(n856), .CO(n52018));
    SB_CARRY add_2794_4 (.CI(n52201), .I0(n3172), .I1(n858), .CO(n52202));
    SB_LUT4 add_2794_3_lut (.I0(n59786), .I1(GND_net), .I2(n538), .I3(n52200), 
            .O(n62059)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2794_3_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_2794_3 (.CI(n52200), .I0(GND_net), .I1(n538), .CO(n52201));
    SB_CARRY add_2794_2 (.CI(VCC_net), .I0(GND_net), .I1(VCC_net), .CO(n52200));
    SB_LUT4 add_2793_23_lut (.I0(GND_net), .I1(n3046), .I2(n3082), .I3(n52199), 
            .O(n8391[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2793_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2793_22_lut (.I0(GND_net), .I1(n3047), .I2(n3188), .I3(n52198), 
            .O(n8391[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2793_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2793_22 (.CI(n52198), .I0(n3047), .I1(n3188), .CO(n52199));
    SB_LUT4 add_2782_3_lut (.I0(GND_net), .I1(n1701), .I2(n698), .I3(n52016), 
            .O(n8105[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2782_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2793_21_lut (.I0(GND_net), .I1(n3048), .I2(n3084), .I3(n52197), 
            .O(n8391[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2793_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2793_21 (.CI(n52197), .I0(n3048), .I1(n3084), .CO(n52198));
    SB_LUT4 add_2793_20_lut (.I0(GND_net), .I1(n3049), .I2(n2977), .I3(n52196), 
            .O(n8391[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2793_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2793_20 (.CI(n52196), .I0(n3049), .I1(n2977), .CO(n52197));
    SB_LUT4 add_2793_19_lut (.I0(GND_net), .I1(n3050), .I2(n2867), .I3(n52195), 
            .O(n8391[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2793_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2782_3 (.CI(n52016), .I0(n1701), .I1(n698), .CO(n52017));
    SB_LUT4 div_37_LessThan_1250_i40_3_lut (.I0(n32_adj_4670), .I1(baudrate[9]), 
            .I2(n43_adj_4668), .I3(GND_net), .O(n40_adj_4671));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1250_i40_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1250_i28_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n1841), .I3(GND_net), .O(n28_adj_4672));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1250_i28_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i53583_3_lut (.I0(n28_adj_4672), .I1(baudrate[5]), .I2(n35_adj_4518), 
            .I3(GND_net), .O(n69277));   // verilog/uart_rx.v(119[33:55])
    defparam i53583_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2793_19 (.CI(n52195), .I0(n3050), .I1(n2867), .CO(n52196));
    SB_LUT4 add_2782_2_lut (.I0(GND_net), .I1(n1702), .I2(n858), .I3(VCC_net), 
            .O(n8105[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2782_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2793_18_lut (.I0(GND_net), .I1(n3051), .I2(n2754), .I3(n52194), 
            .O(n8391[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2793_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2782_2 (.CI(VCC_net), .I0(n1702), .I1(n858), .CO(n52016));
    SB_CARRY add_2793_18 (.CI(n52194), .I0(n3051), .I1(n2754), .CO(n52195));
    SB_LUT4 add_2781_11_lut (.I0(GND_net), .I1(n1552), .I2(n1879), .I3(n52015), 
            .O(n8079[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2781_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i53584_3_lut (.I0(n69277), .I1(baudrate[6]), .I2(n37_adj_4519), 
            .I3(GND_net), .O(n69278));   // verilog/uart_rx.v(119[33:55])
    defparam i53584_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52047_4_lut (.I0(n41_adj_4520), .I1(n39_adj_4521), .I2(n37_adj_4519), 
            .I3(n67745), .O(n67741));
    defparam i52047_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 add_2781_10_lut (.I0(GND_net), .I1(n1553), .I2(n1742), .I3(n52014), 
            .O(n8079[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2781_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2781_10 (.CI(n52014), .I0(n1553), .I1(n1742), .CO(n52015));
    SB_LUT4 add_2781_9_lut (.I0(GND_net), .I1(n1554), .I2(n1602), .I3(n52013), 
            .O(n8079[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2781_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2793_17_lut (.I0(GND_net), .I1(n3052), .I2(n2638), .I3(n52193), 
            .O(n8391[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2793_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2793_17 (.CI(n52193), .I0(n3052), .I1(n2638), .CO(n52194));
    SB_CARRY add_2781_9 (.CI(n52013), .I0(n1554), .I1(n1602), .CO(n52014));
    SB_LUT4 add_2793_16_lut (.I0(GND_net), .I1(n3053), .I2(n2519), .I3(n52192), 
            .O(n8391[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2793_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i54032_4_lut (.I0(n40_adj_4671), .I1(n30_adj_4673), .I2(n43_adj_4668), 
            .I3(n67739), .O(n69726));   // verilog/uart_rx.v(119[33:55])
    defparam i54032_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 add_2781_8_lut (.I0(GND_net), .I1(n1555), .I2(n1459), .I3(n52012), 
            .O(n8079[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2781_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2793_16 (.CI(n52192), .I0(n3053), .I1(n2519), .CO(n52193));
    SB_LUT4 add_2793_15_lut (.I0(GND_net), .I1(n3054), .I2(n2397), .I3(n52191), 
            .O(n8391[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2793_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2793_15 (.CI(n52191), .I0(n3054), .I1(n2397), .CO(n52192));
    SB_CARRY add_2781_8 (.CI(n52012), .I0(n1555), .I1(n1459), .CO(n52013));
    SB_LUT4 add_2793_14_lut (.I0(GND_net), .I1(n3055), .I2(n2272), .I3(n52190), 
            .O(n8391[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2793_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2793_14 (.CI(n52190), .I0(n3055), .I1(n2272), .CO(n52191));
    SB_LUT4 add_2793_13_lut (.I0(GND_net), .I1(n3056), .I2(n2144), .I3(n52189), 
            .O(n8391[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2793_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2781_7_lut (.I0(GND_net), .I1(n1556), .I2(n1460), .I3(n52011), 
            .O(n8079[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2781_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2781_7 (.CI(n52011), .I0(n1556), .I1(n1460), .CO(n52012));
    SB_LUT4 i52777_3_lut (.I0(n69278), .I1(baudrate[7]), .I2(n39_adj_4521), 
            .I3(GND_net), .O(n68471));   // verilog/uart_rx.v(119[33:55])
    defparam i52777_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i54224_4_lut (.I0(n68471), .I1(n69726), .I2(n43_adj_4668), 
            .I3(n67741), .O(n69918));   // verilog/uart_rx.v(119[33:55])
    defparam i54224_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i54225_3_lut (.I0(n69918), .I1(baudrate[10]), .I2(n1832), 
            .I3(GND_net), .O(n69919));   // verilog/uart_rx.v(119[33:55])
    defparam i54225_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i54198_3_lut (.I0(n69919), .I1(baudrate[11]), .I2(n1831), 
            .I3(GND_net), .O(n48_adj_4614));   // verilog/uart_rx.v(119[33:55])
    defparam i54198_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i1_2_lut_adj_1007 (.I0(n62041), .I1(n48_adj_4614), .I2(GND_net), 
            .I3(GND_net), .O(n1977));
    defparam i1_2_lut_adj_1007.LUT_INIT = 16'h2222;
    SB_LUT4 div_37_i1418_3_lut (.I0(n1977), .I1(n8157[12]), .I2(n294[11]), 
            .I3(GND_net), .O(n2109));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1418_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i55124_2_lut_4_lut (.I0(n69030), .I1(baudrate[16]), .I2(n2476), 
            .I3(n63979), .O(n294[7]));   // verilog/uart_rx.v(119[33:55])
    defparam i55124_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_LUT4 div_37_i1505_3_lut (.I0(n2109), .I1(n8183[12]), .I2(n294[10]), 
            .I3(GND_net), .O(n2238));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1505_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1590_3_lut (.I0(n2238), .I1(n8209[12]), .I2(n294[9]), 
            .I3(GND_net), .O(n2364));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1590_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1602_i25_2_lut (.I0(n2364), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_4674));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i942_3_lut (.I0(n1261), .I1(n8027[23]), .I2(n294[16]), 
            .I3(GND_net), .O(n1408));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i942_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1039_3_lut (.I0(n1408), .I1(n8053[23]), .I2(n294[15]), 
            .I3(GND_net), .O(n1552));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1039_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1134_3_lut (.I0(n1552), .I1(n8079[23]), .I2(n294[14]), 
            .I3(GND_net), .O(n1693));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1134_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1227_3_lut (.I0(n1693), .I1(n8105[23]), .I2(n294[13]), 
            .I3(GND_net), .O(n1831));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1227_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1318_3_lut (.I0(n1831), .I1(n8131[23]), .I2(n294[12]), 
            .I3(GND_net), .O(n1966));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1318_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1407_3_lut (.I0(n1966), .I1(n8157[23]), .I2(n294[11]), 
            .I3(GND_net), .O(n2098));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1407_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1494_3_lut (.I0(n2098), .I1(n8183[23]), .I2(n294[10]), 
            .I3(GND_net), .O(n2227));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1494_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1008 (.I0(baudrate[23]), .I1(baudrate[28]), .I2(baudrate[27]), 
            .I3(baudrate[0]), .O(n62363));
    defparam i1_4_lut_adj_1008.LUT_INIT = 16'h0100;
    SB_LUT4 i48517_4_lut (.I0(baudrate[25]), .I1(baudrate[31]), .I2(baudrate[24]), 
            .I3(baudrate[29]), .O(n64202));
    defparam i48517_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1009 (.I0(n59613), .I1(n62363), .I2(n63609), 
            .I3(baudrate[16]), .O(n62391));
    defparam i1_4_lut_adj_1009.LUT_INIT = 16'h0004;
    SB_LUT4 i48589_4_lut (.I0(n64202), .I1(n64124), .I2(n64128), .I3(n63961), 
            .O(n64274));
    defparam i48589_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i54336_4_lut (.I0(n64262), .I1(n67378), .I2(n64274), .I3(n62391), 
            .O(n70030));
    defparam i54336_4_lut.LUT_INIT = 16'hc9cc;
    SB_LUT4 div_37_i535_4_lut (.I0(n70030), .I1(n44_adj_4675), .I2(n294[20]), 
            .I3(baudrate[2]), .O(n803));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i535_4_lut.LUT_INIT = 16'h9565;
    SB_LUT4 div_37_i640_4_lut (.I0(n803), .I1(baudrate[3]), .I2(n294[19]), 
            .I3(n44_adj_4676), .O(n959));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i640_4_lut.LUT_INIT = 16'h6a9a;
    SB_LUT4 i1_2_lut_3_lut (.I0(\r_SM_Main[1] ), .I1(r_SM_Main[0]), .I2(\r_SM_Main[2] ), 
            .I3(GND_net), .O(n4_adj_4559));
    defparam i1_2_lut_3_lut.LUT_INIT = 16'hfdfd;
    SB_LUT4 div_37_i743_4_lut (.I0(n959), .I1(baudrate[4]), .I2(n294[18]), 
            .I3(n44_adj_4677), .O(n1112));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i743_4_lut.LUT_INIT = 16'h6a9a;
    SB_LUT4 div_37_i844_3_lut (.I0(n1112), .I1(n8001[22]), .I2(n294[17]), 
            .I3(GND_net), .O(n1262));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i844_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i943_3_lut (.I0(n1262), .I1(n8027[22]), .I2(n294[16]), 
            .I3(GND_net), .O(n1409));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i943_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1040_3_lut (.I0(n1409), .I1(n8053[22]), .I2(n294[15]), 
            .I3(GND_net), .O(n1553));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1040_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1135_3_lut (.I0(n1553), .I1(n8079[22]), .I2(n294[14]), 
            .I3(GND_net), .O(n1694));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1135_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1228_3_lut (.I0(n1694), .I1(n8105[22]), .I2(n294[13]), 
            .I3(GND_net), .O(n1832));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1228_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1319_3_lut (.I0(n1832), .I1(n8131[22]), .I2(n294[12]), 
            .I3(GND_net), .O(n1967));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1319_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1408_3_lut (.I0(n1967), .I1(n8157[22]), .I2(n294[11]), 
            .I3(GND_net), .O(n2099));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1408_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1495_3_lut (.I0(n2099), .I1(n8183[22]), .I2(n294[10]), 
            .I3(GND_net), .O(n2228));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1495_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1517_i23_2_lut (.I0(n2239), .I1(baudrate[2]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_4678));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i51989_4_lut (.I0(n29_adj_4522), .I1(n27_adj_4524), .I2(n25_adj_4526), 
            .I3(n23_adj_4678), .O(n67683));
    defparam i51989_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i51983_4_lut (.I0(n35_adj_4525), .I1(n33_adj_4530), .I2(n31_adj_4523), 
            .I3(n67683), .O(n67677));
    defparam i51983_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_37_LessThan_1517_i22_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n2240), .I3(GND_net), .O(n22_adj_4679));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i22_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_1517_i30_3_lut (.I0(n28_adj_4680), .I1(baudrate[7]), 
            .I2(n33_adj_4530), .I3(GND_net), .O(n30_adj_4681));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1517_i34_3_lut (.I0(n26_adj_4682), .I1(baudrate[9]), 
            .I2(n37_adj_4527), .I3(GND_net), .O(n34_adj_4683));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i34_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i54060_4_lut (.I0(n34_adj_4683), .I1(n24_adj_4684), .I2(n37_adj_4527), 
            .I3(n67675), .O(n69754));   // verilog/uart_rx.v(119[33:55])
    defparam i54060_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i54061_3_lut (.I0(n69754), .I1(baudrate[10]), .I2(n39_adj_4528), 
            .I3(GND_net), .O(n69755));   // verilog/uart_rx.v(119[33:55])
    defparam i54061_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53880_3_lut (.I0(n69755), .I1(baudrate[11]), .I2(n41_adj_4529), 
            .I3(GND_net), .O(n69574));   // verilog/uart_rx.v(119[33:55])
    defparam i53880_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53754_4_lut (.I0(n41_adj_4529), .I1(n39_adj_4528), .I2(n37_adj_4527), 
            .I3(n67677), .O(n69448));
    defparam i53754_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i53832_4_lut (.I0(n30_adj_4681), .I1(n22_adj_4679), .I2(n33_adj_4530), 
            .I3(n67681), .O(n69526));   // verilog/uart_rx.v(119[33:55])
    defparam i53832_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i52799_3_lut (.I0(n69574), .I1(baudrate[12]), .I2(n43_adj_4531), 
            .I3(GND_net), .O(n68493));   // verilog/uart_rx.v(119[33:55])
    defparam i52799_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i54028_4_lut (.I0(n68493), .I1(n69526), .I2(n43_adj_4531), 
            .I3(n69448), .O(n69722));   // verilog/uart_rx.v(119[33:55])
    defparam i54028_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i54029_3_lut (.I0(n69722), .I1(baudrate[13]), .I2(n2228), 
            .I3(GND_net), .O(n69723));   // verilog/uart_rx.v(119[33:55])
    defparam i54029_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i53952_3_lut (.I0(n69723), .I1(baudrate[14]), .I2(n2227), 
            .I3(GND_net), .O(n48_adj_4685));   // verilog/uart_rx.v(119[33:55])
    defparam i53952_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i1_2_lut_adj_1010 (.I0(n62043), .I1(n48_adj_4685), .I2(GND_net), 
            .I3(GND_net), .O(n2367));
    defparam i1_2_lut_adj_1010.LUT_INIT = 16'h2222;
    SB_LUT4 i1_2_lut_adj_1011 (.I0(baudrate[14]), .I1(baudrate[15]), .I2(GND_net), 
            .I3(GND_net), .O(n63513));
    defparam i1_2_lut_adj_1011.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_1012 (.I0(baudrate[12]), .I1(baudrate[13]), .I2(GND_net), 
            .I3(GND_net), .O(n63369));
    defparam i1_2_lut_adj_1012.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_1013 (.I0(baudrate[10]), .I1(baudrate[11]), .I2(GND_net), 
            .I3(GND_net), .O(n63371));
    defparam i1_2_lut_adj_1013.LUT_INIT = 16'heeee;
    SB_LUT4 i43976_2_lut (.I0(baudrate[2]), .I1(baudrate[3]), .I2(GND_net), 
            .I3(GND_net), .O(n59613));
    defparam i43976_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i48457_2_lut (.I0(baudrate[21]), .I1(baudrate[22]), .I2(GND_net), 
            .I3(GND_net), .O(n64142));
    defparam i48457_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i48577_4_lut (.I0(n64142), .I1(n62687), .I2(n63371), .I3(baudrate[9]), 
            .O(n64262));
    defparam i48577_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1014 (.I0(baudrate[17]), .I1(n64170), .I2(baudrate[2]), 
            .I3(n43066), .O(n61975));
    defparam i1_4_lut_adj_1014.LUT_INIT = 16'h0100;
    SB_LUT4 i1_4_lut_adj_1015 (.I0(n64214), .I1(n61975), .I2(n25574), 
            .I3(n64124), .O(n61167));
    defparam i1_4_lut_adj_1015.LUT_INIT = 16'h0004;
    SB_LUT4 i1_4_lut_adj_1016 (.I0(baudrate[23]), .I1(baudrate[27]), .I2(baudrate[25]), 
            .I3(n43068), .O(n62307));
    defparam i1_4_lut_adj_1016.LUT_INIT = 16'h0100;
    SB_LUT4 i1_4_lut_adj_1017 (.I0(n62307), .I1(baudrate[29]), .I2(baudrate[16]), 
            .I3(baudrate[28]), .O(n62325));
    defparam i1_4_lut_adj_1017.LUT_INIT = 16'h0002;
    SB_LUT4 i48591_4_lut (.I0(n64208), .I1(n64124), .I2(n64128), .I3(n63961), 
            .O(n64276));
    defparam i48591_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1018 (.I0(n64262), .I1(n64276), .I2(n59613), 
            .I3(n62325), .O(n60333));
    defparam i1_4_lut_adj_1018.LUT_INIT = 16'h0100;
    SB_LUT4 i1_2_lut_4_lut_adj_1019 (.I0(n69989), .I1(baudrate[20]), .I2(n2938), 
            .I3(n62055), .O(n3066));   // verilog/uart_rx.v(119[33:55])
    defparam i1_2_lut_4_lut_adj_1019.LUT_INIT = 16'h7100;
    SB_LUT4 i1_4_lut_adj_1020 (.I0(n62545), .I1(n62541), .I2(n62543), 
            .I3(n63961), .O(n62563));
    defparam i1_4_lut_adj_1020.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1021 (.I0(n64170), .I1(n62549), .I2(n62551), 
            .I3(n62547), .O(n62565));
    defparam i1_4_lut_adj_1021.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_3_lut_adj_1022 (.I0(n62565), .I1(n25577), .I2(n62563), 
            .I3(GND_net), .O(n25598));
    defparam i1_3_lut_adj_1022.LUT_INIT = 16'hfefe;
    SB_LUT4 div_37_LessThan_341_i48_3_lut (.I0(n60333), .I1(baudrate[2]), 
            .I2(n61167), .I3(GND_net), .O(n48_adj_4654));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_341_i48_3_lut.LUT_INIT = 16'he8e8;
    SB_LUT4 i48299_2_lut (.I0(baudrate[17]), .I1(n25574), .I2(GND_net), 
            .I3(GND_net), .O(n63979));
    defparam i48299_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i55152_2_lut (.I0(n48_adj_4654), .I1(n25598), .I2(GND_net), 
            .I3(GND_net), .O(n294[21]));
    defparam i55152_2_lut.LUT_INIT = 16'h1111;
    SB_LUT4 i55139_2_lut_4_lut (.I0(n69989), .I1(baudrate[20]), .I2(n2938), 
            .I3(n64248), .O(n294[3]));   // verilog/uart_rx.v(119[33:55])
    defparam i55139_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_LUT4 i54514_2_lut (.I0(n48_adj_4655), .I1(n25608), .I2(GND_net), 
            .I3(GND_net), .O(n294[20]));   // verilog/uart_rx.v(119[33:55])
    defparam i54514_2_lut.LUT_INIT = 16'h1111;
    SB_LUT4 i1_4_lut_adj_1023 (.I0(n63381), .I1(n63513), .I2(baudrate[16]), 
            .I3(n43066), .O(n62629));
    defparam i1_4_lut_adj_1023.LUT_INIT = 16'h0100;
    SB_LUT4 i52416_3_lut (.I0(n60333), .I1(n61167), .I2(baudrate[2]), 
            .I3(GND_net), .O(n67007));   // verilog/uart_rx.v(119[33:55])
    defparam i52416_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i52272_4_lut (.I0(n59613), .I1(n62629), .I2(n63383), .I3(n62683), 
            .O(n67008));   // verilog/uart_rx.v(119[33:55])
    defparam i52272_4_lut.LUT_INIT = 16'h0004;
    SB_LUT4 div_37_i427_4_lut (.I0(n67008), .I1(n67007), .I2(n294[21]), 
            .I3(n63979), .O(n59526));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i427_4_lut.LUT_INIT = 16'hc0ca;
    SB_LUT4 div_37_i534_3_lut (.I0(n59526), .I1(n294[20]), .I2(baudrate[3]), 
            .I3(GND_net), .O(n59528));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i534_3_lut.LUT_INIT = 16'h6a6a;
    SB_LUT4 i54517_2_lut (.I0(n48_adj_4652), .I1(n25605), .I2(GND_net), 
            .I3(GND_net), .O(n294[18]));   // verilog/uart_rx.v(119[33:55])
    defparam i54517_2_lut.LUT_INIT = 16'h1111;
    SB_LUT4 i5581_4_lut (.I0(n803), .I1(baudrate[3]), .I2(n11253), .I3(n20904), 
            .O(n46_adj_4686));   // verilog/uart_rx.v(119[33:55])
    defparam i5581_4_lut.LUT_INIT = 16'hbbb2;
    SB_LUT4 div_37_i639_4_lut (.I0(n59528), .I1(n294[19]), .I2(n46_adj_4686), 
            .I3(baudrate[4]), .O(n59530));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i639_4_lut.LUT_INIT = 16'h6aa6;
    SB_LUT4 i5752_4_lut (.I0(n959), .I1(baudrate[4]), .I2(n11424), .I3(n20914), 
            .O(n46_adj_4687));   // verilog/uart_rx.v(119[33:55])
    defparam i5752_4_lut.LUT_INIT = 16'hbbb2;
    SB_LUT4 div_37_i742_4_lut (.I0(n59530), .I1(n294[18]), .I2(n46_adj_4687), 
            .I3(baudrate[5]), .O(n1111));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i742_4_lut.LUT_INIT = 16'h9559;
    SB_LUT4 div_37_i843_3_lut (.I0(n1111), .I1(n8001[23]), .I2(n294[17]), 
            .I3(GND_net), .O(n1261));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i843_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_866_i36_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n1267), .I3(GND_net), .O(n36_adj_4688));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_866_i36_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_866_i40_3_lut (.I0(n38_adj_4689), .I1(baudrate[4]), 
            .I2(n41_adj_4532), .I3(GND_net), .O(n40_adj_4690));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_866_i40_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i54048_4_lut (.I0(n40_adj_4690), .I1(n36_adj_4688), .I2(n41_adj_4532), 
            .I3(n67786), .O(n69742));   // verilog/uart_rx.v(119[33:55])
    defparam i54048_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i54049_3_lut (.I0(n69742), .I1(baudrate[5]), .I2(n1263), .I3(GND_net), 
            .O(n69743));   // verilog/uart_rx.v(119[33:55])
    defparam i54049_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i53914_3_lut (.I0(n69743), .I1(baudrate[6]), .I2(n1262), .I3(GND_net), 
            .O(n69608));   // verilog/uart_rx.v(119[33:55])
    defparam i53914_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i52755_3_lut (.I0(n69608), .I1(baudrate[7]), .I2(n1261), .I3(GND_net), 
            .O(n48_adj_4691));   // verilog/uart_rx.v(119[33:55])
    defparam i52755_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i54990_4_lut_4_lut (.I0(\r_SM_Main_2__N_3446[1] ), .I1(\r_SM_Main[1] ), 
            .I2(n6_adj_4692), .I3(n61449), .O(n59702));
    defparam i54990_4_lut_4_lut.LUT_INIT = 16'h0703;
    SB_LUT4 i1_2_lut_adj_1024 (.I0(n62037), .I1(n48_adj_4691), .I2(GND_net), 
            .I3(GND_net), .O(n1415));
    defparam i1_2_lut_adj_1024.LUT_INIT = 16'h2222;
    SB_LUT4 div_37_i1046_3_lut (.I0(n1415), .I1(n8053[16]), .I2(n294[15]), 
            .I3(GND_net), .O(n1559));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1046_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1141_3_lut (.I0(n1559), .I1(n8079[16]), .I2(n294[14]), 
            .I3(GND_net), .O(n1700));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1141_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1234_3_lut (.I0(n1700), .I1(n8105[16]), .I2(n294[13]), 
            .I3(GND_net), .O(n1838));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1234_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1325_3_lut (.I0(n1838), .I1(n8131[16]), .I2(n294[12]), 
            .I3(GND_net), .O(n1973));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1325_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1414_3_lut (.I0(n1973), .I1(n8157[16]), .I2(n294[11]), 
            .I3(GND_net), .O(n2105));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1414_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1501_3_lut (.I0(n2105), .I1(n8183[16]), .I2(n294[10]), 
            .I3(GND_net), .O(n2234));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1501_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1586_3_lut (.I0(n2234), .I1(n8209[16]), .I2(n294[9]), 
            .I3(GND_net), .O(n2360));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1586_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1602_i33_2_lut (.I0(n2360), .I1(baudrate[8]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_4693));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1602_i31_2_lut (.I0(n2361), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_4694));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1602_i21_2_lut (.I0(n2366), .I1(baudrate[2]), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_4695));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i51957_4_lut (.I0(n27_adj_4533), .I1(n25_adj_4674), .I2(n23_adj_4660), 
            .I3(n21_adj_4695), .O(n67651));
    defparam i51957_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i51951_4_lut (.I0(n33_adj_4693), .I1(n31_adj_4694), .I2(n29_adj_4534), 
            .I3(n67651), .O(n67645));
    defparam i51951_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_37_LessThan_1602_i28_3_lut (.I0(n26_adj_4696), .I1(baudrate[7]), 
            .I2(n31_adj_4694), .I3(GND_net), .O(n28_adj_4697));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i28_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1602_i32_3_lut (.I0(n24_adj_4698), .I1(baudrate[9]), 
            .I2(n35_adj_4665), .I3(GND_net), .O(n32_adj_4699));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i32_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i54062_4_lut (.I0(n32_adj_4699), .I1(n22_adj_4700), .I2(n35_adj_4665), 
            .I3(n67642), .O(n69756));   // verilog/uart_rx.v(119[33:55])
    defparam i54062_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i54063_3_lut (.I0(n69756), .I1(baudrate[10]), .I2(n37_adj_4653), 
            .I3(GND_net), .O(n69757));   // verilog/uart_rx.v(119[33:55])
    defparam i54063_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53876_3_lut (.I0(n69757), .I1(baudrate[11]), .I2(n39_adj_4659), 
            .I3(GND_net), .O(n69570));   // verilog/uart_rx.v(119[33:55])
    defparam i53876_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53738_4_lut (.I0(n39_adj_4659), .I1(n37_adj_4653), .I2(n35_adj_4665), 
            .I3(n67645), .O(n69432));
    defparam i53738_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i54135_4_lut (.I0(n28_adj_4697), .I1(n20_adj_4701), .I2(n31_adj_4694), 
            .I3(n67649), .O(n69829));   // verilog/uart_rx.v(119[33:55])
    defparam i54135_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i52805_3_lut (.I0(n69570), .I1(baudrate[12]), .I2(n41_adj_4650), 
            .I3(GND_net), .O(n68499));   // verilog/uart_rx.v(119[33:55])
    defparam i52805_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i54228_4_lut (.I0(n68499), .I1(n69829), .I2(n41_adj_4650), 
            .I3(n69432), .O(n69922));   // verilog/uart_rx.v(119[33:55])
    defparam i54228_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i54229_3_lut (.I0(n69922), .I1(baudrate[13]), .I2(n2355), 
            .I3(GND_net), .O(n69923));   // verilog/uart_rx.v(119[33:55])
    defparam i54229_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i54194_3_lut (.I0(n69923), .I1(baudrate[14]), .I2(n2354), 
            .I3(GND_net), .O(n69888));   // verilog/uart_rx.v(119[33:55])
    defparam i54194_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i54115_3_lut (.I0(n69888), .I1(baudrate[15]), .I2(n2353), 
            .I3(GND_net), .O(n48_adj_4566));   // verilog/uart_rx.v(119[33:55])
    defparam i54115_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_i1591_3_lut (.I0(n2239), .I1(n8209[11]), .I2(n294[9]), 
            .I3(GND_net), .O(n2365));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1591_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1674_3_lut (.I0(n2365), .I1(n8235[11]), .I2(n294[8]), 
            .I3(GND_net), .O(n2488));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1674_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1755_3_lut (.I0(n2488), .I1(n8261[11]), .I2(n294[7]), 
            .I3(GND_net), .O(n2608));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1755_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1766_i23_2_lut (.I0(n2608), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_4702));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1766_i25_2_lut (.I0(n2607), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_4703));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1025 (.I0(baudrate[18]), .I1(baudrate[19]), .I2(GND_net), 
            .I3(GND_net), .O(n63509));
    defparam i1_2_lut_adj_1025.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_1026 (.I0(n63519), .I1(n62017), .I2(n62015), 
            .I3(n63509), .O(n25574));
    defparam i1_4_lut_adj_1026.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_LessThan_1766_i17_2_lut (.I0(n2611), .I1(baudrate[2]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_4704));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i51877_4_lut (.I0(n23_adj_4702), .I1(n21_adj_4590), .I2(n19_adj_4589), 
            .I3(n17_adj_4704), .O(n67571));
    defparam i51877_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i51872_4_lut (.I0(n29_adj_4588), .I1(n27_adj_4587), .I2(n25_adj_4703), 
            .I3(n67571), .O(n67566));
    defparam i51872_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i53647_4_lut (.I0(n35_adj_4586), .I1(n33_adj_4585), .I2(n31_adj_4584), 
            .I3(n67566), .O(n69341));
    defparam i53647_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_LessThan_1766_i16_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n2612), .I3(GND_net), .O(n16_adj_4705));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i16_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i53826_3_lut (.I0(n16_adj_4705), .I1(baudrate[13]), .I2(n39_adj_4583), 
            .I3(GND_net), .O(n69520));   // verilog/uart_rx.v(119[33:55])
    defparam i53826_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53827_3_lut (.I0(n69520), .I1(baudrate[14]), .I2(n41_adj_4582), 
            .I3(GND_net), .O(n69521));   // verilog/uart_rx.v(119[33:55])
    defparam i53827_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52745_4_lut (.I0(n41_adj_4582), .I1(n39_adj_4583), .I2(n27_adj_4587), 
            .I3(n67569), .O(n68439));
    defparam i52745_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i53337_3_lut (.I0(n22_adj_4706), .I1(baudrate[7]), .I2(n27_adj_4587), 
            .I3(GND_net), .O(n69031));   // verilog/uart_rx.v(119[33:55])
    defparam i53337_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53680_3_lut (.I0(n69521), .I1(baudrate[15]), .I2(n43_adj_4581), 
            .I3(GND_net), .O(n69374));   // verilog/uart_rx.v(119[33:55])
    defparam i53680_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1766_i28_3_lut (.I0(n20_adj_4707), .I1(baudrate[9]), 
            .I2(n31_adj_4584), .I3(GND_net), .O(n28_adj_4708));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i28_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i54183_4_lut (.I0(n28_adj_4708), .I1(n18_adj_4709), .I2(n31_adj_4584), 
            .I3(n67564), .O(n69877));   // verilog/uart_rx.v(119[33:55])
    defparam i54183_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i54184_3_lut (.I0(n69877), .I1(baudrate[10]), .I2(n33_adj_4585), 
            .I3(GND_net), .O(n69878));   // verilog/uart_rx.v(119[33:55])
    defparam i54184_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i54117_3_lut (.I0(n69878), .I1(baudrate[11]), .I2(n35_adj_4586), 
            .I3(GND_net), .O(n69811));   // verilog/uart_rx.v(119[33:55])
    defparam i54117_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52748_4_lut (.I0(n41_adj_4582), .I1(n39_adj_4583), .I2(n37_adj_4580), 
            .I3(n69341), .O(n68442));
    defparam i52748_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i53824_4_lut (.I0(n69374), .I1(n69031), .I2(n43_adj_4581), 
            .I3(n68439), .O(n69518));   // verilog/uart_rx.v(119[33:55])
    defparam i53824_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i53958_3_lut (.I0(n69811), .I1(baudrate[12]), .I2(n37_adj_4580), 
            .I3(GND_net), .O(n69652));   // verilog/uart_rx.v(119[33:55])
    defparam i53958_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i54155_4_lut (.I0(n69652), .I1(n69518), .I2(n43_adj_4581), 
            .I3(n68442), .O(n69849));   // verilog/uart_rx.v(119[33:55])
    defparam i54155_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i54156_3_lut (.I0(n69849), .I1(baudrate[16]), .I2(n2597), 
            .I3(GND_net), .O(n69850));   // verilog/uart_rx.v(119[33:55])
    defparam i54156_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_1922_i14_3_lut_3_lut (.I0(baudrate[2]), .I1(baudrate[3]), 
            .I2(n2843), .I3(GND_net), .O(n14_adj_4710));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i14_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i51789_2_lut_4_lut (.I0(n2838), .I1(baudrate[8]), .I2(n2842), 
            .I3(baudrate[4]), .O(n67483));
    defparam i51789_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_1922_i16_3_lut_3_lut (.I0(baudrate[4]), .I1(baudrate[8]), 
            .I2(n2838), .I3(GND_net), .O(n16_adj_4711));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i16_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_i1754_3_lut (.I0(n2487), .I1(n8261[12]), .I2(n294[7]), 
            .I3(GND_net), .O(n2607));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1754_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1922_i18_3_lut_3_lut (.I0(baudrate[5]), .I1(baudrate[6]), 
            .I2(n2840), .I3(GND_net), .O(n18_adj_4712));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i18_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i51758_2_lut_4_lut (.I0(n2830), .I1(baudrate[16]), .I2(n2839), 
            .I3(baudrate[7]), .O(n67452));
    defparam i51758_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_i1833_3_lut (.I0(n2607), .I1(n8287[12]), .I2(n294[6]), 
            .I3(GND_net), .O(n2724));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1833_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1835_3_lut (.I0(n2609), .I1(n8287[10]), .I2(n294[6]), 
            .I3(GND_net), .O(n2726));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1835_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1845_i21_2_lut (.I0(n2726), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_4713));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1845_i23_2_lut (.I0(n2725), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_4714));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1845_i25_2_lut (.I0(n2724), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_4715));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1922_i20_3_lut_3_lut (.I0(baudrate[7]), .I1(baudrate[16]), 
            .I2(n2830), .I3(GND_net), .O(n20_adj_4716));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i20_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i1_2_lut_4_lut_adj_1027 (.I0(baudrate[20]), .I1(baudrate[21]), 
            .I2(baudrate[22]), .I3(baudrate[23]), .O(n63519));
    defparam i1_2_lut_4_lut_adj_1027.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_LessThan_1845_i16_3_lut_3_lut (.I0(baudrate[2]), .I1(baudrate[3]), 
            .I2(n2728), .I3(GND_net), .O(n16_adj_4717));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i16_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i51842_2_lut_4_lut (.I0(n2723), .I1(baudrate[8]), .I2(n2727), 
            .I3(baudrate[4]), .O(n67536));
    defparam i51842_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_1845_i18_3_lut_3_lut (.I0(baudrate[4]), .I1(baudrate[8]), 
            .I2(n2723), .I3(GND_net), .O(n18_adj_4718));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i18_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_1845_i37_2_lut (.I0(n2718), .I1(baudrate[13]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_4719));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1845_i20_3_lut_3_lut (.I0(baudrate[5]), .I1(baudrate[6]), 
            .I2(n2725), .I3(GND_net), .O(n20_adj_4720));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i20_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i1_2_lut_adj_1028 (.I0(baudrate[28]), .I1(baudrate[25]), .I2(GND_net), 
            .I3(GND_net), .O(n62569));
    defparam i1_2_lut_adj_1028.LUT_INIT = 16'heeee;
    SB_LUT4 i51818_2_lut_4_lut (.I0(n2715), .I1(baudrate[16]), .I2(n2724), 
            .I3(baudrate[7]), .O(n67512));
    defparam i51818_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_1845_i22_3_lut_3_lut (.I0(baudrate[7]), .I1(baudrate[16]), 
            .I2(n2715), .I3(GND_net), .O(n22_adj_4721));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i22_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i1_2_lut_adj_1029 (.I0(baudrate[27]), .I1(baudrate[30]), .I2(GND_net), 
            .I3(GND_net), .O(n63391));
    defparam i1_2_lut_adj_1029.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_1030 (.I0(baudrate[31]), .I1(baudrate[26]), .I2(GND_net), 
            .I3(GND_net), .O(n63465));
    defparam i1_2_lut_adj_1030.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_1031 (.I0(n63505), .I1(n63391), .I2(n62569), 
            .I3(baudrate[19]), .O(n62589));
    defparam i1_4_lut_adj_1031.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1032 (.I0(n62589), .I1(n63465), .I2(n63507), 
            .I3(n63463), .O(n25577));
    defparam i1_4_lut_adj_1032.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_LessThan_1766_i18_3_lut_3_lut (.I0(baudrate[2]), .I1(baudrate[3]), 
            .I2(n2610), .I3(GND_net), .O(n18_adj_4709));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i18_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i51827_4_lut (.I0(n37_adj_4719), .I1(n25_adj_4715), .I2(n23_adj_4714), 
            .I3(n21_adj_4713), .O(n67521));
    defparam i51827_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i51870_2_lut_4_lut (.I0(n2605), .I1(baudrate[8]), .I2(n2609), 
            .I3(baudrate[4]), .O(n67564));
    defparam i51870_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_1766_i20_3_lut_3_lut (.I0(baudrate[4]), .I1(baudrate[8]), 
            .I2(n2605), .I3(GND_net), .O(n20_adj_4707));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i20_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_1766_i22_3_lut_3_lut (.I0(baudrate[5]), .I1(baudrate[6]), 
            .I2(n2607), .I3(GND_net), .O(n22_adj_4706));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i22_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i52738_4_lut (.I0(n19_adj_4577), .I1(n17_adj_4576), .I2(n2729), 
            .I3(baudrate[2]), .O(n68432));
    defparam i52738_4_lut.LUT_INIT = 16'heffe;
    SB_LUT4 i53318_4_lut (.I0(n25_adj_4715), .I1(n23_adj_4714), .I2(n21_adj_4713), 
            .I3(n68432), .O(n69012));
    defparam i53318_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i53316_4_lut (.I0(n31_adj_4574), .I1(n29_adj_4573), .I2(n27_adj_4572), 
            .I3(n69012), .O(n69010));
    defparam i53316_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i51832_4_lut (.I0(n37_adj_4719), .I1(n35_adj_4579), .I2(n33_adj_4578), 
            .I3(n69010), .O(n67526));
    defparam i51832_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_37_LessThan_1845_i14_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n2730), .I3(GND_net), .O(n14_adj_4722));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i14_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i53820_3_lut (.I0(n14_adj_4722), .I1(baudrate[13]), .I2(n37_adj_4719), 
            .I3(GND_net), .O(n69514));   // verilog/uart_rx.v(119[33:55])
    defparam i53820_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53821_3_lut (.I0(n69514), .I1(baudrate[14]), .I2(n39_adj_4575), 
            .I3(GND_net), .O(n69515));   // verilog/uart_rx.v(119[33:55])
    defparam i53821_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1845_i40_3_lut (.I0(n22_adj_4721), .I1(baudrate[17]), 
            .I2(n45_adj_4570), .I3(GND_net), .O(n40_adj_4723));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i40_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51821_4_lut (.I0(n43_adj_4571), .I1(n41_adj_4569), .I2(n39_adj_4575), 
            .I3(n67521), .O(n67515));
    defparam i51821_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i51875_2_lut_4_lut (.I0(n2607), .I1(baudrate[6]), .I2(n2608), 
            .I3(baudrate[5]), .O(n67569));
    defparam i51875_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i53339_4_lut (.I0(n40_adj_4723), .I1(n20_adj_4720), .I2(n45_adj_4570), 
            .I3(n67512), .O(n69033));   // verilog/uart_rx.v(119[33:55])
    defparam i53339_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i53687_3_lut (.I0(n69515), .I1(baudrate[15]), .I2(n41_adj_4569), 
            .I3(GND_net), .O(n69381));   // verilog/uart_rx.v(119[33:55])
    defparam i53687_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut_4_lut_adj_1033 (.I0(baudrate[28]), .I1(baudrate[25]), 
            .I2(baudrate[26]), .I3(baudrate[29]), .O(n62017));
    defparam i1_3_lut_4_lut_adj_1033.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_LessThan_1845_i26_3_lut (.I0(n18_adj_4718), .I1(baudrate[9]), 
            .I2(n29_adj_4573), .I3(GND_net), .O(n26_adj_4724));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i26_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i54137_4_lut (.I0(n26_adj_4724), .I1(n16_adj_4717), .I2(n29_adj_4573), 
            .I3(n67536), .O(n69831));   // verilog/uart_rx.v(119[33:55])
    defparam i54137_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i54138_3_lut (.I0(n69831), .I1(baudrate[10]), .I2(n31_adj_4574), 
            .I3(GND_net), .O(n69832));   // verilog/uart_rx.v(119[33:55])
    defparam i54138_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i54025_3_lut (.I0(n69832), .I1(baudrate[11]), .I2(n33_adj_4578), 
            .I3(GND_net), .O(n69719));   // verilog/uart_rx.v(119[33:55])
    defparam i54025_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53617_4_lut (.I0(n43_adj_4571), .I1(n41_adj_4569), .I2(n39_adj_4575), 
            .I3(n67526), .O(n69311));
    defparam i53617_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i53961_4_lut (.I0(n69381), .I1(n69033), .I2(n45_adj_4570), 
            .I3(n67515), .O(n69655));   // verilog/uart_rx.v(119[33:55])
    defparam i53961_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i53960_3_lut (.I0(n69719), .I1(baudrate[12]), .I2(n35_adj_4579), 
            .I3(GND_net), .O(n69654));   // verilog/uart_rx.v(119[33:55])
    defparam i53960_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53963_4_lut (.I0(n69654), .I1(n69655), .I2(n45_adj_4570), 
            .I3(n69311), .O(n69657));   // verilog/uart_rx.v(119[33:55])
    defparam i53963_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 div_37_i1834_3_lut (.I0(n2608), .I1(n8287[11]), .I2(n294[6]), 
            .I3(GND_net), .O(n2725));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1834_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1911_3_lut (.I0(n2725), .I1(n8313[11]), .I2(n294[5]), 
            .I3(GND_net), .O(n2839));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1911_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1913_3_lut (.I0(n2727), .I1(n8313[9]), .I2(n294[5]), 
            .I3(GND_net), .O(n2841));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1913_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1922_i19_2_lut (.I0(n2841), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_4725));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1922_i21_2_lut (.I0(n2840), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_4726));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1922_i23_2_lut (.I0(n2839), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_4727));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1922_i35_2_lut (.I0(n2833), .I1(baudrate[13]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_4728));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1034 (.I0(baudrate[22]), .I1(baudrate[23]), .I2(GND_net), 
            .I3(GND_net), .O(n63505));
    defparam i1_2_lut_adj_1034.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_1035 (.I0(baudrate[20]), .I1(baudrate[21]), .I2(GND_net), 
            .I3(GND_net), .O(n63507));
    defparam i1_2_lut_adj_1035.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_1036 (.I0(baudrate[30]), .I1(baudrate[25]), .I2(GND_net), 
            .I3(GND_net), .O(n63459));
    defparam i1_2_lut_adj_1036.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_1037 (.I0(baudrate[29]), .I1(baudrate[24]), .I2(GND_net), 
            .I3(GND_net), .O(n63463));
    defparam i1_2_lut_adj_1037.LUT_INIT = 16'heeee;
    SB_LUT4 div_37_LessThan_1602_i22_3_lut_3_lut (.I0(baudrate[2]), .I1(baudrate[3]), 
            .I2(n2365), .I3(GND_net), .O(n22_adj_4700));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i22_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i1_4_lut_adj_1038 (.I0(baudrate[28]), .I1(baudrate[27]), .I2(baudrate[31]), 
            .I3(baudrate[26]), .O(n62711));
    defparam i1_4_lut_adj_1038.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1039 (.I0(n62711), .I1(n63519), .I2(n63463), 
            .I3(n63459), .O(n25580));
    defparam i1_4_lut_adj_1039.LUT_INIT = 16'hfffe;
    SB_LUT4 i51770_4_lut (.I0(n35_adj_4728), .I1(n23_adj_4727), .I2(n21_adj_4726), 
            .I3(n19_adj_4725), .O(n67464));
    defparam i51770_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i52704_4_lut (.I0(n17_adj_4568), .I1(n15_adj_4567), .I2(n2844), 
            .I3(baudrate[2]), .O(n68398));
    defparam i52704_4_lut.LUT_INIT = 16'heffe;
    SB_LUT4 i51948_2_lut_4_lut (.I0(n2360), .I1(baudrate[8]), .I2(n2364), 
            .I3(baudrate[4]), .O(n67642));
    defparam i51948_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_1602_i24_3_lut_3_lut (.I0(baudrate[4]), .I1(baudrate[8]), 
            .I2(n2360), .I3(GND_net), .O(n24_adj_4698));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i24_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_1602_i20_3_lut_4_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n62043), .I3(n48_adj_4685), .O(n20_adj_4701));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i20_3_lut_4_lut.LUT_INIT = 16'hee8e;
    SB_LUT4 i51955_2_lut_4_lut (.I0(n2362), .I1(baudrate[6]), .I2(n2363), 
            .I3(baudrate[5]), .O(n67649));
    defparam i51955_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_1602_i26_3_lut_3_lut (.I0(baudrate[5]), .I1(baudrate[6]), 
            .I2(n2362), .I3(GND_net), .O(n26_adj_4696));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i26_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i53300_4_lut (.I0(n23_adj_4727), .I1(n21_adj_4726), .I2(n19_adj_4725), 
            .I3(n68398), .O(n68994));
    defparam i53300_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i53290_4_lut (.I0(n29_adj_4565), .I1(n27_adj_4564), .I2(n25_adj_4563), 
            .I3(n68994), .O(n68984));
    defparam i53290_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i51775_4_lut (.I0(n35_adj_4728), .I1(n33_adj_4562), .I2(n31_adj_4561), 
            .I3(n68984), .O(n67469));
    defparam i51775_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_37_LessThan_1922_i12_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n2845), .I3(GND_net), .O(n12_adj_4729));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i12_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i53816_3_lut (.I0(n12_adj_4729), .I1(baudrate[13]), .I2(n35_adj_4728), 
            .I3(GND_net), .O(n69510));   // verilog/uart_rx.v(119[33:55])
    defparam i53816_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1922_i38_3_lut (.I0(n20_adj_4716), .I1(baudrate[17]), 
            .I2(n43_adj_4558), .I3(GND_net), .O(n38_adj_4730));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i38_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53817_3_lut (.I0(n69510), .I1(baudrate[14]), .I2(n37_adj_4557), 
            .I3(GND_net), .O(n69511));   // verilog/uart_rx.v(119[33:55])
    defparam i53817_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51762_4_lut (.I0(n41_adj_4560), .I1(n39_adj_4555), .I2(n37_adj_4557), 
            .I3(n67464), .O(n67456));
    defparam i51762_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i53814_4_lut (.I0(n38_adj_4730), .I1(n18_adj_4712), .I2(n43_adj_4558), 
            .I3(n67452), .O(n69508));   // verilog/uart_rx.v(119[33:55])
    defparam i53814_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i53691_3_lut (.I0(n69511), .I1(baudrate[15]), .I2(n39_adj_4555), 
            .I3(GND_net), .O(n69385));   // verilog/uart_rx.v(119[33:55])
    defparam i53691_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i54619_2_lut_4_lut (.I0(n69866), .I1(baudrate[13]), .I2(n2098), 
            .I3(n25562), .O(n294[10]));   // verilog/uart_rx.v(119[33:55])
    defparam i54619_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_LUT4 div_37_LessThan_1922_i24_3_lut (.I0(n16_adj_4711), .I1(baudrate[9]), 
            .I2(n27_adj_4564), .I3(GND_net), .O(n24_adj_4731));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i54139_4_lut (.I0(n24_adj_4731), .I1(n14_adj_4710), .I2(n27_adj_4564), 
            .I3(n67483), .O(n69833));   // verilog/uart_rx.v(119[33:55])
    defparam i54139_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i54140_3_lut (.I0(n69833), .I1(baudrate[10]), .I2(n29_adj_4565), 
            .I3(GND_net), .O(n69834));   // verilog/uart_rx.v(119[33:55])
    defparam i54140_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i54023_3_lut (.I0(n69834), .I1(baudrate[11]), .I2(n31_adj_4561), 
            .I3(GND_net), .O(n69717));   // verilog/uart_rx.v(119[33:55])
    defparam i54023_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i55115_2_lut_4_lut (.I0(n69870), .I1(baudrate[12]), .I2(n1966), 
            .I3(n64194), .O(n294[11]));
    defparam i55115_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_LUT4 i53609_4_lut (.I0(n41_adj_4560), .I1(n39_adj_4555), .I2(n37_adj_4557), 
            .I3(n67469), .O(n69303));
    defparam i53609_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i54616_2_lut_4_lut (.I0(n69600), .I1(baudrate[10]), .I2(n1693), 
            .I3(n25553), .O(n294[13]));   // verilog/uart_rx.v(119[33:55])
    defparam i54616_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_LUT4 i54127_4_lut (.I0(n69385), .I1(n69508), .I2(n43_adj_4558), 
            .I3(n67456), .O(n69821));   // verilog/uart_rx.v(119[33:55])
    defparam i54127_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i53965_3_lut (.I0(n69717), .I1(baudrate[12]), .I2(n33_adj_4562), 
            .I3(GND_net), .O(n69659));   // verilog/uart_rx.v(119[33:55])
    defparam i53965_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i54282_4_lut (.I0(n69659), .I1(n69821), .I2(n43_adj_4558), 
            .I3(n69303), .O(n69976));   // verilog/uart_rx.v(119[33:55])
    defparam i54282_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i54283_3_lut (.I0(n69976), .I1(baudrate[18]), .I2(n2828), 
            .I3(GND_net), .O(n69977));   // verilog/uart_rx.v(119[33:55])
    defparam i54283_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i55109_2_lut_4_lut (.I0(n69604), .I1(baudrate[9]), .I2(n1552), 
            .I3(n64228), .O(n294[14]));
    defparam i55109_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_LUT4 i54355_2_lut_3_lut_4_lut (.I0(\r_SM_Main_2__N_3446[1] ), .I1(\r_SM_Main[1] ), 
            .I2(r_SM_Main[0]), .I3(\r_SM_Main[2] ), .O(n27901));
    defparam i54355_2_lut_3_lut_4_lut.LUT_INIT = 16'h0007;
    SB_LUT4 div_37_i1909_3_lut (.I0(n2723), .I1(n8313[13]), .I2(n294[5]), 
            .I3(GND_net), .O(n2837));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1909_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1984_3_lut (.I0(n2837), .I1(n8339[13]), .I2(n294[4]), 
            .I3(GND_net), .O(n2948));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1984_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i44144_1_lut (.I0(n25586), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n59790));
    defparam i44144_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_3_lut_4_lut_adj_1040 (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(\r_Bit_Index[0] ), .I3(n4_adj_4559), .O(n62497));   // verilog/uart_rx.v(98[17:39])
    defparam i1_3_lut_4_lut_adj_1040.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_i2164_1_lut (.I0(baudrate[11]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2144));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2164_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i2057_3_lut (.I0(n2948), .I1(n8365[13]), .I2(n294[3]), 
            .I3(GND_net), .O(n3056));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2057_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut_4_lut_adj_1041 (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(\r_Bit_Index[0] ), .I3(n4_adj_4559), .O(n62449));   // verilog/uart_rx.v(98[17:39])
    defparam i1_3_lut_4_lut_adj_1041.LUT_INIT = 16'hffef;
    SB_LUT4 i1_2_lut_4_lut_adj_1042 (.I0(baudrate[12]), .I1(baudrate[13]), 
            .I2(baudrate[14]), .I3(baudrate[15]), .O(n62687));
    defparam i1_2_lut_4_lut_adj_1042.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_LessThan_866_i38_3_lut_3_lut (.I0(n1265), .I1(baudrate[3]), 
            .I2(baudrate[2]), .I3(GND_net), .O(n38_adj_4689));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_866_i38_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 i52092_3_lut_4_lut (.I0(n1265), .I1(baudrate[3]), .I2(baudrate[2]), 
            .I3(n1266), .O(n67786));   // verilog/uart_rx.v(119[33:55])
    defparam i52092_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_765_i40_3_lut_3_lut (.I0(n1114), .I1(baudrate[3]), 
            .I2(baudrate[2]), .I3(GND_net), .O(n40_adj_4663));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_765_i40_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 i52102_3_lut_4_lut (.I0(n1114), .I1(baudrate[3]), .I2(baudrate[2]), 
            .I3(n1115), .O(n67796));   // verilog/uart_rx.v(119[33:55])
    defparam i52102_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_1517_i24_3_lut_3_lut (.I0(baudrate[2]), .I1(baudrate[3]), 
            .I2(n2238), .I3(GND_net), .O(n24_adj_4684));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i24_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i51981_2_lut_4_lut (.I0(n2233), .I1(baudrate[8]), .I2(n2237), 
            .I3(baudrate[4]), .O(n67675));
    defparam i51981_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_1517_i26_3_lut_3_lut (.I0(baudrate[4]), .I1(baudrate[8]), 
            .I2(n2233), .I3(GND_net), .O(n26_adj_4682));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i26_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i51987_2_lut_4_lut (.I0(n2235), .I1(baudrate[6]), .I2(n2236), 
            .I3(baudrate[5]), .O(n67681));
    defparam i51987_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_1517_i28_3_lut_3_lut (.I0(baudrate[5]), .I1(baudrate[6]), 
            .I2(n2235), .I3(GND_net), .O(n28_adj_4680));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i28_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i5574_2_lut_4_lut (.I0(n804), .I1(n43066), .I2(n20902), .I3(baudrate[2]), 
            .O(n44_adj_4676));   // verilog/uart_rx.v(119[33:55])
    defparam i5574_2_lut_4_lut.LUT_INIT = 16'ha2fb;
    SB_LUT4 i52333_4_lut (.I0(\o_Rx_DV_N_3488[8] ), .I1(\o_Rx_DV_N_3488[12] ), 
            .I2(n4935), .I3(n58684), .O(n67033));
    defparam i52333_4_lut.LUT_INIT = 16'h0100;
    SB_LUT4 i52328_4_lut (.I0(n67033), .I1(\o_Rx_DV_N_3488[24] ), .I2(n29), 
            .I3(n23), .O(n67030));
    defparam i52328_4_lut.LUT_INIT = 16'h0002;
    SB_LUT4 i14_4_lut (.I0(\r_SM_Main[1] ), .I1(n67030), .I2(r_SM_Main[0]), 
            .I3(n27), .O(n27661));
    defparam i14_4_lut.LUT_INIT = 16'h05c5;
    SB_LUT4 i52073_3_lut_4_lut (.I0(n1558), .I1(baudrate[3]), .I2(baudrate[2]), 
            .I3(n1559), .O(n67767));   // verilog/uart_rx.v(119[33:55])
    defparam i52073_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_1062_i34_3_lut_3_lut (.I0(n1558), .I1(baudrate[3]), 
            .I2(baudrate[2]), .I3(GND_net), .O(n34_adj_4632));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1062_i34_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 i1_2_lut_4_lut_adj_1043 (.I0(n69404), .I1(baudrate[21]), .I2(n3046), 
            .I3(n62057), .O(n3172));   // verilog/uart_rx.v(119[33:55])
    defparam i1_2_lut_4_lut_adj_1043.LUT_INIT = 16'h7100;
    SB_LUT4 i55149_2_lut_4_lut (.I0(n69404), .I1(baudrate[21]), .I2(n3046), 
            .I3(n25586), .O(n294[2]));   // verilog/uart_rx.v(119[33:55])
    defparam i55149_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_LUT4 i1_3_lut_4_lut_adj_1044 (.I0(n25598), .I1(n48_adj_4654), .I2(baudrate[1]), 
            .I3(baudrate[0]), .O(n44_adj_4675));
    defparam i1_3_lut_4_lut_adj_1044.LUT_INIT = 16'hefff;
    SB_LUT4 i51684_2_lut_3_lut (.I0(baudrate[1]), .I1(n48_adj_4654), .I2(n25598), 
            .I3(GND_net), .O(n67378));   // verilog/uart_rx.v(119[33:55])
    defparam i51684_2_lut_3_lut.LUT_INIT = 16'h0202;
    SB_LUT4 div_37_LessThan_1250_i30_3_lut_3_lut (.I0(baudrate[2]), .I1(baudrate[3]), 
            .I2(n1839), .I3(GND_net), .O(n30_adj_4673));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1250_i30_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i52045_2_lut_4_lut (.I0(n1834), .I1(baudrate[8]), .I2(n1838), 
            .I3(baudrate[4]), .O(n67739));
    defparam i52045_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_1250_i32_3_lut_3_lut (.I0(baudrate[4]), .I1(baudrate[8]), 
            .I2(n1834), .I3(GND_net), .O(n32_adj_4670));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1250_i32_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i51688_2_lut_3_lut (.I0(baudrate[1]), .I1(n48_adj_4655), .I2(n25608), 
            .I3(GND_net), .O(n67382));   // verilog/uart_rx.v(119[33:55])
    defparam i51688_2_lut_3_lut.LUT_INIT = 16'h0202;
    SB_LUT4 i5567_2_lut_3_lut (.I0(n20902), .I1(baudrate[1]), .I2(baudrate[0]), 
            .I3(GND_net), .O(n42_adj_4667));   // verilog/uart_rx.v(119[33:55])
    defparam i5567_2_lut_3_lut.LUT_INIT = 16'habab;
    SB_LUT4 i52349_2_lut (.I0(n58444), .I1(r_Rx_Data), .I2(GND_net), .I3(GND_net), 
            .O(n67056));
    defparam i52349_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i52346_4_lut (.I0(n67056), .I1(n29), .I2(n23), .I3(\o_Rx_DV_N_3488[12] ), 
            .O(n67053));
    defparam i52346_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i51665_4_lut (.I0(n67053), .I1(r_SM_Main[0]), .I2(n27), .I3(\o_Rx_DV_N_3488[24] ), 
            .O(n67050));
    defparam i51665_4_lut.LUT_INIT = 16'hccc8;
    SB_LUT4 i54741_4_lut (.I0(\r_SM_Main[2] ), .I1(n67050), .I2(\r_SM_Main_2__N_3446[1] ), 
            .I3(\r_SM_Main[1] ), .O(n29076));
    defparam i54741_4_lut.LUT_INIT = 16'h0511;
    SB_LUT4 i1_4_lut_adj_1045 (.I0(n58444), .I1(\r_SM_Main[1] ), .I2(r_Rx_Data), 
            .I3(r_SM_Main[0]), .O(n62117));
    defparam i1_4_lut_adj_1045.LUT_INIT = 16'h1000;
    SB_LUT4 i1_4_lut_adj_1046 (.I0(n29), .I1(n23), .I2(\o_Rx_DV_N_3488[12] ), 
            .I3(n62117), .O(n62123));
    defparam i1_4_lut_adj_1046.LUT_INIT = 16'h0100;
    SB_LUT4 i54358_4_lut (.I0(\r_SM_Main[2] ), .I1(\o_Rx_DV_N_3488[24] ), 
            .I2(n27), .I3(n62123), .O(n27701));   // verilog/uart_rx.v(53[7] 144[14])
    defparam i54358_4_lut.LUT_INIT = 16'h5455;
    SB_LUT4 i48505_2_lut_3_lut_4_lut (.I0(baudrate[28]), .I1(baudrate[26]), 
            .I2(baudrate[29]), .I3(baudrate[24]), .O(n64190));
    defparam i48505_2_lut_3_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_3_lut_4_lut (.I0(baudrate[28]), .I1(baudrate[26]), 
            .I2(baudrate[24]), .I3(baudrate[31]), .O(n63401));
    defparam i1_2_lut_3_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i5745_2_lut_4_lut (.I0(n960), .I1(n11417), .I2(n20912), .I3(baudrate[3]), 
            .O(n44_adj_4677));   // verilog/uart_rx.v(119[33:55])
    defparam i5745_2_lut_4_lut.LUT_INIT = 16'ha8fe;
    SB_LUT4 i52353_3_lut_4_lut (.I0(n962), .I1(baudrate[1]), .I2(n48_adj_4652), 
            .I3(n25605), .O(n1115));
    defparam i52353_3_lut_4_lut.LUT_INIT = 16'haaa6;
    SB_LUT4 i52323_2_lut_3_lut (.I0(n25598), .I1(baudrate[1]), .I2(baudrate[0]), 
            .I3(GND_net), .O(n67096));   // verilog/uart_rx.v(119[33:55])
    defparam i52323_2_lut_3_lut.LUT_INIT = 16'h4040;
    SB_LUT4 i1_2_lut_4_lut_adj_1047 (.I0(baudrate[16]), .I1(baudrate[17]), 
            .I2(baudrate[18]), .I3(baudrate[19]), .O(n63521));
    defparam i1_2_lut_4_lut_adj_1047.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_4_lut_adj_1048 (.I0(baudrate[6]), .I1(baudrate[7]), 
            .I2(baudrate[8]), .I3(baudrate[9]), .O(n63383));
    defparam i1_2_lut_4_lut_adj_1048.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_4_lut_adj_1049 (.I0(baudrate[10]), .I1(baudrate[11]), 
            .I2(baudrate[12]), .I3(baudrate[13]), .O(n63381));
    defparam i1_2_lut_4_lut_adj_1049.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_LessThan_965_i34_3_lut_4_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n62037), .I3(n48_adj_4691), .O(n34_adj_4646));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_965_i34_3_lut_4_lut.LUT_INIT = 16'hee8e;
    SB_LUT4 div_37_LessThan_1341_i26_3_lut_4_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n62041), .I3(n48_adj_4614), .O(n26_adj_4639));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1341_i26_3_lut_4_lut.LUT_INIT = 16'hee8e;
    SB_LUT4 div_37_LessThan_1341_i28_3_lut_3_lut (.I0(baudrate[2]), .I1(baudrate[3]), 
            .I2(n1975), .I3(GND_net), .O(n28_adj_4640));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1341_i28_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i52025_2_lut_4_lut (.I0(n1970), .I1(baudrate[8]), .I2(n1974), 
            .I3(baudrate[4]), .O(n67719));
    defparam i52025_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_1341_i30_3_lut_3_lut (.I0(baudrate[4]), .I1(baudrate[8]), 
            .I2(n1970), .I3(GND_net), .O(n30_adj_4637));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1341_i30_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i1_2_lut_4_lut_adj_1050 (.I0(baudrate[30]), .I1(baudrate[25]), 
            .I2(baudrate[31]), .I3(baudrate[26]), .O(n63481));
    defparam i1_2_lut_4_lut_adj_1050.LUT_INIT = 16'hfffe;
    SB_LUT4 i48300_1_lut_2_lut (.I0(baudrate[17]), .I1(n25574), .I2(GND_net), 
            .I3(GND_net), .O(n59810));
    defparam i48300_1_lut_2_lut.LUT_INIT = 16'h1111;
    SB_LUT4 div_37_LessThan_1685_i20_3_lut_3_lut (.I0(baudrate[2]), .I1(baudrate[3]), 
            .I2(n2489), .I3(GND_net), .O(n20_adj_4617));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i20_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i51904_2_lut_4_lut (.I0(n2484), .I1(baudrate[8]), .I2(n2488), 
            .I3(baudrate[4]), .O(n67598));
    defparam i51904_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_1685_i22_3_lut_3_lut (.I0(baudrate[4]), .I1(baudrate[8]), 
            .I2(n2484), .I3(GND_net), .O(n22_adj_4615));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i22_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_1685_i24_3_lut_3_lut (.I0(baudrate[5]), .I1(baudrate[6]), 
            .I2(n2486), .I3(GND_net), .O(n24_adj_4611));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i24_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i2158_3_lut (.I0(r_Bit_Index[2]), .I1(r_Bit_Index[1]), .I2(\r_Bit_Index[0] ), 
            .I3(GND_net), .O(n479[2]));   // verilog/uart_rx.v(103[36:51])
    defparam i2158_3_lut.LUT_INIT = 16'h6a6a;
    SB_LUT4 i2_2_lut (.I0(r_SM_Main[0]), .I1(\r_SM_Main[2] ), .I2(GND_net), 
            .I3(GND_net), .O(n6_adj_4692));
    defparam i2_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 div_37_LessThan_1685_i18_3_lut_4_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n62045), .I3(n48_adj_4566), .O(n18_adj_4610));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i18_3_lut_4_lut.LUT_INIT = 16'hee8e;
    SB_LUT4 i51919_2_lut_4_lut (.I0(n2486), .I1(baudrate[6]), .I2(n2487), 
            .I3(baudrate[5]), .O(n67613));
    defparam i51919_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i48543_2_lut_3_lut_4_lut (.I0(baudrate[12]), .I1(n64194), .I2(baudrate[10]), 
            .I3(baudrate[11]), .O(n64228));
    defparam i48543_2_lut_3_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i2151_2_lut (.I0(r_Bit_Index[1]), .I1(\r_Bit_Index[0] ), .I2(GND_net), 
            .I3(GND_net), .O(n479[1]));   // verilog/uart_rx.v(103[36:51])
    defparam i2151_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i48558_1_lut_2_lut (.I0(baudrate[9]), .I1(n64228), .I2(GND_net), 
            .I3(GND_net), .O(n59836));
    defparam i48558_1_lut_2_lut.LUT_INIT = 16'h1111;
    SB_LUT4 div_37_LessThan_1430_i28_3_lut_3_lut (.I0(baudrate[3]), .I1(baudrate[4]), 
            .I2(n2107), .I3(GND_net), .O(n28));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1430_i28_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i52007_2_lut_4_lut (.I0(n2102), .I1(baudrate[9]), .I2(n2106), 
            .I3(baudrate[5]), .O(n67701));
    defparam i52007_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_1430_i30_3_lut_3_lut (.I0(baudrate[5]), .I1(baudrate[9]), 
            .I2(n2102), .I3(GND_net), .O(n30_adj_4597));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1430_i30_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i55100_2_lut_3_lut_4_lut (.I0(baudrate[8]), .I1(baudrate[9]), 
            .I2(n64228), .I3(n48_adj_4691), .O(n294[16]));
    defparam i55100_2_lut_3_lut_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i48561_2_lut_3_lut_4_lut (.I0(baudrate[8]), .I1(baudrate[9]), 
            .I2(n64228), .I3(baudrate[7]), .O(n64246));
    defparam i48561_2_lut_3_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i48560_1_lut_2_lut_3_lut (.I0(baudrate[8]), .I1(baudrate[9]), 
            .I2(n64228), .I3(GND_net), .O(n59840));
    defparam i48560_1_lut_2_lut_3_lut.LUT_INIT = 16'h0101;
    SB_LUT4 i48439_2_lut_4_lut (.I0(baudrate[5]), .I1(baudrate[6]), .I2(baudrate[7]), 
            .I3(baudrate[8]), .O(n64124));
    defparam i48439_2_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i55094_2_lut_3_lut_4_lut (.I0(baudrate[5]), .I1(baudrate[6]), 
            .I2(n64246), .I3(n48_adj_4556), .O(n294[19]));
    defparam i55094_2_lut_3_lut_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 div_37_LessThan_1997_i12_3_lut_3_lut (.I0(baudrate[2]), .I1(baudrate[3]), 
            .I2(n2955), .I3(GND_net), .O(n12_adj_4554));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i12_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i51726_2_lut_4_lut (.I0(n2950), .I1(baudrate[8]), .I2(n2954), 
            .I3(baudrate[4]), .O(n67420));
    defparam i51726_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_1997_i14_3_lut_3_lut (.I0(baudrate[4]), .I1(baudrate[8]), 
            .I2(n2950), .I3(GND_net), .O(n14_adj_4553));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i14_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_1997_i16_3_lut_3_lut (.I0(baudrate[5]), .I1(baudrate[6]), 
            .I2(n2952), .I3(GND_net), .O(n16_adj_4552));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i16_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i51700_2_lut_4_lut (.I0(n2942), .I1(baudrate[16]), .I2(n2951), 
            .I3(baudrate[7]), .O(n67394));
    defparam i51700_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_1997_i18_3_lut_3_lut (.I0(baudrate[7]), .I1(baudrate[16]), 
            .I2(n2942), .I3(GND_net), .O(n18));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i18_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i1_2_lut_4_lut_adj_1051 (.I0(n69977), .I1(baudrate[19]), .I2(n2827), 
            .I3(n62053), .O(n2957));   // verilog/uart_rx.v(119[33:55])
    defparam i1_2_lut_4_lut_adj_1051.LUT_INIT = 16'h7100;
    SB_LUT4 i55134_2_lut_4_lut (.I0(n69977), .I1(baudrate[19]), .I2(n2827), 
            .I3(n25580), .O(n294[4]));   // verilog/uart_rx.v(119[33:55])
    defparam i55134_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_LUT4 i5743_2_lut_3_lut (.I0(baudrate[3]), .I1(n20912), .I2(n11417), 
            .I3(GND_net), .O(n11424));   // verilog/uart_rx.v(119[33:55])
    defparam i5743_2_lut_3_lut.LUT_INIT = 16'h5454;
    SB_LUT4 i5736_2_lut_3_lut (.I0(baudrate[2]), .I1(n962), .I2(baudrate[1]), 
            .I3(GND_net), .O(n11417));   // verilog/uart_rx.v(119[33:55])
    defparam i5736_2_lut_3_lut.LUT_INIT = 16'h4545;
    SB_LUT4 i7217_2_lut_3_lut (.I0(n805), .I1(baudrate[1]), .I2(baudrate[0]), 
            .I3(GND_net), .O(n20902));   // verilog/uart_rx.v(119[33:55])
    defparam i7217_2_lut_3_lut.LUT_INIT = 16'h2a2a;
    SB_LUT4 i48443_2_lut_3_lut (.I0(baudrate[19]), .I1(baudrate[20]), .I2(baudrate[4]), 
            .I3(GND_net), .O(n64128));
    defparam i48443_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i44140_1_lut_4_lut (.I0(n63613), .I1(n63615), .I2(n63461), 
            .I3(n63611), .O(n59786));
    defparam i44140_1_lut_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i1_2_lut_4_lut_adj_1052 (.I0(n69657), .I1(baudrate[18]), .I2(n2713), 
            .I3(n62051), .O(n2845));   // verilog/uart_rx.v(119[33:55])
    defparam i1_2_lut_4_lut_adj_1052.LUT_INIT = 16'h7100;
    SB_LUT4 i55131_2_lut_4_lut (.I0(n69657), .I1(baudrate[18]), .I2(n2713), 
            .I3(n25577), .O(n294[5]));   // verilog/uart_rx.v(119[33:55])
    defparam i55131_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_LUT4 div_37_LessThan_2070_i10_3_lut_3_lut (.I0(baudrate[2]), .I1(baudrate[3]), 
            .I2(n3064), .I3(GND_net), .O(n10_adj_4505));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i10_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_2070_i14_3_lut_3_lut (.I0(baudrate[5]), .I1(baudrate[6]), 
            .I2(n3061), .I3(GND_net), .O(n14_adj_4504));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i14_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i51635_2_lut_4_lut (.I0(n3051), .I1(baudrate[16]), .I2(n3060), 
            .I3(baudrate[7]), .O(n67329));
    defparam i51635_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_2070_i16_3_lut_3_lut (.I0(baudrate[7]), .I1(baudrate[16]), 
            .I2(n3051), .I3(GND_net), .O(n16_adj_4503));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i16_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_2070_i12_3_lut_3_lut (.I0(baudrate[4]), .I1(baudrate[8]), 
            .I2(n3059), .I3(GND_net), .O(n12_adj_4506));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i12_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i51671_2_lut_4_lut (.I0(n3059), .I1(baudrate[8]), .I2(n3063), 
            .I3(baudrate[4]), .O(n67365));
    defparam i51671_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i55156_2_lut_4_lut (.I0(n69765), .I1(baudrate[22]), .I2(n3151), 
            .I3(n25589), .O(n294[1]));
    defparam i55156_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_LUT4 div_37_LessThan_2141_i8_3_lut_3_lut (.I0(baudrate[2]), .I1(baudrate[3]), 
            .I2(n3170), .I3(GND_net), .O(n8_adj_4485));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i8_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_2141_i12_3_lut_3_lut (.I0(baudrate[5]), .I1(baudrate[6]), 
            .I2(n3167), .I3(GND_net), .O(n12_adj_4484));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i12_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i51589_2_lut_4_lut (.I0(n3157), .I1(baudrate[16]), .I2(n3166), 
            .I3(baudrate[7]), .O(n67283));
    defparam i51589_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i1_2_lut_4_lut_adj_1053 (.I0(n69850), .I1(baudrate[17]), .I2(n2596), 
            .I3(n62049), .O(n2730));   // verilog/uart_rx.v(119[33:55])
    defparam i1_2_lut_4_lut_adj_1053.LUT_INIT = 16'h7100;
    SB_LUT4 div_37_LessThan_2141_i14_3_lut_3_lut (.I0(baudrate[7]), .I1(baudrate[16]), 
            .I2(n3157), .I3(GND_net), .O(n14));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i14_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_2141_i10_3_lut_3_lut (.I0(baudrate[4]), .I1(baudrate[8]), 
            .I2(n3165), .I3(GND_net), .O(n10_adj_4486));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i10_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i55127_2_lut_4_lut (.I0(n69850), .I1(baudrate[17]), .I2(n2596), 
            .I3(n25574), .O(n294[6]));   // verilog/uart_rx.v(119[33:55])
    defparam i55127_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_LUT4 i51613_2_lut_4_lut (.I0(n3165), .I1(baudrate[8]), .I2(n3169), 
            .I3(baudrate[4]), .O(n67307));
    defparam i51613_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i7225_4_lut_4_lut (.I0(n960), .I1(n11417), .I2(n20912), .I3(baudrate[3]), 
            .O(n20914));   // verilog/uart_rx.v(119[33:55])
    defparam i7225_4_lut_4_lut.LUT_INIT = 16'ha8aa;
    SB_LUT4 i48523_3_lut_4_lut (.I0(baudrate[30]), .I1(baudrate[31]), .I2(baudrate[26]), 
            .I3(baudrate[24]), .O(n64208));
    defparam i48523_3_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_3_lut_4_lut_adj_1054 (.I0(baudrate[30]), .I1(baudrate[31]), 
            .I2(baudrate[27]), .I3(baudrate[24]), .O(n62015));
    defparam i1_3_lut_4_lut_adj_1054.LUT_INIT = 16'hfffe;
    SB_LUT4 i55118_2_lut_3_lut_4_lut (.I0(baudrate[16]), .I1(n63979), .I2(n48_adj_4685), 
            .I3(baudrate[15]), .O(n294[9]));
    defparam i55118_2_lut_3_lut_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i48509_2_lut_3_lut_4_lut (.I0(baudrate[16]), .I1(n63979), .I2(n62543), 
            .I3(baudrate[15]), .O(n64194));
    defparam i48509_2_lut_3_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_3_lut_adj_1055 (.I0(baudrate[26]), .I1(baudrate[30]), 
            .I2(baudrate[23]), .I3(GND_net), .O(n63615));
    defparam i1_2_lut_3_lut_adj_1055.LUT_INIT = 16'hfefe;
    
endmodule
//
// Verilog Description of module pwm
//

module pwm (n2873, pwm_out, clk32MHz, reset, \pwm_counter[22] , \pwm_counter[21] , 
            \pwm_counter[12] , pwm_setpoint, GND_net, VCC_net, n25, 
            n45, n43) /* synthesis syn_module_defined=1 */ ;
    input n2873;
    output pwm_out;
    input clk32MHz;
    input reset;
    output \pwm_counter[22] ;
    output \pwm_counter[21] ;
    output \pwm_counter[12] ;
    input [23:0]pwm_setpoint;
    input GND_net;
    input VCC_net;
    input n25;
    input n45;
    input n43;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[16:24])
    
    wire pwm_out_N_577, n58232;
    wire [23:0]pwm_counter;   // verilog/pwm.v(11[19:30])
    
    wire n57282, n57310, n57332, n57360, n57388, n57416, n57442, 
        n57478, n57524, n57556, n57622, n57650, n57674, n57706, 
        n57736, n57764, n57798, n57830, n57988, n58118, n58234, 
        n58236, n58238, n67671, n6, n41, n39, n37, n23, n52262, 
        n48, n52261, n52260, n52259, n29, n52258, n52257, n52256, 
        n52255, n52254, n52253, n52252, n52251, n31, n52250, n52249, 
        n35, n33, n52248, n52247, n52246, n52245, n52244, n52243, 
        n11, n13, n15, n27, n9, n17, n19, n21, n52242, n52241, 
        n52240, n67637, n67628, n12, n30, n68560, n68548, n69680, 
        n69057, n69806, n69430, n69431, n16, n24, n67507, n8, 
        n67498, n68936, n68242, n4, n69047, n69048, n67553, n10, 
        n67534, n69674, n68244, n69902, n69903, n69816, n67509, 
        n69575, n68250, n69786, n61641, n22, n15_adj_4455, n20, 
        n24_adj_4456, n19_adj_4457;
    
    SB_DFFE pwm_out_12 (.Q(pwm_out), .C(clk32MHz), .E(n2873), .D(pwm_out_N_577));   // verilog/pwm.v(16[12] 26[6])
    SB_DFFR pwm_counter_1935__i0 (.Q(pwm_counter[0]), .C(clk32MHz), .D(n58232), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_1935__i23 (.Q(pwm_counter[23]), .C(clk32MHz), .D(n57282), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_1935__i22 (.Q(\pwm_counter[22] ), .C(clk32MHz), 
            .D(n57310), .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_1935__i21 (.Q(\pwm_counter[21] ), .C(clk32MHz), 
            .D(n57332), .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_1935__i20 (.Q(pwm_counter[20]), .C(clk32MHz), .D(n57360), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_1935__i19 (.Q(pwm_counter[19]), .C(clk32MHz), .D(n57388), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_1935__i18 (.Q(pwm_counter[18]), .C(clk32MHz), .D(n57416), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_1935__i17 (.Q(pwm_counter[17]), .C(clk32MHz), .D(n57442), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_1935__i16 (.Q(pwm_counter[16]), .C(clk32MHz), .D(n57478), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_1935__i15 (.Q(pwm_counter[15]), .C(clk32MHz), .D(n57524), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_1935__i14 (.Q(pwm_counter[14]), .C(clk32MHz), .D(n57556), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_1935__i13 (.Q(pwm_counter[13]), .C(clk32MHz), .D(n57622), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_1935__i12 (.Q(\pwm_counter[12] ), .C(clk32MHz), 
            .D(n57650), .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_1935__i11 (.Q(pwm_counter[11]), .C(clk32MHz), .D(n57674), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_1935__i10 (.Q(pwm_counter[10]), .C(clk32MHz), .D(n57706), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_1935__i9 (.Q(pwm_counter[9]), .C(clk32MHz), .D(n57736), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_1935__i8 (.Q(pwm_counter[8]), .C(clk32MHz), .D(n57764), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_1935__i7 (.Q(pwm_counter[7]), .C(clk32MHz), .D(n57798), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_1935__i6 (.Q(pwm_counter[6]), .C(clk32MHz), .D(n57830), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_1935__i5 (.Q(pwm_counter[5]), .C(clk32MHz), .D(n57988), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_1935__i4 (.Q(pwm_counter[4]), .C(clk32MHz), .D(n58118), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_1935__i3 (.Q(pwm_counter[3]), .C(clk32MHz), .D(n58234), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_1935__i2 (.Q(pwm_counter[2]), .C(clk32MHz), .D(n58236), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_1935__i1 (.Q(pwm_counter[1]), .C(clk32MHz), .D(n58238), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_LUT4 i51977_3_lut_4_lut (.I0(pwm_counter[3]), .I1(pwm_setpoint[3]), 
            .I2(pwm_setpoint[2]), .I3(pwm_counter[2]), .O(n67671));   // verilog/pwm.v(21[8:24])
    defparam i51977_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 duty_23__I_0_i6_3_lut_3_lut (.I0(pwm_counter[3]), .I1(pwm_setpoint[3]), 
            .I2(pwm_setpoint[2]), .I3(GND_net), .O(n6));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 duty_23__I_0_i41_2_lut (.I0(pwm_counter[20]), .I1(pwm_setpoint[20]), 
            .I2(GND_net), .I3(GND_net), .O(n41));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i39_2_lut (.I0(pwm_counter[19]), .I1(pwm_setpoint[19]), 
            .I2(GND_net), .I3(GND_net), .O(n39));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i37_2_lut (.I0(pwm_counter[18]), .I1(pwm_setpoint[18]), 
            .I2(GND_net), .I3(GND_net), .O(n37));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i23_2_lut (.I0(pwm_counter[11]), .I1(pwm_setpoint[11]), 
            .I2(GND_net), .I3(GND_net), .O(n23));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 pwm_counter_1935_add_4_25_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[23]), 
            .I3(n52262), .O(n57282)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1935_add_4_25_lut.LUT_INIT = 16'h8228;
    SB_LUT4 pwm_counter_1935_add_4_24_lut (.I0(n48), .I1(GND_net), .I2(\pwm_counter[22] ), 
            .I3(n52261), .O(n57310)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1935_add_4_24_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_1935_add_4_24 (.CI(n52261), .I0(GND_net), .I1(\pwm_counter[22] ), 
            .CO(n52262));
    SB_LUT4 pwm_counter_1935_add_4_23_lut (.I0(n48), .I1(GND_net), .I2(\pwm_counter[21] ), 
            .I3(n52260), .O(n57332)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1935_add_4_23_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_1935_add_4_23 (.CI(n52260), .I0(GND_net), .I1(\pwm_counter[21] ), 
            .CO(n52261));
    SB_LUT4 pwm_counter_1935_add_4_22_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[20]), 
            .I3(n52259), .O(n57360)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1935_add_4_22_lut.LUT_INIT = 16'h8228;
    SB_LUT4 duty_23__I_0_i29_2_lut (.I0(pwm_counter[14]), .I1(pwm_setpoint[14]), 
            .I2(GND_net), .I3(GND_net), .O(n29));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i29_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY pwm_counter_1935_add_4_22 (.CI(n52259), .I0(GND_net), .I1(pwm_counter[20]), 
            .CO(n52260));
    SB_LUT4 pwm_counter_1935_add_4_21_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[19]), 
            .I3(n52258), .O(n57388)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1935_add_4_21_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_1935_add_4_21 (.CI(n52258), .I0(GND_net), .I1(pwm_counter[19]), 
            .CO(n52259));
    SB_LUT4 pwm_counter_1935_add_4_20_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[18]), 
            .I3(n52257), .O(n57416)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1935_add_4_20_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_1935_add_4_20 (.CI(n52257), .I0(GND_net), .I1(pwm_counter[18]), 
            .CO(n52258));
    SB_LUT4 pwm_counter_1935_add_4_19_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[17]), 
            .I3(n52256), .O(n57442)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1935_add_4_19_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_1935_add_4_19 (.CI(n52256), .I0(GND_net), .I1(pwm_counter[17]), 
            .CO(n52257));
    SB_LUT4 pwm_counter_1935_add_4_18_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[16]), 
            .I3(n52255), .O(n57478)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1935_add_4_18_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_1935_add_4_18 (.CI(n52255), .I0(GND_net), .I1(pwm_counter[16]), 
            .CO(n52256));
    SB_LUT4 pwm_counter_1935_add_4_17_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[15]), 
            .I3(n52254), .O(n57524)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1935_add_4_17_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_1935_add_4_17 (.CI(n52254), .I0(GND_net), .I1(pwm_counter[15]), 
            .CO(n52255));
    SB_LUT4 pwm_counter_1935_add_4_16_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[14]), 
            .I3(n52253), .O(n57556)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1935_add_4_16_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_1935_add_4_16 (.CI(n52253), .I0(GND_net), .I1(pwm_counter[14]), 
            .CO(n52254));
    SB_LUT4 pwm_counter_1935_add_4_15_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[13]), 
            .I3(n52252), .O(n57622)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1935_add_4_15_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_1935_add_4_15 (.CI(n52252), .I0(GND_net), .I1(pwm_counter[13]), 
            .CO(n52253));
    SB_LUT4 pwm_counter_1935_add_4_14_lut (.I0(n48), .I1(GND_net), .I2(\pwm_counter[12] ), 
            .I3(n52251), .O(n57650)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1935_add_4_14_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_1935_add_4_14 (.CI(n52251), .I0(GND_net), .I1(\pwm_counter[12] ), 
            .CO(n52252));
    SB_LUT4 duty_23__I_0_i31_2_lut (.I0(pwm_counter[15]), .I1(pwm_setpoint[15]), 
            .I2(GND_net), .I3(GND_net), .O(n31));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 pwm_counter_1935_add_4_13_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[11]), 
            .I3(n52250), .O(n57674)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1935_add_4_13_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_1935_add_4_13 (.CI(n52250), .I0(GND_net), .I1(pwm_counter[11]), 
            .CO(n52251));
    SB_LUT4 pwm_counter_1935_add_4_12_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[10]), 
            .I3(n52249), .O(n57706)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1935_add_4_12_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_1935_add_4_12 (.CI(n52249), .I0(GND_net), .I1(pwm_counter[10]), 
            .CO(n52250));
    SB_LUT4 duty_23__I_0_i35_2_lut (.I0(pwm_counter[17]), .I1(pwm_setpoint[17]), 
            .I2(GND_net), .I3(GND_net), .O(n35));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i33_2_lut (.I0(pwm_counter[16]), .I1(pwm_setpoint[16]), 
            .I2(GND_net), .I3(GND_net), .O(n33));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 pwm_counter_1935_add_4_11_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[9]), 
            .I3(n52248), .O(n57736)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1935_add_4_11_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_1935_add_4_11 (.CI(n52248), .I0(GND_net), .I1(pwm_counter[9]), 
            .CO(n52249));
    SB_LUT4 pwm_counter_1935_add_4_10_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[8]), 
            .I3(n52247), .O(n57764)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1935_add_4_10_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_1935_add_4_10 (.CI(n52247), .I0(GND_net), .I1(pwm_counter[8]), 
            .CO(n52248));
    SB_LUT4 pwm_counter_1935_add_4_9_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[7]), 
            .I3(n52246), .O(n57798)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1935_add_4_9_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_1935_add_4_9 (.CI(n52246), .I0(GND_net), .I1(pwm_counter[7]), 
            .CO(n52247));
    SB_LUT4 pwm_counter_1935_add_4_8_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[6]), 
            .I3(n52245), .O(n57830)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1935_add_4_8_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_1935_add_4_8 (.CI(n52245), .I0(GND_net), .I1(pwm_counter[6]), 
            .CO(n52246));
    SB_LUT4 pwm_counter_1935_add_4_7_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[5]), 
            .I3(n52244), .O(n57988)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1935_add_4_7_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_1935_add_4_7 (.CI(n52244), .I0(GND_net), .I1(pwm_counter[5]), 
            .CO(n52245));
    SB_LUT4 pwm_counter_1935_add_4_6_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[4]), 
            .I3(n52243), .O(n58118)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1935_add_4_6_lut.LUT_INIT = 16'h8228;
    SB_LUT4 duty_23__I_0_i11_2_lut (.I0(pwm_counter[5]), .I1(pwm_setpoint[5]), 
            .I2(GND_net), .I3(GND_net), .O(n11));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i13_2_lut (.I0(pwm_counter[6]), .I1(pwm_setpoint[6]), 
            .I2(GND_net), .I3(GND_net), .O(n13));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i13_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY pwm_counter_1935_add_4_6 (.CI(n52243), .I0(GND_net), .I1(pwm_counter[4]), 
            .CO(n52244));
    SB_LUT4 duty_23__I_0_i15_2_lut (.I0(pwm_counter[7]), .I1(pwm_setpoint[7]), 
            .I2(GND_net), .I3(GND_net), .O(n15));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i27_2_lut (.I0(pwm_counter[13]), .I1(pwm_setpoint[13]), 
            .I2(GND_net), .I3(GND_net), .O(n27));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i9_2_lut (.I0(pwm_counter[4]), .I1(pwm_setpoint[4]), 
            .I2(GND_net), .I3(GND_net), .O(n9));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i17_2_lut (.I0(pwm_counter[8]), .I1(pwm_setpoint[8]), 
            .I2(GND_net), .I3(GND_net), .O(n17));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i19_2_lut (.I0(pwm_counter[9]), .I1(pwm_setpoint[9]), 
            .I2(GND_net), .I3(GND_net), .O(n19));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i21_2_lut (.I0(pwm_counter[10]), .I1(pwm_setpoint[10]), 
            .I2(GND_net), .I3(GND_net), .O(n21));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 pwm_counter_1935_add_4_5_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[3]), 
            .I3(n52242), .O(n58234)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1935_add_4_5_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_1935_add_4_5 (.CI(n52242), .I0(GND_net), .I1(pwm_counter[3]), 
            .CO(n52243));
    SB_LUT4 pwm_counter_1935_add_4_4_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[2]), 
            .I3(n52241), .O(n58236)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1935_add_4_4_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_1935_add_4_4 (.CI(n52241), .I0(GND_net), .I1(pwm_counter[2]), 
            .CO(n52242));
    SB_LUT4 pwm_counter_1935_add_4_3_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[1]), 
            .I3(n52240), .O(n58238)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1935_add_4_3_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_1935_add_4_3 (.CI(n52240), .I0(GND_net), .I1(pwm_counter[1]), 
            .CO(n52241));
    SB_LUT4 i51943_4_lut (.I0(n21), .I1(n19), .I2(n17), .I3(n9), .O(n67637));
    defparam i51943_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i51934_4_lut (.I0(n27), .I1(n15), .I2(n13), .I3(n11), .O(n67628));
    defparam i51934_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 pwm_counter_1935_add_4_2_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[0]), 
            .I3(VCC_net), .O(n58232)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1935_add_4_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_1935_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(pwm_counter[0]), 
            .CO(n52240));
    SB_LUT4 duty_23__I_0_i30_3_lut (.I0(n12), .I1(pwm_setpoint[17]), .I2(n35), 
            .I3(GND_net), .O(n30));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52866_4_lut (.I0(n13), .I1(n11), .I2(n9), .I3(n67671), 
            .O(n68560));
    defparam i52866_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i52854_4_lut (.I0(n19), .I1(n17), .I2(n15), .I3(n68560), 
            .O(n68548));
    defparam i52854_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i53986_4_lut (.I0(n25), .I1(n23), .I2(n21), .I3(n68548), 
            .O(n69680));
    defparam i53986_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i53363_4_lut (.I0(n31), .I1(n29), .I2(n27), .I3(n69680), 
            .O(n69057));
    defparam i53363_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i54112_4_lut (.I0(n37), .I1(n35), .I2(n33), .I3(n69057), 
            .O(n69806));
    defparam i54112_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i53736_3_lut (.I0(n6), .I1(pwm_setpoint[10]), .I2(n21), .I3(GND_net), 
            .O(n69430));   // verilog/pwm.v(21[8:24])
    defparam i53736_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53737_3_lut (.I0(n69430), .I1(pwm_setpoint[11]), .I2(n23), 
            .I3(GND_net), .O(n69431));   // verilog/pwm.v(21[8:24])
    defparam i53737_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i24_3_lut (.I0(n16), .I1(pwm_setpoint[22]), .I2(n45), 
            .I3(GND_net), .O(n24));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51813_4_lut (.I0(n43), .I1(n25), .I2(n23), .I3(n67637), 
            .O(n67507));
    defparam i51813_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i53242_4_lut (.I0(n24), .I1(n8), .I2(n45), .I3(n67498), 
            .O(n68936));   // verilog/pwm.v(21[8:24])
    defparam i53242_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i52548_3_lut (.I0(n69431), .I1(pwm_setpoint[12]), .I2(n25), 
            .I3(GND_net), .O(n68242));   // verilog/pwm.v(21[8:24])
    defparam i52548_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i4_4_lut (.I0(pwm_counter[0]), .I1(pwm_setpoint[1]), 
            .I2(pwm_counter[1]), .I3(pwm_setpoint[0]), .O(n4));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i4_4_lut.LUT_INIT = 16'h4d0c;
    SB_LUT4 i53353_3_lut (.I0(n4), .I1(pwm_setpoint[13]), .I2(n27), .I3(GND_net), 
            .O(n69047));   // verilog/pwm.v(21[8:24])
    defparam i53353_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53354_3_lut (.I0(n69047), .I1(pwm_setpoint[14]), .I2(n29), 
            .I3(GND_net), .O(n69048));   // verilog/pwm.v(21[8:24])
    defparam i53354_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51859_4_lut (.I0(n33), .I1(n31), .I2(n29), .I3(n67628), 
            .O(n67553));
    defparam i51859_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i53980_4_lut (.I0(n30), .I1(n10), .I2(n35), .I3(n67534), 
            .O(n69674));   // verilog/pwm.v(21[8:24])
    defparam i53980_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i52550_3_lut (.I0(n69048), .I1(pwm_setpoint[15]), .I2(n31), 
            .I3(GND_net), .O(n68244));   // verilog/pwm.v(21[8:24])
    defparam i52550_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i54208_4_lut (.I0(n68244), .I1(n69674), .I2(n35), .I3(n67553), 
            .O(n69902));   // verilog/pwm.v(21[8:24])
    defparam i54208_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i54209_3_lut (.I0(n69902), .I1(pwm_setpoint[18]), .I2(n37), 
            .I3(GND_net), .O(n69903));   // verilog/pwm.v(21[8:24])
    defparam i54209_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i54122_3_lut (.I0(n69903), .I1(pwm_setpoint[19]), .I2(n39), 
            .I3(GND_net), .O(n69816));   // verilog/pwm.v(21[8:24])
    defparam i54122_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51815_4_lut (.I0(n43), .I1(n41), .I2(n39), .I3(n69806), 
            .O(n67509));
    defparam i51815_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i53881_4_lut (.I0(n68242), .I1(n68936), .I2(n45), .I3(n67507), 
            .O(n69575));   // verilog/pwm.v(21[8:24])
    defparam i53881_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i52556_3_lut (.I0(n69816), .I1(pwm_setpoint[20]), .I2(n41), 
            .I3(GND_net), .O(n68250));   // verilog/pwm.v(21[8:24])
    defparam i52556_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i54092_4_lut (.I0(n68250), .I1(n69575), .I2(n45), .I3(n67509), 
            .O(n69786));   // verilog/pwm.v(21[8:24])
    defparam i54092_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i54093_3_lut (.I0(n69786), .I1(pwm_counter[23]), .I2(pwm_setpoint[23]), 
            .I3(GND_net), .O(pwm_out_N_577));   // verilog/pwm.v(21[8:24])
    defparam i54093_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i2_3_lut (.I0(pwm_counter[6]), .I1(pwm_counter[8]), .I2(pwm_counter[7]), 
            .I3(GND_net), .O(n61641));
    defparam i2_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i9_4_lut (.I0(pwm_counter[15]), .I1(pwm_counter[16]), .I2(pwm_counter[20]), 
            .I3(pwm_counter[19]), .O(n22));
    defparam i9_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_4_lut (.I0(n61641), .I1(\pwm_counter[21] ), .I2(pwm_counter[10]), 
            .I3(pwm_counter[9]), .O(n15_adj_4455));
    defparam i2_4_lut.LUT_INIT = 16'heccc;
    SB_LUT4 i7_3_lut (.I0(pwm_counter[13]), .I1(\pwm_counter[22] ), .I2(pwm_counter[11]), 
            .I3(GND_net), .O(n20));
    defparam i7_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i11_4_lut (.I0(n15_adj_4455), .I1(n22), .I2(\pwm_counter[12] ), 
            .I3(pwm_counter[18]), .O(n24_adj_4456));
    defparam i11_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i6_2_lut (.I0(pwm_counter[14]), .I1(pwm_counter[17]), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_4457));
    defparam i6_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut (.I0(pwm_counter[23]), .I1(n19_adj_4457), .I2(n24_adj_4456), 
            .I3(n20), .O(n48));   // verilog/pwm.v(17[20:33])
    defparam i1_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 duty_23__I_0_i8_3_lut_3_lut (.I0(pwm_setpoint[4]), .I1(pwm_setpoint[8]), 
            .I2(pwm_counter[8]), .I3(GND_net), .O(n8));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i8_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i51804_2_lut_4_lut (.I0(pwm_setpoint[21]), .I1(\pwm_counter[21] ), 
            .I2(pwm_counter[9]), .I3(pwm_setpoint[9]), .O(n67498));
    defparam i51804_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 duty_23__I_0_i16_3_lut_3_lut (.I0(pwm_setpoint[9]), .I1(pwm_setpoint[21]), 
            .I2(\pwm_counter[21] ), .I3(GND_net), .O(n16));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i16_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 duty_23__I_0_i10_3_lut_3_lut (.I0(pwm_setpoint[5]), .I1(pwm_setpoint[6]), 
            .I2(pwm_counter[6]), .I3(GND_net), .O(n10));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i10_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i51840_2_lut_4_lut (.I0(pwm_counter[16]), .I1(pwm_setpoint[16]), 
            .I2(pwm_counter[7]), .I3(pwm_setpoint[7]), .O(n67534));
    defparam i51840_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 duty_23__I_0_i12_3_lut_3_lut (.I0(pwm_setpoint[7]), .I1(pwm_setpoint[16]), 
            .I2(pwm_counter[16]), .I3(GND_net), .O(n12));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i12_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    
endmodule
//
// Verilog Description of module pll32MHz
//

module pll32MHz (GND_net, clk16MHz, VCC_net, clk32MHz) /* synthesis syn_module_defined=1 */ ;
    input GND_net;
    input clk16MHz;
    input VCC_net;
    output clk32MHz;
    
    wire clk16MHz /* synthesis SET_AS_NETWORK=clk16MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[16:24])
    
    SB_PLL40_CORE pll32MHz_inst (.REFERENCECLK(clk16MHz), .PLLOUTCORE(clk32MHz), 
            .BYPASS(GND_net), .RESETB(VCC_net)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=52, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=34, LSE_RLINE=38 */ ;   // verilog/TinyFPGA_B.v(34[10] 38[2])
    defparam pll32MHz_inst.FEEDBACK_PATH = "PHASE_AND_DELAY";
    defparam pll32MHz_inst.DELAY_ADJUSTMENT_MODE_FEEDBACK = "FIXED";
    defparam pll32MHz_inst.DELAY_ADJUSTMENT_MODE_RELATIVE = "FIXED";
    defparam pll32MHz_inst.SHIFTREG_DIV_MODE = 2'b00;
    defparam pll32MHz_inst.FDA_FEEDBACK = 4'b0000;
    defparam pll32MHz_inst.FDA_RELATIVE = 4'b0000;
    defparam pll32MHz_inst.PLLOUT_SELECT = "SHIFTREG_0deg";
    defparam pll32MHz_inst.DIVR = 4'b0000;
    defparam pll32MHz_inst.DIVF = 7'b0000001;
    defparam pll32MHz_inst.DIVQ = 3'b011;
    defparam pll32MHz_inst.FILTER_RANGE = 3'b001;
    defparam pll32MHz_inst.ENABLE_ICEGATE = 1'b0;
    defparam pll32MHz_inst.TEST_MODE = 1'b0;
    defparam pll32MHz_inst.EXTERNAL_DIVIDE_FACTOR = 1;
    
endmodule
//
// Verilog Description of module \quadrature_decoder(0)_U0 
//

module \quadrature_decoder(0)_U0  (n1744, GND_net, \encoder0_position[30] , 
            \encoder0_position[29] , ENCODER0_B_N_keep, n1779, ENCODER0_A_N_keep, 
            \encoder0_position[28] , \encoder0_position[27] , \encoder0_position[26] , 
            \encoder0_position[25] , \encoder0_position[24] , b_prev, 
            \a_new[1] , \encoder0_position[23] , \encoder0_position[22] , 
            \encoder0_position[21] , \encoder0_position[20] , \encoder0_position[19] , 
            \encoder0_position[18] , \encoder0_position[17] , \encoder0_position[16] , 
            \encoder0_position[15] , \encoder0_position[14] , \encoder0_position[13] , 
            \encoder0_position[12] , \encoder0_position[11] , \encoder0_position[10] , 
            \encoder0_position[9] , \encoder0_position[8] , \encoder0_position[7] , 
            \encoder0_position[6] , \encoder0_position[5] , \encoder0_position[4] , 
            \encoder0_position[3] , \encoder0_position[2] , \encoder0_position[1] , 
            \encoder0_position[0] , VCC_net, n29648, a_prev, n29647, 
            n29628, n1742, position_31__N_3836, \b_new[1] , debounce_cnt_N_3833) /* synthesis lattice_noprune=1 */ ;
    output n1744;
    input GND_net;
    output \encoder0_position[30] ;
    output \encoder0_position[29] ;
    input ENCODER0_B_N_keep;
    input n1779;
    input ENCODER0_A_N_keep;
    output \encoder0_position[28] ;
    output \encoder0_position[27] ;
    output \encoder0_position[26] ;
    output \encoder0_position[25] ;
    output \encoder0_position[24] ;
    output b_prev;
    output \a_new[1] ;
    output \encoder0_position[23] ;
    output \encoder0_position[22] ;
    output \encoder0_position[21] ;
    output \encoder0_position[20] ;
    output \encoder0_position[19] ;
    output \encoder0_position[18] ;
    output \encoder0_position[17] ;
    output \encoder0_position[16] ;
    output \encoder0_position[15] ;
    output \encoder0_position[14] ;
    output \encoder0_position[13] ;
    output \encoder0_position[12] ;
    output \encoder0_position[11] ;
    output \encoder0_position[10] ;
    output \encoder0_position[9] ;
    output \encoder0_position[8] ;
    output \encoder0_position[7] ;
    output \encoder0_position[6] ;
    output \encoder0_position[5] ;
    output \encoder0_position[4] ;
    output \encoder0_position[3] ;
    output \encoder0_position[2] ;
    output \encoder0_position[1] ;
    output \encoder0_position[0] ;
    input VCC_net;
    input n29648;
    output a_prev;
    input n29647;
    input n29628;
    output n1742;
    output position_31__N_3836;
    output \b_new[1] ;
    output debounce_cnt_N_3833;
    
    wire [31:0]n133;
    
    wire direction_N_3840, n52426, n52425, n52424;
    wire [1:0]b_new;   // vhdl/quadrature_decoder.vhd(40[9:14])
    wire [1:0]a_new;   // vhdl/quadrature_decoder.vhd(39[9:14])
    
    wire n52423, n52422, n52421, n52420, n52419, n52418, n52417, 
        n52416, n52415, n52414, n52413, n52412, n52411, n52410, 
        n52409, n52408, n52407, n52406, n52405, n52404, n52403, 
        n52402, n52401, n52400, n52399, n52398, n52397, n52396;
    
    SB_LUT4 position_1952_add_4_33_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(n1744), .I3(n52426), .O(n133[31])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1952_add_4_33_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 position_1952_add_4_32_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder0_position[30] ), .I3(n52425), .O(n133[30])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1952_add_4_32_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1952_add_4_32 (.CI(n52425), .I0(direction_N_3840), 
            .I1(\encoder0_position[30] ), .CO(n52426));
    SB_LUT4 position_1952_add_4_31_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder0_position[29] ), .I3(n52424), .O(n133[29])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1952_add_4_31_lut.LUT_INIT = 16'hC33C;
    SB_DFF b_new_i0 (.Q(b_new[0]), .C(n1779), .D(ENCODER0_B_N_keep));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_DFF a_new_i0 (.Q(a_new[0]), .C(n1779), .D(ENCODER0_A_N_keep));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_CARRY position_1952_add_4_31 (.CI(n52424), .I0(direction_N_3840), 
            .I1(\encoder0_position[29] ), .CO(n52425));
    SB_LUT4 position_1952_add_4_30_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder0_position[28] ), .I3(n52423), .O(n133[28])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1952_add_4_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1952_add_4_30 (.CI(n52423), .I0(direction_N_3840), 
            .I1(\encoder0_position[28] ), .CO(n52424));
    SB_LUT4 position_1952_add_4_29_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder0_position[27] ), .I3(n52422), .O(n133[27])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1952_add_4_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1952_add_4_29 (.CI(n52422), .I0(direction_N_3840), 
            .I1(\encoder0_position[27] ), .CO(n52423));
    SB_LUT4 position_1952_add_4_28_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder0_position[26] ), .I3(n52421), .O(n133[26])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1952_add_4_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1952_add_4_28 (.CI(n52421), .I0(direction_N_3840), 
            .I1(\encoder0_position[26] ), .CO(n52422));
    SB_LUT4 position_1952_add_4_27_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder0_position[25] ), .I3(n52420), .O(n133[25])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1952_add_4_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1952_add_4_27 (.CI(n52420), .I0(direction_N_3840), 
            .I1(\encoder0_position[25] ), .CO(n52421));
    SB_LUT4 position_1952_add_4_26_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder0_position[24] ), .I3(n52419), .O(n133[24])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1952_add_4_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1952_add_4_26 (.CI(n52419), .I0(direction_N_3840), 
            .I1(\encoder0_position[24] ), .CO(n52420));
    SB_LUT4 b_prev_I_0_48_2_lut (.I0(b_prev), .I1(\a_new[1] ), .I2(GND_net), 
            .I3(GND_net), .O(direction_N_3840));   // vhdl/quadrature_decoder.vhd(64[18:37])
    defparam b_prev_I_0_48_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 position_1952_add_4_25_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder0_position[23] ), .I3(n52418), .O(n133[23])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1952_add_4_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1952_add_4_25 (.CI(n52418), .I0(direction_N_3840), 
            .I1(\encoder0_position[23] ), .CO(n52419));
    SB_LUT4 position_1952_add_4_24_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder0_position[22] ), .I3(n52417), .O(n133[22])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1952_add_4_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1952_add_4_24 (.CI(n52417), .I0(direction_N_3840), 
            .I1(\encoder0_position[22] ), .CO(n52418));
    SB_LUT4 position_1952_add_4_23_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder0_position[21] ), .I3(n52416), .O(n133[21])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1952_add_4_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1952_add_4_23 (.CI(n52416), .I0(direction_N_3840), 
            .I1(\encoder0_position[21] ), .CO(n52417));
    SB_LUT4 position_1952_add_4_22_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder0_position[20] ), .I3(n52415), .O(n133[20])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1952_add_4_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1952_add_4_22 (.CI(n52415), .I0(direction_N_3840), 
            .I1(\encoder0_position[20] ), .CO(n52416));
    SB_LUT4 position_1952_add_4_21_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder0_position[19] ), .I3(n52414), .O(n133[19])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1952_add_4_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1952_add_4_21 (.CI(n52414), .I0(direction_N_3840), 
            .I1(\encoder0_position[19] ), .CO(n52415));
    SB_LUT4 position_1952_add_4_20_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder0_position[18] ), .I3(n52413), .O(n133[18])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1952_add_4_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1952_add_4_20 (.CI(n52413), .I0(direction_N_3840), 
            .I1(\encoder0_position[18] ), .CO(n52414));
    SB_LUT4 position_1952_add_4_19_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder0_position[17] ), .I3(n52412), .O(n133[17])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1952_add_4_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1952_add_4_19 (.CI(n52412), .I0(direction_N_3840), 
            .I1(\encoder0_position[17] ), .CO(n52413));
    SB_LUT4 position_1952_add_4_18_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder0_position[16] ), .I3(n52411), .O(n133[16])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1952_add_4_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1952_add_4_18 (.CI(n52411), .I0(direction_N_3840), 
            .I1(\encoder0_position[16] ), .CO(n52412));
    SB_LUT4 position_1952_add_4_17_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder0_position[15] ), .I3(n52410), .O(n133[15])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1952_add_4_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1952_add_4_17 (.CI(n52410), .I0(direction_N_3840), 
            .I1(\encoder0_position[15] ), .CO(n52411));
    SB_LUT4 position_1952_add_4_16_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder0_position[14] ), .I3(n52409), .O(n133[14])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1952_add_4_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1952_add_4_16 (.CI(n52409), .I0(direction_N_3840), 
            .I1(\encoder0_position[14] ), .CO(n52410));
    SB_LUT4 position_1952_add_4_15_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder0_position[13] ), .I3(n52408), .O(n133[13])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1952_add_4_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1952_add_4_15 (.CI(n52408), .I0(direction_N_3840), 
            .I1(\encoder0_position[13] ), .CO(n52409));
    SB_LUT4 position_1952_add_4_14_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder0_position[12] ), .I3(n52407), .O(n133[12])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1952_add_4_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1952_add_4_14 (.CI(n52407), .I0(direction_N_3840), 
            .I1(\encoder0_position[12] ), .CO(n52408));
    SB_LUT4 position_1952_add_4_13_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder0_position[11] ), .I3(n52406), .O(n133[11])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1952_add_4_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1952_add_4_13 (.CI(n52406), .I0(direction_N_3840), 
            .I1(\encoder0_position[11] ), .CO(n52407));
    SB_LUT4 position_1952_add_4_12_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder0_position[10] ), .I3(n52405), .O(n133[10])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1952_add_4_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1952_add_4_12 (.CI(n52405), .I0(direction_N_3840), 
            .I1(\encoder0_position[10] ), .CO(n52406));
    SB_LUT4 position_1952_add_4_11_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder0_position[9] ), .I3(n52404), .O(n133[9])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1952_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1952_add_4_11 (.CI(n52404), .I0(direction_N_3840), 
            .I1(\encoder0_position[9] ), .CO(n52405));
    SB_LUT4 position_1952_add_4_10_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder0_position[8] ), .I3(n52403), .O(n133[8])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1952_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1952_add_4_10 (.CI(n52403), .I0(direction_N_3840), 
            .I1(\encoder0_position[8] ), .CO(n52404));
    SB_LUT4 position_1952_add_4_9_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder0_position[7] ), .I3(n52402), .O(n133[7])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1952_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1952_add_4_9 (.CI(n52402), .I0(direction_N_3840), 
            .I1(\encoder0_position[7] ), .CO(n52403));
    SB_LUT4 position_1952_add_4_8_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder0_position[6] ), .I3(n52401), .O(n133[6])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1952_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1952_add_4_8 (.CI(n52401), .I0(direction_N_3840), 
            .I1(\encoder0_position[6] ), .CO(n52402));
    SB_LUT4 position_1952_add_4_7_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder0_position[5] ), .I3(n52400), .O(n133[5])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1952_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1952_add_4_7 (.CI(n52400), .I0(direction_N_3840), 
            .I1(\encoder0_position[5] ), .CO(n52401));
    SB_LUT4 position_1952_add_4_6_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder0_position[4] ), .I3(n52399), .O(n133[4])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1952_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1952_add_4_6 (.CI(n52399), .I0(direction_N_3840), 
            .I1(\encoder0_position[4] ), .CO(n52400));
    SB_LUT4 position_1952_add_4_5_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder0_position[3] ), .I3(n52398), .O(n133[3])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1952_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1952_add_4_5 (.CI(n52398), .I0(direction_N_3840), 
            .I1(\encoder0_position[3] ), .CO(n52399));
    SB_LUT4 position_1952_add_4_4_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder0_position[2] ), .I3(n52397), .O(n133[2])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1952_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1952_add_4_4 (.CI(n52397), .I0(direction_N_3840), 
            .I1(\encoder0_position[2] ), .CO(n52398));
    SB_LUT4 position_1952_add_4_3_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder0_position[1] ), .I3(n52396), .O(n133[1])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1952_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1952_add_4_3 (.CI(n52396), .I0(direction_N_3840), 
            .I1(\encoder0_position[1] ), .CO(n52397));
    SB_LUT4 position_1952_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(\encoder0_position[0] ), 
            .I3(VCC_net), .O(n133[0])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1952_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1952_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(\encoder0_position[0] ), 
            .CO(n52396));
    SB_DFF a_prev_40 (.Q(a_prev), .C(n1779), .D(n29648));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_DFF b_prev_41 (.Q(b_prev), .C(n1779), .D(n29647));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_DFF direction_42 (.Q(n1742), .C(n1779), .D(n29628));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_DFFE position_1952__i31 (.Q(n1744), .C(n1779), .E(position_31__N_3836), 
            .D(n133[31]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1952__i30 (.Q(\encoder0_position[30] ), .C(n1779), 
            .E(position_31__N_3836), .D(n133[30]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1952__i29 (.Q(\encoder0_position[29] ), .C(n1779), 
            .E(position_31__N_3836), .D(n133[29]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1952__i28 (.Q(\encoder0_position[28] ), .C(n1779), 
            .E(position_31__N_3836), .D(n133[28]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1952__i27 (.Q(\encoder0_position[27] ), .C(n1779), 
            .E(position_31__N_3836), .D(n133[27]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1952__i26 (.Q(\encoder0_position[26] ), .C(n1779), 
            .E(position_31__N_3836), .D(n133[26]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1952__i25 (.Q(\encoder0_position[25] ), .C(n1779), 
            .E(position_31__N_3836), .D(n133[25]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1952__i24 (.Q(\encoder0_position[24] ), .C(n1779), 
            .E(position_31__N_3836), .D(n133[24]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1952__i23 (.Q(\encoder0_position[23] ), .C(n1779), 
            .E(position_31__N_3836), .D(n133[23]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1952__i22 (.Q(\encoder0_position[22] ), .C(n1779), 
            .E(position_31__N_3836), .D(n133[22]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1952__i21 (.Q(\encoder0_position[21] ), .C(n1779), 
            .E(position_31__N_3836), .D(n133[21]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1952__i20 (.Q(\encoder0_position[20] ), .C(n1779), 
            .E(position_31__N_3836), .D(n133[20]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1952__i19 (.Q(\encoder0_position[19] ), .C(n1779), 
            .E(position_31__N_3836), .D(n133[19]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1952__i18 (.Q(\encoder0_position[18] ), .C(n1779), 
            .E(position_31__N_3836), .D(n133[18]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1952__i17 (.Q(\encoder0_position[17] ), .C(n1779), 
            .E(position_31__N_3836), .D(n133[17]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1952__i16 (.Q(\encoder0_position[16] ), .C(n1779), 
            .E(position_31__N_3836), .D(n133[16]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1952__i15 (.Q(\encoder0_position[15] ), .C(n1779), 
            .E(position_31__N_3836), .D(n133[15]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1952__i14 (.Q(\encoder0_position[14] ), .C(n1779), 
            .E(position_31__N_3836), .D(n133[14]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1952__i13 (.Q(\encoder0_position[13] ), .C(n1779), 
            .E(position_31__N_3836), .D(n133[13]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1952__i12 (.Q(\encoder0_position[12] ), .C(n1779), 
            .E(position_31__N_3836), .D(n133[12]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1952__i11 (.Q(\encoder0_position[11] ), .C(n1779), 
            .E(position_31__N_3836), .D(n133[11]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1952__i10 (.Q(\encoder0_position[10] ), .C(n1779), 
            .E(position_31__N_3836), .D(n133[10]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1952__i9 (.Q(\encoder0_position[9] ), .C(n1779), .E(position_31__N_3836), 
            .D(n133[9]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1952__i8 (.Q(\encoder0_position[8] ), .C(n1779), .E(position_31__N_3836), 
            .D(n133[8]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1952__i7 (.Q(\encoder0_position[7] ), .C(n1779), .E(position_31__N_3836), 
            .D(n133[7]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1952__i6 (.Q(\encoder0_position[6] ), .C(n1779), .E(position_31__N_3836), 
            .D(n133[6]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1952__i5 (.Q(\encoder0_position[5] ), .C(n1779), .E(position_31__N_3836), 
            .D(n133[5]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1952__i4 (.Q(\encoder0_position[4] ), .C(n1779), .E(position_31__N_3836), 
            .D(n133[4]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1952__i3 (.Q(\encoder0_position[3] ), .C(n1779), .E(position_31__N_3836), 
            .D(n133[3]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1952__i2 (.Q(\encoder0_position[2] ), .C(n1779), .E(position_31__N_3836), 
            .D(n133[2]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1952__i1 (.Q(\encoder0_position[1] ), .C(n1779), .E(position_31__N_3836), 
            .D(n133[1]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1952__i0 (.Q(\encoder0_position[0] ), .C(n1779), .E(position_31__N_3836), 
            .D(n133[0]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFF a_new_i1 (.Q(\a_new[1] ), .C(n1779), .D(a_new[0]));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_DFF b_new_i1 (.Q(\b_new[1] ), .C(n1779), .D(b_new[0]));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_LUT4 position_31__I_938_4_lut (.I0(a_prev), .I1(b_prev), .I2(\a_new[1] ), 
            .I3(\b_new[1] ), .O(position_31__N_3836));   // vhdl/quadrature_decoder.vhd(63[11:57])
    defparam position_31__I_938_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 debounce_cnt_I_937_4_lut (.I0(a_new[0]), .I1(b_new[0]), .I2(\a_new[1] ), 
            .I3(\b_new[1] ), .O(debounce_cnt_N_3833));   // vhdl/quadrature_decoder.vhd(53[8:58])
    defparam debounce_cnt_I_937_4_lut.LUT_INIT = 16'h7bde;
    
endmodule
//
// Verilog Description of module TLI4970
//

module TLI4970 (\state[1] , GND_net, clk16MHz, VCC_net, n6, n5, 
            n11, n15, \state[0] , \data[12] , n29622, \data[15] , 
            clk_out, CS_c, CS_CLK_c, n29602, n9, n29567, n29565, 
            \current[0] , n29563, \data[11] , n29562, \data[10] , 
            n29550, \data[9] , n29549, \data[8] , n29548, \data[7] , 
            n29547, \data[6] , n29546, \data[5] , n29545, \data[4] , 
            n29538, \data[3] , n29530, \data[2] , n29529, \data[1] , 
            n25499, n4, n25508, n30424, \data[0] , n30319, \current[1] , 
            n30318, \current[2] , n30317, \current[3] , n30316, \current[4] , 
            n30315, \current[5] , n30313, \current[6] , n30312, \current[7] , 
            n30311, \current[8] , n30310, \current[9] , n30309, \current[10] , 
            n30308, \current[11] , n25504, n25512, n27643, \current[15] , 
            n6_adj_7, n5_adj_8, n5_adj_9, n6_adj_10, state_7__N_4319, 
            n42981) /* synthesis syn_noprune=1, syn_module_defined=1 */ ;
    output \state[1] ;
    input GND_net;
    input clk16MHz;
    input VCC_net;
    output n6;
    output n5;
    output n11;
    output n15;
    output \state[0] ;
    output \data[12] ;
    input n29622;
    output \data[15] ;
    output clk_out;
    output CS_c;
    output CS_CLK_c;
    input n29602;
    input n9;
    input n29567;
    input n29565;
    output \current[0] ;
    input n29563;
    output \data[11] ;
    input n29562;
    output \data[10] ;
    input n29550;
    output \data[9] ;
    input n29549;
    output \data[8] ;
    input n29548;
    output \data[7] ;
    input n29547;
    output \data[6] ;
    input n29546;
    output \data[5] ;
    input n29545;
    output \data[4] ;
    input n29538;
    output \data[3] ;
    input n29530;
    output \data[2] ;
    input n29529;
    output \data[1] ;
    output n25499;
    output n4;
    output n25508;
    input n30424;
    output \data[0] ;
    input n30319;
    output \current[1] ;
    input n30318;
    output \current[2] ;
    input n30317;
    output \current[3] ;
    input n30316;
    output \current[4] ;
    input n30315;
    output \current[5] ;
    input n30313;
    output \current[6] ;
    input n30312;
    output \current[7] ;
    input n30311;
    output \current[8] ;
    input n30310;
    output \current[9] ;
    input n30309;
    output \current[10] ;
    input n30308;
    output \current[11] ;
    output n25504;
    output n25512;
    output n27643;
    output \current[15] ;
    output n6_adj_7;
    output n5_adj_8;
    output n5_adj_9;
    output n6_adj_10;
    output state_7__N_4319;
    output n42981;
    
    wire clk_slow /* synthesis is_clock=1, SET_AS_NETWORK=\tli/clk_slow */ ;   // verilog/tli4970.v(11[7:15])
    wire clk16MHz /* synthesis SET_AS_NETWORK=clk16MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    
    wire n12167, n27924, n28816;
    wire [7:0]counter;   // verilog/tli4970.v(12[13:20])
    
    wire clk_slow_N_4233, clk_slow_N_4232;
    wire [2:0]n17;
    
    wire n52375, n52374;
    wire [11:0]n53;
    wire [15:0]delay_counter;   // verilog/tli4970.v(28[14:27])
    
    wire n52373, n52372, n52371, n52370, n52369, n52368, n52367, 
        n52366, n52365, n52364, n52363;
    wire [7:0]bit_counter;   // verilog/tli4970.v(26[13:24])
    
    wire n6_adj_4450, n8, n12, n10, delay_counter_15__N_4314;
    wire [1:0]n1859;
    
    wire n22550, n27696;
    wire [7:0]n37;
    
    wire n29087, n22552, n22554, n22556, n43529, n52269, n52268, 
        n52267, n52266, n67045, n52265, n2, n67041, n52264, n67039, 
        n52263, n67046;
    
    SB_DFFNESR state_i1 (.Q(\state[1] ), .C(clk_slow), .E(n27924), .D(n12167), 
            .R(n28816));   // verilog/tli4970.v(35[10] 68[6])
    SB_LUT4 i2061_3_lut (.I0(counter[0]), .I1(counter[2]), .I2(counter[1]), 
            .I3(GND_net), .O(clk_slow_N_4233));
    defparam i2061_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 clk_slow_I_0_72_2_lut (.I0(clk_slow), .I1(clk_slow_N_4233), 
            .I2(GND_net), .I3(GND_net), .O(clk_slow_N_4232));   // verilog/tli4970.v(15[5] 18[8])
    defparam clk_slow_I_0_72_2_lut.LUT_INIT = 16'h6666;
    SB_DFF clk_slow_63 (.Q(clk_slow), .C(clk16MHz), .D(clk_slow_N_4232));   // verilog/tli4970.v(13[10] 19[6])
    SB_LUT4 counter_1944_1945_add_4_4_lut (.I0(GND_net), .I1(GND_net), .I2(counter[2]), 
            .I3(n52375), .O(n17[2])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1944_1945_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 counter_1944_1945_add_4_3_lut (.I0(GND_net), .I1(GND_net), .I2(counter[1]), 
            .I3(n52374), .O(n17[1])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1944_1945_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_1944_1945_add_4_3 (.CI(n52374), .I0(GND_net), .I1(counter[1]), 
            .CO(n52375));
    SB_LUT4 counter_1944_1945_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(counter[0]), 
            .I3(VCC_net), .O(n17[0])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1944_1945_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_1944_1945_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(counter[0]), 
            .CO(n52374));
    SB_LUT4 delay_counter_1942_1943_add_4_13_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[11]), .I3(n52373), .O(n53[11])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_1942_1943_add_4_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 delay_counter_1942_1943_add_4_12_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[10]), .I3(n52372), .O(n53[10])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_1942_1943_add_4_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_1942_1943_add_4_12 (.CI(n52372), .I0(GND_net), 
            .I1(delay_counter[10]), .CO(n52373));
    SB_LUT4 delay_counter_1942_1943_add_4_11_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[9]), .I3(n52371), .O(n53[9])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_1942_1943_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_1942_1943_add_4_11 (.CI(n52371), .I0(GND_net), 
            .I1(delay_counter[9]), .CO(n52372));
    SB_LUT4 delay_counter_1942_1943_add_4_10_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[8]), .I3(n52370), .O(n53[8])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_1942_1943_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_1942_1943_add_4_10 (.CI(n52370), .I0(GND_net), 
            .I1(delay_counter[8]), .CO(n52371));
    SB_LUT4 delay_counter_1942_1943_add_4_9_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[7]), .I3(n52369), .O(n53[7])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_1942_1943_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_1942_1943_add_4_9 (.CI(n52369), .I0(GND_net), 
            .I1(delay_counter[7]), .CO(n52370));
    SB_LUT4 delay_counter_1942_1943_add_4_8_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[6]), .I3(n52368), .O(n53[6])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_1942_1943_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_1942_1943_add_4_8 (.CI(n52368), .I0(GND_net), 
            .I1(delay_counter[6]), .CO(n52369));
    SB_LUT4 delay_counter_1942_1943_add_4_7_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[5]), .I3(n52367), .O(n53[5])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_1942_1943_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_1942_1943_add_4_7 (.CI(n52367), .I0(GND_net), 
            .I1(delay_counter[5]), .CO(n52368));
    SB_LUT4 delay_counter_1942_1943_add_4_6_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[4]), .I3(n52366), .O(n53[4])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_1942_1943_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_1942_1943_add_4_6 (.CI(n52366), .I0(GND_net), 
            .I1(delay_counter[4]), .CO(n52367));
    SB_LUT4 delay_counter_1942_1943_add_4_5_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[3]), .I3(n52365), .O(n53[3])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_1942_1943_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_1942_1943_add_4_5 (.CI(n52365), .I0(GND_net), 
            .I1(delay_counter[3]), .CO(n52366));
    SB_LUT4 delay_counter_1942_1943_add_4_4_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[2]), .I3(n52364), .O(n53[2])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_1942_1943_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_1942_1943_add_4_4 (.CI(n52364), .I0(GND_net), 
            .I1(delay_counter[2]), .CO(n52365));
    SB_LUT4 delay_counter_1942_1943_add_4_3_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[1]), .I3(n52363), .O(n53[1])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_1942_1943_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_1942_1943_add_4_3 (.CI(n52363), .I0(GND_net), 
            .I1(delay_counter[1]), .CO(n52364));
    SB_LUT4 delay_counter_1942_1943_add_4_2_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[0]), .I3(VCC_net), .O(n53[0])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_1942_1943_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_1942_1943_add_4_2 (.CI(VCC_net), .I0(GND_net), 
            .I1(delay_counter[0]), .CO(n52363));
    SB_LUT4 equal_335_i6_2_lut (.I0(bit_counter[2]), .I1(bit_counter[3]), 
            .I2(GND_net), .I3(GND_net), .O(n6));   // verilog/tli4970.v(54[9:26])
    defparam equal_335_i6_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 equal_326_i5_2_lut (.I0(bit_counter[0]), .I1(bit_counter[1]), 
            .I2(GND_net), .I3(GND_net), .O(n5));   // verilog/tli4970.v(54[9:26])
    defparam equal_326_i5_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut (.I0(bit_counter[5]), .I1(bit_counter[4]), .I2(GND_net), 
            .I3(GND_net), .O(n6_adj_4450));   // verilog/tli4970.v(56[12:26])
    defparam i1_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i4_4_lut (.I0(bit_counter[6]), .I1(n11), .I2(bit_counter[7]), 
            .I3(n6_adj_4450), .O(n15));   // verilog/tli4970.v(56[12:26])
    defparam i4_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i3_3_lut (.I0(delay_counter[1]), .I1(delay_counter[2]), .I2(delay_counter[4]), 
            .I3(GND_net), .O(n8));
    defparam i3_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i2062_4_lut (.I0(delay_counter[3]), .I1(delay_counter[5]), .I2(n8), 
            .I3(delay_counter[0]), .O(n12));
    defparam i2062_4_lut.LUT_INIT = 16'hccc8;
    SB_LUT4 i4_4_lut_adj_958 (.I0(delay_counter[11]), .I1(delay_counter[7]), 
            .I2(delay_counter[8]), .I3(delay_counter[9]), .O(n10));
    defparam i4_4_lut_adj_958.LUT_INIT = 16'h8000;
    SB_LUT4 i5_4_lut (.I0(delay_counter[10]), .I1(n10), .I2(n12), .I3(delay_counter[6]), 
            .O(delay_counter_15__N_4314));
    defparam i5_4_lut.LUT_INIT = 16'h8880;
    SB_LUT4 mux_2029_i2_3_lut (.I0(n15), .I1(\state[1] ), .I2(\state[0] ), 
            .I3(GND_net), .O(n12167));
    defparam mux_2029_i2_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i2117_1_lut (.I0(\data[12] ), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1859[0]));
    defparam i2117_1_lut.LUT_INIT = 16'h5555;
    SB_DFFN data_i15 (.Q(\data[15] ), .C(clk_slow), .D(n29622));   // verilog/tli4970.v(35[10] 68[6])
    SB_LUT4 spi_clk_I_0_i1_3_lut (.I0(clk_slow), .I1(clk_out), .I2(CS_c), 
            .I3(GND_net), .O(CS_CLK_c));   // verilog/tli4970.v(23[20:53])
    defparam spi_clk_I_0_i1_3_lut.LUT_INIT = 16'hc8c8;
    SB_DFFN data_i12 (.Q(\data[12] ), .C(clk_slow), .D(n29602));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN clk_out_67 (.Q(clk_out), .C(clk_slow), .D(n9));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN slave_select_66 (.Q(CS_c), .C(clk_slow), .D(n29567));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i1 (.Q(\current[0] ), .C(clk_slow), .D(n29565));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i11 (.Q(\data[11] ), .C(clk_slow), .D(n29563));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i10 (.Q(\data[10] ), .C(clk_slow), .D(n29562));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i9 (.Q(\data[9] ), .C(clk_slow), .D(n29550));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i8 (.Q(\data[8] ), .C(clk_slow), .D(n29549));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i7 (.Q(\data[7] ), .C(clk_slow), .D(n29548));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i6 (.Q(\data[6] ), .C(clk_slow), .D(n29547));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i5 (.Q(\data[5] ), .C(clk_slow), .D(n29546));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i4 (.Q(\data[4] ), .C(clk_slow), .D(n29545));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i3 (.Q(\data[3] ), .C(clk_slow), .D(n29538));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i2 (.Q(\data[2] ), .C(clk_slow), .D(n29530));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i1 (.Q(\data[1] ), .C(clk_slow), .D(n29529));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFNE bit_counter_1936__i0 (.Q(bit_counter[0]), .C(clk_slow), .E(n27696), 
            .D(n22550));   // verilog/tli4970.v(55[24:39])
    SB_DFFNSR delay_counter_1942_1943__i1 (.Q(delay_counter[0]), .C(clk_slow), 
            .D(n53[0]), .R(delay_counter_15__N_4314));   // verilog/tli4970.v(40[24:39])
    SB_DFFSR counter_1944_1945__i1 (.Q(counter[0]), .C(clk16MHz), .D(n17[0]), 
            .R(clk_slow_N_4233));   // verilog/tli4970.v(14[16:27])
    SB_DFFSR counter_1944_1945__i3 (.Q(counter[2]), .C(clk16MHz), .D(n17[2]), 
            .R(clk_slow_N_4233));   // verilog/tli4970.v(14[16:27])
    SB_DFFSR counter_1944_1945__i2 (.Q(counter[1]), .C(clk16MHz), .D(n17[1]), 
            .R(clk_slow_N_4233));   // verilog/tli4970.v(14[16:27])
    SB_DFFNSR delay_counter_1942_1943__i12 (.Q(delay_counter[11]), .C(clk_slow), 
            .D(n53[11]), .R(delay_counter_15__N_4314));   // verilog/tli4970.v(40[24:39])
    SB_DFFNSR delay_counter_1942_1943__i11 (.Q(delay_counter[10]), .C(clk_slow), 
            .D(n53[10]), .R(delay_counter_15__N_4314));   // verilog/tli4970.v(40[24:39])
    SB_DFFNSR delay_counter_1942_1943__i10 (.Q(delay_counter[9]), .C(clk_slow), 
            .D(n53[9]), .R(delay_counter_15__N_4314));   // verilog/tli4970.v(40[24:39])
    SB_DFFNSR delay_counter_1942_1943__i9 (.Q(delay_counter[8]), .C(clk_slow), 
            .D(n53[8]), .R(delay_counter_15__N_4314));   // verilog/tli4970.v(40[24:39])
    SB_DFFNSR delay_counter_1942_1943__i8 (.Q(delay_counter[7]), .C(clk_slow), 
            .D(n53[7]), .R(delay_counter_15__N_4314));   // verilog/tli4970.v(40[24:39])
    SB_DFFNSR delay_counter_1942_1943__i7 (.Q(delay_counter[6]), .C(clk_slow), 
            .D(n53[6]), .R(delay_counter_15__N_4314));   // verilog/tli4970.v(40[24:39])
    SB_DFFNSR delay_counter_1942_1943__i6 (.Q(delay_counter[5]), .C(clk_slow), 
            .D(n53[5]), .R(delay_counter_15__N_4314));   // verilog/tli4970.v(40[24:39])
    SB_DFFNSR delay_counter_1942_1943__i5 (.Q(delay_counter[4]), .C(clk_slow), 
            .D(n53[4]), .R(delay_counter_15__N_4314));   // verilog/tli4970.v(40[24:39])
    SB_DFFNSR delay_counter_1942_1943__i4 (.Q(delay_counter[3]), .C(clk_slow), 
            .D(n53[3]), .R(delay_counter_15__N_4314));   // verilog/tli4970.v(40[24:39])
    SB_DFFNSR delay_counter_1942_1943__i3 (.Q(delay_counter[2]), .C(clk_slow), 
            .D(n53[2]), .R(delay_counter_15__N_4314));   // verilog/tli4970.v(40[24:39])
    SB_DFFNSR delay_counter_1942_1943__i2 (.Q(delay_counter[1]), .C(clk_slow), 
            .D(n53[1]), .R(delay_counter_15__N_4314));   // verilog/tli4970.v(40[24:39])
    SB_DFFNESR bit_counter_1936__i4 (.Q(bit_counter[4]), .C(clk_slow), .E(n27696), 
            .D(n37[4]), .R(n29087));   // verilog/tli4970.v(55[24:39])
    SB_DFFNESR bit_counter_1936__i5 (.Q(bit_counter[5]), .C(clk_slow), .E(n27696), 
            .D(n37[5]), .R(n29087));   // verilog/tli4970.v(55[24:39])
    SB_DFFNESR bit_counter_1936__i6 (.Q(bit_counter[6]), .C(clk_slow), .E(n27696), 
            .D(n37[6]), .R(n29087));   // verilog/tli4970.v(55[24:39])
    SB_DFFNESR bit_counter_1936__i7 (.Q(bit_counter[7]), .C(clk_slow), .E(n27696), 
            .D(n37[7]), .R(n29087));   // verilog/tli4970.v(55[24:39])
    SB_DFFNE bit_counter_1936__i3 (.Q(bit_counter[3]), .C(clk_slow), .E(n27696), 
            .D(n22552));   // verilog/tli4970.v(55[24:39])
    SB_DFFNE bit_counter_1936__i2 (.Q(bit_counter[2]), .C(clk_slow), .E(n27696), 
            .D(n22554));   // verilog/tli4970.v(55[24:39])
    SB_DFFNE bit_counter_1936__i1 (.Q(bit_counter[1]), .C(clk_slow), .E(n27696), 
            .D(n22556));   // verilog/tli4970.v(55[24:39])
    SB_LUT4 i2_3_lut_4_lut (.I0(bit_counter[0]), .I1(bit_counter[1]), .I2(\state[0] ), 
            .I3(\state[1] ), .O(n25499));
    defparam i2_3_lut_4_lut.LUT_INIT = 16'hf7ff;
    SB_LUT4 i1_2_lut_4_lut (.I0(\state[0] ), .I1(\state[1] ), .I2(bit_counter[2]), 
            .I3(bit_counter[3]), .O(n4));   // verilog/tli4970.v(43[5] 67[12])
    defparam i1_2_lut_4_lut.LUT_INIT = 16'hbfff;
    SB_LUT4 i1_2_lut_4_lut_adj_959 (.I0(\state[0] ), .I1(\state[1] ), .I2(bit_counter[2]), 
            .I3(bit_counter[3]), .O(n25508));   // verilog/tli4970.v(43[5] 67[12])
    defparam i1_2_lut_4_lut_adj_959.LUT_INIT = 16'hfbff;
    SB_DFFN data_i0 (.Q(\data[0] ), .C(clk_slow), .D(n30424));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i2 (.Q(\current[1] ), .C(clk_slow), .D(n30319));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i3 (.Q(\current[2] ), .C(clk_slow), .D(n30318));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i4 (.Q(\current[3] ), .C(clk_slow), .D(n30317));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i5 (.Q(\current[4] ), .C(clk_slow), .D(n30316));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i6 (.Q(\current[5] ), .C(clk_slow), .D(n30315));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i7 (.Q(\current[6] ), .C(clk_slow), .D(n30313));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i8 (.Q(\current[7] ), .C(clk_slow), .D(n30312));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i9 (.Q(\current[8] ), .C(clk_slow), .D(n30311));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i10 (.Q(\current[9] ), .C(clk_slow), .D(n30310));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i11 (.Q(\current[10] ), .C(clk_slow), .D(n30309));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i12 (.Q(\current[11] ), .C(clk_slow), .D(n30308));   // verilog/tli4970.v(35[10] 68[6])
    SB_LUT4 i1_2_lut_4_lut_adj_960 (.I0(\state[0] ), .I1(\state[1] ), .I2(bit_counter[2]), 
            .I3(bit_counter[3]), .O(n25504));   // verilog/tli4970.v(43[5] 67[12])
    defparam i1_2_lut_4_lut_adj_960.LUT_INIT = 16'hffbf;
    SB_LUT4 i1_2_lut_4_lut_adj_961 (.I0(\state[0] ), .I1(\state[1] ), .I2(bit_counter[2]), 
            .I3(bit_counter[3]), .O(n25512));   // verilog/tli4970.v(43[5] 67[12])
    defparam i1_2_lut_4_lut_adj_961.LUT_INIT = 16'hfffb;
    SB_DFFNE current__i13 (.Q(\current[15] ), .C(clk_slow), .E(n27643), 
            .D(n1859[0]));   // verilog/tli4970.v(35[10] 68[6])
    SB_LUT4 i15082_2_lut_2_lut (.I0(\state[1] ), .I1(\state[0] ), .I2(GND_net), 
            .I3(GND_net), .O(n29087));   // verilog/tli4970.v(55[24:39])
    defparam i15082_2_lut_2_lut.LUT_INIT = 16'h4444;
    SB_DFFNESS state_i0 (.Q(\state[0] ), .C(clk_slow), .E(n27924), .D(n43529), 
            .S(n28816));   // verilog/tli4970.v(35[10] 68[6])
    SB_LUT4 bit_counter_1936_add_4_9_lut (.I0(GND_net), .I1(VCC_net), .I2(bit_counter[7]), 
            .I3(n52269), .O(n37[7])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_counter_1936_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 bit_counter_1936_add_4_8_lut (.I0(GND_net), .I1(VCC_net), .I2(bit_counter[6]), 
            .I3(n52268), .O(n37[6])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_counter_1936_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY bit_counter_1936_add_4_8 (.CI(n52268), .I0(VCC_net), .I1(bit_counter[6]), 
            .CO(n52269));
    SB_LUT4 bit_counter_1936_add_4_7_lut (.I0(GND_net), .I1(VCC_net), .I2(bit_counter[5]), 
            .I3(n52267), .O(n37[5])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_counter_1936_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY bit_counter_1936_add_4_7 (.CI(n52267), .I0(VCC_net), .I1(bit_counter[5]), 
            .CO(n52268));
    SB_LUT4 bit_counter_1936_add_4_6_lut (.I0(GND_net), .I1(VCC_net), .I2(bit_counter[4]), 
            .I3(n52266), .O(n37[4])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_counter_1936_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY bit_counter_1936_add_4_6 (.CI(n52266), .I0(VCC_net), .I1(bit_counter[4]), 
            .CO(n52267));
    SB_LUT4 bit_counter_1936_add_4_5_lut (.I0(n2), .I1(VCC_net), .I2(bit_counter[3]), 
            .I3(n52265), .O(n67045)) /* synthesis syn_instantiated=1 */ ;
    defparam bit_counter_1936_add_4_5_lut.LUT_INIT = 16'h8228;
    SB_CARRY bit_counter_1936_add_4_5 (.CI(n52265), .I0(VCC_net), .I1(bit_counter[3]), 
            .CO(n52266));
    SB_LUT4 bit_counter_1936_add_4_4_lut (.I0(n2), .I1(VCC_net), .I2(bit_counter[2]), 
            .I3(n52264), .O(n67041)) /* synthesis syn_instantiated=1 */ ;
    defparam bit_counter_1936_add_4_4_lut.LUT_INIT = 16'h8228;
    SB_CARRY bit_counter_1936_add_4_4 (.CI(n52264), .I0(VCC_net), .I1(bit_counter[2]), 
            .CO(n52265));
    SB_LUT4 bit_counter_1936_add_4_3_lut (.I0(n2), .I1(VCC_net), .I2(bit_counter[1]), 
            .I3(n52263), .O(n67039)) /* synthesis syn_instantiated=1 */ ;
    defparam bit_counter_1936_add_4_3_lut.LUT_INIT = 16'h8228;
    SB_CARRY bit_counter_1936_add_4_3 (.CI(n52263), .I0(VCC_net), .I1(bit_counter[1]), 
            .CO(n52264));
    SB_LUT4 bit_counter_1936_add_4_2_lut (.I0(n2), .I1(GND_net), .I2(bit_counter[0]), 
            .I3(VCC_net), .O(n67046)) /* synthesis syn_instantiated=1 */ ;
    defparam bit_counter_1936_add_4_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY bit_counter_1936_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(bit_counter[0]), 
            .CO(n52263));
    SB_LUT4 i2389_1_lut (.I0(\state[0] ), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2));
    defparam i2389_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_2_lut_4_lut_adj_962 (.I0(n15), .I1(\state[0] ), .I2(\state[1] ), 
            .I3(delay_counter_15__N_4314), .O(n27924));
    defparam i1_2_lut_4_lut_adj_962.LUT_INIT = 16'hffdc;
    SB_LUT4 i14810_2_lut_4_lut (.I0(n15), .I1(\state[0] ), .I2(\state[1] ), 
            .I3(delay_counter_15__N_4314), .O(n28816));
    defparam i14810_2_lut_4_lut.LUT_INIT = 16'h2300;
    SB_LUT4 i8813_3_lut (.I0(\state[0] ), .I1(n67039), .I2(\state[1] ), 
            .I3(GND_net), .O(n22556));   // verilog/tli4970.v(55[24:39])
    defparam i8813_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8811_3_lut (.I0(\state[0] ), .I1(n67041), .I2(\state[1] ), 
            .I3(GND_net), .O(n22554));   // verilog/tli4970.v(55[24:39])
    defparam i8811_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8809_3_lut (.I0(\state[0] ), .I1(n67045), .I2(\state[1] ), 
            .I3(GND_net), .O(n22552));   // verilog/tli4970.v(55[24:39])
    defparam i8809_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13957_2_lut (.I0(\state[1] ), .I1(\state[0] ), .I2(GND_net), 
            .I3(GND_net), .O(n27696));
    defparam i13957_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i8807_3_lut (.I0(\state[0] ), .I1(n67046), .I2(\state[1] ), 
            .I3(GND_net), .O(n22550));   // verilog/tli4970.v(55[24:39])
    defparam i8807_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 equal_333_i6_2_lut (.I0(bit_counter[2]), .I1(bit_counter[3]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_7));   // verilog/tli4970.v(54[9:26])
    defparam equal_333_i6_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 equal_325_i5_2_lut (.I0(bit_counter[0]), .I1(bit_counter[1]), 
            .I2(GND_net), .I3(GND_net), .O(n5_adj_8));   // verilog/tli4970.v(54[9:26])
    defparam equal_325_i5_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 equal_264_i11_2_lut_4_lut (.I0(bit_counter[0]), .I1(bit_counter[1]), 
            .I2(bit_counter[2]), .I3(bit_counter[3]), .O(n11));   // verilog/tli4970.v(56[12:26])
    defparam equal_264_i11_2_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 equal_324_i5_2_lut (.I0(bit_counter[0]), .I1(bit_counter[1]), 
            .I2(GND_net), .I3(GND_net), .O(n5_adj_9));   // verilog/tli4970.v(54[9:26])
    defparam equal_324_i5_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 equal_328_i6_2_lut (.I0(bit_counter[2]), .I1(bit_counter[3]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_10));   // verilog/tli4970.v(54[9:26])
    defparam equal_328_i6_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 i54366_3_lut (.I0(\data[15] ), .I1(\state[1] ), .I2(\state[0] ), 
            .I3(GND_net), .O(n27643));
    defparam i54366_3_lut.LUT_INIT = 16'h4040;
    SB_LUT4 state_7__I_0_77_i9_2_lut (.I0(\state[0] ), .I1(\state[1] ), 
            .I2(GND_net), .I3(GND_net), .O(state_7__N_4319));   // verilog/tli4970.v(53[7:17])
    defparam state_7__I_0_77_i9_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 i29089_2_lut (.I0(bit_counter[2]), .I1(bit_counter[3]), .I2(GND_net), 
            .I3(GND_net), .O(n42981));
    defparam i29089_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i54383_2_lut (.I0(n15), .I1(\state[0] ), .I2(GND_net), .I3(GND_net), 
            .O(n43529));
    defparam i54383_2_lut.LUT_INIT = 16'h1111;
    
endmodule
//
// Verilog Description of module EEPROM
//

module EEPROM (n25391, \state[0] , \state[1] , enable_slow_N_4213, n5771, 
            ready_prev, clk16MHz, \state[2] , GND_net, n43543, \state_7__N_3918[0] , 
            n42885, n29566, rw, n58190, data_ready, ID, n57800, 
            n58002, baudrate, n30330, n30329, n30328, n30327, n30326, 
            n30325, n30324, n30323, \state[0]_adj_3 , n58751, n4, 
            data, n61888, n25490, scl_enable, \state_7__N_4110[0] , 
            VCC_net, scl, sda_enable, sda_out, n29573, \saved_addr[0] , 
            n6426, n30410, n8, n30134, n30133, n30132, n30131, 
            n30130, n30129, n30128, n4_adj_4, n4_adj_5, n42994, 
            n6, \state_7__N_4126[3] , n10, n25522, n25517, n10_adj_6) /* synthesis syn_noprune=1, syn_module_defined=1 */ ;
    output n25391;
    output \state[0] ;
    output \state[1] ;
    output enable_slow_N_4213;
    output [0:0]n5771;
    output ready_prev;
    input clk16MHz;
    output \state[2] ;
    input GND_net;
    output n43543;
    input \state_7__N_3918[0] ;
    output n42885;
    input n29566;
    output rw;
    input n58190;
    output data_ready;
    output [7:0]ID;
    input n57800;
    input n58002;
    output [31:0]baudrate;
    input n30330;
    input n30329;
    input n30328;
    input n30327;
    input n30326;
    input n30325;
    input n30324;
    input n30323;
    output \state[0]_adj_3 ;
    output n58751;
    output n4;
    output [7:0]data;
    output n61888;
    output n25490;
    output scl_enable;
    output \state_7__N_4110[0] ;
    input VCC_net;
    output scl;
    output sda_enable;
    output sda_out;
    input n29573;
    output \saved_addr[0] ;
    output n6426;
    input n30410;
    input n8;
    input n30134;
    input n30133;
    input n30132;
    input n30131;
    input n30130;
    input n30129;
    input n30128;
    output n4_adj_4;
    output n4_adj_5;
    output n42994;
    output n6;
    input \state_7__N_4126[3] ;
    output n10;
    output n25522;
    output n25517;
    output n10_adj_6;
    
    wire clk16MHz /* synthesis SET_AS_NETWORK=clk16MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    wire [15:0]delay_counter;   // verilog/eeprom.v(28[12:25])
    
    wire n28, n26, n27, n25, enable;
    wire [15:0]delay_counter_15__N_3956;
    wire [15:0]n5111;
    
    wire n51261, n51260, n51259, n51258, n51257, n6685, n51256, 
        n43433, n6684, n51255, n6683, n51254, n6682, n51253, n6681, 
        n51252, n51251, n6679, n51250, n51249, n51248, n51247;
    wire [2:0]byte_counter;   // verilog/eeprom.v(30[11:23])
    
    wire n4_c, n63957;
    wire [7:0]state;   // verilog/i2c_controller.v(33[12:17])
    
    wire n67179, n61588;
    wire [7:0]state_7__N_3885;
    
    wire n29561;
    wire [2:0]n17;
    
    wire n27703, n29084, n53631, n30362, n30361, n30360, n30359, 
        n30358, n30357, n30356, n30355, n30354, n30353, n30352, 
        n30351, n30350, n30348, n30347, n30346, n30345, n30344, 
        n30343, n30342, n30341, n30340, n30339, n30338, n30337, 
        n30336, n30335, n30334, n30333, n30332, n30331, n27634, 
        n28835, n58746, n52727, n58743, n6_c;
    
    SB_LUT4 i12_4_lut (.I0(delay_counter[6]), .I1(delay_counter[10]), .I2(delay_counter[12]), 
            .I3(delay_counter[8]), .O(n28));   // verilog/eeprom.v(55[12:28])
    defparam i12_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i10_4_lut (.I0(delay_counter[11]), .I1(delay_counter[2]), .I2(delay_counter[7]), 
            .I3(delay_counter[5]), .O(n26));   // verilog/eeprom.v(55[12:28])
    defparam i10_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i11_4_lut (.I0(delay_counter[15]), .I1(delay_counter[3]), .I2(delay_counter[14]), 
            .I3(delay_counter[1]), .O(n27));   // verilog/eeprom.v(55[12:28])
    defparam i11_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i9_4_lut (.I0(delay_counter[4]), .I1(delay_counter[9]), .I2(delay_counter[13]), 
            .I3(delay_counter[0]), .O(n25));   // verilog/eeprom.v(55[12:28])
    defparam i9_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut (.I0(n25), .I1(n27), .I2(n26), .I3(n28), .O(n25391));   // verilog/eeprom.v(55[12:28])
    defparam i15_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 mux_1448_Mux_0_i3_4_lut (.I0(\state[0] ), .I1(n25391), .I2(\state[1] ), 
            .I3(enable_slow_N_4213), .O(n5771[0]));   // verilog/eeprom.v(38[3] 80[10])
    defparam mux_1448_Mux_0_i3_4_lut.LUT_INIT = 16'h1a0a;
    SB_DFF ready_prev_59 (.Q(ready_prev), .C(clk16MHz), .D(enable_slow_N_4213));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFSR enable_58 (.Q(enable), .C(clk16MHz), .D(n5771[0]), .R(\state[2] ));   // verilog/eeprom.v(35[8] 81[4])
    SB_LUT4 add_1101_17_lut (.I0(GND_net), .I1(delay_counter[15]), .I2(n5111[11]), 
            .I3(n51261), .O(delay_counter_15__N_3956[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1101_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_1101_16_lut (.I0(GND_net), .I1(delay_counter[14]), .I2(n5111[11]), 
            .I3(n51260), .O(delay_counter_15__N_3956[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1101_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1101_16 (.CI(n51260), .I0(delay_counter[14]), .I1(n5111[11]), 
            .CO(n51261));
    SB_LUT4 add_1101_15_lut (.I0(GND_net), .I1(delay_counter[13]), .I2(n5111[11]), 
            .I3(n51259), .O(delay_counter_15__N_3956[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1101_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1101_15 (.CI(n51259), .I0(delay_counter[13]), .I1(n5111[11]), 
            .CO(n51260));
    SB_LUT4 add_1101_14_lut (.I0(GND_net), .I1(delay_counter[12]), .I2(n5111[11]), 
            .I3(n51258), .O(delay_counter_15__N_3956[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1101_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1101_14 (.CI(n51258), .I0(delay_counter[12]), .I1(n5111[11]), 
            .CO(n51259));
    SB_LUT4 add_1101_13_lut (.I0(GND_net), .I1(delay_counter[11]), .I2(n5111[11]), 
            .I3(n51257), .O(delay_counter_15__N_3956[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1101_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1101_13 (.CI(n51257), .I0(delay_counter[11]), .I1(n5111[11]), 
            .CO(n51258));
    SB_LUT4 add_1101_12_lut (.I0(n43433), .I1(delay_counter[10]), .I2(n5111[11]), 
            .I3(n51256), .O(n6685)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1101_12_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_1101_12 (.CI(n51256), .I0(delay_counter[10]), .I1(n5111[11]), 
            .CO(n51257));
    SB_LUT4 add_1101_11_lut (.I0(n43433), .I1(delay_counter[9]), .I2(n5111[11]), 
            .I3(n51255), .O(n6684)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1101_11_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_1101_11 (.CI(n51255), .I0(delay_counter[9]), .I1(n5111[11]), 
            .CO(n51256));
    SB_LUT4 add_1101_10_lut (.I0(n43433), .I1(delay_counter[8]), .I2(n5111[11]), 
            .I3(n51254), .O(n6683)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1101_10_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_1101_10 (.CI(n51254), .I0(delay_counter[8]), .I1(n5111[11]), 
            .CO(n51255));
    SB_LUT4 add_1101_9_lut (.I0(n43433), .I1(delay_counter[7]), .I2(n5111[11]), 
            .I3(n51253), .O(n6682)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1101_9_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_1101_9 (.CI(n51253), .I0(delay_counter[7]), .I1(n5111[11]), 
            .CO(n51254));
    SB_LUT4 add_1101_8_lut (.I0(n43433), .I1(delay_counter[6]), .I2(n5111[11]), 
            .I3(n51252), .O(n6681)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1101_8_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_1101_8 (.CI(n51252), .I0(delay_counter[6]), .I1(n5111[11]), 
            .CO(n51253));
    SB_LUT4 add_1101_7_lut (.I0(GND_net), .I1(delay_counter[5]), .I2(n5111[11]), 
            .I3(n51251), .O(delay_counter_15__N_3956[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1101_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1101_7 (.CI(n51251), .I0(delay_counter[5]), .I1(n5111[11]), 
            .CO(n51252));
    SB_LUT4 add_1101_6_lut (.I0(n43433), .I1(delay_counter[4]), .I2(n5111[11]), 
            .I3(n51250), .O(n6679)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1101_6_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_1101_6 (.CI(n51250), .I0(delay_counter[4]), .I1(n5111[11]), 
            .CO(n51251));
    SB_LUT4 add_1101_5_lut (.I0(GND_net), .I1(delay_counter[3]), .I2(n5111[11]), 
            .I3(n51249), .O(delay_counter_15__N_3956[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1101_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1101_5 (.CI(n51249), .I0(delay_counter[3]), .I1(n5111[11]), 
            .CO(n51250));
    SB_LUT4 add_1101_4_lut (.I0(GND_net), .I1(delay_counter[2]), .I2(n5111[11]), 
            .I3(n51248), .O(delay_counter_15__N_3956[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1101_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1101_4 (.CI(n51248), .I0(delay_counter[2]), .I1(n5111[11]), 
            .CO(n51249));
    SB_LUT4 add_1101_3_lut (.I0(GND_net), .I1(delay_counter[1]), .I2(n5111[11]), 
            .I3(n51247), .O(delay_counter_15__N_3956[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1101_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1101_3 (.CI(n51247), .I0(delay_counter[1]), .I1(n5111[11]), 
            .CO(n51248));
    SB_LUT4 add_1101_2_lut (.I0(GND_net), .I1(delay_counter[0]), .I2(n5111[11]), 
            .I3(GND_net), .O(delay_counter_15__N_3956[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1101_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1101_2 (.CI(GND_net), .I0(delay_counter[0]), .I1(n5111[11]), 
            .CO(n51247));
    SB_LUT4 i29649_3_lut (.I0(byte_counter[0]), .I1(byte_counter[2]), .I2(byte_counter[1]), 
            .I3(GND_net), .O(n43543));
    defparam i29649_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i54385_2_lut (.I0(n25391), .I1(enable_slow_N_4213), .I2(GND_net), 
            .I3(GND_net), .O(n5111[11]));   // verilog/eeprom.v(59[18] 61[12])
    defparam i54385_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut (.I0(\state[2] ), .I1(\state[1] ), .I2(\state_7__N_3918[0] ), 
            .I3(\state[0] ), .O(n4_c));
    defparam i1_4_lut.LUT_INIT = 16'hbbba;
    SB_LUT4 i52344_4_lut (.I0(n63957), .I1(n25391), .I2(\state[1] ), .I3(state[3]), 
            .O(n67179));
    defparam i52344_4_lut.LUT_INIT = 16'h0010;
    SB_LUT4 i2_4_lut (.I0(n67179), .I1(n4_c), .I2(n42885), .I3(\state[0] ), 
            .O(n61588));
    defparam i2_4_lut.LUT_INIT = 16'hcfee;
    SB_LUT4 i8907_4_lut (.I0(\state[1] ), .I1(n43543), .I2(\state[2] ), 
            .I3(\state[0] ), .O(state_7__N_3885[1]));   // verilog/eeprom.v(38[3] 80[10])
    defparam i8907_4_lut.LUT_INIT = 16'ha5ba;
    SB_DFF rw_64 (.Q(rw), .C(clk16MHz), .D(n29566));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF data_ready_61 (.Q(data_ready), .C(clk16MHz), .D(n58190));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i1 (.Q(ID[0]), .C(clk16MHz), .D(n29561));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF state_i2 (.Q(\state[2] ), .C(clk16MHz), .D(n57800));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESR byte_counter_1941__i1 (.Q(byte_counter[1]), .C(clk16MHz), 
            .E(n27703), .D(n17[1]), .R(n29084));   // verilog/eeprom.v(68[25:39])
    SB_DFFESR byte_counter_1941__i2 (.Q(byte_counter[2]), .C(clk16MHz), 
            .E(n27703), .D(n17[2]), .R(n29084));   // verilog/eeprom.v(68[25:39])
    SB_DFFESR byte_counter_1941__i0 (.Q(byte_counter[0]), .C(clk16MHz), 
            .E(n27703), .D(n53631), .R(n29084));   // verilog/eeprom.v(68[25:39])
    SB_DFF state_i0 (.Q(\state[0] ), .C(clk16MHz), .D(n58002));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i2 (.Q(ID[1]), .C(clk16MHz), .D(n30362));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i3 (.Q(ID[2]), .C(clk16MHz), .D(n30361));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i4 (.Q(ID[3]), .C(clk16MHz), .D(n30360));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i5 (.Q(ID[4]), .C(clk16MHz), .D(n30359));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i6 (.Q(ID[5]), .C(clk16MHz), .D(n30358));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i7 (.Q(ID[6]), .C(clk16MHz), .D(n30357));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i8 (.Q(ID[7]), .C(clk16MHz), .D(n30356));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i9 (.Q(baudrate[0]), .C(clk16MHz), .D(n30355));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i10 (.Q(baudrate[1]), .C(clk16MHz), .D(n30354));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i11 (.Q(baudrate[2]), .C(clk16MHz), .D(n30353));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i12 (.Q(baudrate[3]), .C(clk16MHz), .D(n30352));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i13 (.Q(baudrate[4]), .C(clk16MHz), .D(n30351));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i14 (.Q(baudrate[5]), .C(clk16MHz), .D(n30350));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i15 (.Q(baudrate[6]), .C(clk16MHz), .D(n30348));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i16 (.Q(baudrate[7]), .C(clk16MHz), .D(n30347));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i17 (.Q(baudrate[8]), .C(clk16MHz), .D(n30346));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i18 (.Q(baudrate[9]), .C(clk16MHz), .D(n30345));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i19 (.Q(baudrate[10]), .C(clk16MHz), .D(n30344));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i20 (.Q(baudrate[11]), .C(clk16MHz), .D(n30343));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i21 (.Q(baudrate[12]), .C(clk16MHz), .D(n30342));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i22 (.Q(baudrate[13]), .C(clk16MHz), .D(n30341));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i23 (.Q(baudrate[14]), .C(clk16MHz), .D(n30340));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i24 (.Q(baudrate[15]), .C(clk16MHz), .D(n30339));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i25 (.Q(baudrate[16]), .C(clk16MHz), .D(n30338));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i26 (.Q(baudrate[17]), .C(clk16MHz), .D(n30337));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i27 (.Q(baudrate[18]), .C(clk16MHz), .D(n30336));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i28 (.Q(baudrate[19]), .C(clk16MHz), .D(n30335));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i29 (.Q(baudrate[20]), .C(clk16MHz), .D(n30334));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i30 (.Q(baudrate[21]), .C(clk16MHz), .D(n30333));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i31 (.Q(baudrate[22]), .C(clk16MHz), .D(n30332));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i32 (.Q(baudrate[23]), .C(clk16MHz), .D(n30331));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i33 (.Q(baudrate[24]), .C(clk16MHz), .D(n30330));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i34 (.Q(baudrate[25]), .C(clk16MHz), .D(n30329));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i35 (.Q(baudrate[26]), .C(clk16MHz), .D(n30328));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i36 (.Q(baudrate[27]), .C(clk16MHz), .D(n30327));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i37 (.Q(baudrate[28]), .C(clk16MHz), .D(n30326));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i38 (.Q(baudrate[29]), .C(clk16MHz), .D(n30325));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i39 (.Q(baudrate[30]), .C(clk16MHz), .D(n30324));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i40 (.Q(baudrate[31]), .C(clk16MHz), .D(n30323));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFE state_i1 (.Q(\state[1] ), .C(clk16MHz), .E(n61588), .D(state_7__N_3885[1]));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESR delay_counter_i0_i15 (.Q(delay_counter[15]), .C(clk16MHz), 
            .E(n27634), .D(delay_counter_15__N_3956[15]), .R(n28835));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESR delay_counter_i0_i14 (.Q(delay_counter[14]), .C(clk16MHz), 
            .E(n27634), .D(delay_counter_15__N_3956[14]), .R(n28835));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESR delay_counter_i0_i13 (.Q(delay_counter[13]), .C(clk16MHz), 
            .E(n27634), .D(delay_counter_15__N_3956[13]), .R(n28835));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESR delay_counter_i0_i12 (.Q(delay_counter[12]), .C(clk16MHz), 
            .E(n27634), .D(delay_counter_15__N_3956[12]), .R(n28835));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESR delay_counter_i0_i11 (.Q(delay_counter[11]), .C(clk16MHz), 
            .E(n27634), .D(delay_counter_15__N_3956[11]), .R(n28835));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESS delay_counter_i0_i10 (.Q(delay_counter[10]), .C(clk16MHz), 
            .E(n27634), .D(n6685), .S(n28835));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESS delay_counter_i0_i9 (.Q(delay_counter[9]), .C(clk16MHz), .E(n27634), 
            .D(n6684), .S(n28835));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESS delay_counter_i0_i8 (.Q(delay_counter[8]), .C(clk16MHz), .E(n27634), 
            .D(n6683), .S(n28835));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESS delay_counter_i0_i7 (.Q(delay_counter[7]), .C(clk16MHz), .E(n27634), 
            .D(n6682), .S(n28835));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESS delay_counter_i0_i6 (.Q(delay_counter[6]), .C(clk16MHz), .E(n27634), 
            .D(n6681), .S(n28835));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESR delay_counter_i0_i5 (.Q(delay_counter[5]), .C(clk16MHz), .E(n27634), 
            .D(delay_counter_15__N_3956[5]), .R(n28835));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESS delay_counter_i0_i4 (.Q(delay_counter[4]), .C(clk16MHz), .E(n27634), 
            .D(n6679), .S(n28835));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESR delay_counter_i0_i3 (.Q(delay_counter[3]), .C(clk16MHz), .E(n27634), 
            .D(delay_counter_15__N_3956[3]), .R(n28835));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESR delay_counter_i0_i2 (.Q(delay_counter[2]), .C(clk16MHz), .E(n27634), 
            .D(delay_counter_15__N_3956[2]), .R(n28835));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESR delay_counter_i0_i1 (.Q(delay_counter[1]), .C(clk16MHz), .E(n27634), 
            .D(delay_counter_15__N_3956[1]), .R(n28835));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESR delay_counter_i0_i0 (.Q(delay_counter[0]), .C(clk16MHz), .E(n27634), 
            .D(delay_counter_15__N_3956[0]), .R(n28835));   // verilog/eeprom.v(35[8] 81[4])
    SB_LUT4 i1_2_lut_3_lut (.I0(enable_slow_N_4213), .I1(ready_prev), .I2(byte_counter[0]), 
            .I3(GND_net), .O(n53631));
    defparam i1_2_lut_3_lut.LUT_INIT = 16'hd2d2;
    SB_LUT4 i2_3_lut_4_lut (.I0(\state[0]_adj_3 ), .I1(state[3]), .I2(state[2]), 
            .I3(state[1]), .O(n58751));   // verilog/eeprom.v(55[12:28])
    defparam i2_3_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_3_lut_4_lut (.I0(\state[0]_adj_3 ), .I1(state[3]), 
            .I2(state[1]), .I3(state[2]), .O(n4));   // verilog/eeprom.v(55[12:28])
    defparam i1_2_lut_3_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i16350_3_lut_4_lut (.I0(byte_counter[0]), .I1(n58746), .I2(data[7]), 
            .I3(ID[7]), .O(n30356));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16350_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16351_3_lut_4_lut (.I0(byte_counter[0]), .I1(n58746), .I2(data[6]), 
            .I3(ID[6]), .O(n30357));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16351_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16352_3_lut_4_lut (.I0(byte_counter[0]), .I1(n58746), .I2(data[5]), 
            .I3(ID[5]), .O(n30358));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16352_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16353_3_lut_4_lut (.I0(byte_counter[0]), .I1(n58746), .I2(data[4]), 
            .I3(ID[4]), .O(n30359));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16353_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16354_3_lut_4_lut (.I0(byte_counter[0]), .I1(n58746), .I2(data[3]), 
            .I3(ID[3]), .O(n30360));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16354_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16355_3_lut_4_lut (.I0(byte_counter[0]), .I1(n58746), .I2(data[2]), 
            .I3(ID[2]), .O(n30361));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16355_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16356_3_lut_4_lut (.I0(byte_counter[0]), .I1(n58746), .I2(data[1]), 
            .I3(ID[1]), .O(n30362));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16356_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15555_3_lut_4_lut (.I0(byte_counter[0]), .I1(n58746), .I2(data[0]), 
            .I3(ID[0]), .O(n29561));   // verilog/eeprom.v(35[8] 81[4])
    defparam i15555_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i3_3_lut_4_lut (.I0(byte_counter[1]), .I1(n52727), .I2(byte_counter[0]), 
            .I3(byte_counter[2]), .O(n61888));
    defparam i3_3_lut_4_lut.LUT_INIT = 16'hfbff;
    SB_LUT4 i2_2_lut_3_lut (.I0(byte_counter[1]), .I1(n52727), .I2(byte_counter[2]), 
            .I3(GND_net), .O(n58746));
    defparam i2_2_lut_3_lut.LUT_INIT = 16'hfbfb;
    SB_LUT4 i54371_3_lut_4_lut_4_lut (.I0(\state[2] ), .I1(n43543), .I2(\state[0] ), 
            .I3(\state[1] ), .O(n27634));
    defparam i54371_3_lut_4_lut_4_lut.LUT_INIT = 16'h0552;
    SB_LUT4 i36978_2_lut_3_lut_4_lut (.I0(enable_slow_N_4213), .I1(ready_prev), 
            .I2(byte_counter[0]), .I3(byte_counter[1]), .O(n17[1]));   // verilog/eeprom.v(68[25:39])
    defparam i36978_2_lut_3_lut_4_lut.LUT_INIT = 16'hdf20;
    SB_LUT4 i2_3_lut_4_lut_adj_956 (.I0(\state_7__N_3918[0] ), .I1(\state[1] ), 
            .I2(\state[0] ), .I3(\state[2] ), .O(n29084));   // verilog/eeprom.v(68[25:39])
    defparam i2_3_lut_4_lut_adj_956.LUT_INIT = 16'h0002;
    SB_LUT4 i1_4_lut_4_lut (.I0(\state_7__N_3918[0] ), .I1(\state[1] ), 
            .I2(\state[0] ), .I3(\state[2] ), .O(n27703));   // verilog/eeprom.v(68[25:39])
    defparam i1_4_lut_4_lut.LUT_INIT = 16'h00c2;
    SB_LUT4 i36985_3_lut_4_lut (.I0(n42885), .I1(byte_counter[0]), .I2(byte_counter[1]), 
            .I3(byte_counter[2]), .O(n17[2]));   // verilog/eeprom.v(68[25:39])
    defparam i36985_3_lut_4_lut.LUT_INIT = 16'hbf40;
    SB_LUT4 i2_3_lut (.I0(byte_counter[2]), .I1(n52727), .I2(byte_counter[1]), 
            .I3(GND_net), .O(n58743));   // verilog/eeprom.v(66[9:28])
    defparam i2_3_lut.LUT_INIT = 16'hbfbf;
    SB_LUT4 i16341_3_lut_4_lut (.I0(byte_counter[0]), .I1(n58746), .I2(data[7]), 
            .I3(baudrate[7]), .O(n30347));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16341_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i16342_3_lut_4_lut (.I0(byte_counter[0]), .I1(n58746), .I2(data[6]), 
            .I3(baudrate[6]), .O(n30348));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16342_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i16344_3_lut_4_lut (.I0(byte_counter[0]), .I1(n58746), .I2(data[5]), 
            .I3(baudrate[5]), .O(n30350));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16344_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i16345_3_lut_4_lut (.I0(byte_counter[0]), .I1(n58746), .I2(data[4]), 
            .I3(baudrate[4]), .O(n30351));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16345_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i16346_3_lut_4_lut (.I0(byte_counter[0]), .I1(n58746), .I2(data[3]), 
            .I3(baudrate[3]), .O(n30352));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16346_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i16347_3_lut_4_lut (.I0(byte_counter[0]), .I1(n58746), .I2(data[2]), 
            .I3(baudrate[2]), .O(n30353));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16347_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i16348_3_lut_4_lut (.I0(byte_counter[0]), .I1(n58746), .I2(data[1]), 
            .I3(baudrate[1]), .O(n30354));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16348_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i16349_3_lut_4_lut (.I0(byte_counter[0]), .I1(n58746), .I2(data[0]), 
            .I3(baudrate[0]), .O(n30355));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16349_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i29540_1_lut_2_lut (.I0(\state[2] ), .I1(n43543), .I2(GND_net), 
            .I3(GND_net), .O(n43433));
    defparam i29540_1_lut_2_lut.LUT_INIT = 16'h7777;
    SB_LUT4 i28993_2_lut (.I0(enable_slow_N_4213), .I1(ready_prev), .I2(GND_net), 
            .I3(GND_net), .O(n42885));
    defparam i28993_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 i16333_3_lut_4_lut (.I0(byte_counter[0]), .I1(n58743), .I2(data[7]), 
            .I3(baudrate[15]), .O(n30339));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16333_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16334_3_lut_4_lut (.I0(byte_counter[0]), .I1(n58743), .I2(data[6]), 
            .I3(baudrate[14]), .O(n30340));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16334_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16335_3_lut_4_lut (.I0(byte_counter[0]), .I1(n58743), .I2(data[5]), 
            .I3(baudrate[13]), .O(n30341));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16335_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16336_3_lut_4_lut (.I0(byte_counter[0]), .I1(n58743), .I2(data[4]), 
            .I3(baudrate[12]), .O(n30342));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16336_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16337_3_lut_4_lut (.I0(byte_counter[0]), .I1(n58743), .I2(data[3]), 
            .I3(baudrate[11]), .O(n30343));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16337_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16338_3_lut_4_lut (.I0(byte_counter[0]), .I1(n58743), .I2(data[2]), 
            .I3(baudrate[10]), .O(n30344));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16338_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16339_3_lut_4_lut (.I0(byte_counter[0]), .I1(n58743), .I2(data[1]), 
            .I3(baudrate[9]), .O(n30345));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16339_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16340_3_lut_4_lut (.I0(byte_counter[0]), .I1(n58743), .I2(data[0]), 
            .I3(baudrate[8]), .O(n30346));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16340_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16325_3_lut_4_lut (.I0(byte_counter[0]), .I1(n58743), .I2(data[7]), 
            .I3(baudrate[23]), .O(n30331));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16325_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i16326_3_lut_4_lut (.I0(byte_counter[0]), .I1(n58743), .I2(data[6]), 
            .I3(baudrate[22]), .O(n30332));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16326_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i16327_3_lut_4_lut (.I0(byte_counter[0]), .I1(n58743), .I2(data[5]), 
            .I3(baudrate[21]), .O(n30333));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16327_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i16328_3_lut_4_lut (.I0(byte_counter[0]), .I1(n58743), .I2(data[4]), 
            .I3(baudrate[20]), .O(n30334));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16328_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i16329_3_lut_4_lut (.I0(byte_counter[0]), .I1(n58743), .I2(data[3]), 
            .I3(baudrate[19]), .O(n30335));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16329_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i16330_3_lut_4_lut (.I0(byte_counter[0]), .I1(n58743), .I2(data[2]), 
            .I3(baudrate[18]), .O(n30336));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16330_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i16331_3_lut_4_lut (.I0(byte_counter[0]), .I1(n58743), .I2(data[1]), 
            .I3(baudrate[17]), .O(n30337));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16331_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i16332_3_lut_4_lut (.I0(byte_counter[0]), .I1(n58743), .I2(data[0]), 
            .I3(baudrate[16]), .O(n30338));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16332_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut (.I0(\state[0] ), .I1(\state[1] ), .I2(GND_net), 
            .I3(GND_net), .O(n6_c));
    defparam i1_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i4_4_lut (.I0(ready_prev), .I1(n58751), .I2(\state[2] ), .I3(n6_c), 
            .O(n52727));
    defparam i4_4_lut.LUT_INIT = 16'h0100;
    SB_LUT4 i1_2_lut_adj_957 (.I0(\state[0] ), .I1(\state[1] ), .I2(GND_net), 
            .I3(GND_net), .O(n25490));   // verilog/eeprom.v(38[3] 80[10])
    defparam i1_2_lut_adj_957.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_4_lut (.I0(\state[2] ), .I1(\state[1] ), .I2(\state[0] ), 
            .I3(n43543), .O(n28835));   // verilog/eeprom.v(35[8] 81[4])
    defparam i1_2_lut_4_lut.LUT_INIT = 16'h1012;
    i2c_controller i2c (.clk16MHz(clk16MHz), .scl_enable(scl_enable), .\state[2] (state[2]), 
            .\state[3] (state[3]), .\state[0] (\state[0]_adj_3 ), .GND_net(GND_net), 
            .\state_7__N_4110[0] (\state_7__N_4110[0] ), .VCC_net(VCC_net), 
            .scl(scl), .\state[1] (state[1]), .enable_slow_N_4213(enable_slow_N_4213), 
            .sda_enable(sda_enable), .sda_out(sda_out), .n29573(n29573), 
            .\saved_addr[0] (\saved_addr[0] ), .n6426(n6426), .n30410(n30410), 
            .data({data}), .n8(n8), .n30134(n30134), .n30133(n30133), 
            .n30132(n30132), .n30131(n30131), .n30130(n30130), .n30129(n30129), 
            .n30128(n30128), .n4(n4_adj_4), .n4_adj_1(n4_adj_5), .n42994(n42994), 
            .n6(n6), .n63957(n63957), .\state_7__N_4126[3] (\state_7__N_4126[3] ), 
            .n10(n10), .n25522(n25522), .n25517(n25517), .enable(enable), 
            .n10_adj_2(n10_adj_6)) /* synthesis syn_noprune=1, syn_module_defined=1 */ ;   // verilog/eeprom.v(83[16] 97[4])
    
endmodule
//
// Verilog Description of module i2c_controller
//

module i2c_controller (clk16MHz, scl_enable, \state[2] , \state[3] , 
            \state[0] , GND_net, \state_7__N_4110[0] , VCC_net, scl, 
            \state[1] , enable_slow_N_4213, sda_enable, sda_out, n29573, 
            \saved_addr[0] , n6426, n30410, data, n8, n30134, n30133, 
            n30132, n30131, n30130, n30129, n30128, n4, n4_adj_1, 
            n42994, n6, n63957, \state_7__N_4126[3] , n10, n25522, 
            n25517, enable, n10_adj_2) /* synthesis syn_noprune=1, syn_module_defined=1 */ ;
    input clk16MHz;
    output scl_enable;
    output \state[2] ;
    output \state[3] ;
    output \state[0] ;
    input GND_net;
    output \state_7__N_4110[0] ;
    input VCC_net;
    output scl;
    output \state[1] ;
    output enable_slow_N_4213;
    output sda_enable;
    output sda_out;
    input n29573;
    output \saved_addr[0] ;
    output n6426;
    input n30410;
    output [7:0]data;
    input n8;
    input n30134;
    input n30133;
    input n30132;
    input n30131;
    input n30130;
    input n30129;
    input n30128;
    output n4;
    output n4_adj_1;
    output n42994;
    output n6;
    output n63957;
    input \state_7__N_4126[3] ;
    output n10;
    output n25522;
    output n25517;
    input enable;
    output n10_adj_2;
    
    wire i2c_clk /* synthesis is_clock=1, SET_AS_NETWORK=\eeprom/i2c/i2c_clk */ ;   // verilog/i2c_controller.v(41[6:13])
    wire clk16MHz /* synthesis SET_AS_NETWORK=clk16MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    
    wire i2c_clk_N_4199, scl_enable_N_4200, n6754, enable_slow_N_4212, 
        n27694;
    wire [5:0]n29;
    wire [7:0]counter2;   // verilog/i2c_controller.v(37[12:20])
    
    wire n52395, n52394, n52393, n52392, n52391, sda_out_adj_4430;
    wire [7:0]n119;
    wire [7:0]counter;   // verilog/i2c_controller.v(36[12:19])
    
    wire n51268, n51267, n51266, n51265, n51264, n51263, n51262, 
        n29067, n61820, n59742, n4_c, n27887, n28826, n5, n61950, 
        n43152, n43440, n52718, n60756, n27558, n42860, n11, n27689, 
        n58048, n60892, n27687, n4_adj_4433, n11_adj_4434, n67181, 
        n9, n52714, n11_adj_4435, n10_adj_4436, n66964, n42883, 
        n11_adj_4437, n4_adj_4438, n6419, n11_adj_4439, n12, n28, 
        n70034, n59642, n28_adj_4441;
    
    SB_DFF i2c_clk_122 (.Q(i2c_clk), .C(clk16MHz), .D(i2c_clk_N_4199));   // verilog/i2c_controller.v(58[9] 71[5])
    SB_DFFN i2c_scl_enable_124 (.Q(scl_enable), .C(i2c_clk), .D(scl_enable_N_4200));   // verilog/i2c_controller.v(76[12] 82[6])
    SB_LUT4 i1_2_lut_3_lut (.I0(\state[2] ), .I1(\state[3] ), .I2(\state[0] ), 
            .I3(GND_net), .O(n6754));   // verilog/i2c_controller.v(44[32:47])
    defparam i1_2_lut_3_lut.LUT_INIT = 16'h1010;
    SB_DFFE enable_slow_121 (.Q(\state_7__N_4110[0] ), .C(clk16MHz), .E(n27694), 
            .D(enable_slow_N_4212));   // verilog/i2c_controller.v(58[9] 71[5])
    SB_LUT4 counter2_1950_1951_add_4_7_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter2[5]), .I3(n52395), .O(n29[5])) /* synthesis syn_instantiated=1 */ ;
    defparam counter2_1950_1951_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 counter2_1950_1951_add_4_6_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter2[4]), .I3(n52394), .O(n29[4])) /* synthesis syn_instantiated=1 */ ;
    defparam counter2_1950_1951_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter2_1950_1951_add_4_6 (.CI(n52394), .I0(GND_net), .I1(counter2[4]), 
            .CO(n52395));
    SB_LUT4 counter2_1950_1951_add_4_5_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter2[3]), .I3(n52393), .O(n29[3])) /* synthesis syn_instantiated=1 */ ;
    defparam counter2_1950_1951_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter2_1950_1951_add_4_5 (.CI(n52393), .I0(GND_net), .I1(counter2[3]), 
            .CO(n52394));
    SB_LUT4 counter2_1950_1951_add_4_4_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter2[2]), .I3(n52392), .O(n29[2])) /* synthesis syn_instantiated=1 */ ;
    defparam counter2_1950_1951_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter2_1950_1951_add_4_4 (.CI(n52392), .I0(GND_net), .I1(counter2[2]), 
            .CO(n52393));
    SB_LUT4 counter2_1950_1951_add_4_3_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter2[1]), .I3(n52391), .O(n29[1])) /* synthesis syn_instantiated=1 */ ;
    defparam counter2_1950_1951_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter2_1950_1951_add_4_3 (.CI(n52391), .I0(GND_net), .I1(counter2[1]), 
            .CO(n52392));
    SB_LUT4 counter2_1950_1951_add_4_2_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter2[0]), .I3(VCC_net), .O(n29[0])) /* synthesis syn_instantiated=1 */ ;
    defparam counter2_1950_1951_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter2_1950_1951_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(counter2[0]), 
            .CO(n52391));
    SB_LUT4 i29013_2_lut (.I0(i2c_clk), .I1(scl_enable), .I2(GND_net), 
            .I3(GND_net), .O(scl));   // verilog/i2c_controller.v(45[19:61])
    defparam i29013_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 i54392_3_lut_4_lut (.I0(\state[2] ), .I1(\state[3] ), .I2(\state[0] ), 
            .I3(\state[1] ), .O(enable_slow_N_4213));   // verilog/i2c_controller.v(44[32:47])
    defparam i54392_3_lut_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i2423_2_lut (.I0(sda_out_adj_4430), .I1(sda_enable), .I2(GND_net), 
            .I3(GND_net), .O(sda_out));   // verilog/i2c_controller.v(46[9:20])
    defparam i2423_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 sub_39_add_2_9_lut (.I0(GND_net), .I1(counter[7]), .I2(VCC_net), 
            .I3(n51268), .O(n119[7])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_39_add_2_8_lut (.I0(GND_net), .I1(counter[6]), .I2(VCC_net), 
            .I3(n51267), .O(n119[6])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_39_add_2_8 (.CI(n51267), .I0(counter[6]), .I1(VCC_net), 
            .CO(n51268));
    SB_LUT4 sub_39_add_2_7_lut (.I0(GND_net), .I1(counter[5]), .I2(VCC_net), 
            .I3(n51266), .O(n119[5])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_39_add_2_7 (.CI(n51266), .I0(counter[5]), .I1(VCC_net), 
            .CO(n51267));
    SB_LUT4 sub_39_add_2_6_lut (.I0(GND_net), .I1(counter[4]), .I2(VCC_net), 
            .I3(n51265), .O(n119[4])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_39_add_2_6 (.CI(n51265), .I0(counter[4]), .I1(VCC_net), 
            .CO(n51266));
    SB_LUT4 sub_39_add_2_5_lut (.I0(GND_net), .I1(counter[3]), .I2(VCC_net), 
            .I3(n51264), .O(n119[3])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_39_add_2_5 (.CI(n51264), .I0(counter[3]), .I1(VCC_net), 
            .CO(n51265));
    SB_LUT4 sub_39_add_2_4_lut (.I0(GND_net), .I1(counter[2]), .I2(VCC_net), 
            .I3(n51263), .O(n119[2])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_39_add_2_4 (.CI(n51263), .I0(counter[2]), .I1(VCC_net), 
            .CO(n51264));
    SB_LUT4 sub_39_add_2_3_lut (.I0(GND_net), .I1(counter[1]), .I2(VCC_net), 
            .I3(n51262), .O(n119[1])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_39_add_2_3 (.CI(n51262), .I0(counter[1]), .I1(VCC_net), 
            .CO(n51263));
    SB_LUT4 sub_39_add_2_2_lut (.I0(GND_net), .I1(counter[0]), .I2(GND_net), 
            .I3(VCC_net), .O(n119[0])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_39_add_2_2 (.CI(VCC_net), .I0(counter[0]), .I1(GND_net), 
            .CO(n51262));
    SB_DFF saved_addr__i1 (.Q(\saved_addr[0] ), .C(i2c_clk), .D(n29573));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFSR counter2_1950_1951__i6 (.Q(counter2[5]), .C(clk16MHz), .D(n29[5]), 
            .R(n29067));   // verilog/i2c_controller.v(69[20:35])
    SB_DFFSR counter2_1950_1951__i5 (.Q(counter2[4]), .C(clk16MHz), .D(n29[4]), 
            .R(n29067));   // verilog/i2c_controller.v(69[20:35])
    SB_DFFSR counter2_1950_1951__i4 (.Q(counter2[3]), .C(clk16MHz), .D(n29[3]), 
            .R(n29067));   // verilog/i2c_controller.v(69[20:35])
    SB_DFFSR counter2_1950_1951__i3 (.Q(counter2[2]), .C(clk16MHz), .D(n29[2]), 
            .R(n29067));   // verilog/i2c_controller.v(69[20:35])
    SB_DFFSR counter2_1950_1951__i2 (.Q(counter2[1]), .C(clk16MHz), .D(n29[1]), 
            .R(n29067));   // verilog/i2c_controller.v(69[20:35])
    SB_LUT4 i2_2_lut_4_lut (.I0(\state[1] ), .I1(\state[2] ), .I2(\state[0] ), 
            .I3(\state[3] ), .O(n61820));
    defparam i2_2_lut_4_lut.LUT_INIT = 16'h0054;
    SB_LUT4 i44102_2_lut_3_lut (.I0(\state[2] ), .I1(\state[0] ), .I2(\state[3] ), 
            .I3(GND_net), .O(n59742));
    defparam i44102_2_lut_3_lut.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_945 (.I0(\state[2] ), .I1(\state[0] ), .I2(\state[3] ), 
            .I3(GND_net), .O(n4_c));
    defparam i1_2_lut_3_lut_adj_945.LUT_INIT = 16'h0e0e;
    SB_DFFESS counter_i1 (.Q(counter[1]), .C(i2c_clk), .E(n27887), .D(n119[1]), 
            .S(n28826));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESS counter_i2 (.Q(counter[2]), .C(i2c_clk), .E(n27887), .D(n119[2]), 
            .S(n28826));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESR counter_i3 (.Q(counter[3]), .C(i2c_clk), .E(n27887), .D(n119[3]), 
            .R(n28826));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESR counter_i4 (.Q(counter[4]), .C(i2c_clk), .E(n27887), .D(n119[4]), 
            .R(n28826));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESR counter_i5 (.Q(counter[5]), .C(i2c_clk), .E(n27887), .D(n119[5]), 
            .R(n28826));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESR counter_i6 (.Q(counter[6]), .C(i2c_clk), .E(n27887), .D(n119[6]), 
            .R(n28826));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESR counter_i7 (.Q(counter[7]), .C(i2c_clk), .E(n27887), .D(n119[7]), 
            .R(n28826));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESS state_i0_i1 (.Q(\state[1] ), .C(i2c_clk), .E(n6426), .D(n5), 
            .S(n61950));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESS state_i0_i2 (.Q(\state[2] ), .C(i2c_clk), .E(n6426), .D(n43152), 
            .S(n43440));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESS state_i0_i3 (.Q(\state[3] ), .C(i2c_clk), .E(n6426), .D(n52718), 
            .S(n60756));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFSR counter2_1950_1951__i1 (.Q(counter2[0]), .C(clk16MHz), .D(n29[0]), 
            .R(n29067));   // verilog/i2c_controller.v(69[20:35])
    SB_DFF data_out_i0_i0 (.Q(data[0]), .C(i2c_clk), .D(n30410));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFE state_i0_i0 (.Q(\state[0] ), .C(i2c_clk), .E(VCC_net), .D(n8));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFF data_out_i0_i7 (.Q(data[7]), .C(i2c_clk), .D(n30134));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFF data_out_i0_i6 (.Q(data[6]), .C(i2c_clk), .D(n30133));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFF data_out_i0_i5 (.Q(data[5]), .C(i2c_clk), .D(n30132));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFF data_out_i0_i4 (.Q(data[4]), .C(i2c_clk), .D(n30131));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFF data_out_i0_i3 (.Q(data[3]), .C(i2c_clk), .D(n30130));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFF data_out_i0_i2 (.Q(data[2]), .C(i2c_clk), .D(n30129));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFF data_out_i0_i1 (.Q(data[1]), .C(i2c_clk), .D(n30128));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_LUT4 i54378_2_lut (.I0(\state_7__N_4110[0] ), .I1(enable_slow_N_4213), 
            .I2(GND_net), .I3(GND_net), .O(enable_slow_N_4212));   // verilog/i2c_controller.v(62[6:32])
    defparam i54378_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 i14820_2_lut_4_lut (.I0(n27887), .I1(\state[2] ), .I2(\state[3] ), 
            .I3(\state[0] ), .O(n28826));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i14820_2_lut_4_lut.LUT_INIT = 16'h0200;
    SB_LUT4 i1_3_lut_4_lut (.I0(\state[3] ), .I1(\state[2] ), .I2(\state[1] ), 
            .I3(\state[0] ), .O(n27558));
    defparam i1_3_lut_4_lut.LUT_INIT = 16'ha888;
    SB_LUT4 i29148_2_lut_3_lut (.I0(\state[2] ), .I1(\state[3] ), .I2(\state[0] ), 
            .I3(GND_net), .O(n42860));
    defparam i29148_2_lut_3_lut.LUT_INIT = 16'hfdfd;
    SB_LUT4 i54952_3_lut_4_lut (.I0(\state[2] ), .I1(\state[3] ), .I2(\state[1] ), 
            .I3(n6426), .O(n60756));
    defparam i54952_3_lut_4_lut.LUT_INIT = 16'h0200;
    SB_LUT4 equal_1515_i11_2_lut_4_lut (.I0(\state[1] ), .I1(\state[0] ), 
            .I2(\state[2] ), .I3(\state[3] ), .O(n11));   // verilog/i2c_controller.v(181[4] 217[11])
    defparam equal_1515_i11_2_lut_4_lut.LUT_INIT = 16'hff7f;
    SB_DFFNESS write_enable_132 (.Q(sda_enable), .C(i2c_clk), .E(n27689), 
            .D(n61820), .S(n58048));   // verilog/i2c_controller.v(180[12] 218[6])
    SB_DFFNESS sda_out_133 (.Q(sda_out_adj_4430), .C(i2c_clk), .E(n27687), 
            .D(n60892), .S(n58048));   // verilog/i2c_controller.v(180[12] 218[6])
    SB_DFFESS counter_i0 (.Q(counter[0]), .C(i2c_clk), .E(n27887), .D(n119[0]), 
            .S(n28826));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_LUT4 i1_2_lut (.I0(counter[2]), .I1(counter[1]), .I2(GND_net), 
            .I3(GND_net), .O(n4));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i1_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 equal_349_i4_2_lut (.I0(counter[1]), .I1(counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n4_adj_1));   // verilog/i2c_controller.v(153[6:23])
    defparam equal_349_i4_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 i29102_2_lut (.I0(counter[1]), .I1(counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n42994));
    defparam i29102_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_2_lut_4_lut_adj_946 (.I0(\state[2] ), .I1(\state[3] ), .I2(\state[0] ), 
            .I3(\state[1] ), .O(n6));
    defparam i2_2_lut_4_lut_adj_946.LUT_INIT = 16'hfebf;
    SB_LUT4 i48279_2_lut_3_lut (.I0(\state[2] ), .I1(\state[1] ), .I2(\state[0] ), 
            .I3(GND_net), .O(n63957));
    defparam i48279_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_4_lut_4_lut (.I0(\state[2] ), .I1(\state[1] ), .I2(\state[0] ), 
            .I3(\state[3] ), .O(n4_adj_4433));
    defparam i1_4_lut_4_lut.LUT_INIT = 16'hffa1;
    SB_LUT4 state_7__I_0_142_i11_2_lut_3_lut_4_lut (.I0(\state[0] ), .I1(\state[1] ), 
            .I2(\state[2] ), .I3(\state[3] ), .O(n11_adj_4434));   // verilog/i2c_controller.v(77[27:43])
    defparam state_7__I_0_142_i11_2_lut_3_lut_4_lut.LUT_INIT = 16'hfdff;
    SB_LUT4 i52079_2_lut_3_lut (.I0(\state[0] ), .I1(\state[1] ), .I2(\state_7__N_4126[3] ), 
            .I3(GND_net), .O(n67181));   // verilog/i2c_controller.v(77[27:43])
    defparam i52079_2_lut_3_lut.LUT_INIT = 16'hd0d0;
    SB_LUT4 i1_2_lut_3_lut_adj_947 (.I0(n9), .I1(n10), .I2(counter[0]), 
            .I3(GND_net), .O(n25522));   // verilog/i2c_controller.v(151[5:14])
    defparam i1_2_lut_3_lut_adj_947.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_2_lut_3_lut_adj_948 (.I0(n9), .I1(n10), .I2(counter[0]), 
            .I3(GND_net), .O(n25517));   // verilog/i2c_controller.v(151[5:14])
    defparam i1_2_lut_3_lut_adj_948.LUT_INIT = 16'hefef;
    SB_LUT4 i54962_3_lut_4_lut (.I0(n9), .I1(n10), .I2(n11_adj_4434), 
            .I3(n6426), .O(n43440));   // verilog/i2c_controller.v(151[5:14])
    defparam i54962_3_lut_4_lut.LUT_INIT = 16'h1f00;
    SB_LUT4 i54397_3_lut_4_lut (.I0(\state[3] ), .I1(\state[2] ), .I2(n52714), 
            .I3(n9), .O(n52718));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i54397_3_lut_4_lut.LUT_INIT = 16'h0f2f;
    SB_LUT4 state_7__I_0_145_i11_2_lut_3_lut_4_lut (.I0(\state[0] ), .I1(\state[1] ), 
            .I2(\state[2] ), .I3(\state[3] ), .O(n11_adj_4435));   // verilog/i2c_controller.v(77[27:43])
    defparam state_7__I_0_145_i11_2_lut_3_lut_4_lut.LUT_INIT = 16'hffdf;
    SB_LUT4 i2_4_lut (.I0(\state[1] ), .I1(\state[0] ), .I2(\state[2] ), 
            .I3(\state[3] ), .O(scl_enable_N_4200));
    defparam i2_4_lut.LUT_INIT = 16'hfefa;
    SB_LUT4 i4_4_lut (.I0(counter2[3]), .I1(counter2[5]), .I2(counter2[2]), 
            .I3(counter2[4]), .O(n10_adj_4436));
    defparam i4_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i5_3_lut (.I0(counter2[1]), .I1(n10_adj_4436), .I2(counter2[0]), 
            .I3(GND_net), .O(n29067));
    defparam i5_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i1_2_lut_adj_949 (.I0(i2c_clk), .I1(n29067), .I2(GND_net), 
            .I3(GND_net), .O(i2c_clk_N_4199));
    defparam i1_2_lut_adj_949.LUT_INIT = 16'h6666;
    SB_LUT4 i51673_2_lut (.I0(enable), .I1(n11), .I2(GND_net), .I3(GND_net), 
            .O(n66964));   // verilog/i2c_controller.v(33[12:17])
    defparam i51673_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i38_4_lut (.I0(n66964), .I1(n42883), .I2(\state_7__N_4126[3] ), 
            .I3(\state[3] ), .O(n52714));   // verilog/i2c_controller.v(33[12:17])
    defparam i38_4_lut.LUT_INIT = 16'hfa3a;
    SB_LUT4 i54866_2_lut (.I0(\state_7__N_4126[3] ), .I1(n11_adj_4437), 
            .I2(GND_net), .I3(GND_net), .O(n43152));
    defparam i54866_2_lut.LUT_INIT = 16'h1111;
    SB_LUT4 state_7__I_0_141_i10_2_lut (.I0(\state[2] ), .I1(\state[3] ), 
            .I2(GND_net), .I3(GND_net), .O(n10));   // verilog/i2c_controller.v(130[5:15])
    defparam state_7__I_0_141_i10_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 i1_2_lut_adj_950 (.I0(\state[0] ), .I1(\state[1] ), .I2(GND_net), 
            .I3(GND_net), .O(n9));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i1_2_lut_adj_950.LUT_INIT = 16'hbbbb;
    SB_LUT4 i28991_2_lut (.I0(\state[1] ), .I1(\state[0] ), .I2(GND_net), 
            .I3(GND_net), .O(n42883));
    defparam i28991_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_951 (.I0(n6426), .I1(\state[2] ), .I2(GND_net), 
            .I3(GND_net), .O(n4_adj_4438));
    defparam i1_2_lut_adj_951.LUT_INIT = 16'hdddd;
    SB_LUT4 i54964_4_lut (.I0(\state[3] ), .I1(n4_adj_4438), .I2(\state[0] ), 
            .I3(\state[1] ), .O(n61950));
    defparam i54964_4_lut.LUT_INIT = 16'h0130;
    SB_LUT4 i54364_4_lut (.I0(n27558), .I1(n6419), .I2(n11_adj_4439), 
            .I3(n42860), .O(n6426));
    defparam i54364_4_lut.LUT_INIT = 16'h5111;
    SB_LUT4 i1_4_lut (.I0(\state_7__N_4126[3] ), .I1(n11_adj_4435), .I2(\saved_addr[0] ), 
            .I3(n11_adj_4437), .O(n5));   // verilog/i2c_controller.v(33[12:17])
    defparam i1_4_lut.LUT_INIT = 16'h3373;
    SB_LUT4 i1_2_lut_3_lut_adj_952 (.I0(enable), .I1(\state_7__N_4110[0] ), 
            .I2(enable_slow_N_4213), .I3(GND_net), .O(n27694));
    defparam i1_2_lut_3_lut_adj_952.LUT_INIT = 16'haeae;
    SB_LUT4 i2_2_lut (.I0(counter[2]), .I1(counter[1]), .I2(GND_net), 
            .I3(GND_net), .O(n10_adj_2));   // verilog/i2c_controller.v(110[10:22])
    defparam i2_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i5_4_lut (.I0(counter[3]), .I1(counter[4]), .I2(counter[0]), 
            .I3(counter[6]), .O(n12));   // verilog/i2c_controller.v(110[10:22])
    defparam i5_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i6_4_lut (.I0(counter[5]), .I1(n12), .I2(counter[7]), .I3(n10_adj_2), 
            .O(n6419));   // verilog/i2c_controller.v(110[10:22])
    defparam i6_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i14_4_lut (.I0(n6419), .I1(n67181), .I2(n6754), .I3(n4_adj_4433), 
            .O(n27887));
    defparam i14_4_lut.LUT_INIT = 16'h303a;
    SB_LUT4 state_7__I_0_139_i11_2_lut_3_lut_4_lut (.I0(\state[2] ), .I1(\state[3] ), 
            .I2(\state[0] ), .I3(\state[1] ), .O(n11_adj_4439));   // verilog/i2c_controller.v(44[32:47])
    defparam state_7__I_0_139_i11_2_lut_3_lut_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i1_4_lut_adj_953 (.I0(\state[3] ), .I1(\state[2] ), .I2(\state[0] ), 
            .I3(\state[1] ), .O(n28));
    defparam i1_4_lut_adj_953.LUT_INIT = 16'h4054;
    SB_LUT4 i54340_2_lut (.I0(\state[3] ), .I1(\state[1] ), .I2(GND_net), 
            .I3(GND_net), .O(n70034));
    defparam i54340_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 state_7__I_0_140_i11_2_lut_3_lut_4_lut (.I0(\state[2] ), .I1(\state[3] ), 
            .I2(\state[1] ), .I3(\state[0] ), .O(n11_adj_4437));   // verilog/i2c_controller.v(44[32:47])
    defparam state_7__I_0_140_i11_2_lut_3_lut_4_lut.LUT_INIT = 16'hefff;
    SB_LUT4 i1_4_lut_adj_954 (.I0(n11), .I1(n70034), .I2(n28), .I3(n59642), 
            .O(n27687));
    defparam i1_4_lut_adj_954.LUT_INIT = 16'ha0a8;
    SB_LUT4 i35_4_lut (.I0(counter[1]), .I1(counter[0]), .I2(counter[2]), 
            .I3(\saved_addr[0] ), .O(n28_adj_4441));   // verilog/i2c_controller.v(36[12:19])
    defparam i35_4_lut.LUT_INIT = 16'hc1c0;
    SB_LUT4 i44004_2_lut (.I0(\state[2] ), .I1(\state[0] ), .I2(GND_net), 
            .I3(GND_net), .O(n59642));
    defparam i44004_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i3_4_lut (.I0(\state[3] ), .I1(n11), .I2(\state[1] ), .I3(n59642), 
            .O(n58048));
    defparam i3_4_lut.LUT_INIT = 16'h0008;
    SB_LUT4 i1_4_lut_adj_955 (.I0(n11), .I1(\state[1] ), .I2(n4_c), .I3(n59742), 
            .O(n27689));
    defparam i1_4_lut_adj_955.LUT_INIT = 16'ha0a2;
    SB_LUT4 i2_3_lut_4_lut (.I0(\state[2] ), .I1(\state[3] ), .I2(\state[1] ), 
            .I3(n28_adj_4441), .O(n60892));   // verilog/i2c_controller.v(44[32:47])
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h1000;
    
endmodule
