// ******************************************************************************

// iCEcube Netlister

// Version:            2017.08.27940

// Build Date:         Sep 12 2017 08:25:46

// File Generated:     Jan 29 2020 19:23:48

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "TinyFPGA_B" view "INTERFACE"

module TinyFPGA_B (
    USBPU,
    TX,
    SDA,
    SCL,
    RX,
    NEOPXL,
    LED,
    INLC,
    INLB,
    INLA,
    INHC,
    INHB,
    INHA,
    HALL3,
    HALL2,
    HALL1,
    FAULT_N,
    ENCODER1_B,
    ENCODER1_A,
    ENCODER0_B,
    ENCODER0_A,
    DE,
    CS_MISO,
    CS_CLK,
    CS,
    CLK);

    output USBPU;
    output TX;
    inout SDA;
    inout SCL;
    input RX;
    output NEOPXL;
    output LED;
    output INLC;
    output INLB;
    output INLA;
    output INHC;
    output INHB;
    output INHA;
    input HALL3;
    input HALL2;
    input HALL1;
    input FAULT_N;
    input ENCODER1_B;
    input ENCODER1_A;
    input ENCODER0_B;
    input ENCODER0_A;
    output DE;
    input CS_MISO;
    output CS_CLK;
    output CS;
    input CLK;

    wire N__5901;
    wire N__5900;
    wire N__5899;
    wire N__5892;
    wire N__5891;
    wire N__5890;
    wire N__5883;
    wire N__5882;
    wire N__5881;
    wire N__5874;
    wire N__5873;
    wire N__5872;
    wire N__5865;
    wire N__5864;
    wire N__5863;
    wire N__5856;
    wire N__5855;
    wire N__5854;
    wire N__5847;
    wire N__5846;
    wire N__5845;
    wire N__5838;
    wire N__5837;
    wire N__5836;
    wire N__5829;
    wire N__5828;
    wire N__5827;
    wire N__5820;
    wire N__5819;
    wire N__5818;
    wire N__5811;
    wire N__5810;
    wire N__5809;
    wire N__5802;
    wire N__5801;
    wire N__5800;
    wire N__5793;
    wire N__5792;
    wire N__5791;
    wire N__5784;
    wire N__5783;
    wire N__5782;
    wire N__5775;
    wire N__5774;
    wire N__5773;
    wire N__5766;
    wire N__5765;
    wire N__5764;
    wire N__5747;
    wire N__5746;
    wire N__5743;
    wire N__5740;
    wire N__5737;
    wire N__5732;
    wire N__5731;
    wire N__5728;
    wire N__5725;
    wire N__5720;
    wire N__5717;
    wire N__5714;
    wire N__5713;
    wire N__5710;
    wire N__5707;
    wire N__5706;
    wire N__5705;
    wire N__5702;
    wire N__5699;
    wire N__5696;
    wire N__5693;
    wire N__5684;
    wire N__5683;
    wire N__5682;
    wire N__5679;
    wire N__5676;
    wire N__5673;
    wire N__5670;
    wire N__5667;
    wire N__5664;
    wire N__5657;
    wire N__5654;
    wire N__5651;
    wire N__5650;
    wire N__5649;
    wire N__5646;
    wire N__5643;
    wire N__5640;
    wire N__5633;
    wire N__5632;
    wire N__5631;
    wire N__5630;
    wire N__5627;
    wire N__5626;
    wire N__5625;
    wire N__5622;
    wire N__5619;
    wire N__5616;
    wire N__5613;
    wire N__5608;
    wire N__5597;
    wire N__5594;
    wire N__5591;
    wire N__5588;
    wire N__5585;
    wire N__5582;
    wire N__5579;
    wire N__5578;
    wire N__5575;
    wire N__5574;
    wire N__5573;
    wire N__5570;
    wire N__5569;
    wire N__5568;
    wire N__5567;
    wire N__5566;
    wire N__5565;
    wire N__5564;
    wire N__5563;
    wire N__5562;
    wire N__5559;
    wire N__5556;
    wire N__5553;
    wire N__5550;
    wire N__5547;
    wire N__5546;
    wire N__5539;
    wire N__5536;
    wire N__5535;
    wire N__5532;
    wire N__5531;
    wire N__5530;
    wire N__5527;
    wire N__5526;
    wire N__5525;
    wire N__5524;
    wire N__5521;
    wire N__5514;
    wire N__5509;
    wire N__5506;
    wire N__5501;
    wire N__5500;
    wire N__5499;
    wire N__5498;
    wire N__5497;
    wire N__5496;
    wire N__5493;
    wire N__5490;
    wire N__5483;
    wire N__5476;
    wire N__5473;
    wire N__5466;
    wire N__5463;
    wire N__5456;
    wire N__5451;
    wire N__5448;
    wire N__5429;
    wire N__5428;
    wire N__5425;
    wire N__5424;
    wire N__5423;
    wire N__5422;
    wire N__5421;
    wire N__5420;
    wire N__5419;
    wire N__5416;
    wire N__5415;
    wire N__5414;
    wire N__5411;
    wire N__5408;
    wire N__5405;
    wire N__5402;
    wire N__5401;
    wire N__5400;
    wire N__5399;
    wire N__5398;
    wire N__5397;
    wire N__5396;
    wire N__5395;
    wire N__5392;
    wire N__5389;
    wire N__5384;
    wire N__5381;
    wire N__5378;
    wire N__5373;
    wire N__5368;
    wire N__5367;
    wire N__5366;
    wire N__5365;
    wire N__5364;
    wire N__5361;
    wire N__5360;
    wire N__5357;
    wire N__5356;
    wire N__5353;
    wire N__5350;
    wire N__5347;
    wire N__5342;
    wire N__5335;
    wire N__5328;
    wire N__5325;
    wire N__5316;
    wire N__5313;
    wire N__5310;
    wire N__5305;
    wire N__5282;
    wire N__5281;
    wire N__5280;
    wire N__5279;
    wire N__5278;
    wire N__5277;
    wire N__5274;
    wire N__5271;
    wire N__5270;
    wire N__5267;
    wire N__5266;
    wire N__5263;
    wire N__5262;
    wire N__5261;
    wire N__5260;
    wire N__5259;
    wire N__5258;
    wire N__5257;
    wire N__5254;
    wire N__5249;
    wire N__5246;
    wire N__5241;
    wire N__5238;
    wire N__5237;
    wire N__5236;
    wire N__5233;
    wire N__5230;
    wire N__5227;
    wire N__5222;
    wire N__5217;
    wire N__5214;
    wire N__5211;
    wire N__5204;
    wire N__5201;
    wire N__5200;
    wire N__5199;
    wire N__5196;
    wire N__5195;
    wire N__5194;
    wire N__5193;
    wire N__5192;
    wire N__5189;
    wire N__5186;
    wire N__5179;
    wire N__5172;
    wire N__5169;
    wire N__5162;
    wire N__5159;
    wire N__5152;
    wire N__5135;
    wire N__5134;
    wire N__5133;
    wire N__5132;
    wire N__5131;
    wire N__5130;
    wire N__5129;
    wire N__5128;
    wire N__5127;
    wire N__5126;
    wire N__5125;
    wire N__5124;
    wire N__5123;
    wire N__5120;
    wire N__5119;
    wire N__5114;
    wire N__5111;
    wire N__5108;
    wire N__5101;
    wire N__5098;
    wire N__5097;
    wire N__5094;
    wire N__5087;
    wire N__5086;
    wire N__5083;
    wire N__5080;
    wire N__5071;
    wire N__5070;
    wire N__5069;
    wire N__5068;
    wire N__5067;
    wire N__5066;
    wire N__5065;
    wire N__5064;
    wire N__5061;
    wire N__5058;
    wire N__5055;
    wire N__5052;
    wire N__5049;
    wire N__5042;
    wire N__5035;
    wire N__5026;
    wire N__5009;
    wire N__5006;
    wire N__5003;
    wire N__5000;
    wire N__4997;
    wire N__4994;
    wire N__4991;
    wire N__4990;
    wire N__4987;
    wire N__4984;
    wire N__4979;
    wire N__4976;
    wire N__4975;
    wire N__4974;
    wire N__4973;
    wire N__4972;
    wire N__4969;
    wire N__4966;
    wire N__4963;
    wire N__4960;
    wire N__4957;
    wire N__4956;
    wire N__4955;
    wire N__4954;
    wire N__4953;
    wire N__4950;
    wire N__4947;
    wire N__4946;
    wire N__4941;
    wire N__4938;
    wire N__4935;
    wire N__4932;
    wire N__4929;
    wire N__4926;
    wire N__4921;
    wire N__4918;
    wire N__4915;
    wire N__4912;
    wire N__4907;
    wire N__4904;
    wire N__4897;
    wire N__4896;
    wire N__4895;
    wire N__4894;
    wire N__4891;
    wire N__4886;
    wire N__4883;
    wire N__4880;
    wire N__4877;
    wire N__4872;
    wire N__4859;
    wire N__4856;
    wire N__4853;
    wire N__4850;
    wire N__4847;
    wire N__4844;
    wire N__4841;
    wire N__4840;
    wire N__4837;
    wire N__4834;
    wire N__4829;
    wire N__4826;
    wire N__4825;
    wire N__4822;
    wire N__4821;
    wire N__4820;
    wire N__4817;
    wire N__4814;
    wire N__4809;
    wire N__4802;
    wire N__4799;
    wire N__4796;
    wire N__4795;
    wire N__4792;
    wire N__4791;
    wire N__4790;
    wire N__4789;
    wire N__4786;
    wire N__4783;
    wire N__4776;
    wire N__4769;
    wire N__4766;
    wire N__4763;
    wire N__4760;
    wire N__4757;
    wire N__4754;
    wire N__4751;
    wire N__4748;
    wire N__4747;
    wire N__4746;
    wire N__4739;
    wire N__4736;
    wire N__4733;
    wire N__4730;
    wire N__4727;
    wire N__4724;
    wire N__4721;
    wire N__4718;
    wire N__4715;
    wire N__4714;
    wire N__4713;
    wire N__4710;
    wire N__4707;
    wire N__4704;
    wire N__4697;
    wire N__4694;
    wire N__4691;
    wire N__4688;
    wire N__4687;
    wire N__4684;
    wire N__4681;
    wire N__4678;
    wire N__4675;
    wire N__4670;
    wire N__4669;
    wire N__4666;
    wire N__4663;
    wire N__4660;
    wire N__4657;
    wire N__4652;
    wire N__4649;
    wire N__4648;
    wire N__4645;
    wire N__4642;
    wire N__4639;
    wire N__4634;
    wire N__4633;
    wire N__4630;
    wire N__4627;
    wire N__4624;
    wire N__4619;
    wire N__4618;
    wire N__4615;
    wire N__4612;
    wire N__4609;
    wire N__4604;
    wire N__4601;
    wire N__4600;
    wire N__4597;
    wire N__4596;
    wire N__4593;
    wire N__4590;
    wire N__4587;
    wire N__4584;
    wire N__4577;
    wire N__4574;
    wire N__4571;
    wire N__4568;
    wire N__4565;
    wire N__4562;
    wire N__4559;
    wire N__4556;
    wire N__4553;
    wire N__4550;
    wire N__4547;
    wire N__4544;
    wire N__4541;
    wire N__4538;
    wire N__4535;
    wire N__4532;
    wire N__4531;
    wire N__4530;
    wire N__4527;
    wire N__4522;
    wire N__4517;
    wire N__4516;
    wire N__4511;
    wire N__4508;
    wire N__4505;
    wire N__4502;
    wire N__4499;
    wire N__4496;
    wire N__4493;
    wire N__4490;
    wire N__4487;
    wire N__4486;
    wire N__4483;
    wire N__4480;
    wire N__4479;
    wire N__4476;
    wire N__4473;
    wire N__4470;
    wire N__4463;
    wire N__4460;
    wire N__4457;
    wire N__4454;
    wire N__4451;
    wire N__4448;
    wire N__4445;
    wire N__4444;
    wire N__4443;
    wire N__4440;
    wire N__4437;
    wire N__4434;
    wire N__4427;
    wire N__4424;
    wire N__4421;
    wire N__4418;
    wire N__4415;
    wire N__4414;
    wire N__4413;
    wire N__4412;
    wire N__4411;
    wire N__4408;
    wire N__4407;
    wire N__4404;
    wire N__4403;
    wire N__4400;
    wire N__4385;
    wire N__4382;
    wire N__4379;
    wire N__4376;
    wire N__4373;
    wire N__4370;
    wire N__4367;
    wire N__4364;
    wire N__4361;
    wire N__4358;
    wire N__4355;
    wire N__4352;
    wire N__4351;
    wire N__4348;
    wire N__4345;
    wire N__4342;
    wire N__4341;
    wire N__4338;
    wire N__4335;
    wire N__4332;
    wire N__4329;
    wire N__4324;
    wire N__4319;
    wire N__4316;
    wire N__4313;
    wire N__4310;
    wire N__4307;
    wire N__4304;
    wire N__4301;
    wire N__4298;
    wire N__4295;
    wire N__4292;
    wire N__4289;
    wire N__4286;
    wire N__4283;
    wire N__4280;
    wire N__4277;
    wire N__4274;
    wire N__4271;
    wire N__4268;
    wire N__4265;
    wire N__4262;
    wire N__4259;
    wire N__4256;
    wire N__4253;
    wire N__4250;
    wire N__4247;
    wire N__4244;
    wire N__4241;
    wire N__4238;
    wire N__4235;
    wire N__4232;
    wire N__4231;
    wire N__4228;
    wire N__4225;
    wire N__4220;
    wire N__4219;
    wire N__4218;
    wire N__4217;
    wire N__4216;
    wire N__4211;
    wire N__4208;
    wire N__4205;
    wire N__4202;
    wire N__4197;
    wire N__4194;
    wire N__4191;
    wire N__4188;
    wire N__4185;
    wire N__4184;
    wire N__4181;
    wire N__4176;
    wire N__4173;
    wire N__4166;
    wire N__4165;
    wire N__4160;
    wire N__4157;
    wire N__4156;
    wire N__4153;
    wire N__4150;
    wire N__4145;
    wire N__4142;
    wire N__4141;
    wire N__4138;
    wire N__4135;
    wire N__4130;
    wire N__4127;
    wire N__4126;
    wire N__4123;
    wire N__4120;
    wire N__4115;
    wire N__4112;
    wire N__4111;
    wire N__4108;
    wire N__4105;
    wire N__4100;
    wire N__4097;
    wire N__4094;
    wire N__4093;
    wire N__4090;
    wire N__4087;
    wire N__4082;
    wire N__4079;
    wire N__4076;
    wire N__4075;
    wire N__4074;
    wire N__4071;
    wire N__4068;
    wire N__4065;
    wire N__4058;
    wire N__4057;
    wire N__4056;
    wire N__4053;
    wire N__4052;
    wire N__4051;
    wire N__4046;
    wire N__4043;
    wire N__4040;
    wire N__4037;
    wire N__4034;
    wire N__4029;
    wire N__4026;
    wire N__4021;
    wire N__4018;
    wire N__4015;
    wire N__4010;
    wire N__4007;
    wire N__4006;
    wire N__4005;
    wire N__4004;
    wire N__4003;
    wire N__4002;
    wire N__4001;
    wire N__4000;
    wire N__3999;
    wire N__3998;
    wire N__3995;
    wire N__3992;
    wire N__3987;
    wire N__3978;
    wire N__3973;
    wire N__3962;
    wire N__3961;
    wire N__3960;
    wire N__3957;
    wire N__3954;
    wire N__3951;
    wire N__3948;
    wire N__3941;
    wire N__3940;
    wire N__3939;
    wire N__3938;
    wire N__3937;
    wire N__3936;
    wire N__3935;
    wire N__3934;
    wire N__3933;
    wire N__3932;
    wire N__3931;
    wire N__3930;
    wire N__3929;
    wire N__3928;
    wire N__3927;
    wire N__3926;
    wire N__3925;
    wire N__3890;
    wire N__3887;
    wire N__3884;
    wire N__3881;
    wire N__3878;
    wire N__3877;
    wire N__3876;
    wire N__3875;
    wire N__3874;
    wire N__3873;
    wire N__3870;
    wire N__3865;
    wire N__3860;
    wire N__3857;
    wire N__3848;
    wire N__3845;
    wire N__3842;
    wire N__3841;
    wire N__3838;
    wire N__3835;
    wire N__3830;
    wire N__3829;
    wire N__3826;
    wire N__3823;
    wire N__3818;
    wire N__3817;
    wire N__3814;
    wire N__3811;
    wire N__3808;
    wire N__3803;
    wire N__3802;
    wire N__3799;
    wire N__3796;
    wire N__3791;
    wire N__3790;
    wire N__3787;
    wire N__3784;
    wire N__3779;
    wire N__3778;
    wire N__3775;
    wire N__3772;
    wire N__3767;
    wire N__3764;
    wire N__3763;
    wire N__3760;
    wire N__3757;
    wire N__3752;
    wire N__3749;
    wire N__3746;
    wire N__3745;
    wire N__3742;
    wire N__3739;
    wire N__3734;
    wire N__3731;
    wire N__3730;
    wire N__3727;
    wire N__3724;
    wire N__3719;
    wire N__3716;
    wire N__3715;
    wire N__3712;
    wire N__3709;
    wire N__3704;
    wire N__3701;
    wire N__3698;
    wire N__3695;
    wire N__3692;
    wire N__3689;
    wire N__3686;
    wire N__3683;
    wire N__3680;
    wire N__3679;
    wire N__3678;
    wire N__3675;
    wire N__3670;
    wire N__3665;
    wire N__3662;
    wire N__3661;
    wire N__3658;
    wire N__3655;
    wire N__3650;
    wire N__3649;
    wire N__3646;
    wire N__3643;
    wire N__3640;
    wire N__3637;
    wire N__3632;
    wire N__3631;
    wire N__3628;
    wire N__3625;
    wire N__3620;
    wire N__3617;
    wire N__3616;
    wire N__3613;
    wire N__3610;
    wire N__3605;
    wire N__3602;
    wire N__3599;
    wire N__3598;
    wire N__3597;
    wire N__3596;
    wire N__3595;
    wire N__3594;
    wire N__3593;
    wire N__3592;
    wire N__3591;
    wire N__3590;
    wire N__3587;
    wire N__3586;
    wire N__3583;
    wire N__3582;
    wire N__3579;
    wire N__3578;
    wire N__3575;
    wire N__3572;
    wire N__3569;
    wire N__3568;
    wire N__3565;
    wire N__3564;
    wire N__3561;
    wire N__3560;
    wire N__3543;
    wire N__3540;
    wire N__3525;
    wire N__3518;
    wire N__3517;
    wire N__3514;
    wire N__3511;
    wire N__3506;
    wire N__3503;
    wire N__3502;
    wire N__3499;
    wire N__3496;
    wire N__3493;
    wire N__3488;
    wire N__3487;
    wire N__3484;
    wire N__3481;
    wire N__3476;
    wire N__3473;
    wire N__3472;
    wire N__3469;
    wire N__3466;
    wire N__3461;
    wire N__3458;
    wire N__3455;
    wire N__3452;
    wire N__3449;
    wire N__3446;
    wire N__3443;
    wire N__3440;
    wire N__3437;
    wire N__3434;
    wire N__3431;
    wire N__3428;
    wire N__3425;
    wire N__3422;
    wire N__3419;
    wire N__3416;
    wire N__3413;
    wire N__3410;
    wire N__3407;
    wire N__3404;
    wire N__3401;
    wire N__3400;
    wire N__3397;
    wire N__3394;
    wire N__3389;
    wire N__3386;
    wire N__3385;
    wire N__3382;
    wire N__3379;
    wire N__3374;
    wire N__3371;
    wire N__3370;
    wire N__3367;
    wire N__3364;
    wire N__3359;
    wire N__3358;
    wire N__3355;
    wire N__3352;
    wire N__3347;
    wire N__3346;
    wire N__3343;
    wire N__3340;
    wire N__3335;
    wire N__3332;
    wire N__3331;
    wire N__3328;
    wire N__3325;
    wire N__3322;
    wire N__3317;
    wire N__3316;
    wire N__3313;
    wire N__3310;
    wire N__3305;
    wire N__3304;
    wire N__3301;
    wire N__3298;
    wire N__3293;
    wire N__3290;
    wire N__3289;
    wire N__3286;
    wire N__3283;
    wire N__3278;
    wire N__3275;
    wire N__3272;
    wire N__3269;
    wire N__3268;
    wire N__3267;
    wire N__3266;
    wire N__3263;
    wire N__3260;
    wire N__3257;
    wire N__3254;
    wire N__3245;
    wire N__3244;
    wire N__3243;
    wire N__3240;
    wire N__3237;
    wire N__3234;
    wire N__3227;
    wire N__3224;
    wire N__3221;
    wire N__3220;
    wire N__3217;
    wire N__3214;
    wire N__3209;
    wire N__3208;
    wire N__3205;
    wire N__3202;
    wire N__3197;
    wire N__3196;
    wire N__3193;
    wire N__3190;
    wire N__3187;
    wire N__3182;
    wire N__3181;
    wire N__3178;
    wire N__3175;
    wire N__3170;
    wire N__3169;
    wire N__3164;
    wire N__3161;
    wire N__3158;
    wire N__3155;
    wire N__3154;
    wire N__3151;
    wire N__3148;
    wire N__3143;
    wire N__3142;
    wire N__3139;
    wire N__3136;
    wire N__3131;
    wire N__3130;
    wire N__3127;
    wire N__3124;
    wire N__3121;
    wire N__3116;
    wire N__3115;
    wire N__3112;
    wire N__3109;
    wire N__3104;
    wire N__3103;
    wire N__3100;
    wire N__3097;
    wire N__3092;
    wire N__3091;
    wire N__3088;
    wire N__3085;
    wire N__3080;
    wire N__3079;
    wire N__3076;
    wire N__3073;
    wire N__3070;
    wire N__3065;
    wire N__3064;
    wire N__3061;
    wire N__3058;
    wire N__3053;
    wire N__3052;
    wire N__3049;
    wire N__3046;
    wire N__3041;
    wire N__3040;
    wire N__3037;
    wire N__3034;
    wire N__3029;
    wire N__3026;
    wire N__3023;
    wire N__3020;
    wire N__3017;
    wire N__3014;
    wire N__3011;
    wire N__3010;
    wire N__3007;
    wire N__3004;
    wire N__2999;
    wire N__2998;
    wire N__2995;
    wire N__2992;
    wire N__2987;
    wire N__2984;
    wire N__2983;
    wire N__2980;
    wire N__2977;
    wire N__2972;
    wire N__2971;
    wire N__2968;
    wire N__2965;
    wire N__2962;
    wire N__2957;
    wire N__2956;
    wire N__2953;
    wire N__2950;
    wire N__2945;
    wire N__2944;
    wire N__2941;
    wire N__2938;
    wire N__2933;
    wire N__2930;
    wire N__2927;
    wire N__2926;
    wire N__2923;
    wire N__2920;
    wire N__2915;
    wire N__2914;
    wire N__2911;
    wire N__2908;
    wire N__2905;
    wire N__2900;
    wire N__2897;
    wire N__2894;
    wire N__2891;
    wire N__2888;
    wire N__2885;
    wire N__2882;
    wire N__2879;
    wire N__2876;
    wire N__2873;
    wire N__2870;
    wire N__2867;
    wire N__2864;
    wire N__2861;
    wire N__2858;
    wire N__2855;
    wire N__2852;
    wire N__2849;
    wire N__2846;
    wire N__2843;
    wire N__2840;
    wire N__2837;
    wire N__2834;
    wire N__2831;
    wire N__2828;
    wire N__2825;
    wire N__2822;
    wire N__2819;
    wire N__2816;
    wire N__2813;
    wire N__2810;
    wire N__2807;
    wire N__2804;
    wire N__2803;
    wire N__2802;
    wire N__2797;
    wire N__2794;
    wire N__2789;
    wire N__2788;
    wire N__2787;
    wire N__2780;
    wire N__2777;
    wire N__2776;
    wire N__2773;
    wire N__2770;
    wire N__2769;
    wire N__2764;
    wire N__2761;
    wire N__2756;
    wire N__2755;
    wire N__2754;
    wire N__2749;
    wire N__2746;
    wire N__2741;
    wire N__2738;
    wire N__2735;
    wire N__2732;
    wire N__2731;
    wire N__2726;
    wire N__2723;
    wire N__2720;
    wire N__2717;
    wire N__2714;
    wire N__2711;
    wire N__2708;
    wire N__2705;
    wire N__2702;
    wire N__2699;
    wire N__2696;
    wire N__2693;
    wire N__2690;
    wire N__2687;
    wire N__2684;
    wire N__2681;
    wire N__2678;
    wire N__2675;
    wire N__2672;
    wire N__2669;
    wire N__2666;
    wire N__2663;
    wire N__2660;
    wire N__2657;
    wire N__2654;
    wire N__2651;
    wire N__2648;
    wire N__2645;
    wire N__2642;
    wire N__2639;
    wire N__2636;
    wire N__2633;
    wire N__2630;
    wire N__2627;
    wire N__2624;
    wire N__2621;
    wire N__2618;
    wire N__2615;
    wire N__2612;
    wire N__2609;
    wire N__2606;
    wire N__2603;
    wire N__2600;
    wire N__2597;
    wire N__2594;
    wire N__2591;
    wire N__2588;
    wire N__2585;
    wire N__2582;
    wire N__2579;
    wire N__2576;
    wire N__2573;
    wire N__2570;
    wire N__2567;
    wire N__2564;
    wire N__2561;
    wire N__2558;
    wire N__2555;
    wire N__2552;
    wire N__2549;
    wire N__2546;
    wire N__2543;
    wire N__2540;
    wire N__2537;
    wire N__2534;
    wire N__2531;
    wire N__2528;
    wire N__2525;
    wire N__2522;
    wire N__2519;
    wire N__2516;
    wire N__2513;
    wire N__2510;
    wire N__2507;
    wire N__2504;
    wire N__2501;
    wire N__2498;
    wire N__2495;
    wire N__2492;
    wire N__2489;
    wire N__2486;
    wire N__2483;
    wire CLK_pad_gb_input;
    wire VCCG0;
    wire GNDG0;
    wire n26;
    wire bfn_13_21_0_;
    wire n25;
    wire n2535;
    wire n24;
    wire n2536;
    wire n23;
    wire n2537;
    wire n22;
    wire n2538;
    wire n21;
    wire n2539;
    wire n20;
    wire n2540;
    wire n19;
    wire n2541;
    wire n2542;
    wire n18;
    wire bfn_13_22_0_;
    wire n17_adj_394;
    wire n2543;
    wire n16_adj_393;
    wire n2544;
    wire n15_adj_392;
    wire n2545;
    wire n14_adj_391;
    wire n2546;
    wire n13_adj_390;
    wire n2547;
    wire n12_adj_389;
    wire n2548;
    wire n11;
    wire n2549;
    wire n2550;
    wire n10;
    wire bfn_13_23_0_;
    wire n9;
    wire n2551;
    wire n8_adj_388;
    wire n2552;
    wire n7_adj_387;
    wire n2553;
    wire n6;
    wire n2554;
    wire n2555;
    wire n2556;
    wire n2557;
    wire n2558;
    wire bfn_13_24_0_;
    wire n2559;
    wire blink_counter_21;
    wire blink_counter_24;
    wire blink_counter_23;
    wire blink_counter_22;
    wire n2730;
    wire n2731_cascade_;
    wire blink_counter_25;
    wire LED_c;
    wire bfn_14_21_0_;
    wire n2478;
    wire n2479;
    wire n2480;
    wire n2481;
    wire n2482;
    wire n2483;
    wire n2484;
    wire n2485;
    wire bfn_14_22_0_;
    wire n2486;
    wire n2487;
    wire n2488;
    wire n2489;
    wire n2490;
    wire n2491;
    wire n2492;
    wire n2493;
    wire bfn_14_23_0_;
    wire n2494;
    wire n2495;
    wire n2496;
    wire n2497;
    wire n2498;
    wire n2499;
    wire n2500;
    wire n2501;
    wire bfn_14_24_0_;
    wire n2502;
    wire n2503;
    wire n2504;
    wire n2505;
    wire n2506;
    wire n2507;
    wire n2508;
    wire delay_counter_6;
    wire delay_counter_0;
    wire delay_counter_9;
    wire delay_counter_4;
    wire delay_counter_2;
    wire delay_counter_7;
    wire delay_counter_5;
    wire delay_counter_3;
    wire delay_counter_8;
    wire delay_counter_1;
    wire n17;
    wire n16;
    wire delay_counter_11;
    wire delay_counter_10;
    wire n2722_cascade_;
    wire delay_counter_12;
    wire delay_counter_17;
    wire delay_counter_15;
    wire delay_counter_14;
    wire n8;
    wire delay_counter_16;
    wire delay_counter_13;
    wire n2715;
    wire delay_counter_18;
    wire delay_counter_19;
    wire n2721_cascade_;
    wire delay_counter_22;
    wire delay_counter_21;
    wire delay_counter_23;
    wire n7_cascade_;
    wire delay_counter_20;
    wire delay_counter_29;
    wire delay_counter_25;
    wire n2695_cascade_;
    wire delay_counter_28;
    wire n13_cascade_;
    wire addr_10__N_70;
    wire delay_counter_31;
    wire n13;
    wire delay_counter_26;
    wire delay_counter_30;
    wire delay_counter_27;
    wire delay_counter_24;
    wire n14;
    wire n2077_cascade_;
    wire n2077;
    wire n12_cascade_;
    wire bfn_17_19_0_;
    wire \eeprom.n2516 ;
    wire \eeprom.n2517 ;
    wire \eeprom.n2518 ;
    wire \eeprom.n2519 ;
    wire \eeprom.n2520 ;
    wire \eeprom.n2521 ;
    wire \eeprom.n2522 ;
    wire \eeprom.n2523 ;
    wire bfn_17_20_0_;
    wire \eeprom.n2524 ;
    wire \eeprom.n2525 ;
    wire \eeprom.n2526 ;
    wire \eeprom.n2527 ;
    wire \eeprom.n2528 ;
    wire \eeprom.n2529 ;
    wire \eeprom.n2530 ;
    wire n6_adj_397_cascade_;
    wire n2662_cascade_;
    wire n2668;
    wire \eeprom.delay_counter_0 ;
    wire \eeprom.delay_counter_2 ;
    wire \eeprom.delay_counter_5 ;
    wire \eeprom.delay_counter_10 ;
    wire \eeprom.n24_cascade_ ;
    wire \eeprom.n1338_cascade_ ;
    wire \eeprom.n575 ;
    wire \eeprom.n1435 ;
    wire \eeprom.n1435_cascade_ ;
    wire \eeprom.n1503 ;
    wire \eeprom.delay_counter_6 ;
    wire \eeprom.delay_counter_12 ;
    wire \eeprom.n16 ;
    wire n624_cascade_;
    wire \eeprom.delay_counter_14 ;
    wire \eeprom.delay_counter_11 ;
    wire \eeprom.delay_counter_15 ;
    wire \eeprom.delay_counter_9 ;
    wire \eeprom.delay_counter_1 ;
    wire \eeprom.delay_counter_7 ;
    wire \eeprom.n2685_cascade_ ;
    wire \eeprom.delay_counter_3 ;
    wire \eeprom.n22 ;
    wire \eeprom.delay_counter_13 ;
    wire \eeprom.delay_counter_8 ;
    wire \eeprom.delay_counter_4 ;
    wire \eeprom.n20 ;
    wire \eeprom.i2c.n6_cascade_ ;
    wire \eeprom.i2c.counter2_7__N_256_cascade_ ;
    wire \eeprom.i2c.n1384 ;
    wire \eeprom.i2c.counter2_0 ;
    wire bfn_19_17_0_;
    wire \eeprom.i2c.counter2_1 ;
    wire \eeprom.i2c.n2531 ;
    wire \eeprom.i2c.counter2_2 ;
    wire \eeprom.i2c.n2532 ;
    wire \eeprom.i2c.counter2_3 ;
    wire \eeprom.i2c.n2533 ;
    wire \eeprom.i2c.n2534 ;
    wire \eeprom.i2c.counter2_4 ;
    wire \eeprom.i2c.counter2_7__N_256 ;
    wire read;
    wire state_0;
    wire \eeprom.n1338 ;
    wire CLK_c;
    wire state_1;
    wire \eeprom.i2c.n2740_cascade_ ;
    wire \eeprom.i2c.n970 ;
    wire \eeprom.i2c.n2747_cascade_ ;
    wire \eeprom.i2c.n15_adj_381_cascade_ ;
    wire \eeprom.i2c.n2671 ;
    wire \eeprom.i2c.n2671_cascade_ ;
    wire rw;
    wire n15;
    wire state_7_N_269_0;
    wire n15_cascade_;
    wire \eeprom.i2c.n37 ;
    wire n7_adj_385;
    wire bfn_21_14_0_;
    wire \eeprom.i2c.n2509 ;
    wire \eeprom.i2c.n2510 ;
    wire \eeprom.i2c.n2511 ;
    wire \eeprom.i2c.n2512 ;
    wire \eeprom.i2c.n2513 ;
    wire \eeprom.i2c.n2514 ;
    wire CONSTANT_ONE_NET;
    wire \eeprom.i2c.n2515 ;
    wire \eeprom.i2c.n1413 ;
    wire \eeprom.i2c.n1495 ;
    wire \eeprom.i2c.n2734 ;
    wire \INVeeprom.i2c.sda_out_133C_net ;
    wire \eeprom.enable ;
    wire \INVeeprom.i2c.write_enable_132C_net ;
    wire \eeprom.i2c.n2736 ;
    wire \eeprom.i2c.n2664 ;
    wire \eeprom.i2c.n39_cascade_ ;
    wire \eeprom.i2c.n952 ;
    wire \eeprom.i2c.n33_cascade_ ;
    wire \eeprom.i2c.n16 ;
    wire \eeprom.i2c.n34_cascade_ ;
    wire \eeprom.i2c.n2616 ;
    wire \eeprom.i2c.n36 ;
    wire \eeprom.i2c.n33 ;
    wire \eeprom.i2c.n36_cascade_ ;
    wire \eeprom.i2c.n1493 ;
    wire state_7_N_285_3;
    wire \eeprom.i2c.n11 ;
    wire saved_addr_0;
    wire \eeprom.i2c.n11_adj_377 ;
    wire \eeprom.i2c.n11_adj_378 ;
    wire \eeprom.i2c.counter_4 ;
    wire \eeprom.i2c.counter_6 ;
    wire \eeprom.i2c.counter_7 ;
    wire \eeprom.i2c.counter_5 ;
    wire \eeprom.i2c.counter_3 ;
    wire \eeprom.i2c.n10_adj_380_cascade_ ;
    wire \eeprom.i2c.counter_2 ;
    wire \eeprom.i2c.n2706 ;
    wire \eeprom.i2c.n2654 ;
    wire \eeprom.i2c.counter_1 ;
    wire \eeprom.i2c.n2063_cascade_ ;
    wire \eeprom.i2c.counter_0 ;
    wire \eeprom.i2c.n1358_cascade_ ;
    wire \eeprom.i2c.n2726 ;
    wire \eeprom.i2c.n876_cascade_ ;
    wire \eeprom.i2c.n2078 ;
    wire \eeprom.i2c.n11_adj_376 ;
    wire \eeprom.i2c.n21 ;
    wire \eeprom.i2c.n2714 ;
    wire \eeprom.i2c.n2741_cascade_ ;
    wire \eeprom.i2c.n10_adj_379 ;
    wire \eeprom.i2c.n2018 ;
    wire sda_enable;
    wire \eeprom.i2c.n10 ;
    wire \eeprom.i2c.sda_out ;
    wire \eeprom.i2c.n876 ;
    wire \eeprom.i2c.n2008 ;
    wire \INVeeprom.i2c.i2c_scl_enable_124C_net ;
    wire \eeprom.i2c.n9 ;
    wire \eeprom.state_3 ;
    wire state_0_adj_386;
    wire \eeprom.state_1_adj_383 ;
    wire \eeprom.state_2 ;
    wire \eeprom.i2c.n11_adj_382 ;
    wire scl_enable;
    wire \eeprom.i2c.i2c_clk ;
    wire scl_c;
    wire _gnd_net_;

    defparam CS_CLK_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam CS_CLK_pad_iopad.PULLUP=1'b0;
    IO_PAD CS_CLK_pad_iopad (
            .OE(N__5901),
            .DIN(N__5900),
            .DOUT(N__5899),
            .PACKAGEPIN(CS_CLK));
    defparam CS_CLK_pad_preio.PIN_TYPE=6'b011001;
    defparam CS_CLK_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO CS_CLK_pad_preio (
            .PADOEN(N__5901),
            .PADOUT(N__5900),
            .PADIN(N__5899),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam CS_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam CS_pad_iopad.PULLUP=1'b0;
    IO_PAD CS_pad_iopad (
            .OE(N__5892),
            .DIN(N__5891),
            .DOUT(N__5890),
            .PACKAGEPIN(CS));
    defparam CS_pad_preio.PIN_TYPE=6'b011001;
    defparam CS_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO CS_pad_preio (
            .PADOEN(N__5892),
            .PADOUT(N__5891),
            .PADIN(N__5890),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam DE_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam DE_pad_iopad.PULLUP=1'b0;
    IO_PAD DE_pad_iopad (
            .OE(N__5883),
            .DIN(N__5882),
            .DOUT(N__5881),
            .PACKAGEPIN(DE));
    defparam DE_pad_preio.PIN_TYPE=6'b011001;
    defparam DE_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO DE_pad_preio (
            .PADOEN(N__5883),
            .PADOUT(N__5882),
            .PADIN(N__5881),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam INHA_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam INHA_pad_iopad.PULLUP=1'b0;
    IO_PAD INHA_pad_iopad (
            .OE(N__5874),
            .DIN(N__5873),
            .DOUT(N__5872),
            .PACKAGEPIN(INHA));
    defparam INHA_pad_preio.PIN_TYPE=6'b011001;
    defparam INHA_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO INHA_pad_preio (
            .PADOEN(N__5874),
            .PADOUT(N__5873),
            .PADIN(N__5872),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam INHB_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam INHB_pad_iopad.PULLUP=1'b0;
    IO_PAD INHB_pad_iopad (
            .OE(N__5865),
            .DIN(N__5864),
            .DOUT(N__5863),
            .PACKAGEPIN(INHB));
    defparam INHB_pad_preio.PIN_TYPE=6'b011001;
    defparam INHB_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO INHB_pad_preio (
            .PADOEN(N__5865),
            .PADOUT(N__5864),
            .PADIN(N__5863),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam INHC_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam INHC_pad_iopad.PULLUP=1'b0;
    IO_PAD INHC_pad_iopad (
            .OE(N__5856),
            .DIN(N__5855),
            .DOUT(N__5854),
            .PACKAGEPIN(INHC));
    defparam INHC_pad_preio.PIN_TYPE=6'b011001;
    defparam INHC_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO INHC_pad_preio (
            .PADOEN(N__5856),
            .PADOUT(N__5855),
            .PADIN(N__5854),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam INLA_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam INLA_pad_iopad.PULLUP=1'b0;
    IO_PAD INLA_pad_iopad (
            .OE(N__5847),
            .DIN(N__5846),
            .DOUT(N__5845),
            .PACKAGEPIN(INLA));
    defparam INLA_pad_preio.PIN_TYPE=6'b011001;
    defparam INLA_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO INLA_pad_preio (
            .PADOEN(N__5847),
            .PADOUT(N__5846),
            .PADIN(N__5845),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam INLB_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam INLB_pad_iopad.PULLUP=1'b0;
    IO_PAD INLB_pad_iopad (
            .OE(N__5838),
            .DIN(N__5837),
            .DOUT(N__5836),
            .PACKAGEPIN(INLB));
    defparam INLB_pad_preio.PIN_TYPE=6'b011001;
    defparam INLB_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO INLB_pad_preio (
            .PADOEN(N__5838),
            .PADOUT(N__5837),
            .PADIN(N__5836),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam INLC_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam INLC_pad_iopad.PULLUP=1'b0;
    IO_PAD INLC_pad_iopad (
            .OE(N__5829),
            .DIN(N__5828),
            .DOUT(N__5827),
            .PACKAGEPIN(INLC));
    defparam INLC_pad_preio.PIN_TYPE=6'b011001;
    defparam INLC_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO INLC_pad_preio (
            .PADOEN(N__5829),
            .PADOUT(N__5828),
            .PADIN(N__5827),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam LED_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam LED_pad_iopad.PULLUP=1'b0;
    IO_PAD LED_pad_iopad (
            .OE(N__5820),
            .DIN(N__5819),
            .DOUT(N__5818),
            .PACKAGEPIN(LED));
    defparam LED_pad_preio.PIN_TYPE=6'b011001;
    defparam LED_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO LED_pad_preio (
            .PADOEN(N__5820),
            .PADOUT(N__5819),
            .PADIN(N__5818),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__2723),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam NEOPXL_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam NEOPXL_pad_iopad.PULLUP=1'b0;
    IO_PAD NEOPXL_pad_iopad (
            .OE(N__5811),
            .DIN(N__5810),
            .DOUT(N__5809),
            .PACKAGEPIN(NEOPXL));
    defparam NEOPXL_pad_preio.PIN_TYPE=6'b011001;
    defparam NEOPXL_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO NEOPXL_pad_preio (
            .PADOEN(N__5811),
            .PADOUT(N__5810),
            .PADIN(N__5809),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam TX_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam TX_pad_iopad.PULLUP=1'b0;
    IO_PAD TX_pad_iopad (
            .OE(N__5802),
            .DIN(N__5801),
            .DOUT(N__5800),
            .PACKAGEPIN(TX));
    defparam TX_pad_preio.PIN_TYPE=6'b011001;
    defparam TX_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO TX_pad_preio (
            .PADOEN(N__5802),
            .PADOUT(N__5801),
            .PADIN(N__5800),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam USBPU_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam USBPU_pad_iopad.PULLUP=1'b0;
    IO_PAD USBPU_pad_iopad (
            .OE(N__5793),
            .DIN(N__5792),
            .DOUT(N__5791),
            .PACKAGEPIN(USBPU));
    defparam USBPU_pad_preio.PIN_TYPE=6'b011001;
    defparam USBPU_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO USBPU_pad_preio (
            .PADOEN(N__5793),
            .PADOUT(N__5792),
            .PADIN(N__5791),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam scl_output_iopad.IO_STANDARD="SB_LVCMOS";
    defparam scl_output_iopad.PULLUP=1'b1;
    IO_PAD scl_output_iopad (
            .OE(N__5784),
            .DIN(N__5783),
            .DOUT(N__5782),
            .PACKAGEPIN(SCL));
    defparam scl_output_preio.PIN_TYPE=6'b101001;
    defparam scl_output_preio.NEG_TRIGGER=1'b0;
    PRE_IO scl_output_preio (
            .PADOEN(N__5784),
            .PADOUT(N__5783),
            .PADIN(N__5782),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__4859),
            .DOUT1(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__5000));
    defparam sda_output_iopad.IO_STANDARD="SB_LVCMOS";
    defparam sda_output_iopad.PULLUP=1'b1;
    IO_PAD sda_output_iopad (
            .OE(N__5775),
            .DIN(N__5774),
            .DOUT(N__5773),
            .PACKAGEPIN(SDA));
    defparam sda_output_preio.PIN_TYPE=6'b101001;
    defparam sda_output_preio.NEG_TRIGGER=1'b0;
    PRE_IO sda_output_preio (
            .PADOEN(N__5775),
            .PADOUT(N__5774),
            .PADIN(N__5773),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__4493),
            .DOUT1(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__5717));
    defparam CLK_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam CLK_pad_iopad.PULLUP=1'b0;
    IO_PAD CLK_pad_iopad (
            .OE(N__5766),
            .DIN(N__5765),
            .DOUT(N__5764),
            .PACKAGEPIN(CLK));
    defparam CLK_pad_preio.PIN_TYPE=6'b000001;
    defparam CLK_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO CLK_pad_preio (
            .PADOEN(N__5766),
            .PADOUT(N__5765),
            .PADIN(N__5764),
            .CLOCKENABLE(),
            .DIN0(CLK_pad_gb_input),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    InMux I__1302 (
            .O(N__5747),
            .I(N__5743));
    InMux I__1301 (
            .O(N__5746),
            .I(N__5740));
    LocalMux I__1300 (
            .O(N__5743),
            .I(N__5737));
    LocalMux I__1299 (
            .O(N__5740),
            .I(\eeprom.i2c.n10_adj_379 ));
    Odrv4 I__1298 (
            .O(N__5737),
            .I(\eeprom.i2c.n10_adj_379 ));
    InMux I__1297 (
            .O(N__5732),
            .I(N__5728));
    InMux I__1296 (
            .O(N__5731),
            .I(N__5725));
    LocalMux I__1295 (
            .O(N__5728),
            .I(N__5720));
    LocalMux I__1294 (
            .O(N__5725),
            .I(N__5720));
    Odrv4 I__1293 (
            .O(N__5720),
            .I(\eeprom.i2c.n2018 ));
    IoInMux I__1292 (
            .O(N__5717),
            .I(N__5714));
    LocalMux I__1291 (
            .O(N__5714),
            .I(N__5710));
    InMux I__1290 (
            .O(N__5713),
            .I(N__5707));
    Span12Mux_s11_h I__1289 (
            .O(N__5710),
            .I(N__5702));
    LocalMux I__1288 (
            .O(N__5707),
            .I(N__5699));
    InMux I__1287 (
            .O(N__5706),
            .I(N__5696));
    InMux I__1286 (
            .O(N__5705),
            .I(N__5693));
    Odrv12 I__1285 (
            .O(N__5702),
            .I(sda_enable));
    Odrv4 I__1284 (
            .O(N__5699),
            .I(sda_enable));
    LocalMux I__1283 (
            .O(N__5696),
            .I(sda_enable));
    LocalMux I__1282 (
            .O(N__5693),
            .I(sda_enable));
    CascadeMux I__1281 (
            .O(N__5684),
            .I(N__5679));
    InMux I__1280 (
            .O(N__5683),
            .I(N__5676));
    InMux I__1279 (
            .O(N__5682),
            .I(N__5673));
    InMux I__1278 (
            .O(N__5679),
            .I(N__5670));
    LocalMux I__1277 (
            .O(N__5676),
            .I(N__5667));
    LocalMux I__1276 (
            .O(N__5673),
            .I(N__5664));
    LocalMux I__1275 (
            .O(N__5670),
            .I(\eeprom.i2c.n10 ));
    Odrv4 I__1274 (
            .O(N__5667),
            .I(\eeprom.i2c.n10 ));
    Odrv4 I__1273 (
            .O(N__5664),
            .I(\eeprom.i2c.n10 ));
    InMux I__1272 (
            .O(N__5657),
            .I(N__5654));
    LocalMux I__1271 (
            .O(N__5654),
            .I(N__5651));
    Span4Mux_h I__1270 (
            .O(N__5651),
            .I(N__5646));
    InMux I__1269 (
            .O(N__5650),
            .I(N__5643));
    InMux I__1268 (
            .O(N__5649),
            .I(N__5640));
    Odrv4 I__1267 (
            .O(N__5646),
            .I(\eeprom.i2c.sda_out ));
    LocalMux I__1266 (
            .O(N__5643),
            .I(\eeprom.i2c.sda_out ));
    LocalMux I__1265 (
            .O(N__5640),
            .I(\eeprom.i2c.sda_out ));
    CascadeMux I__1264 (
            .O(N__5633),
            .I(N__5627));
    CEMux I__1263 (
            .O(N__5632),
            .I(N__5622));
    CEMux I__1262 (
            .O(N__5631),
            .I(N__5619));
    CEMux I__1261 (
            .O(N__5630),
            .I(N__5616));
    InMux I__1260 (
            .O(N__5627),
            .I(N__5613));
    InMux I__1259 (
            .O(N__5626),
            .I(N__5608));
    InMux I__1258 (
            .O(N__5625),
            .I(N__5608));
    LocalMux I__1257 (
            .O(N__5622),
            .I(\eeprom.i2c.n876 ));
    LocalMux I__1256 (
            .O(N__5619),
            .I(\eeprom.i2c.n876 ));
    LocalMux I__1255 (
            .O(N__5616),
            .I(\eeprom.i2c.n876 ));
    LocalMux I__1254 (
            .O(N__5613),
            .I(\eeprom.i2c.n876 ));
    LocalMux I__1253 (
            .O(N__5608),
            .I(\eeprom.i2c.n876 ));
    SRMux I__1252 (
            .O(N__5597),
            .I(N__5594));
    LocalMux I__1251 (
            .O(N__5594),
            .I(N__5591));
    Odrv4 I__1250 (
            .O(N__5591),
            .I(\eeprom.i2c.n2008 ));
    CascadeMux I__1249 (
            .O(N__5588),
            .I(N__5585));
    InMux I__1248 (
            .O(N__5585),
            .I(N__5582));
    LocalMux I__1247 (
            .O(N__5582),
            .I(\eeprom.i2c.n9 ));
    InMux I__1246 (
            .O(N__5579),
            .I(N__5575));
    InMux I__1245 (
            .O(N__5578),
            .I(N__5570));
    LocalMux I__1244 (
            .O(N__5575),
            .I(N__5559));
    InMux I__1243 (
            .O(N__5574),
            .I(N__5556));
    InMux I__1242 (
            .O(N__5573),
            .I(N__5553));
    LocalMux I__1241 (
            .O(N__5570),
            .I(N__5550));
    InMux I__1240 (
            .O(N__5569),
            .I(N__5547));
    InMux I__1239 (
            .O(N__5568),
            .I(N__5539));
    InMux I__1238 (
            .O(N__5567),
            .I(N__5539));
    InMux I__1237 (
            .O(N__5566),
            .I(N__5539));
    InMux I__1236 (
            .O(N__5565),
            .I(N__5536));
    InMux I__1235 (
            .O(N__5564),
            .I(N__5532));
    CascadeMux I__1234 (
            .O(N__5563),
            .I(N__5527));
    InMux I__1233 (
            .O(N__5562),
            .I(N__5521));
    Span4Mux_h I__1232 (
            .O(N__5559),
            .I(N__5514));
    LocalMux I__1231 (
            .O(N__5556),
            .I(N__5514));
    LocalMux I__1230 (
            .O(N__5553),
            .I(N__5514));
    Span4Mux_h I__1229 (
            .O(N__5550),
            .I(N__5509));
    LocalMux I__1228 (
            .O(N__5547),
            .I(N__5509));
    InMux I__1227 (
            .O(N__5546),
            .I(N__5506));
    LocalMux I__1226 (
            .O(N__5539),
            .I(N__5501));
    LocalMux I__1225 (
            .O(N__5536),
            .I(N__5501));
    InMux I__1224 (
            .O(N__5535),
            .I(N__5493));
    LocalMux I__1223 (
            .O(N__5532),
            .I(N__5490));
    InMux I__1222 (
            .O(N__5531),
            .I(N__5483));
    InMux I__1221 (
            .O(N__5530),
            .I(N__5483));
    InMux I__1220 (
            .O(N__5527),
            .I(N__5483));
    InMux I__1219 (
            .O(N__5526),
            .I(N__5476));
    InMux I__1218 (
            .O(N__5525),
            .I(N__5476));
    InMux I__1217 (
            .O(N__5524),
            .I(N__5476));
    LocalMux I__1216 (
            .O(N__5521),
            .I(N__5473));
    Span4Mux_v I__1215 (
            .O(N__5514),
            .I(N__5466));
    Span4Mux_v I__1214 (
            .O(N__5509),
            .I(N__5466));
    LocalMux I__1213 (
            .O(N__5506),
            .I(N__5466));
    Span4Mux_h I__1212 (
            .O(N__5501),
            .I(N__5463));
    InMux I__1211 (
            .O(N__5500),
            .I(N__5456));
    InMux I__1210 (
            .O(N__5499),
            .I(N__5456));
    InMux I__1209 (
            .O(N__5498),
            .I(N__5456));
    InMux I__1208 (
            .O(N__5497),
            .I(N__5451));
    InMux I__1207 (
            .O(N__5496),
            .I(N__5451));
    LocalMux I__1206 (
            .O(N__5493),
            .I(N__5448));
    Odrv4 I__1205 (
            .O(N__5490),
            .I(\eeprom.state_3 ));
    LocalMux I__1204 (
            .O(N__5483),
            .I(\eeprom.state_3 ));
    LocalMux I__1203 (
            .O(N__5476),
            .I(\eeprom.state_3 ));
    Odrv12 I__1202 (
            .O(N__5473),
            .I(\eeprom.state_3 ));
    Odrv4 I__1201 (
            .O(N__5466),
            .I(\eeprom.state_3 ));
    Odrv4 I__1200 (
            .O(N__5463),
            .I(\eeprom.state_3 ));
    LocalMux I__1199 (
            .O(N__5456),
            .I(\eeprom.state_3 ));
    LocalMux I__1198 (
            .O(N__5451),
            .I(\eeprom.state_3 ));
    Odrv4 I__1197 (
            .O(N__5448),
            .I(\eeprom.state_3 ));
    InMux I__1196 (
            .O(N__5429),
            .I(N__5425));
    CascadeMux I__1195 (
            .O(N__5428),
            .I(N__5416));
    LocalMux I__1194 (
            .O(N__5425),
            .I(N__5411));
    InMux I__1193 (
            .O(N__5424),
            .I(N__5408));
    InMux I__1192 (
            .O(N__5423),
            .I(N__5405));
    InMux I__1191 (
            .O(N__5422),
            .I(N__5402));
    InMux I__1190 (
            .O(N__5421),
            .I(N__5392));
    InMux I__1189 (
            .O(N__5420),
            .I(N__5389));
    InMux I__1188 (
            .O(N__5419),
            .I(N__5384));
    InMux I__1187 (
            .O(N__5416),
            .I(N__5384));
    InMux I__1186 (
            .O(N__5415),
            .I(N__5381));
    InMux I__1185 (
            .O(N__5414),
            .I(N__5378));
    Span4Mux_v I__1184 (
            .O(N__5411),
            .I(N__5373));
    LocalMux I__1183 (
            .O(N__5408),
            .I(N__5373));
    LocalMux I__1182 (
            .O(N__5405),
            .I(N__5368));
    LocalMux I__1181 (
            .O(N__5402),
            .I(N__5368));
    CascadeMux I__1180 (
            .O(N__5401),
            .I(N__5361));
    CascadeMux I__1179 (
            .O(N__5400),
            .I(N__5357));
    InMux I__1178 (
            .O(N__5399),
            .I(N__5353));
    InMux I__1177 (
            .O(N__5398),
            .I(N__5350));
    InMux I__1176 (
            .O(N__5397),
            .I(N__5347));
    InMux I__1175 (
            .O(N__5396),
            .I(N__5342));
    InMux I__1174 (
            .O(N__5395),
            .I(N__5342));
    LocalMux I__1173 (
            .O(N__5392),
            .I(N__5335));
    LocalMux I__1172 (
            .O(N__5389),
            .I(N__5335));
    LocalMux I__1171 (
            .O(N__5384),
            .I(N__5335));
    LocalMux I__1170 (
            .O(N__5381),
            .I(N__5328));
    LocalMux I__1169 (
            .O(N__5378),
            .I(N__5328));
    Span4Mux_h I__1168 (
            .O(N__5373),
            .I(N__5328));
    Span4Mux_h I__1167 (
            .O(N__5368),
            .I(N__5325));
    InMux I__1166 (
            .O(N__5367),
            .I(N__5316));
    InMux I__1165 (
            .O(N__5366),
            .I(N__5316));
    InMux I__1164 (
            .O(N__5365),
            .I(N__5316));
    InMux I__1163 (
            .O(N__5364),
            .I(N__5316));
    InMux I__1162 (
            .O(N__5361),
            .I(N__5313));
    InMux I__1161 (
            .O(N__5360),
            .I(N__5310));
    InMux I__1160 (
            .O(N__5357),
            .I(N__5305));
    InMux I__1159 (
            .O(N__5356),
            .I(N__5305));
    LocalMux I__1158 (
            .O(N__5353),
            .I(state_0_adj_386));
    LocalMux I__1157 (
            .O(N__5350),
            .I(state_0_adj_386));
    LocalMux I__1156 (
            .O(N__5347),
            .I(state_0_adj_386));
    LocalMux I__1155 (
            .O(N__5342),
            .I(state_0_adj_386));
    Odrv4 I__1154 (
            .O(N__5335),
            .I(state_0_adj_386));
    Odrv4 I__1153 (
            .O(N__5328),
            .I(state_0_adj_386));
    Odrv4 I__1152 (
            .O(N__5325),
            .I(state_0_adj_386));
    LocalMux I__1151 (
            .O(N__5316),
            .I(state_0_adj_386));
    LocalMux I__1150 (
            .O(N__5313),
            .I(state_0_adj_386));
    LocalMux I__1149 (
            .O(N__5310),
            .I(state_0_adj_386));
    LocalMux I__1148 (
            .O(N__5305),
            .I(state_0_adj_386));
    CascadeMux I__1147 (
            .O(N__5282),
            .I(N__5274));
    CascadeMux I__1146 (
            .O(N__5281),
            .I(N__5271));
    CascadeMux I__1145 (
            .O(N__5280),
            .I(N__5267));
    CascadeMux I__1144 (
            .O(N__5279),
            .I(N__5263));
    InMux I__1143 (
            .O(N__5278),
            .I(N__5254));
    InMux I__1142 (
            .O(N__5277),
            .I(N__5249));
    InMux I__1141 (
            .O(N__5274),
            .I(N__5249));
    InMux I__1140 (
            .O(N__5271),
            .I(N__5246));
    InMux I__1139 (
            .O(N__5270),
            .I(N__5241));
    InMux I__1138 (
            .O(N__5267),
            .I(N__5241));
    InMux I__1137 (
            .O(N__5266),
            .I(N__5238));
    InMux I__1136 (
            .O(N__5263),
            .I(N__5233));
    CascadeMux I__1135 (
            .O(N__5262),
            .I(N__5230));
    InMux I__1134 (
            .O(N__5261),
            .I(N__5227));
    InMux I__1133 (
            .O(N__5260),
            .I(N__5222));
    InMux I__1132 (
            .O(N__5259),
            .I(N__5222));
    InMux I__1131 (
            .O(N__5258),
            .I(N__5217));
    InMux I__1130 (
            .O(N__5257),
            .I(N__5217));
    LocalMux I__1129 (
            .O(N__5254),
            .I(N__5214));
    LocalMux I__1128 (
            .O(N__5249),
            .I(N__5211));
    LocalMux I__1127 (
            .O(N__5246),
            .I(N__5204));
    LocalMux I__1126 (
            .O(N__5241),
            .I(N__5204));
    LocalMux I__1125 (
            .O(N__5238),
            .I(N__5204));
    CascadeMux I__1124 (
            .O(N__5237),
            .I(N__5201));
    CascadeMux I__1123 (
            .O(N__5236),
            .I(N__5196));
    LocalMux I__1122 (
            .O(N__5233),
            .I(N__5189));
    InMux I__1121 (
            .O(N__5230),
            .I(N__5186));
    LocalMux I__1120 (
            .O(N__5227),
            .I(N__5179));
    LocalMux I__1119 (
            .O(N__5222),
            .I(N__5179));
    LocalMux I__1118 (
            .O(N__5217),
            .I(N__5179));
    Span4Mux_v I__1117 (
            .O(N__5214),
            .I(N__5172));
    Span4Mux_v I__1116 (
            .O(N__5211),
            .I(N__5172));
    Span4Mux_v I__1115 (
            .O(N__5204),
            .I(N__5172));
    InMux I__1114 (
            .O(N__5201),
            .I(N__5169));
    InMux I__1113 (
            .O(N__5200),
            .I(N__5162));
    InMux I__1112 (
            .O(N__5199),
            .I(N__5162));
    InMux I__1111 (
            .O(N__5196),
            .I(N__5162));
    InMux I__1110 (
            .O(N__5195),
            .I(N__5159));
    InMux I__1109 (
            .O(N__5194),
            .I(N__5152));
    InMux I__1108 (
            .O(N__5193),
            .I(N__5152));
    InMux I__1107 (
            .O(N__5192),
            .I(N__5152));
    Odrv4 I__1106 (
            .O(N__5189),
            .I(\eeprom.state_1_adj_383 ));
    LocalMux I__1105 (
            .O(N__5186),
            .I(\eeprom.state_1_adj_383 ));
    Odrv4 I__1104 (
            .O(N__5179),
            .I(\eeprom.state_1_adj_383 ));
    Odrv4 I__1103 (
            .O(N__5172),
            .I(\eeprom.state_1_adj_383 ));
    LocalMux I__1102 (
            .O(N__5169),
            .I(\eeprom.state_1_adj_383 ));
    LocalMux I__1101 (
            .O(N__5162),
            .I(\eeprom.state_1_adj_383 ));
    LocalMux I__1100 (
            .O(N__5159),
            .I(\eeprom.state_1_adj_383 ));
    LocalMux I__1099 (
            .O(N__5152),
            .I(\eeprom.state_1_adj_383 ));
    InMux I__1098 (
            .O(N__5135),
            .I(N__5120));
    InMux I__1097 (
            .O(N__5134),
            .I(N__5114));
    InMux I__1096 (
            .O(N__5133),
            .I(N__5114));
    InMux I__1095 (
            .O(N__5132),
            .I(N__5111));
    InMux I__1094 (
            .O(N__5131),
            .I(N__5108));
    InMux I__1093 (
            .O(N__5130),
            .I(N__5101));
    InMux I__1092 (
            .O(N__5129),
            .I(N__5101));
    InMux I__1091 (
            .O(N__5128),
            .I(N__5101));
    InMux I__1090 (
            .O(N__5127),
            .I(N__5098));
    InMux I__1089 (
            .O(N__5126),
            .I(N__5094));
    InMux I__1088 (
            .O(N__5125),
            .I(N__5087));
    InMux I__1087 (
            .O(N__5124),
            .I(N__5087));
    InMux I__1086 (
            .O(N__5123),
            .I(N__5087));
    LocalMux I__1085 (
            .O(N__5120),
            .I(N__5083));
    InMux I__1084 (
            .O(N__5119),
            .I(N__5080));
    LocalMux I__1083 (
            .O(N__5114),
            .I(N__5071));
    LocalMux I__1082 (
            .O(N__5111),
            .I(N__5071));
    LocalMux I__1081 (
            .O(N__5108),
            .I(N__5071));
    LocalMux I__1080 (
            .O(N__5101),
            .I(N__5071));
    LocalMux I__1079 (
            .O(N__5098),
            .I(N__5061));
    InMux I__1078 (
            .O(N__5097),
            .I(N__5058));
    LocalMux I__1077 (
            .O(N__5094),
            .I(N__5055));
    LocalMux I__1076 (
            .O(N__5087),
            .I(N__5052));
    InMux I__1075 (
            .O(N__5086),
            .I(N__5049));
    Span4Mux_v I__1074 (
            .O(N__5083),
            .I(N__5042));
    LocalMux I__1073 (
            .O(N__5080),
            .I(N__5042));
    Span4Mux_v I__1072 (
            .O(N__5071),
            .I(N__5042));
    InMux I__1071 (
            .O(N__5070),
            .I(N__5035));
    InMux I__1070 (
            .O(N__5069),
            .I(N__5035));
    InMux I__1069 (
            .O(N__5068),
            .I(N__5035));
    InMux I__1068 (
            .O(N__5067),
            .I(N__5026));
    InMux I__1067 (
            .O(N__5066),
            .I(N__5026));
    InMux I__1066 (
            .O(N__5065),
            .I(N__5026));
    InMux I__1065 (
            .O(N__5064),
            .I(N__5026));
    Odrv4 I__1064 (
            .O(N__5061),
            .I(\eeprom.state_2 ));
    LocalMux I__1063 (
            .O(N__5058),
            .I(\eeprom.state_2 ));
    Odrv4 I__1062 (
            .O(N__5055),
            .I(\eeprom.state_2 ));
    Odrv4 I__1061 (
            .O(N__5052),
            .I(\eeprom.state_2 ));
    LocalMux I__1060 (
            .O(N__5049),
            .I(\eeprom.state_2 ));
    Odrv4 I__1059 (
            .O(N__5042),
            .I(\eeprom.state_2 ));
    LocalMux I__1058 (
            .O(N__5035),
            .I(\eeprom.state_2 ));
    LocalMux I__1057 (
            .O(N__5026),
            .I(\eeprom.state_2 ));
    CascadeMux I__1056 (
            .O(N__5009),
            .I(N__5006));
    InMux I__1055 (
            .O(N__5006),
            .I(N__5003));
    LocalMux I__1054 (
            .O(N__5003),
            .I(\eeprom.i2c.n11_adj_382 ));
    IoInMux I__1053 (
            .O(N__5000),
            .I(N__4997));
    LocalMux I__1052 (
            .O(N__4997),
            .I(N__4994));
    Span4Mux_s2_h I__1051 (
            .O(N__4994),
            .I(N__4991));
    Span4Mux_v I__1050 (
            .O(N__4991),
            .I(N__4987));
    InMux I__1049 (
            .O(N__4990),
            .I(N__4984));
    Sp12to4 I__1048 (
            .O(N__4987),
            .I(N__4979));
    LocalMux I__1047 (
            .O(N__4984),
            .I(N__4979));
    Odrv12 I__1046 (
            .O(N__4979),
            .I(scl_enable));
    ClkMux I__1045 (
            .O(N__4976),
            .I(N__4969));
    ClkMux I__1044 (
            .O(N__4975),
            .I(N__4966));
    ClkMux I__1043 (
            .O(N__4974),
            .I(N__4963));
    ClkMux I__1042 (
            .O(N__4973),
            .I(N__4960));
    InMux I__1041 (
            .O(N__4972),
            .I(N__4957));
    LocalMux I__1040 (
            .O(N__4969),
            .I(N__4950));
    LocalMux I__1039 (
            .O(N__4966),
            .I(N__4947));
    LocalMux I__1038 (
            .O(N__4963),
            .I(N__4941));
    LocalMux I__1037 (
            .O(N__4960),
            .I(N__4941));
    LocalMux I__1036 (
            .O(N__4957),
            .I(N__4938));
    ClkMux I__1035 (
            .O(N__4956),
            .I(N__4935));
    ClkMux I__1034 (
            .O(N__4955),
            .I(N__4932));
    ClkMux I__1033 (
            .O(N__4954),
            .I(N__4929));
    ClkMux I__1032 (
            .O(N__4953),
            .I(N__4926));
    Span4Mux_h I__1031 (
            .O(N__4950),
            .I(N__4921));
    Span4Mux_v I__1030 (
            .O(N__4947),
            .I(N__4921));
    ClkMux I__1029 (
            .O(N__4946),
            .I(N__4918));
    Span4Mux_v I__1028 (
            .O(N__4941),
            .I(N__4915));
    Span4Mux_v I__1027 (
            .O(N__4938),
            .I(N__4912));
    LocalMux I__1026 (
            .O(N__4935),
            .I(N__4907));
    LocalMux I__1025 (
            .O(N__4932),
            .I(N__4907));
    LocalMux I__1024 (
            .O(N__4929),
            .I(N__4904));
    LocalMux I__1023 (
            .O(N__4926),
            .I(N__4897));
    Span4Mux_h I__1022 (
            .O(N__4921),
            .I(N__4897));
    LocalMux I__1021 (
            .O(N__4918),
            .I(N__4897));
    Span4Mux_h I__1020 (
            .O(N__4915),
            .I(N__4891));
    Span4Mux_h I__1019 (
            .O(N__4912),
            .I(N__4886));
    Span4Mux_v I__1018 (
            .O(N__4907),
            .I(N__4886));
    Span4Mux_v I__1017 (
            .O(N__4904),
            .I(N__4883));
    Span4Mux_v I__1016 (
            .O(N__4897),
            .I(N__4880));
    InMux I__1015 (
            .O(N__4896),
            .I(N__4877));
    InMux I__1014 (
            .O(N__4895),
            .I(N__4872));
    InMux I__1013 (
            .O(N__4894),
            .I(N__4872));
    Odrv4 I__1012 (
            .O(N__4891),
            .I(\eeprom.i2c.i2c_clk ));
    Odrv4 I__1011 (
            .O(N__4886),
            .I(\eeprom.i2c.i2c_clk ));
    Odrv4 I__1010 (
            .O(N__4883),
            .I(\eeprom.i2c.i2c_clk ));
    Odrv4 I__1009 (
            .O(N__4880),
            .I(\eeprom.i2c.i2c_clk ));
    LocalMux I__1008 (
            .O(N__4877),
            .I(\eeprom.i2c.i2c_clk ));
    LocalMux I__1007 (
            .O(N__4872),
            .I(\eeprom.i2c.i2c_clk ));
    IoInMux I__1006 (
            .O(N__4859),
            .I(N__4856));
    LocalMux I__1005 (
            .O(N__4856),
            .I(N__4853));
    Span4Mux_s3_h I__1004 (
            .O(N__4853),
            .I(N__4850));
    Span4Mux_v I__1003 (
            .O(N__4850),
            .I(N__4847));
    Odrv4 I__1002 (
            .O(N__4847),
            .I(scl_c));
    InMux I__1001 (
            .O(N__4844),
            .I(N__4841));
    LocalMux I__1000 (
            .O(N__4841),
            .I(N__4837));
    InMux I__999 (
            .O(N__4840),
            .I(N__4834));
    Odrv12 I__998 (
            .O(N__4837),
            .I(\eeprom.i2c.n2654 ));
    LocalMux I__997 (
            .O(N__4834),
            .I(\eeprom.i2c.n2654 ));
    InMux I__996 (
            .O(N__4829),
            .I(N__4826));
    LocalMux I__995 (
            .O(N__4826),
            .I(N__4822));
    InMux I__994 (
            .O(N__4825),
            .I(N__4817));
    Span4Mux_h I__993 (
            .O(N__4822),
            .I(N__4814));
    InMux I__992 (
            .O(N__4821),
            .I(N__4809));
    InMux I__991 (
            .O(N__4820),
            .I(N__4809));
    LocalMux I__990 (
            .O(N__4817),
            .I(\eeprom.i2c.counter_1 ));
    Odrv4 I__989 (
            .O(N__4814),
            .I(\eeprom.i2c.counter_1 ));
    LocalMux I__988 (
            .O(N__4809),
            .I(\eeprom.i2c.counter_1 ));
    CascadeMux I__987 (
            .O(N__4802),
            .I(\eeprom.i2c.n2063_cascade_ ));
    InMux I__986 (
            .O(N__4799),
            .I(N__4796));
    LocalMux I__985 (
            .O(N__4796),
            .I(N__4792));
    InMux I__984 (
            .O(N__4795),
            .I(N__4786));
    Span4Mux_h I__983 (
            .O(N__4792),
            .I(N__4783));
    InMux I__982 (
            .O(N__4791),
            .I(N__4776));
    InMux I__981 (
            .O(N__4790),
            .I(N__4776));
    InMux I__980 (
            .O(N__4789),
            .I(N__4776));
    LocalMux I__979 (
            .O(N__4786),
            .I(\eeprom.i2c.counter_0 ));
    Odrv4 I__978 (
            .O(N__4783),
            .I(\eeprom.i2c.counter_0 ));
    LocalMux I__977 (
            .O(N__4776),
            .I(\eeprom.i2c.counter_0 ));
    CascadeMux I__976 (
            .O(N__4769),
            .I(\eeprom.i2c.n1358_cascade_ ));
    InMux I__975 (
            .O(N__4766),
            .I(N__4763));
    LocalMux I__974 (
            .O(N__4763),
            .I(N__4760));
    Odrv4 I__973 (
            .O(N__4760),
            .I(\eeprom.i2c.n2726 ));
    CascadeMux I__972 (
            .O(N__4757),
            .I(\eeprom.i2c.n876_cascade_ ));
    SRMux I__971 (
            .O(N__4754),
            .I(N__4751));
    LocalMux I__970 (
            .O(N__4751),
            .I(\eeprom.i2c.n2078 ));
    InMux I__969 (
            .O(N__4748),
            .I(N__4739));
    InMux I__968 (
            .O(N__4747),
            .I(N__4739));
    InMux I__967 (
            .O(N__4746),
            .I(N__4739));
    LocalMux I__966 (
            .O(N__4739),
            .I(\eeprom.i2c.n11_adj_376 ));
    InMux I__965 (
            .O(N__4736),
            .I(N__4733));
    LocalMux I__964 (
            .O(N__4733),
            .I(\eeprom.i2c.n21 ));
    InMux I__963 (
            .O(N__4730),
            .I(N__4727));
    LocalMux I__962 (
            .O(N__4727),
            .I(N__4724));
    Odrv12 I__961 (
            .O(N__4724),
            .I(\eeprom.i2c.n2714 ));
    CascadeMux I__960 (
            .O(N__4721),
            .I(\eeprom.i2c.n2741_cascade_ ));
    CascadeMux I__959 (
            .O(N__4718),
            .I(N__4715));
    InMux I__958 (
            .O(N__4715),
            .I(N__4710));
    InMux I__957 (
            .O(N__4714),
            .I(N__4707));
    InMux I__956 (
            .O(N__4713),
            .I(N__4704));
    LocalMux I__955 (
            .O(N__4710),
            .I(\eeprom.i2c.n11_adj_377 ));
    LocalMux I__954 (
            .O(N__4707),
            .I(\eeprom.i2c.n11_adj_377 ));
    LocalMux I__953 (
            .O(N__4704),
            .I(\eeprom.i2c.n11_adj_377 ));
    InMux I__952 (
            .O(N__4697),
            .I(N__4694));
    LocalMux I__951 (
            .O(N__4694),
            .I(N__4691));
    Odrv4 I__950 (
            .O(N__4691),
            .I(\eeprom.i2c.n11_adj_378 ));
    CascadeMux I__949 (
            .O(N__4688),
            .I(N__4684));
    InMux I__948 (
            .O(N__4687),
            .I(N__4681));
    InMux I__947 (
            .O(N__4684),
            .I(N__4678));
    LocalMux I__946 (
            .O(N__4681),
            .I(N__4675));
    LocalMux I__945 (
            .O(N__4678),
            .I(\eeprom.i2c.counter_4 ));
    Odrv4 I__944 (
            .O(N__4675),
            .I(\eeprom.i2c.counter_4 ));
    CascadeMux I__943 (
            .O(N__4670),
            .I(N__4666));
    InMux I__942 (
            .O(N__4669),
            .I(N__4663));
    InMux I__941 (
            .O(N__4666),
            .I(N__4660));
    LocalMux I__940 (
            .O(N__4663),
            .I(N__4657));
    LocalMux I__939 (
            .O(N__4660),
            .I(\eeprom.i2c.counter_6 ));
    Odrv12 I__938 (
            .O(N__4657),
            .I(\eeprom.i2c.counter_6 ));
    CascadeMux I__937 (
            .O(N__4652),
            .I(N__4649));
    InMux I__936 (
            .O(N__4649),
            .I(N__4645));
    InMux I__935 (
            .O(N__4648),
            .I(N__4642));
    LocalMux I__934 (
            .O(N__4645),
            .I(N__4639));
    LocalMux I__933 (
            .O(N__4642),
            .I(\eeprom.i2c.counter_7 ));
    Odrv4 I__932 (
            .O(N__4639),
            .I(\eeprom.i2c.counter_7 ));
    InMux I__931 (
            .O(N__4634),
            .I(N__4630));
    InMux I__930 (
            .O(N__4633),
            .I(N__4627));
    LocalMux I__929 (
            .O(N__4630),
            .I(N__4624));
    LocalMux I__928 (
            .O(N__4627),
            .I(\eeprom.i2c.counter_5 ));
    Odrv4 I__927 (
            .O(N__4624),
            .I(\eeprom.i2c.counter_5 ));
    InMux I__926 (
            .O(N__4619),
            .I(N__4615));
    InMux I__925 (
            .O(N__4618),
            .I(N__4612));
    LocalMux I__924 (
            .O(N__4615),
            .I(N__4609));
    LocalMux I__923 (
            .O(N__4612),
            .I(\eeprom.i2c.counter_3 ));
    Odrv4 I__922 (
            .O(N__4609),
            .I(\eeprom.i2c.counter_3 ));
    CascadeMux I__921 (
            .O(N__4604),
            .I(\eeprom.i2c.n10_adj_380_cascade_ ));
    CascadeMux I__920 (
            .O(N__4601),
            .I(N__4597));
    InMux I__919 (
            .O(N__4600),
            .I(N__4593));
    InMux I__918 (
            .O(N__4597),
            .I(N__4590));
    InMux I__917 (
            .O(N__4596),
            .I(N__4587));
    LocalMux I__916 (
            .O(N__4593),
            .I(N__4584));
    LocalMux I__915 (
            .O(N__4590),
            .I(\eeprom.i2c.counter_2 ));
    LocalMux I__914 (
            .O(N__4587),
            .I(\eeprom.i2c.counter_2 ));
    Odrv4 I__913 (
            .O(N__4584),
            .I(\eeprom.i2c.counter_2 ));
    SRMux I__912 (
            .O(N__4577),
            .I(N__4574));
    LocalMux I__911 (
            .O(N__4574),
            .I(\eeprom.i2c.n2706 ));
    CascadeMux I__910 (
            .O(N__4571),
            .I(\eeprom.i2c.n39_cascade_ ));
    CEMux I__909 (
            .O(N__4568),
            .I(N__4565));
    LocalMux I__908 (
            .O(N__4565),
            .I(N__4562));
    Span4Mux_h I__907 (
            .O(N__4562),
            .I(N__4559));
    Odrv4 I__906 (
            .O(N__4559),
            .I(\eeprom.i2c.n952 ));
    CascadeMux I__905 (
            .O(N__4556),
            .I(\eeprom.i2c.n33_cascade_ ));
    InMux I__904 (
            .O(N__4553),
            .I(N__4550));
    LocalMux I__903 (
            .O(N__4550),
            .I(\eeprom.i2c.n16 ));
    CascadeMux I__902 (
            .O(N__4547),
            .I(\eeprom.i2c.n34_cascade_ ));
    CEMux I__901 (
            .O(N__4544),
            .I(N__4541));
    LocalMux I__900 (
            .O(N__4541),
            .I(N__4538));
    Odrv4 I__899 (
            .O(N__4538),
            .I(\eeprom.i2c.n2616 ));
    InMux I__898 (
            .O(N__4535),
            .I(N__4532));
    LocalMux I__897 (
            .O(N__4532),
            .I(N__4527));
    InMux I__896 (
            .O(N__4531),
            .I(N__4522));
    InMux I__895 (
            .O(N__4530),
            .I(N__4522));
    Odrv4 I__894 (
            .O(N__4527),
            .I(\eeprom.i2c.n36 ));
    LocalMux I__893 (
            .O(N__4522),
            .I(\eeprom.i2c.n36 ));
    InMux I__892 (
            .O(N__4517),
            .I(N__4511));
    InMux I__891 (
            .O(N__4516),
            .I(N__4511));
    LocalMux I__890 (
            .O(N__4511),
            .I(\eeprom.i2c.n33 ));
    CascadeMux I__889 (
            .O(N__4508),
            .I(\eeprom.i2c.n36_cascade_ ));
    SRMux I__888 (
            .O(N__4505),
            .I(N__4502));
    LocalMux I__887 (
            .O(N__4502),
            .I(N__4499));
    Span4Mux_h I__886 (
            .O(N__4499),
            .I(N__4496));
    Odrv4 I__885 (
            .O(N__4496),
            .I(\eeprom.i2c.n1493 ));
    IoInMux I__884 (
            .O(N__4493),
            .I(N__4490));
    LocalMux I__883 (
            .O(N__4490),
            .I(N__4487));
    Span12Mux_s6_h I__882 (
            .O(N__4487),
            .I(N__4483));
    InMux I__881 (
            .O(N__4486),
            .I(N__4480));
    Span12Mux_v I__880 (
            .O(N__4483),
            .I(N__4476));
    LocalMux I__879 (
            .O(N__4480),
            .I(N__4473));
    InMux I__878 (
            .O(N__4479),
            .I(N__4470));
    Odrv12 I__877 (
            .O(N__4476),
            .I(state_7_N_285_3));
    Odrv4 I__876 (
            .O(N__4473),
            .I(state_7_N_285_3));
    LocalMux I__875 (
            .O(N__4470),
            .I(state_7_N_285_3));
    CascadeMux I__874 (
            .O(N__4463),
            .I(N__4460));
    InMux I__873 (
            .O(N__4460),
            .I(N__4457));
    LocalMux I__872 (
            .O(N__4457),
            .I(N__4454));
    Odrv12 I__871 (
            .O(N__4454),
            .I(\eeprom.i2c.n11 ));
    InMux I__870 (
            .O(N__4451),
            .I(N__4448));
    LocalMux I__869 (
            .O(N__4448),
            .I(N__4445));
    Span4Mux_v I__868 (
            .O(N__4445),
            .I(N__4440));
    InMux I__867 (
            .O(N__4444),
            .I(N__4437));
    InMux I__866 (
            .O(N__4443),
            .I(N__4434));
    Odrv4 I__865 (
            .O(N__4440),
            .I(saved_addr_0));
    LocalMux I__864 (
            .O(N__4437),
            .I(saved_addr_0));
    LocalMux I__863 (
            .O(N__4434),
            .I(saved_addr_0));
    InMux I__862 (
            .O(N__4427),
            .I(\eeprom.i2c.n2511 ));
    InMux I__861 (
            .O(N__4424),
            .I(\eeprom.i2c.n2512 ));
    InMux I__860 (
            .O(N__4421),
            .I(\eeprom.i2c.n2513 ));
    InMux I__859 (
            .O(N__4418),
            .I(\eeprom.i2c.n2514 ));
    CascadeMux I__858 (
            .O(N__4415),
            .I(N__4408));
    CascadeMux I__857 (
            .O(N__4414),
            .I(N__4404));
    CascadeMux I__856 (
            .O(N__4413),
            .I(N__4400));
    InMux I__855 (
            .O(N__4412),
            .I(N__4385));
    InMux I__854 (
            .O(N__4411),
            .I(N__4385));
    InMux I__853 (
            .O(N__4408),
            .I(N__4385));
    InMux I__852 (
            .O(N__4407),
            .I(N__4385));
    InMux I__851 (
            .O(N__4404),
            .I(N__4385));
    InMux I__850 (
            .O(N__4403),
            .I(N__4385));
    InMux I__849 (
            .O(N__4400),
            .I(N__4385));
    LocalMux I__848 (
            .O(N__4385),
            .I(CONSTANT_ONE_NET));
    InMux I__847 (
            .O(N__4382),
            .I(\eeprom.i2c.n2515 ));
    CEMux I__846 (
            .O(N__4379),
            .I(N__4376));
    LocalMux I__845 (
            .O(N__4376),
            .I(N__4373));
    Odrv4 I__844 (
            .O(N__4373),
            .I(\eeprom.i2c.n1413 ));
    SRMux I__843 (
            .O(N__4370),
            .I(N__4367));
    LocalMux I__842 (
            .O(N__4367),
            .I(N__4364));
    Span4Mux_h I__841 (
            .O(N__4364),
            .I(N__4361));
    Odrv4 I__840 (
            .O(N__4361),
            .I(\eeprom.i2c.n1495 ));
    InMux I__839 (
            .O(N__4358),
            .I(N__4355));
    LocalMux I__838 (
            .O(N__4355),
            .I(\eeprom.i2c.n2734 ));
    CascadeMux I__837 (
            .O(N__4352),
            .I(N__4348));
    SRMux I__836 (
            .O(N__4351),
            .I(N__4345));
    InMux I__835 (
            .O(N__4348),
            .I(N__4342));
    LocalMux I__834 (
            .O(N__4345),
            .I(N__4338));
    LocalMux I__833 (
            .O(N__4342),
            .I(N__4335));
    InMux I__832 (
            .O(N__4341),
            .I(N__4332));
    Span4Mux_h I__831 (
            .O(N__4338),
            .I(N__4329));
    Span4Mux_h I__830 (
            .O(N__4335),
            .I(N__4324));
    LocalMux I__829 (
            .O(N__4332),
            .I(N__4324));
    Odrv4 I__828 (
            .O(N__4329),
            .I(\eeprom.enable ));
    Odrv4 I__827 (
            .O(N__4324),
            .I(\eeprom.enable ));
    InMux I__826 (
            .O(N__4319),
            .I(N__4316));
    LocalMux I__825 (
            .O(N__4316),
            .I(\eeprom.i2c.n2736 ));
    CascadeMux I__824 (
            .O(N__4313),
            .I(N__4310));
    InMux I__823 (
            .O(N__4310),
            .I(N__4307));
    LocalMux I__822 (
            .O(N__4307),
            .I(N__4304));
    Span4Mux_v I__821 (
            .O(N__4304),
            .I(N__4301));
    Odrv4 I__820 (
            .O(N__4301),
            .I(\eeprom.i2c.n2664 ));
    CascadeMux I__819 (
            .O(N__4298),
            .I(n15_cascade_));
    InMux I__818 (
            .O(N__4295),
            .I(N__4292));
    LocalMux I__817 (
            .O(N__4292),
            .I(N__4289));
    Odrv4 I__816 (
            .O(N__4289),
            .I(\eeprom.i2c.n37 ));
    InMux I__815 (
            .O(N__4286),
            .I(N__4283));
    LocalMux I__814 (
            .O(N__4283),
            .I(N__4280));
    Odrv12 I__813 (
            .O(N__4280),
            .I(n7_adj_385));
    InMux I__812 (
            .O(N__4277),
            .I(bfn_21_14_0_));
    InMux I__811 (
            .O(N__4274),
            .I(\eeprom.i2c.n2509 ));
    InMux I__810 (
            .O(N__4271),
            .I(\eeprom.i2c.n2510 ));
    CascadeMux I__809 (
            .O(N__4268),
            .I(\eeprom.i2c.n2740_cascade_ ));
    InMux I__808 (
            .O(N__4265),
            .I(N__4262));
    LocalMux I__807 (
            .O(N__4262),
            .I(\eeprom.i2c.n970 ));
    CascadeMux I__806 (
            .O(N__4259),
            .I(\eeprom.i2c.n2747_cascade_ ));
    CascadeMux I__805 (
            .O(N__4256),
            .I(\eeprom.i2c.n15_adj_381_cascade_ ));
    InMux I__804 (
            .O(N__4253),
            .I(N__4250));
    LocalMux I__803 (
            .O(N__4250),
            .I(\eeprom.i2c.n2671 ));
    CascadeMux I__802 (
            .O(N__4247),
            .I(\eeprom.i2c.n2671_cascade_ ));
    CascadeMux I__801 (
            .O(N__4244),
            .I(N__4241));
    InMux I__800 (
            .O(N__4241),
            .I(N__4238));
    LocalMux I__799 (
            .O(N__4238),
            .I(N__4235));
    Span4Mux_h I__798 (
            .O(N__4235),
            .I(N__4232));
    Span4Mux_v I__797 (
            .O(N__4232),
            .I(N__4228));
    InMux I__796 (
            .O(N__4231),
            .I(N__4225));
    Odrv4 I__795 (
            .O(N__4228),
            .I(rw));
    LocalMux I__794 (
            .O(N__4225),
            .I(rw));
    InMux I__793 (
            .O(N__4220),
            .I(N__4211));
    InMux I__792 (
            .O(N__4219),
            .I(N__4211));
    InMux I__791 (
            .O(N__4218),
            .I(N__4208));
    CascadeMux I__790 (
            .O(N__4217),
            .I(N__4205));
    InMux I__789 (
            .O(N__4216),
            .I(N__4202));
    LocalMux I__788 (
            .O(N__4211),
            .I(N__4197));
    LocalMux I__787 (
            .O(N__4208),
            .I(N__4197));
    InMux I__786 (
            .O(N__4205),
            .I(N__4194));
    LocalMux I__785 (
            .O(N__4202),
            .I(N__4191));
    Span4Mux_v I__784 (
            .O(N__4197),
            .I(N__4188));
    LocalMux I__783 (
            .O(N__4194),
            .I(N__4185));
    Span4Mux_v I__782 (
            .O(N__4191),
            .I(N__4181));
    Sp12to4 I__781 (
            .O(N__4188),
            .I(N__4176));
    Span12Mux_v I__780 (
            .O(N__4185),
            .I(N__4176));
    InMux I__779 (
            .O(N__4184),
            .I(N__4173));
    Odrv4 I__778 (
            .O(N__4181),
            .I(n15));
    Odrv12 I__777 (
            .O(N__4176),
            .I(n15));
    LocalMux I__776 (
            .O(N__4173),
            .I(n15));
    InMux I__775 (
            .O(N__4166),
            .I(N__4160));
    InMux I__774 (
            .O(N__4165),
            .I(N__4160));
    LocalMux I__773 (
            .O(N__4160),
            .I(state_7_N_269_0));
    InMux I__772 (
            .O(N__4157),
            .I(N__4153));
    InMux I__771 (
            .O(N__4156),
            .I(N__4150));
    LocalMux I__770 (
            .O(N__4153),
            .I(\eeprom.i2c.counter2_0 ));
    LocalMux I__769 (
            .O(N__4150),
            .I(\eeprom.i2c.counter2_0 ));
    InMux I__768 (
            .O(N__4145),
            .I(bfn_19_17_0_));
    InMux I__767 (
            .O(N__4142),
            .I(N__4138));
    InMux I__766 (
            .O(N__4141),
            .I(N__4135));
    LocalMux I__765 (
            .O(N__4138),
            .I(\eeprom.i2c.counter2_1 ));
    LocalMux I__764 (
            .O(N__4135),
            .I(\eeprom.i2c.counter2_1 ));
    InMux I__763 (
            .O(N__4130),
            .I(\eeprom.i2c.n2531 ));
    InMux I__762 (
            .O(N__4127),
            .I(N__4123));
    InMux I__761 (
            .O(N__4126),
            .I(N__4120));
    LocalMux I__760 (
            .O(N__4123),
            .I(\eeprom.i2c.counter2_2 ));
    LocalMux I__759 (
            .O(N__4120),
            .I(\eeprom.i2c.counter2_2 ));
    InMux I__758 (
            .O(N__4115),
            .I(\eeprom.i2c.n2532 ));
    InMux I__757 (
            .O(N__4112),
            .I(N__4108));
    InMux I__756 (
            .O(N__4111),
            .I(N__4105));
    LocalMux I__755 (
            .O(N__4108),
            .I(\eeprom.i2c.counter2_3 ));
    LocalMux I__754 (
            .O(N__4105),
            .I(\eeprom.i2c.counter2_3 ));
    InMux I__753 (
            .O(N__4100),
            .I(\eeprom.i2c.n2533 ));
    InMux I__752 (
            .O(N__4097),
            .I(\eeprom.i2c.n2534 ));
    InMux I__751 (
            .O(N__4094),
            .I(N__4090));
    InMux I__750 (
            .O(N__4093),
            .I(N__4087));
    LocalMux I__749 (
            .O(N__4090),
            .I(\eeprom.i2c.counter2_4 ));
    LocalMux I__748 (
            .O(N__4087),
            .I(\eeprom.i2c.counter2_4 ));
    SRMux I__747 (
            .O(N__4082),
            .I(N__4079));
    LocalMux I__746 (
            .O(N__4079),
            .I(N__4076));
    Span4Mux_h I__745 (
            .O(N__4076),
            .I(N__4071));
    InMux I__744 (
            .O(N__4075),
            .I(N__4068));
    InMux I__743 (
            .O(N__4074),
            .I(N__4065));
    Odrv4 I__742 (
            .O(N__4071),
            .I(\eeprom.i2c.counter2_7__N_256 ));
    LocalMux I__741 (
            .O(N__4068),
            .I(\eeprom.i2c.counter2_7__N_256 ));
    LocalMux I__740 (
            .O(N__4065),
            .I(\eeprom.i2c.counter2_7__N_256 ));
    CascadeMux I__739 (
            .O(N__4058),
            .I(N__4053));
    InMux I__738 (
            .O(N__4057),
            .I(N__4046));
    InMux I__737 (
            .O(N__4056),
            .I(N__4046));
    InMux I__736 (
            .O(N__4053),
            .I(N__4043));
    InMux I__735 (
            .O(N__4052),
            .I(N__4040));
    InMux I__734 (
            .O(N__4051),
            .I(N__4037));
    LocalMux I__733 (
            .O(N__4046),
            .I(N__4034));
    LocalMux I__732 (
            .O(N__4043),
            .I(N__4029));
    LocalMux I__731 (
            .O(N__4040),
            .I(N__4029));
    LocalMux I__730 (
            .O(N__4037),
            .I(N__4026));
    Span4Mux_v I__729 (
            .O(N__4034),
            .I(N__4021));
    Span4Mux_h I__728 (
            .O(N__4029),
            .I(N__4021));
    Span12Mux_h I__727 (
            .O(N__4026),
            .I(N__4018));
    Span4Mux_v I__726 (
            .O(N__4021),
            .I(N__4015));
    Odrv12 I__725 (
            .O(N__4018),
            .I(read));
    Odrv4 I__724 (
            .O(N__4015),
            .I(read));
    InMux I__723 (
            .O(N__4010),
            .I(N__4007));
    LocalMux I__722 (
            .O(N__4007),
            .I(N__3995));
    InMux I__721 (
            .O(N__4006),
            .I(N__3992));
    InMux I__720 (
            .O(N__4005),
            .I(N__3987));
    InMux I__719 (
            .O(N__4004),
            .I(N__3987));
    InMux I__718 (
            .O(N__4003),
            .I(N__3978));
    InMux I__717 (
            .O(N__4002),
            .I(N__3978));
    InMux I__716 (
            .O(N__4001),
            .I(N__3978));
    InMux I__715 (
            .O(N__4000),
            .I(N__3978));
    InMux I__714 (
            .O(N__3999),
            .I(N__3973));
    InMux I__713 (
            .O(N__3998),
            .I(N__3973));
    Odrv4 I__712 (
            .O(N__3995),
            .I(state_0));
    LocalMux I__711 (
            .O(N__3992),
            .I(state_0));
    LocalMux I__710 (
            .O(N__3987),
            .I(state_0));
    LocalMux I__709 (
            .O(N__3978),
            .I(state_0));
    LocalMux I__708 (
            .O(N__3973),
            .I(state_0));
    CascadeMux I__707 (
            .O(N__3962),
            .I(N__3957));
    InMux I__706 (
            .O(N__3961),
            .I(N__3954));
    InMux I__705 (
            .O(N__3960),
            .I(N__3951));
    InMux I__704 (
            .O(N__3957),
            .I(N__3948));
    LocalMux I__703 (
            .O(N__3954),
            .I(\eeprom.n1338 ));
    LocalMux I__702 (
            .O(N__3951),
            .I(\eeprom.n1338 ));
    LocalMux I__701 (
            .O(N__3948),
            .I(\eeprom.n1338 ));
    ClkMux I__700 (
            .O(N__3941),
            .I(N__3890));
    ClkMux I__699 (
            .O(N__3940),
            .I(N__3890));
    ClkMux I__698 (
            .O(N__3939),
            .I(N__3890));
    ClkMux I__697 (
            .O(N__3938),
            .I(N__3890));
    ClkMux I__696 (
            .O(N__3937),
            .I(N__3890));
    ClkMux I__695 (
            .O(N__3936),
            .I(N__3890));
    ClkMux I__694 (
            .O(N__3935),
            .I(N__3890));
    ClkMux I__693 (
            .O(N__3934),
            .I(N__3890));
    ClkMux I__692 (
            .O(N__3933),
            .I(N__3890));
    ClkMux I__691 (
            .O(N__3932),
            .I(N__3890));
    ClkMux I__690 (
            .O(N__3931),
            .I(N__3890));
    ClkMux I__689 (
            .O(N__3930),
            .I(N__3890));
    ClkMux I__688 (
            .O(N__3929),
            .I(N__3890));
    ClkMux I__687 (
            .O(N__3928),
            .I(N__3890));
    ClkMux I__686 (
            .O(N__3927),
            .I(N__3890));
    ClkMux I__685 (
            .O(N__3926),
            .I(N__3890));
    ClkMux I__684 (
            .O(N__3925),
            .I(N__3890));
    GlobalMux I__683 (
            .O(N__3890),
            .I(N__3887));
    gio2CtrlBuf I__682 (
            .O(N__3887),
            .I(CLK_c));
    SRMux I__681 (
            .O(N__3884),
            .I(N__3881));
    LocalMux I__680 (
            .O(N__3881),
            .I(N__3878));
    Span4Mux_h I__679 (
            .O(N__3878),
            .I(N__3870));
    InMux I__678 (
            .O(N__3877),
            .I(N__3865));
    InMux I__677 (
            .O(N__3876),
            .I(N__3865));
    InMux I__676 (
            .O(N__3875),
            .I(N__3860));
    InMux I__675 (
            .O(N__3874),
            .I(N__3860));
    InMux I__674 (
            .O(N__3873),
            .I(N__3857));
    Odrv4 I__673 (
            .O(N__3870),
            .I(state_1));
    LocalMux I__672 (
            .O(N__3865),
            .I(state_1));
    LocalMux I__671 (
            .O(N__3860),
            .I(state_1));
    LocalMux I__670 (
            .O(N__3857),
            .I(state_1));
    CascadeMux I__669 (
            .O(N__3848),
            .I(n624_cascade_));
    CascadeMux I__668 (
            .O(N__3845),
            .I(N__3842));
    InMux I__667 (
            .O(N__3842),
            .I(N__3838));
    InMux I__666 (
            .O(N__3841),
            .I(N__3835));
    LocalMux I__665 (
            .O(N__3838),
            .I(\eeprom.delay_counter_14 ));
    LocalMux I__664 (
            .O(N__3835),
            .I(\eeprom.delay_counter_14 ));
    InMux I__663 (
            .O(N__3830),
            .I(N__3826));
    InMux I__662 (
            .O(N__3829),
            .I(N__3823));
    LocalMux I__661 (
            .O(N__3826),
            .I(\eeprom.delay_counter_11 ));
    LocalMux I__660 (
            .O(N__3823),
            .I(\eeprom.delay_counter_11 ));
    CascadeMux I__659 (
            .O(N__3818),
            .I(N__3814));
    InMux I__658 (
            .O(N__3817),
            .I(N__3811));
    InMux I__657 (
            .O(N__3814),
            .I(N__3808));
    LocalMux I__656 (
            .O(N__3811),
            .I(\eeprom.delay_counter_15 ));
    LocalMux I__655 (
            .O(N__3808),
            .I(\eeprom.delay_counter_15 ));
    InMux I__654 (
            .O(N__3803),
            .I(N__3799));
    InMux I__653 (
            .O(N__3802),
            .I(N__3796));
    LocalMux I__652 (
            .O(N__3799),
            .I(\eeprom.delay_counter_9 ));
    LocalMux I__651 (
            .O(N__3796),
            .I(\eeprom.delay_counter_9 ));
    InMux I__650 (
            .O(N__3791),
            .I(N__3787));
    InMux I__649 (
            .O(N__3790),
            .I(N__3784));
    LocalMux I__648 (
            .O(N__3787),
            .I(\eeprom.delay_counter_1 ));
    LocalMux I__647 (
            .O(N__3784),
            .I(\eeprom.delay_counter_1 ));
    InMux I__646 (
            .O(N__3779),
            .I(N__3775));
    InMux I__645 (
            .O(N__3778),
            .I(N__3772));
    LocalMux I__644 (
            .O(N__3775),
            .I(\eeprom.delay_counter_7 ));
    LocalMux I__643 (
            .O(N__3772),
            .I(\eeprom.delay_counter_7 ));
    CascadeMux I__642 (
            .O(N__3767),
            .I(\eeprom.n2685_cascade_ ));
    InMux I__641 (
            .O(N__3764),
            .I(N__3760));
    InMux I__640 (
            .O(N__3763),
            .I(N__3757));
    LocalMux I__639 (
            .O(N__3760),
            .I(\eeprom.delay_counter_3 ));
    LocalMux I__638 (
            .O(N__3757),
            .I(\eeprom.delay_counter_3 ));
    InMux I__637 (
            .O(N__3752),
            .I(N__3749));
    LocalMux I__636 (
            .O(N__3749),
            .I(\eeprom.n22 ));
    InMux I__635 (
            .O(N__3746),
            .I(N__3742));
    InMux I__634 (
            .O(N__3745),
            .I(N__3739));
    LocalMux I__633 (
            .O(N__3742),
            .I(\eeprom.delay_counter_13 ));
    LocalMux I__632 (
            .O(N__3739),
            .I(\eeprom.delay_counter_13 ));
    CascadeMux I__631 (
            .O(N__3734),
            .I(N__3731));
    InMux I__630 (
            .O(N__3731),
            .I(N__3727));
    InMux I__629 (
            .O(N__3730),
            .I(N__3724));
    LocalMux I__628 (
            .O(N__3727),
            .I(\eeprom.delay_counter_8 ));
    LocalMux I__627 (
            .O(N__3724),
            .I(\eeprom.delay_counter_8 ));
    CascadeMux I__626 (
            .O(N__3719),
            .I(N__3716));
    InMux I__625 (
            .O(N__3716),
            .I(N__3712));
    InMux I__624 (
            .O(N__3715),
            .I(N__3709));
    LocalMux I__623 (
            .O(N__3712),
            .I(\eeprom.delay_counter_4 ));
    LocalMux I__622 (
            .O(N__3709),
            .I(\eeprom.delay_counter_4 ));
    InMux I__621 (
            .O(N__3704),
            .I(N__3701));
    LocalMux I__620 (
            .O(N__3701),
            .I(\eeprom.n20 ));
    CascadeMux I__619 (
            .O(N__3698),
            .I(\eeprom.i2c.n6_cascade_ ));
    CascadeMux I__618 (
            .O(N__3695),
            .I(\eeprom.i2c.counter2_7__N_256_cascade_ ));
    CEMux I__617 (
            .O(N__3692),
            .I(N__3689));
    LocalMux I__616 (
            .O(N__3689),
            .I(\eeprom.i2c.n1384 ));
    CascadeMux I__615 (
            .O(N__3686),
            .I(n6_adj_397_cascade_));
    CascadeMux I__614 (
            .O(N__3683),
            .I(n2662_cascade_));
    InMux I__613 (
            .O(N__3680),
            .I(N__3675));
    InMux I__612 (
            .O(N__3679),
            .I(N__3670));
    InMux I__611 (
            .O(N__3678),
            .I(N__3670));
    LocalMux I__610 (
            .O(N__3675),
            .I(n2668));
    LocalMux I__609 (
            .O(N__3670),
            .I(n2668));
    CascadeMux I__608 (
            .O(N__3665),
            .I(N__3662));
    InMux I__607 (
            .O(N__3662),
            .I(N__3658));
    InMux I__606 (
            .O(N__3661),
            .I(N__3655));
    LocalMux I__605 (
            .O(N__3658),
            .I(\eeprom.delay_counter_0 ));
    LocalMux I__604 (
            .O(N__3655),
            .I(\eeprom.delay_counter_0 ));
    CascadeMux I__603 (
            .O(N__3650),
            .I(N__3646));
    CascadeMux I__602 (
            .O(N__3649),
            .I(N__3643));
    InMux I__601 (
            .O(N__3646),
            .I(N__3640));
    InMux I__600 (
            .O(N__3643),
            .I(N__3637));
    LocalMux I__599 (
            .O(N__3640),
            .I(\eeprom.delay_counter_2 ));
    LocalMux I__598 (
            .O(N__3637),
            .I(\eeprom.delay_counter_2 ));
    InMux I__597 (
            .O(N__3632),
            .I(N__3628));
    InMux I__596 (
            .O(N__3631),
            .I(N__3625));
    LocalMux I__595 (
            .O(N__3628),
            .I(\eeprom.delay_counter_5 ));
    LocalMux I__594 (
            .O(N__3625),
            .I(\eeprom.delay_counter_5 ));
    CascadeMux I__593 (
            .O(N__3620),
            .I(N__3617));
    InMux I__592 (
            .O(N__3617),
            .I(N__3613));
    InMux I__591 (
            .O(N__3616),
            .I(N__3610));
    LocalMux I__590 (
            .O(N__3613),
            .I(\eeprom.delay_counter_10 ));
    LocalMux I__589 (
            .O(N__3610),
            .I(\eeprom.delay_counter_10 ));
    CascadeMux I__588 (
            .O(N__3605),
            .I(\eeprom.n24_cascade_ ));
    CascadeMux I__587 (
            .O(N__3602),
            .I(\eeprom.n1338_cascade_ ));
    CascadeMux I__586 (
            .O(N__3599),
            .I(N__3587));
    CascadeMux I__585 (
            .O(N__3598),
            .I(N__3583));
    CascadeMux I__584 (
            .O(N__3597),
            .I(N__3579));
    CascadeMux I__583 (
            .O(N__3596),
            .I(N__3575));
    CascadeMux I__582 (
            .O(N__3595),
            .I(N__3572));
    CascadeMux I__581 (
            .O(N__3594),
            .I(N__3569));
    CascadeMux I__580 (
            .O(N__3593),
            .I(N__3565));
    CascadeMux I__579 (
            .O(N__3592),
            .I(N__3561));
    InMux I__578 (
            .O(N__3591),
            .I(N__3543));
    InMux I__577 (
            .O(N__3590),
            .I(N__3543));
    InMux I__576 (
            .O(N__3587),
            .I(N__3543));
    InMux I__575 (
            .O(N__3586),
            .I(N__3543));
    InMux I__574 (
            .O(N__3583),
            .I(N__3543));
    InMux I__573 (
            .O(N__3582),
            .I(N__3543));
    InMux I__572 (
            .O(N__3579),
            .I(N__3543));
    InMux I__571 (
            .O(N__3578),
            .I(N__3543));
    InMux I__570 (
            .O(N__3575),
            .I(N__3540));
    InMux I__569 (
            .O(N__3572),
            .I(N__3525));
    InMux I__568 (
            .O(N__3569),
            .I(N__3525));
    InMux I__567 (
            .O(N__3568),
            .I(N__3525));
    InMux I__566 (
            .O(N__3565),
            .I(N__3525));
    InMux I__565 (
            .O(N__3564),
            .I(N__3525));
    InMux I__564 (
            .O(N__3561),
            .I(N__3525));
    InMux I__563 (
            .O(N__3560),
            .I(N__3525));
    LocalMux I__562 (
            .O(N__3543),
            .I(\eeprom.n575 ));
    LocalMux I__561 (
            .O(N__3540),
            .I(\eeprom.n575 ));
    LocalMux I__560 (
            .O(N__3525),
            .I(\eeprom.n575 ));
    CEMux I__559 (
            .O(N__3518),
            .I(N__3514));
    CEMux I__558 (
            .O(N__3517),
            .I(N__3511));
    LocalMux I__557 (
            .O(N__3514),
            .I(\eeprom.n1435 ));
    LocalMux I__556 (
            .O(N__3511),
            .I(\eeprom.n1435 ));
    CascadeMux I__555 (
            .O(N__3506),
            .I(\eeprom.n1435_cascade_ ));
    SRMux I__554 (
            .O(N__3503),
            .I(N__3499));
    SRMux I__553 (
            .O(N__3502),
            .I(N__3496));
    LocalMux I__552 (
            .O(N__3499),
            .I(N__3493));
    LocalMux I__551 (
            .O(N__3496),
            .I(\eeprom.n1503 ));
    Odrv4 I__550 (
            .O(N__3493),
            .I(\eeprom.n1503 ));
    InMux I__549 (
            .O(N__3488),
            .I(N__3484));
    InMux I__548 (
            .O(N__3487),
            .I(N__3481));
    LocalMux I__547 (
            .O(N__3484),
            .I(\eeprom.delay_counter_6 ));
    LocalMux I__546 (
            .O(N__3481),
            .I(\eeprom.delay_counter_6 ));
    CascadeMux I__545 (
            .O(N__3476),
            .I(N__3473));
    InMux I__544 (
            .O(N__3473),
            .I(N__3469));
    InMux I__543 (
            .O(N__3472),
            .I(N__3466));
    LocalMux I__542 (
            .O(N__3469),
            .I(\eeprom.delay_counter_12 ));
    LocalMux I__541 (
            .O(N__3466),
            .I(\eeprom.delay_counter_12 ));
    InMux I__540 (
            .O(N__3461),
            .I(N__3458));
    LocalMux I__539 (
            .O(N__3458),
            .I(\eeprom.n16 ));
    InMux I__538 (
            .O(N__3455),
            .I(bfn_17_20_0_));
    InMux I__537 (
            .O(N__3452),
            .I(\eeprom.n2524 ));
    InMux I__536 (
            .O(N__3449),
            .I(\eeprom.n2525 ));
    InMux I__535 (
            .O(N__3446),
            .I(\eeprom.n2526 ));
    InMux I__534 (
            .O(N__3443),
            .I(\eeprom.n2527 ));
    InMux I__533 (
            .O(N__3440),
            .I(\eeprom.n2528 ));
    InMux I__532 (
            .O(N__3437),
            .I(\eeprom.n2529 ));
    InMux I__531 (
            .O(N__3434),
            .I(\eeprom.n2530 ));
    InMux I__530 (
            .O(N__3431),
            .I(N__3428));
    LocalMux I__529 (
            .O(N__3428),
            .I(n2077));
    CascadeMux I__528 (
            .O(N__3425),
            .I(n12_cascade_));
    InMux I__527 (
            .O(N__3422),
            .I(\eeprom.n2516 ));
    InMux I__526 (
            .O(N__3419),
            .I(\eeprom.n2517 ));
    InMux I__525 (
            .O(N__3416),
            .I(\eeprom.n2518 ));
    InMux I__524 (
            .O(N__3413),
            .I(\eeprom.n2519 ));
    InMux I__523 (
            .O(N__3410),
            .I(\eeprom.n2520 ));
    InMux I__522 (
            .O(N__3407),
            .I(\eeprom.n2521 ));
    InMux I__521 (
            .O(N__3404),
            .I(\eeprom.n2522 ));
    InMux I__520 (
            .O(N__3401),
            .I(N__3397));
    InMux I__519 (
            .O(N__3400),
            .I(N__3394));
    LocalMux I__518 (
            .O(N__3397),
            .I(N__3389));
    LocalMux I__517 (
            .O(N__3394),
            .I(N__3389));
    Odrv4 I__516 (
            .O(N__3389),
            .I(delay_counter_18));
    InMux I__515 (
            .O(N__3386),
            .I(N__3382));
    InMux I__514 (
            .O(N__3385),
            .I(N__3379));
    LocalMux I__513 (
            .O(N__3382),
            .I(delay_counter_19));
    LocalMux I__512 (
            .O(N__3379),
            .I(delay_counter_19));
    CascadeMux I__511 (
            .O(N__3374),
            .I(n2721_cascade_));
    InMux I__510 (
            .O(N__3371),
            .I(N__3367));
    InMux I__509 (
            .O(N__3370),
            .I(N__3364));
    LocalMux I__508 (
            .O(N__3367),
            .I(delay_counter_22));
    LocalMux I__507 (
            .O(N__3364),
            .I(delay_counter_22));
    InMux I__506 (
            .O(N__3359),
            .I(N__3355));
    InMux I__505 (
            .O(N__3358),
            .I(N__3352));
    LocalMux I__504 (
            .O(N__3355),
            .I(delay_counter_21));
    LocalMux I__503 (
            .O(N__3352),
            .I(delay_counter_21));
    InMux I__502 (
            .O(N__3347),
            .I(N__3343));
    InMux I__501 (
            .O(N__3346),
            .I(N__3340));
    LocalMux I__500 (
            .O(N__3343),
            .I(delay_counter_23));
    LocalMux I__499 (
            .O(N__3340),
            .I(delay_counter_23));
    CascadeMux I__498 (
            .O(N__3335),
            .I(n7_cascade_));
    InMux I__497 (
            .O(N__3332),
            .I(N__3328));
    InMux I__496 (
            .O(N__3331),
            .I(N__3325));
    LocalMux I__495 (
            .O(N__3328),
            .I(N__3322));
    LocalMux I__494 (
            .O(N__3325),
            .I(delay_counter_20));
    Odrv4 I__493 (
            .O(N__3322),
            .I(delay_counter_20));
    InMux I__492 (
            .O(N__3317),
            .I(N__3313));
    InMux I__491 (
            .O(N__3316),
            .I(N__3310));
    LocalMux I__490 (
            .O(N__3313),
            .I(delay_counter_29));
    LocalMux I__489 (
            .O(N__3310),
            .I(delay_counter_29));
    InMux I__488 (
            .O(N__3305),
            .I(N__3301));
    InMux I__487 (
            .O(N__3304),
            .I(N__3298));
    LocalMux I__486 (
            .O(N__3301),
            .I(delay_counter_25));
    LocalMux I__485 (
            .O(N__3298),
            .I(delay_counter_25));
    CascadeMux I__484 (
            .O(N__3293),
            .I(n2695_cascade_));
    InMux I__483 (
            .O(N__3290),
            .I(N__3286));
    InMux I__482 (
            .O(N__3289),
            .I(N__3283));
    LocalMux I__481 (
            .O(N__3286),
            .I(delay_counter_28));
    LocalMux I__480 (
            .O(N__3283),
            .I(delay_counter_28));
    CascadeMux I__479 (
            .O(N__3278),
            .I(n13_cascade_));
    SRMux I__478 (
            .O(N__3275),
            .I(N__3272));
    LocalMux I__477 (
            .O(N__3272),
            .I(N__3269));
    Span4Mux_h I__476 (
            .O(N__3269),
            .I(N__3263));
    SRMux I__475 (
            .O(N__3268),
            .I(N__3260));
    SRMux I__474 (
            .O(N__3267),
            .I(N__3257));
    SRMux I__473 (
            .O(N__3266),
            .I(N__3254));
    Odrv4 I__472 (
            .O(N__3263),
            .I(addr_10__N_70));
    LocalMux I__471 (
            .O(N__3260),
            .I(addr_10__N_70));
    LocalMux I__470 (
            .O(N__3257),
            .I(addr_10__N_70));
    LocalMux I__469 (
            .O(N__3254),
            .I(addr_10__N_70));
    InMux I__468 (
            .O(N__3245),
            .I(N__3240));
    InMux I__467 (
            .O(N__3244),
            .I(N__3237));
    InMux I__466 (
            .O(N__3243),
            .I(N__3234));
    LocalMux I__465 (
            .O(N__3240),
            .I(delay_counter_31));
    LocalMux I__464 (
            .O(N__3237),
            .I(delay_counter_31));
    LocalMux I__463 (
            .O(N__3234),
            .I(delay_counter_31));
    InMux I__462 (
            .O(N__3227),
            .I(N__3224));
    LocalMux I__461 (
            .O(N__3224),
            .I(n13));
    InMux I__460 (
            .O(N__3221),
            .I(N__3217));
    InMux I__459 (
            .O(N__3220),
            .I(N__3214));
    LocalMux I__458 (
            .O(N__3217),
            .I(delay_counter_26));
    LocalMux I__457 (
            .O(N__3214),
            .I(delay_counter_26));
    InMux I__456 (
            .O(N__3209),
            .I(N__3205));
    InMux I__455 (
            .O(N__3208),
            .I(N__3202));
    LocalMux I__454 (
            .O(N__3205),
            .I(delay_counter_30));
    LocalMux I__453 (
            .O(N__3202),
            .I(delay_counter_30));
    CascadeMux I__452 (
            .O(N__3197),
            .I(N__3193));
    InMux I__451 (
            .O(N__3196),
            .I(N__3190));
    InMux I__450 (
            .O(N__3193),
            .I(N__3187));
    LocalMux I__449 (
            .O(N__3190),
            .I(delay_counter_27));
    LocalMux I__448 (
            .O(N__3187),
            .I(delay_counter_27));
    InMux I__447 (
            .O(N__3182),
            .I(N__3178));
    InMux I__446 (
            .O(N__3181),
            .I(N__3175));
    LocalMux I__445 (
            .O(N__3178),
            .I(delay_counter_24));
    LocalMux I__444 (
            .O(N__3175),
            .I(delay_counter_24));
    InMux I__443 (
            .O(N__3170),
            .I(N__3164));
    InMux I__442 (
            .O(N__3169),
            .I(N__3164));
    LocalMux I__441 (
            .O(N__3164),
            .I(n14));
    CascadeMux I__440 (
            .O(N__3161),
            .I(n2077_cascade_));
    InMux I__439 (
            .O(N__3158),
            .I(n2508));
    InMux I__438 (
            .O(N__3155),
            .I(N__3151));
    InMux I__437 (
            .O(N__3154),
            .I(N__3148));
    LocalMux I__436 (
            .O(N__3151),
            .I(delay_counter_6));
    LocalMux I__435 (
            .O(N__3148),
            .I(delay_counter_6));
    InMux I__434 (
            .O(N__3143),
            .I(N__3139));
    InMux I__433 (
            .O(N__3142),
            .I(N__3136));
    LocalMux I__432 (
            .O(N__3139),
            .I(delay_counter_0));
    LocalMux I__431 (
            .O(N__3136),
            .I(delay_counter_0));
    CascadeMux I__430 (
            .O(N__3131),
            .I(N__3127));
    InMux I__429 (
            .O(N__3130),
            .I(N__3124));
    InMux I__428 (
            .O(N__3127),
            .I(N__3121));
    LocalMux I__427 (
            .O(N__3124),
            .I(delay_counter_9));
    LocalMux I__426 (
            .O(N__3121),
            .I(delay_counter_9));
    InMux I__425 (
            .O(N__3116),
            .I(N__3112));
    InMux I__424 (
            .O(N__3115),
            .I(N__3109));
    LocalMux I__423 (
            .O(N__3112),
            .I(delay_counter_4));
    LocalMux I__422 (
            .O(N__3109),
            .I(delay_counter_4));
    InMux I__421 (
            .O(N__3104),
            .I(N__3100));
    InMux I__420 (
            .O(N__3103),
            .I(N__3097));
    LocalMux I__419 (
            .O(N__3100),
            .I(delay_counter_2));
    LocalMux I__418 (
            .O(N__3097),
            .I(delay_counter_2));
    InMux I__417 (
            .O(N__3092),
            .I(N__3088));
    InMux I__416 (
            .O(N__3091),
            .I(N__3085));
    LocalMux I__415 (
            .O(N__3088),
            .I(delay_counter_7));
    LocalMux I__414 (
            .O(N__3085),
            .I(delay_counter_7));
    CascadeMux I__413 (
            .O(N__3080),
            .I(N__3076));
    InMux I__412 (
            .O(N__3079),
            .I(N__3073));
    InMux I__411 (
            .O(N__3076),
            .I(N__3070));
    LocalMux I__410 (
            .O(N__3073),
            .I(delay_counter_5));
    LocalMux I__409 (
            .O(N__3070),
            .I(delay_counter_5));
    InMux I__408 (
            .O(N__3065),
            .I(N__3061));
    InMux I__407 (
            .O(N__3064),
            .I(N__3058));
    LocalMux I__406 (
            .O(N__3061),
            .I(delay_counter_3));
    LocalMux I__405 (
            .O(N__3058),
            .I(delay_counter_3));
    InMux I__404 (
            .O(N__3053),
            .I(N__3049));
    InMux I__403 (
            .O(N__3052),
            .I(N__3046));
    LocalMux I__402 (
            .O(N__3049),
            .I(delay_counter_8));
    LocalMux I__401 (
            .O(N__3046),
            .I(delay_counter_8));
    InMux I__400 (
            .O(N__3041),
            .I(N__3037));
    InMux I__399 (
            .O(N__3040),
            .I(N__3034));
    LocalMux I__398 (
            .O(N__3037),
            .I(delay_counter_1));
    LocalMux I__397 (
            .O(N__3034),
            .I(delay_counter_1));
    CascadeMux I__396 (
            .O(N__3029),
            .I(N__3026));
    InMux I__395 (
            .O(N__3026),
            .I(N__3023));
    LocalMux I__394 (
            .O(N__3023),
            .I(N__3020));
    Odrv4 I__393 (
            .O(N__3020),
            .I(n17));
    InMux I__392 (
            .O(N__3017),
            .I(N__3014));
    LocalMux I__391 (
            .O(N__3014),
            .I(n16));
    InMux I__390 (
            .O(N__3011),
            .I(N__3007));
    InMux I__389 (
            .O(N__3010),
            .I(N__3004));
    LocalMux I__388 (
            .O(N__3007),
            .I(delay_counter_11));
    LocalMux I__387 (
            .O(N__3004),
            .I(delay_counter_11));
    InMux I__386 (
            .O(N__2999),
            .I(N__2995));
    InMux I__385 (
            .O(N__2998),
            .I(N__2992));
    LocalMux I__384 (
            .O(N__2995),
            .I(delay_counter_10));
    LocalMux I__383 (
            .O(N__2992),
            .I(delay_counter_10));
    CascadeMux I__382 (
            .O(N__2987),
            .I(n2722_cascade_));
    InMux I__381 (
            .O(N__2984),
            .I(N__2980));
    InMux I__380 (
            .O(N__2983),
            .I(N__2977));
    LocalMux I__379 (
            .O(N__2980),
            .I(delay_counter_12));
    LocalMux I__378 (
            .O(N__2977),
            .I(delay_counter_12));
    InMux I__377 (
            .O(N__2972),
            .I(N__2968));
    InMux I__376 (
            .O(N__2971),
            .I(N__2965));
    LocalMux I__375 (
            .O(N__2968),
            .I(N__2962));
    LocalMux I__374 (
            .O(N__2965),
            .I(delay_counter_17));
    Odrv4 I__373 (
            .O(N__2962),
            .I(delay_counter_17));
    InMux I__372 (
            .O(N__2957),
            .I(N__2953));
    InMux I__371 (
            .O(N__2956),
            .I(N__2950));
    LocalMux I__370 (
            .O(N__2953),
            .I(delay_counter_15));
    LocalMux I__369 (
            .O(N__2950),
            .I(delay_counter_15));
    InMux I__368 (
            .O(N__2945),
            .I(N__2941));
    InMux I__367 (
            .O(N__2944),
            .I(N__2938));
    LocalMux I__366 (
            .O(N__2941),
            .I(delay_counter_14));
    LocalMux I__365 (
            .O(N__2938),
            .I(delay_counter_14));
    InMux I__364 (
            .O(N__2933),
            .I(N__2930));
    LocalMux I__363 (
            .O(N__2930),
            .I(n8));
    InMux I__362 (
            .O(N__2927),
            .I(N__2923));
    InMux I__361 (
            .O(N__2926),
            .I(N__2920));
    LocalMux I__360 (
            .O(N__2923),
            .I(delay_counter_16));
    LocalMux I__359 (
            .O(N__2920),
            .I(delay_counter_16));
    CascadeMux I__358 (
            .O(N__2915),
            .I(N__2911));
    InMux I__357 (
            .O(N__2914),
            .I(N__2908));
    InMux I__356 (
            .O(N__2911),
            .I(N__2905));
    LocalMux I__355 (
            .O(N__2908),
            .I(delay_counter_13));
    LocalMux I__354 (
            .O(N__2905),
            .I(delay_counter_13));
    InMux I__353 (
            .O(N__2900),
            .I(N__2897));
    LocalMux I__352 (
            .O(N__2897),
            .I(n2715));
    InMux I__351 (
            .O(N__2894),
            .I(n2499));
    InMux I__350 (
            .O(N__2891),
            .I(n2500));
    InMux I__349 (
            .O(N__2888),
            .I(bfn_14_24_0_));
    InMux I__348 (
            .O(N__2885),
            .I(n2502));
    InMux I__347 (
            .O(N__2882),
            .I(n2503));
    InMux I__346 (
            .O(N__2879),
            .I(n2504));
    InMux I__345 (
            .O(N__2876),
            .I(n2505));
    InMux I__344 (
            .O(N__2873),
            .I(n2506));
    InMux I__343 (
            .O(N__2870),
            .I(n2507));
    InMux I__342 (
            .O(N__2867),
            .I(n2490));
    InMux I__341 (
            .O(N__2864),
            .I(n2491));
    InMux I__340 (
            .O(N__2861),
            .I(n2492));
    InMux I__339 (
            .O(N__2858),
            .I(bfn_14_23_0_));
    InMux I__338 (
            .O(N__2855),
            .I(n2494));
    InMux I__337 (
            .O(N__2852),
            .I(n2495));
    InMux I__336 (
            .O(N__2849),
            .I(n2496));
    InMux I__335 (
            .O(N__2846),
            .I(n2497));
    InMux I__334 (
            .O(N__2843),
            .I(n2498));
    InMux I__333 (
            .O(N__2840),
            .I(n2480));
    InMux I__332 (
            .O(N__2837),
            .I(n2481));
    InMux I__331 (
            .O(N__2834),
            .I(n2482));
    InMux I__330 (
            .O(N__2831),
            .I(n2483));
    InMux I__329 (
            .O(N__2828),
            .I(n2484));
    InMux I__328 (
            .O(N__2825),
            .I(bfn_14_22_0_));
    InMux I__327 (
            .O(N__2822),
            .I(n2486));
    InMux I__326 (
            .O(N__2819),
            .I(n2487));
    InMux I__325 (
            .O(N__2816),
            .I(n2488));
    InMux I__324 (
            .O(N__2813),
            .I(n2489));
    InMux I__323 (
            .O(N__2810),
            .I(bfn_13_24_0_));
    InMux I__322 (
            .O(N__2807),
            .I(n2559));
    InMux I__321 (
            .O(N__2804),
            .I(N__2797));
    InMux I__320 (
            .O(N__2803),
            .I(N__2797));
    InMux I__319 (
            .O(N__2802),
            .I(N__2794));
    LocalMux I__318 (
            .O(N__2797),
            .I(blink_counter_21));
    LocalMux I__317 (
            .O(N__2794),
            .I(blink_counter_21));
    InMux I__316 (
            .O(N__2789),
            .I(N__2780));
    InMux I__315 (
            .O(N__2788),
            .I(N__2780));
    InMux I__314 (
            .O(N__2787),
            .I(N__2780));
    LocalMux I__313 (
            .O(N__2780),
            .I(blink_counter_24));
    CascadeMux I__312 (
            .O(N__2777),
            .I(N__2773));
    CascadeMux I__311 (
            .O(N__2776),
            .I(N__2770));
    InMux I__310 (
            .O(N__2773),
            .I(N__2764));
    InMux I__309 (
            .O(N__2770),
            .I(N__2764));
    InMux I__308 (
            .O(N__2769),
            .I(N__2761));
    LocalMux I__307 (
            .O(N__2764),
            .I(blink_counter_23));
    LocalMux I__306 (
            .O(N__2761),
            .I(blink_counter_23));
    InMux I__305 (
            .O(N__2756),
            .I(N__2749));
    InMux I__304 (
            .O(N__2755),
            .I(N__2749));
    InMux I__303 (
            .O(N__2754),
            .I(N__2746));
    LocalMux I__302 (
            .O(N__2749),
            .I(blink_counter_22));
    LocalMux I__301 (
            .O(N__2746),
            .I(blink_counter_22));
    InMux I__300 (
            .O(N__2741),
            .I(N__2738));
    LocalMux I__299 (
            .O(N__2738),
            .I(n2730));
    CascadeMux I__298 (
            .O(N__2735),
            .I(n2731_cascade_));
    InMux I__297 (
            .O(N__2732),
            .I(N__2726));
    InMux I__296 (
            .O(N__2731),
            .I(N__2726));
    LocalMux I__295 (
            .O(N__2726),
            .I(blink_counter_25));
    IoInMux I__294 (
            .O(N__2723),
            .I(N__2720));
    LocalMux I__293 (
            .O(N__2720),
            .I(N__2717));
    Span4Mux_s3_v I__292 (
            .O(N__2717),
            .I(N__2714));
    Sp12to4 I__291 (
            .O(N__2714),
            .I(N__2711));
    Span12Mux_h I__290 (
            .O(N__2711),
            .I(N__2708));
    Odrv12 I__289 (
            .O(N__2708),
            .I(LED_c));
    InMux I__288 (
            .O(N__2705),
            .I(bfn_14_21_0_));
    InMux I__287 (
            .O(N__2702),
            .I(n2478));
    InMux I__286 (
            .O(N__2699),
            .I(n2479));
    InMux I__285 (
            .O(N__2696),
            .I(N__2693));
    LocalMux I__284 (
            .O(N__2693),
            .I(n11));
    InMux I__283 (
            .O(N__2690),
            .I(n2549));
    InMux I__282 (
            .O(N__2687),
            .I(N__2684));
    LocalMux I__281 (
            .O(N__2684),
            .I(n10));
    InMux I__280 (
            .O(N__2681),
            .I(bfn_13_23_0_));
    InMux I__279 (
            .O(N__2678),
            .I(N__2675));
    LocalMux I__278 (
            .O(N__2675),
            .I(n9));
    InMux I__277 (
            .O(N__2672),
            .I(n2551));
    InMux I__276 (
            .O(N__2669),
            .I(N__2666));
    LocalMux I__275 (
            .O(N__2666),
            .I(n8_adj_388));
    InMux I__274 (
            .O(N__2663),
            .I(n2552));
    InMux I__273 (
            .O(N__2660),
            .I(N__2657));
    LocalMux I__272 (
            .O(N__2657),
            .I(n7_adj_387));
    InMux I__271 (
            .O(N__2654),
            .I(n2553));
    InMux I__270 (
            .O(N__2651),
            .I(N__2648));
    LocalMux I__269 (
            .O(N__2648),
            .I(n6));
    InMux I__268 (
            .O(N__2645),
            .I(n2554));
    InMux I__267 (
            .O(N__2642),
            .I(n2555));
    InMux I__266 (
            .O(N__2639),
            .I(n2556));
    InMux I__265 (
            .O(N__2636),
            .I(n2557));
    InMux I__264 (
            .O(N__2633),
            .I(N__2630));
    LocalMux I__263 (
            .O(N__2630),
            .I(n19));
    InMux I__262 (
            .O(N__2627),
            .I(n2541));
    InMux I__261 (
            .O(N__2624),
            .I(N__2621));
    LocalMux I__260 (
            .O(N__2621),
            .I(n18));
    InMux I__259 (
            .O(N__2618),
            .I(bfn_13_22_0_));
    InMux I__258 (
            .O(N__2615),
            .I(N__2612));
    LocalMux I__257 (
            .O(N__2612),
            .I(n17_adj_394));
    InMux I__256 (
            .O(N__2609),
            .I(n2543));
    InMux I__255 (
            .O(N__2606),
            .I(N__2603));
    LocalMux I__254 (
            .O(N__2603),
            .I(n16_adj_393));
    InMux I__253 (
            .O(N__2600),
            .I(n2544));
    InMux I__252 (
            .O(N__2597),
            .I(N__2594));
    LocalMux I__251 (
            .O(N__2594),
            .I(n15_adj_392));
    InMux I__250 (
            .O(N__2591),
            .I(n2545));
    InMux I__249 (
            .O(N__2588),
            .I(N__2585));
    LocalMux I__248 (
            .O(N__2585),
            .I(n14_adj_391));
    InMux I__247 (
            .O(N__2582),
            .I(n2546));
    InMux I__246 (
            .O(N__2579),
            .I(N__2576));
    LocalMux I__245 (
            .O(N__2576),
            .I(n13_adj_390));
    InMux I__244 (
            .O(N__2573),
            .I(n2547));
    InMux I__243 (
            .O(N__2570),
            .I(N__2567));
    LocalMux I__242 (
            .O(N__2567),
            .I(n12_adj_389));
    InMux I__241 (
            .O(N__2564),
            .I(n2548));
    InMux I__240 (
            .O(N__2561),
            .I(N__2558));
    LocalMux I__239 (
            .O(N__2558),
            .I(n26));
    InMux I__238 (
            .O(N__2555),
            .I(bfn_13_21_0_));
    InMux I__237 (
            .O(N__2552),
            .I(N__2549));
    LocalMux I__236 (
            .O(N__2549),
            .I(n25));
    InMux I__235 (
            .O(N__2546),
            .I(n2535));
    InMux I__234 (
            .O(N__2543),
            .I(N__2540));
    LocalMux I__233 (
            .O(N__2540),
            .I(n24));
    InMux I__232 (
            .O(N__2537),
            .I(n2536));
    InMux I__231 (
            .O(N__2534),
            .I(N__2531));
    LocalMux I__230 (
            .O(N__2531),
            .I(n23));
    InMux I__229 (
            .O(N__2528),
            .I(n2537));
    InMux I__228 (
            .O(N__2525),
            .I(N__2522));
    LocalMux I__227 (
            .O(N__2522),
            .I(n22));
    InMux I__226 (
            .O(N__2519),
            .I(n2538));
    InMux I__225 (
            .O(N__2516),
            .I(N__2513));
    LocalMux I__224 (
            .O(N__2513),
            .I(n21));
    InMux I__223 (
            .O(N__2510),
            .I(n2539));
    InMux I__222 (
            .O(N__2507),
            .I(N__2504));
    LocalMux I__221 (
            .O(N__2504),
            .I(n20));
    InMux I__220 (
            .O(N__2501),
            .I(n2540));
    IoInMux I__219 (
            .O(N__2498),
            .I(N__2495));
    LocalMux I__218 (
            .O(N__2495),
            .I(N__2492));
    IoSpan4Mux I__217 (
            .O(N__2492),
            .I(N__2489));
    IoSpan4Mux I__216 (
            .O(N__2489),
            .I(N__2486));
    IoSpan4Mux I__215 (
            .O(N__2486),
            .I(N__2483));
    Odrv4 I__214 (
            .O(N__2483),
            .I(CLK_pad_gb_input));
    INV \INVeeprom.i2c.i2c_scl_enable_124C  (
            .O(\INVeeprom.i2c.i2c_scl_enable_124C_net ),
            .I(N__4974));
    INV \INVeeprom.i2c.write_enable_132C  (
            .O(\INVeeprom.i2c.write_enable_132C_net ),
            .I(N__4946));
    INV \INVeeprom.i2c.sda_out_133C  (
            .O(\INVeeprom.i2c.sda_out_133C_net ),
            .I(N__4975));
    defparam IN_MUX_bfv_21_14_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_21_14_0_ (
            .carryinitin(),
            .carryinitout(bfn_21_14_0_));
    defparam IN_MUX_bfv_19_17_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_19_17_0_ (
            .carryinitin(),
            .carryinitout(bfn_19_17_0_));
    defparam IN_MUX_bfv_17_19_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_19_0_ (
            .carryinitin(),
            .carryinitout(bfn_17_19_0_));
    defparam IN_MUX_bfv_17_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_20_0_ (
            .carryinitin(\eeprom.n2523 ),
            .carryinitout(bfn_17_20_0_));
    defparam IN_MUX_bfv_14_21_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_21_0_ (
            .carryinitin(),
            .carryinitout(bfn_14_21_0_));
    defparam IN_MUX_bfv_14_22_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_22_0_ (
            .carryinitin(n2485),
            .carryinitout(bfn_14_22_0_));
    defparam IN_MUX_bfv_14_23_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_23_0_ (
            .carryinitin(n2493),
            .carryinitout(bfn_14_23_0_));
    defparam IN_MUX_bfv_14_24_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_24_0_ (
            .carryinitin(n2501),
            .carryinitout(bfn_14_24_0_));
    defparam IN_MUX_bfv_13_21_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_21_0_ (
            .carryinitin(),
            .carryinitout(bfn_13_21_0_));
    defparam IN_MUX_bfv_13_22_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_22_0_ (
            .carryinitin(n2542),
            .carryinitout(bfn_13_22_0_));
    defparam IN_MUX_bfv_13_23_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_23_0_ (
            .carryinitin(n2550),
            .carryinitout(bfn_13_23_0_));
    defparam IN_MUX_bfv_13_24_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_24_0_ (
            .carryinitin(n2558),
            .carryinitout(bfn_13_24_0_));
    ICE_GB CLK_pad_gb (
            .USERSIGNALTOGLOBALBUFFER(N__2498),
            .GLOBALBUFFEROUTPUT(CLK_c));
    VCC VCC (
            .Y(VCCG0));
    GND GND (
            .Y(GNDG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam blink_counter_332__i0_LC_13_21_0.C_ON=1'b1;
    defparam blink_counter_332__i0_LC_13_21_0.SEQ_MODE=4'b1000;
    defparam blink_counter_332__i0_LC_13_21_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_332__i0_LC_13_21_0 (
            .in0(_gnd_net_),
            .in1(N__2561),
            .in2(_gnd_net_),
            .in3(N__2555),
            .lcout(n26),
            .ltout(),
            .carryin(bfn_13_21_0_),
            .carryout(n2535),
            .clk(N__3925),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_332__i1_LC_13_21_1.C_ON=1'b1;
    defparam blink_counter_332__i1_LC_13_21_1.SEQ_MODE=4'b1000;
    defparam blink_counter_332__i1_LC_13_21_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_332__i1_LC_13_21_1 (
            .in0(_gnd_net_),
            .in1(N__2552),
            .in2(_gnd_net_),
            .in3(N__2546),
            .lcout(n25),
            .ltout(),
            .carryin(n2535),
            .carryout(n2536),
            .clk(N__3925),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_332__i2_LC_13_21_2.C_ON=1'b1;
    defparam blink_counter_332__i2_LC_13_21_2.SEQ_MODE=4'b1000;
    defparam blink_counter_332__i2_LC_13_21_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_332__i2_LC_13_21_2 (
            .in0(_gnd_net_),
            .in1(N__2543),
            .in2(_gnd_net_),
            .in3(N__2537),
            .lcout(n24),
            .ltout(),
            .carryin(n2536),
            .carryout(n2537),
            .clk(N__3925),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_332__i3_LC_13_21_3.C_ON=1'b1;
    defparam blink_counter_332__i3_LC_13_21_3.SEQ_MODE=4'b1000;
    defparam blink_counter_332__i3_LC_13_21_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_332__i3_LC_13_21_3 (
            .in0(_gnd_net_),
            .in1(N__2534),
            .in2(_gnd_net_),
            .in3(N__2528),
            .lcout(n23),
            .ltout(),
            .carryin(n2537),
            .carryout(n2538),
            .clk(N__3925),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_332__i4_LC_13_21_4.C_ON=1'b1;
    defparam blink_counter_332__i4_LC_13_21_4.SEQ_MODE=4'b1000;
    defparam blink_counter_332__i4_LC_13_21_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_332__i4_LC_13_21_4 (
            .in0(_gnd_net_),
            .in1(N__2525),
            .in2(_gnd_net_),
            .in3(N__2519),
            .lcout(n22),
            .ltout(),
            .carryin(n2538),
            .carryout(n2539),
            .clk(N__3925),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_332__i5_LC_13_21_5.C_ON=1'b1;
    defparam blink_counter_332__i5_LC_13_21_5.SEQ_MODE=4'b1000;
    defparam blink_counter_332__i5_LC_13_21_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_332__i5_LC_13_21_5 (
            .in0(_gnd_net_),
            .in1(N__2516),
            .in2(_gnd_net_),
            .in3(N__2510),
            .lcout(n21),
            .ltout(),
            .carryin(n2539),
            .carryout(n2540),
            .clk(N__3925),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_332__i6_LC_13_21_6.C_ON=1'b1;
    defparam blink_counter_332__i6_LC_13_21_6.SEQ_MODE=4'b1000;
    defparam blink_counter_332__i6_LC_13_21_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_332__i6_LC_13_21_6 (
            .in0(_gnd_net_),
            .in1(N__2507),
            .in2(_gnd_net_),
            .in3(N__2501),
            .lcout(n20),
            .ltout(),
            .carryin(n2540),
            .carryout(n2541),
            .clk(N__3925),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_332__i7_LC_13_21_7.C_ON=1'b1;
    defparam blink_counter_332__i7_LC_13_21_7.SEQ_MODE=4'b1000;
    defparam blink_counter_332__i7_LC_13_21_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_332__i7_LC_13_21_7 (
            .in0(_gnd_net_),
            .in1(N__2633),
            .in2(_gnd_net_),
            .in3(N__2627),
            .lcout(n19),
            .ltout(),
            .carryin(n2541),
            .carryout(n2542),
            .clk(N__3925),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_332__i8_LC_13_22_0.C_ON=1'b1;
    defparam blink_counter_332__i8_LC_13_22_0.SEQ_MODE=4'b1000;
    defparam blink_counter_332__i8_LC_13_22_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_332__i8_LC_13_22_0 (
            .in0(_gnd_net_),
            .in1(N__2624),
            .in2(_gnd_net_),
            .in3(N__2618),
            .lcout(n18),
            .ltout(),
            .carryin(bfn_13_22_0_),
            .carryout(n2543),
            .clk(N__3926),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_332__i9_LC_13_22_1.C_ON=1'b1;
    defparam blink_counter_332__i9_LC_13_22_1.SEQ_MODE=4'b1000;
    defparam blink_counter_332__i9_LC_13_22_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_332__i9_LC_13_22_1 (
            .in0(_gnd_net_),
            .in1(N__2615),
            .in2(_gnd_net_),
            .in3(N__2609),
            .lcout(n17_adj_394),
            .ltout(),
            .carryin(n2543),
            .carryout(n2544),
            .clk(N__3926),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_332__i10_LC_13_22_2.C_ON=1'b1;
    defparam blink_counter_332__i10_LC_13_22_2.SEQ_MODE=4'b1000;
    defparam blink_counter_332__i10_LC_13_22_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_332__i10_LC_13_22_2 (
            .in0(_gnd_net_),
            .in1(N__2606),
            .in2(_gnd_net_),
            .in3(N__2600),
            .lcout(n16_adj_393),
            .ltout(),
            .carryin(n2544),
            .carryout(n2545),
            .clk(N__3926),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_332__i11_LC_13_22_3.C_ON=1'b1;
    defparam blink_counter_332__i11_LC_13_22_3.SEQ_MODE=4'b1000;
    defparam blink_counter_332__i11_LC_13_22_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_332__i11_LC_13_22_3 (
            .in0(_gnd_net_),
            .in1(N__2597),
            .in2(_gnd_net_),
            .in3(N__2591),
            .lcout(n15_adj_392),
            .ltout(),
            .carryin(n2545),
            .carryout(n2546),
            .clk(N__3926),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_332__i12_LC_13_22_4.C_ON=1'b1;
    defparam blink_counter_332__i12_LC_13_22_4.SEQ_MODE=4'b1000;
    defparam blink_counter_332__i12_LC_13_22_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_332__i12_LC_13_22_4 (
            .in0(_gnd_net_),
            .in1(N__2588),
            .in2(_gnd_net_),
            .in3(N__2582),
            .lcout(n14_adj_391),
            .ltout(),
            .carryin(n2546),
            .carryout(n2547),
            .clk(N__3926),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_332__i13_LC_13_22_5.C_ON=1'b1;
    defparam blink_counter_332__i13_LC_13_22_5.SEQ_MODE=4'b1000;
    defparam blink_counter_332__i13_LC_13_22_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_332__i13_LC_13_22_5 (
            .in0(_gnd_net_),
            .in1(N__2579),
            .in2(_gnd_net_),
            .in3(N__2573),
            .lcout(n13_adj_390),
            .ltout(),
            .carryin(n2547),
            .carryout(n2548),
            .clk(N__3926),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_332__i14_LC_13_22_6.C_ON=1'b1;
    defparam blink_counter_332__i14_LC_13_22_6.SEQ_MODE=4'b1000;
    defparam blink_counter_332__i14_LC_13_22_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_332__i14_LC_13_22_6 (
            .in0(_gnd_net_),
            .in1(N__2570),
            .in2(_gnd_net_),
            .in3(N__2564),
            .lcout(n12_adj_389),
            .ltout(),
            .carryin(n2548),
            .carryout(n2549),
            .clk(N__3926),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_332__i15_LC_13_22_7.C_ON=1'b1;
    defparam blink_counter_332__i15_LC_13_22_7.SEQ_MODE=4'b1000;
    defparam blink_counter_332__i15_LC_13_22_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_332__i15_LC_13_22_7 (
            .in0(_gnd_net_),
            .in1(N__2696),
            .in2(_gnd_net_),
            .in3(N__2690),
            .lcout(n11),
            .ltout(),
            .carryin(n2549),
            .carryout(n2550),
            .clk(N__3926),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_332__i16_LC_13_23_0.C_ON=1'b1;
    defparam blink_counter_332__i16_LC_13_23_0.SEQ_MODE=4'b1000;
    defparam blink_counter_332__i16_LC_13_23_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_332__i16_LC_13_23_0 (
            .in0(_gnd_net_),
            .in1(N__2687),
            .in2(_gnd_net_),
            .in3(N__2681),
            .lcout(n10),
            .ltout(),
            .carryin(bfn_13_23_0_),
            .carryout(n2551),
            .clk(N__3930),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_332__i17_LC_13_23_1.C_ON=1'b1;
    defparam blink_counter_332__i17_LC_13_23_1.SEQ_MODE=4'b1000;
    defparam blink_counter_332__i17_LC_13_23_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_332__i17_LC_13_23_1 (
            .in0(_gnd_net_),
            .in1(N__2678),
            .in2(_gnd_net_),
            .in3(N__2672),
            .lcout(n9),
            .ltout(),
            .carryin(n2551),
            .carryout(n2552),
            .clk(N__3930),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_332__i18_LC_13_23_2.C_ON=1'b1;
    defparam blink_counter_332__i18_LC_13_23_2.SEQ_MODE=4'b1000;
    defparam blink_counter_332__i18_LC_13_23_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_332__i18_LC_13_23_2 (
            .in0(_gnd_net_),
            .in1(N__2669),
            .in2(_gnd_net_),
            .in3(N__2663),
            .lcout(n8_adj_388),
            .ltout(),
            .carryin(n2552),
            .carryout(n2553),
            .clk(N__3930),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_332__i19_LC_13_23_3.C_ON=1'b1;
    defparam blink_counter_332__i19_LC_13_23_3.SEQ_MODE=4'b1000;
    defparam blink_counter_332__i19_LC_13_23_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_332__i19_LC_13_23_3 (
            .in0(_gnd_net_),
            .in1(N__2660),
            .in2(_gnd_net_),
            .in3(N__2654),
            .lcout(n7_adj_387),
            .ltout(),
            .carryin(n2553),
            .carryout(n2554),
            .clk(N__3930),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_332__i20_LC_13_23_4.C_ON=1'b1;
    defparam blink_counter_332__i20_LC_13_23_4.SEQ_MODE=4'b1000;
    defparam blink_counter_332__i20_LC_13_23_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_332__i20_LC_13_23_4 (
            .in0(_gnd_net_),
            .in1(N__2651),
            .in2(_gnd_net_),
            .in3(N__2645),
            .lcout(n6),
            .ltout(),
            .carryin(n2554),
            .carryout(n2555),
            .clk(N__3930),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_332__i21_LC_13_23_5.C_ON=1'b1;
    defparam blink_counter_332__i21_LC_13_23_5.SEQ_MODE=4'b1000;
    defparam blink_counter_332__i21_LC_13_23_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_332__i21_LC_13_23_5 (
            .in0(_gnd_net_),
            .in1(N__2802),
            .in2(_gnd_net_),
            .in3(N__2642),
            .lcout(blink_counter_21),
            .ltout(),
            .carryin(n2555),
            .carryout(n2556),
            .clk(N__3930),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_332__i22_LC_13_23_6.C_ON=1'b1;
    defparam blink_counter_332__i22_LC_13_23_6.SEQ_MODE=4'b1000;
    defparam blink_counter_332__i22_LC_13_23_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_332__i22_LC_13_23_6 (
            .in0(_gnd_net_),
            .in1(N__2754),
            .in2(_gnd_net_),
            .in3(N__2639),
            .lcout(blink_counter_22),
            .ltout(),
            .carryin(n2556),
            .carryout(n2557),
            .clk(N__3930),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_332__i23_LC_13_23_7.C_ON=1'b1;
    defparam blink_counter_332__i23_LC_13_23_7.SEQ_MODE=4'b1000;
    defparam blink_counter_332__i23_LC_13_23_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_332__i23_LC_13_23_7 (
            .in0(_gnd_net_),
            .in1(N__2769),
            .in2(_gnd_net_),
            .in3(N__2636),
            .lcout(blink_counter_23),
            .ltout(),
            .carryin(n2557),
            .carryout(n2558),
            .clk(N__3930),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_332__i24_LC_13_24_0.C_ON=1'b1;
    defparam blink_counter_332__i24_LC_13_24_0.SEQ_MODE=4'b1000;
    defparam blink_counter_332__i24_LC_13_24_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_332__i24_LC_13_24_0 (
            .in0(_gnd_net_),
            .in1(N__2787),
            .in2(_gnd_net_),
            .in3(N__2810),
            .lcout(blink_counter_24),
            .ltout(),
            .carryin(bfn_13_24_0_),
            .carryout(n2559),
            .clk(N__3933),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_332__i25_LC_13_24_1.C_ON=1'b0;
    defparam blink_counter_332__i25_LC_13_24_1.SEQ_MODE=4'b1000;
    defparam blink_counter_332__i25_LC_13_24_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_332__i25_LC_13_24_1 (
            .in0(_gnd_net_),
            .in1(N__2731),
            .in2(_gnd_net_),
            .in3(N__2807),
            .lcout(blink_counter_25),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3933),
            .ce(),
            .sr(_gnd_net_));
    defparam i1846_4_lut_LC_13_24_2.C_ON=1'b0;
    defparam i1846_4_lut_LC_13_24_2.SEQ_MODE=4'b0000;
    defparam i1846_4_lut_LC_13_24_2.LUT_INIT=16'b1011101000100010;
    LogicCell40 i1846_4_lut_LC_13_24_2 (
            .in0(N__2803),
            .in1(N__2788),
            .in2(N__2776),
            .in3(N__2755),
            .lcout(n2730),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1847_4_lut_LC_13_24_4.C_ON=1'b0;
    defparam i1847_4_lut_LC_13_24_4.SEQ_MODE=4'b0000;
    defparam i1847_4_lut_LC_13_24_4.LUT_INIT=16'b1110101011111000;
    LogicCell40 i1847_4_lut_LC_13_24_4 (
            .in0(N__2804),
            .in1(N__2789),
            .in2(N__2777),
            .in3(N__2756),
            .lcout(),
            .ltout(n2731_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1848_3_lut_LC_13_24_5.C_ON=1'b0;
    defparam i1848_3_lut_LC_13_24_5.SEQ_MODE=4'b0000;
    defparam i1848_3_lut_LC_13_24_5.LUT_INIT=16'b0000111101010101;
    LogicCell40 i1848_3_lut_LC_13_24_5 (
            .in0(N__2741),
            .in1(_gnd_net_),
            .in2(N__2735),
            .in3(N__2732),
            .lcout(LED_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam delay_counter_331__i0_LC_14_21_0.C_ON=1'b1;
    defparam delay_counter_331__i0_LC_14_21_0.SEQ_MODE=4'b1000;
    defparam delay_counter_331__i0_LC_14_21_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 delay_counter_331__i0_LC_14_21_0 (
            .in0(_gnd_net_),
            .in1(N__3143),
            .in2(_gnd_net_),
            .in3(N__2705),
            .lcout(delay_counter_0),
            .ltout(),
            .carryin(bfn_14_21_0_),
            .carryout(n2478),
            .clk(N__3927),
            .ce(),
            .sr(N__3275));
    defparam delay_counter_331__i1_LC_14_21_1.C_ON=1'b1;
    defparam delay_counter_331__i1_LC_14_21_1.SEQ_MODE=4'b1000;
    defparam delay_counter_331__i1_LC_14_21_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 delay_counter_331__i1_LC_14_21_1 (
            .in0(_gnd_net_),
            .in1(N__3041),
            .in2(_gnd_net_),
            .in3(N__2702),
            .lcout(delay_counter_1),
            .ltout(),
            .carryin(n2478),
            .carryout(n2479),
            .clk(N__3927),
            .ce(),
            .sr(N__3275));
    defparam delay_counter_331__i2_LC_14_21_2.C_ON=1'b1;
    defparam delay_counter_331__i2_LC_14_21_2.SEQ_MODE=4'b1000;
    defparam delay_counter_331__i2_LC_14_21_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 delay_counter_331__i2_LC_14_21_2 (
            .in0(_gnd_net_),
            .in1(N__3104),
            .in2(_gnd_net_),
            .in3(N__2699),
            .lcout(delay_counter_2),
            .ltout(),
            .carryin(n2479),
            .carryout(n2480),
            .clk(N__3927),
            .ce(),
            .sr(N__3275));
    defparam delay_counter_331__i3_LC_14_21_3.C_ON=1'b1;
    defparam delay_counter_331__i3_LC_14_21_3.SEQ_MODE=4'b1000;
    defparam delay_counter_331__i3_LC_14_21_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 delay_counter_331__i3_LC_14_21_3 (
            .in0(_gnd_net_),
            .in1(N__3065),
            .in2(_gnd_net_),
            .in3(N__2840),
            .lcout(delay_counter_3),
            .ltout(),
            .carryin(n2480),
            .carryout(n2481),
            .clk(N__3927),
            .ce(),
            .sr(N__3275));
    defparam delay_counter_331__i4_LC_14_21_4.C_ON=1'b1;
    defparam delay_counter_331__i4_LC_14_21_4.SEQ_MODE=4'b1000;
    defparam delay_counter_331__i4_LC_14_21_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 delay_counter_331__i4_LC_14_21_4 (
            .in0(_gnd_net_),
            .in1(N__3116),
            .in2(_gnd_net_),
            .in3(N__2837),
            .lcout(delay_counter_4),
            .ltout(),
            .carryin(n2481),
            .carryout(n2482),
            .clk(N__3927),
            .ce(),
            .sr(N__3275));
    defparam delay_counter_331__i5_LC_14_21_5.C_ON=1'b1;
    defparam delay_counter_331__i5_LC_14_21_5.SEQ_MODE=4'b1000;
    defparam delay_counter_331__i5_LC_14_21_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 delay_counter_331__i5_LC_14_21_5 (
            .in0(_gnd_net_),
            .in1(N__3079),
            .in2(_gnd_net_),
            .in3(N__2834),
            .lcout(delay_counter_5),
            .ltout(),
            .carryin(n2482),
            .carryout(n2483),
            .clk(N__3927),
            .ce(),
            .sr(N__3275));
    defparam delay_counter_331__i6_LC_14_21_6.C_ON=1'b1;
    defparam delay_counter_331__i6_LC_14_21_6.SEQ_MODE=4'b1000;
    defparam delay_counter_331__i6_LC_14_21_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 delay_counter_331__i6_LC_14_21_6 (
            .in0(_gnd_net_),
            .in1(N__3155),
            .in2(_gnd_net_),
            .in3(N__2831),
            .lcout(delay_counter_6),
            .ltout(),
            .carryin(n2483),
            .carryout(n2484),
            .clk(N__3927),
            .ce(),
            .sr(N__3275));
    defparam delay_counter_331__i7_LC_14_21_7.C_ON=1'b1;
    defparam delay_counter_331__i7_LC_14_21_7.SEQ_MODE=4'b1000;
    defparam delay_counter_331__i7_LC_14_21_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 delay_counter_331__i7_LC_14_21_7 (
            .in0(_gnd_net_),
            .in1(N__3092),
            .in2(_gnd_net_),
            .in3(N__2828),
            .lcout(delay_counter_7),
            .ltout(),
            .carryin(n2484),
            .carryout(n2485),
            .clk(N__3927),
            .ce(),
            .sr(N__3275));
    defparam delay_counter_331__i8_LC_14_22_0.C_ON=1'b1;
    defparam delay_counter_331__i8_LC_14_22_0.SEQ_MODE=4'b1000;
    defparam delay_counter_331__i8_LC_14_22_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 delay_counter_331__i8_LC_14_22_0 (
            .in0(_gnd_net_),
            .in1(N__3053),
            .in2(_gnd_net_),
            .in3(N__2825),
            .lcout(delay_counter_8),
            .ltout(),
            .carryin(bfn_14_22_0_),
            .carryout(n2486),
            .clk(N__3931),
            .ce(),
            .sr(N__3267));
    defparam delay_counter_331__i9_LC_14_22_1.C_ON=1'b1;
    defparam delay_counter_331__i9_LC_14_22_1.SEQ_MODE=4'b1000;
    defparam delay_counter_331__i9_LC_14_22_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 delay_counter_331__i9_LC_14_22_1 (
            .in0(_gnd_net_),
            .in1(N__3130),
            .in2(_gnd_net_),
            .in3(N__2822),
            .lcout(delay_counter_9),
            .ltout(),
            .carryin(n2486),
            .carryout(n2487),
            .clk(N__3931),
            .ce(),
            .sr(N__3267));
    defparam delay_counter_331__i10_LC_14_22_2.C_ON=1'b1;
    defparam delay_counter_331__i10_LC_14_22_2.SEQ_MODE=4'b1000;
    defparam delay_counter_331__i10_LC_14_22_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 delay_counter_331__i10_LC_14_22_2 (
            .in0(_gnd_net_),
            .in1(N__2999),
            .in2(_gnd_net_),
            .in3(N__2819),
            .lcout(delay_counter_10),
            .ltout(),
            .carryin(n2487),
            .carryout(n2488),
            .clk(N__3931),
            .ce(),
            .sr(N__3267));
    defparam delay_counter_331__i11_LC_14_22_3.C_ON=1'b1;
    defparam delay_counter_331__i11_LC_14_22_3.SEQ_MODE=4'b1000;
    defparam delay_counter_331__i11_LC_14_22_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 delay_counter_331__i11_LC_14_22_3 (
            .in0(_gnd_net_),
            .in1(N__3011),
            .in2(_gnd_net_),
            .in3(N__2816),
            .lcout(delay_counter_11),
            .ltout(),
            .carryin(n2488),
            .carryout(n2489),
            .clk(N__3931),
            .ce(),
            .sr(N__3267));
    defparam delay_counter_331__i12_LC_14_22_4.C_ON=1'b1;
    defparam delay_counter_331__i12_LC_14_22_4.SEQ_MODE=4'b1000;
    defparam delay_counter_331__i12_LC_14_22_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 delay_counter_331__i12_LC_14_22_4 (
            .in0(_gnd_net_),
            .in1(N__2984),
            .in2(_gnd_net_),
            .in3(N__2813),
            .lcout(delay_counter_12),
            .ltout(),
            .carryin(n2489),
            .carryout(n2490),
            .clk(N__3931),
            .ce(),
            .sr(N__3267));
    defparam delay_counter_331__i13_LC_14_22_5.C_ON=1'b1;
    defparam delay_counter_331__i13_LC_14_22_5.SEQ_MODE=4'b1000;
    defparam delay_counter_331__i13_LC_14_22_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 delay_counter_331__i13_LC_14_22_5 (
            .in0(_gnd_net_),
            .in1(N__2914),
            .in2(_gnd_net_),
            .in3(N__2867),
            .lcout(delay_counter_13),
            .ltout(),
            .carryin(n2490),
            .carryout(n2491),
            .clk(N__3931),
            .ce(),
            .sr(N__3267));
    defparam delay_counter_331__i14_LC_14_22_6.C_ON=1'b1;
    defparam delay_counter_331__i14_LC_14_22_6.SEQ_MODE=4'b1000;
    defparam delay_counter_331__i14_LC_14_22_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 delay_counter_331__i14_LC_14_22_6 (
            .in0(_gnd_net_),
            .in1(N__2945),
            .in2(_gnd_net_),
            .in3(N__2864),
            .lcout(delay_counter_14),
            .ltout(),
            .carryin(n2491),
            .carryout(n2492),
            .clk(N__3931),
            .ce(),
            .sr(N__3267));
    defparam delay_counter_331__i15_LC_14_22_7.C_ON=1'b1;
    defparam delay_counter_331__i15_LC_14_22_7.SEQ_MODE=4'b1000;
    defparam delay_counter_331__i15_LC_14_22_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 delay_counter_331__i15_LC_14_22_7 (
            .in0(_gnd_net_),
            .in1(N__2957),
            .in2(_gnd_net_),
            .in3(N__2861),
            .lcout(delay_counter_15),
            .ltout(),
            .carryin(n2492),
            .carryout(n2493),
            .clk(N__3931),
            .ce(),
            .sr(N__3267));
    defparam delay_counter_331__i16_LC_14_23_0.C_ON=1'b1;
    defparam delay_counter_331__i16_LC_14_23_0.SEQ_MODE=4'b1000;
    defparam delay_counter_331__i16_LC_14_23_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 delay_counter_331__i16_LC_14_23_0 (
            .in0(_gnd_net_),
            .in1(N__2927),
            .in2(_gnd_net_),
            .in3(N__2858),
            .lcout(delay_counter_16),
            .ltout(),
            .carryin(bfn_14_23_0_),
            .carryout(n2494),
            .clk(N__3934),
            .ce(),
            .sr(N__3266));
    defparam delay_counter_331__i17_LC_14_23_1.C_ON=1'b1;
    defparam delay_counter_331__i17_LC_14_23_1.SEQ_MODE=4'b1000;
    defparam delay_counter_331__i17_LC_14_23_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 delay_counter_331__i17_LC_14_23_1 (
            .in0(_gnd_net_),
            .in1(N__2971),
            .in2(_gnd_net_),
            .in3(N__2855),
            .lcout(delay_counter_17),
            .ltout(),
            .carryin(n2494),
            .carryout(n2495),
            .clk(N__3934),
            .ce(),
            .sr(N__3266));
    defparam delay_counter_331__i18_LC_14_23_2.C_ON=1'b1;
    defparam delay_counter_331__i18_LC_14_23_2.SEQ_MODE=4'b1000;
    defparam delay_counter_331__i18_LC_14_23_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 delay_counter_331__i18_LC_14_23_2 (
            .in0(_gnd_net_),
            .in1(N__3401),
            .in2(_gnd_net_),
            .in3(N__2852),
            .lcout(delay_counter_18),
            .ltout(),
            .carryin(n2495),
            .carryout(n2496),
            .clk(N__3934),
            .ce(),
            .sr(N__3266));
    defparam delay_counter_331__i19_LC_14_23_3.C_ON=1'b1;
    defparam delay_counter_331__i19_LC_14_23_3.SEQ_MODE=4'b1000;
    defparam delay_counter_331__i19_LC_14_23_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 delay_counter_331__i19_LC_14_23_3 (
            .in0(_gnd_net_),
            .in1(N__3386),
            .in2(_gnd_net_),
            .in3(N__2849),
            .lcout(delay_counter_19),
            .ltout(),
            .carryin(n2496),
            .carryout(n2497),
            .clk(N__3934),
            .ce(),
            .sr(N__3266));
    defparam delay_counter_331__i20_LC_14_23_4.C_ON=1'b1;
    defparam delay_counter_331__i20_LC_14_23_4.SEQ_MODE=4'b1000;
    defparam delay_counter_331__i20_LC_14_23_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 delay_counter_331__i20_LC_14_23_4 (
            .in0(_gnd_net_),
            .in1(N__3331),
            .in2(_gnd_net_),
            .in3(N__2846),
            .lcout(delay_counter_20),
            .ltout(),
            .carryin(n2497),
            .carryout(n2498),
            .clk(N__3934),
            .ce(),
            .sr(N__3266));
    defparam delay_counter_331__i21_LC_14_23_5.C_ON=1'b1;
    defparam delay_counter_331__i21_LC_14_23_5.SEQ_MODE=4'b1000;
    defparam delay_counter_331__i21_LC_14_23_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 delay_counter_331__i21_LC_14_23_5 (
            .in0(_gnd_net_),
            .in1(N__3359),
            .in2(_gnd_net_),
            .in3(N__2843),
            .lcout(delay_counter_21),
            .ltout(),
            .carryin(n2498),
            .carryout(n2499),
            .clk(N__3934),
            .ce(),
            .sr(N__3266));
    defparam delay_counter_331__i22_LC_14_23_6.C_ON=1'b1;
    defparam delay_counter_331__i22_LC_14_23_6.SEQ_MODE=4'b1000;
    defparam delay_counter_331__i22_LC_14_23_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 delay_counter_331__i22_LC_14_23_6 (
            .in0(_gnd_net_),
            .in1(N__3371),
            .in2(_gnd_net_),
            .in3(N__2894),
            .lcout(delay_counter_22),
            .ltout(),
            .carryin(n2499),
            .carryout(n2500),
            .clk(N__3934),
            .ce(),
            .sr(N__3266));
    defparam delay_counter_331__i23_LC_14_23_7.C_ON=1'b1;
    defparam delay_counter_331__i23_LC_14_23_7.SEQ_MODE=4'b1000;
    defparam delay_counter_331__i23_LC_14_23_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 delay_counter_331__i23_LC_14_23_7 (
            .in0(_gnd_net_),
            .in1(N__3347),
            .in2(_gnd_net_),
            .in3(N__2891),
            .lcout(delay_counter_23),
            .ltout(),
            .carryin(n2500),
            .carryout(n2501),
            .clk(N__3934),
            .ce(),
            .sr(N__3266));
    defparam delay_counter_331__i24_LC_14_24_0.C_ON=1'b1;
    defparam delay_counter_331__i24_LC_14_24_0.SEQ_MODE=4'b1000;
    defparam delay_counter_331__i24_LC_14_24_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 delay_counter_331__i24_LC_14_24_0 (
            .in0(_gnd_net_),
            .in1(N__3182),
            .in2(_gnd_net_),
            .in3(N__2888),
            .lcout(delay_counter_24),
            .ltout(),
            .carryin(bfn_14_24_0_),
            .carryout(n2502),
            .clk(N__3939),
            .ce(),
            .sr(N__3268));
    defparam delay_counter_331__i25_LC_14_24_1.C_ON=1'b1;
    defparam delay_counter_331__i25_LC_14_24_1.SEQ_MODE=4'b1000;
    defparam delay_counter_331__i25_LC_14_24_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 delay_counter_331__i25_LC_14_24_1 (
            .in0(_gnd_net_),
            .in1(N__3305),
            .in2(_gnd_net_),
            .in3(N__2885),
            .lcout(delay_counter_25),
            .ltout(),
            .carryin(n2502),
            .carryout(n2503),
            .clk(N__3939),
            .ce(),
            .sr(N__3268));
    defparam delay_counter_331__i26_LC_14_24_2.C_ON=1'b1;
    defparam delay_counter_331__i26_LC_14_24_2.SEQ_MODE=4'b1000;
    defparam delay_counter_331__i26_LC_14_24_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 delay_counter_331__i26_LC_14_24_2 (
            .in0(_gnd_net_),
            .in1(N__3221),
            .in2(_gnd_net_),
            .in3(N__2882),
            .lcout(delay_counter_26),
            .ltout(),
            .carryin(n2503),
            .carryout(n2504),
            .clk(N__3939),
            .ce(),
            .sr(N__3268));
    defparam delay_counter_331__i27_LC_14_24_3.C_ON=1'b1;
    defparam delay_counter_331__i27_LC_14_24_3.SEQ_MODE=4'b1000;
    defparam delay_counter_331__i27_LC_14_24_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 delay_counter_331__i27_LC_14_24_3 (
            .in0(_gnd_net_),
            .in1(N__3196),
            .in2(_gnd_net_),
            .in3(N__2879),
            .lcout(delay_counter_27),
            .ltout(),
            .carryin(n2504),
            .carryout(n2505),
            .clk(N__3939),
            .ce(),
            .sr(N__3268));
    defparam delay_counter_331__i28_LC_14_24_4.C_ON=1'b1;
    defparam delay_counter_331__i28_LC_14_24_4.SEQ_MODE=4'b1000;
    defparam delay_counter_331__i28_LC_14_24_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 delay_counter_331__i28_LC_14_24_4 (
            .in0(_gnd_net_),
            .in1(N__3290),
            .in2(_gnd_net_),
            .in3(N__2876),
            .lcout(delay_counter_28),
            .ltout(),
            .carryin(n2505),
            .carryout(n2506),
            .clk(N__3939),
            .ce(),
            .sr(N__3268));
    defparam delay_counter_331__i29_LC_14_24_5.C_ON=1'b1;
    defparam delay_counter_331__i29_LC_14_24_5.SEQ_MODE=4'b1000;
    defparam delay_counter_331__i29_LC_14_24_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 delay_counter_331__i29_LC_14_24_5 (
            .in0(_gnd_net_),
            .in1(N__3317),
            .in2(_gnd_net_),
            .in3(N__2873),
            .lcout(delay_counter_29),
            .ltout(),
            .carryin(n2506),
            .carryout(n2507),
            .clk(N__3939),
            .ce(),
            .sr(N__3268));
    defparam delay_counter_331__i30_LC_14_24_6.C_ON=1'b1;
    defparam delay_counter_331__i30_LC_14_24_6.SEQ_MODE=4'b1000;
    defparam delay_counter_331__i30_LC_14_24_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 delay_counter_331__i30_LC_14_24_6 (
            .in0(_gnd_net_),
            .in1(N__3209),
            .in2(_gnd_net_),
            .in3(N__2870),
            .lcout(delay_counter_30),
            .ltout(),
            .carryin(n2507),
            .carryout(n2508),
            .clk(N__3939),
            .ce(),
            .sr(N__3268));
    defparam delay_counter_331__i31_LC_14_24_7.C_ON=1'b0;
    defparam delay_counter_331__i31_LC_14_24_7.SEQ_MODE=4'b1000;
    defparam delay_counter_331__i31_LC_14_24_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 delay_counter_331__i31_LC_14_24_7 (
            .in0(_gnd_net_),
            .in1(N__3245),
            .in2(_gnd_net_),
            .in3(N__3158),
            .lcout(delay_counter_31),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3939),
            .ce(),
            .sr(N__3268));
    defparam i6_4_lut_adj_15_LC_15_21_4.C_ON=1'b0;
    defparam i6_4_lut_adj_15_LC_15_21_4.SEQ_MODE=4'b0000;
    defparam i6_4_lut_adj_15_LC_15_21_4.LUT_INIT=16'b1111111111111110;
    LogicCell40 i6_4_lut_adj_15_LC_15_21_4 (
            .in0(N__3154),
            .in1(N__3142),
            .in2(N__3131),
            .in3(N__3115),
            .lcout(n16),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i7_4_lut_LC_15_21_6.C_ON=1'b0;
    defparam i7_4_lut_LC_15_21_6.SEQ_MODE=4'b0000;
    defparam i7_4_lut_LC_15_21_6.LUT_INIT=16'b1111111111111110;
    LogicCell40 i7_4_lut_LC_15_21_6 (
            .in0(N__3103),
            .in1(N__3091),
            .in2(N__3080),
            .in3(N__3064),
            .lcout(n17),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i9_4_lut_LC_15_22_1.C_ON=1'b0;
    defparam i9_4_lut_LC_15_22_1.SEQ_MODE=4'b0000;
    defparam i9_4_lut_LC_15_22_1.LUT_INIT=16'b1111111111111110;
    LogicCell40 i9_4_lut_LC_15_22_1 (
            .in0(N__3052),
            .in1(N__3040),
            .in2(N__3029),
            .in3(N__3017),
            .lcout(),
            .ltout(n2722_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i2_4_lut_adj_17_LC_15_22_2.C_ON=1'b0;
    defparam i2_4_lut_adj_17_LC_15_22_2.SEQ_MODE=4'b0000;
    defparam i2_4_lut_adj_17_LC_15_22_2.LUT_INIT=16'b1111111111101010;
    LogicCell40 i2_4_lut_adj_17_LC_15_22_2 (
            .in0(N__3010),
            .in1(N__2998),
            .in2(N__2987),
            .in3(N__2983),
            .lcout(n2715),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i3_3_lut_LC_15_22_4.C_ON=1'b0;
    defparam i3_3_lut_LC_15_22_4.SEQ_MODE=4'b0000;
    defparam i3_3_lut_LC_15_22_4.LUT_INIT=16'b1111111111101110;
    LogicCell40 i3_3_lut_LC_15_22_4 (
            .in0(N__2972),
            .in1(N__2956),
            .in2(_gnd_net_),
            .in3(N__2944),
            .lcout(n8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i4_4_lut_adj_18_LC_15_23_1.C_ON=1'b0;
    defparam i4_4_lut_adj_18_LC_15_23_1.SEQ_MODE=4'b0000;
    defparam i4_4_lut_adj_18_LC_15_23_1.LUT_INIT=16'b1111111011101110;
    LogicCell40 i4_4_lut_adj_18_LC_15_23_1 (
            .in0(N__2933),
            .in1(N__2926),
            .in2(N__2915),
            .in3(N__2900),
            .lcout(),
            .ltout(n2721_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i2_4_lut_LC_15_23_2.C_ON=1'b0;
    defparam i2_4_lut_LC_15_23_2.SEQ_MODE=4'b0000;
    defparam i2_4_lut_LC_15_23_2.LUT_INIT=16'b1110110000000000;
    LogicCell40 i2_4_lut_LC_15_23_2 (
            .in0(N__3400),
            .in1(N__3385),
            .in2(N__3374),
            .in3(N__3370),
            .lcout(),
            .ltout(n7_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i4_4_lut_LC_15_23_3.C_ON=1'b0;
    defparam i4_4_lut_LC_15_23_3.SEQ_MODE=4'b0000;
    defparam i4_4_lut_LC_15_23_3.LUT_INIT=16'b1000000000000000;
    LogicCell40 i4_4_lut_LC_15_23_3 (
            .in0(N__3358),
            .in1(N__3346),
            .in2(N__3335),
            .in3(N__3332),
            .lcout(),
            .ltout(n2695_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i5_4_lut_LC_15_23_4.C_ON=1'b0;
    defparam i5_4_lut_LC_15_23_4.SEQ_MODE=4'b0000;
    defparam i5_4_lut_LC_15_23_4.LUT_INIT=16'b1111111111111110;
    LogicCell40 i5_4_lut_LC_15_23_4 (
            .in0(N__3316),
            .in1(N__3304),
            .in2(N__3293),
            .in3(N__3289),
            .lcout(n13),
            .ltout(n13_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1200_3_lut_LC_15_23_5.C_ON=1'b0;
    defparam i1200_3_lut_LC_15_23_5.SEQ_MODE=4'b0000;
    defparam i1200_3_lut_LC_15_23_5.LUT_INIT=16'b0011001100110000;
    LogicCell40 i1200_3_lut_LC_15_23_5 (
            .in0(_gnd_net_),
            .in1(N__3243),
            .in2(N__3278),
            .in3(N__3169),
            .lcout(addr_10__N_70),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam read_15_LC_15_23_7.C_ON=1'b0;
    defparam read_15_LC_15_23_7.SEQ_MODE=4'b1000;
    defparam read_15_LC_15_23_7.LUT_INIT=16'b0101010101000100;
    LogicCell40 read_15_LC_15_23_7 (
            .in0(N__3244),
            .in1(N__3170),
            .in2(_gnd_net_),
            .in3(N__3227),
            .lcout(read),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3940),
            .ce(),
            .sr(_gnd_net_));
    defparam i6_4_lut_LC_15_24_6.C_ON=1'b0;
    defparam i6_4_lut_LC_15_24_6.SEQ_MODE=4'b0000;
    defparam i6_4_lut_LC_15_24_6.LUT_INIT=16'b1111111111111110;
    LogicCell40 i6_4_lut_LC_15_24_6 (
            .in0(N__3220),
            .in1(N__3208),
            .in2(N__3197),
            .in3(N__3181),
            .lcout(n14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i1275_2_lut_3_lut_LC_17_18_0 .C_ON=1'b0;
    defparam \eeprom.i1275_2_lut_3_lut_LC_17_18_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.i1275_2_lut_3_lut_LC_17_18_0 .LUT_INIT=16'b1111111110111011;
    LogicCell40 \eeprom.i1275_2_lut_3_lut_LC_17_18_0  (
            .in0(N__4216),
            .in1(N__3876),
            .in2(_gnd_net_),
            .in3(N__4004),
            .lcout(n2077),
            .ltout(n2077_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.state__i0_LC_17_18_1 .C_ON=1'b0;
    defparam \eeprom.state__i0_LC_17_18_1 .SEQ_MODE=4'b1000;
    defparam \eeprom.state__i0_LC_17_18_1 .LUT_INIT=16'b1001000010000000;
    LogicCell40 \eeprom.state__i0_LC_17_18_1  (
            .in0(N__4005),
            .in1(N__3680),
            .in2(N__3161),
            .in3(N__4057),
            .lcout(state_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3928),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_3_lut_LC_17_18_4.C_ON=1'b0;
    defparam i1_3_lut_LC_17_18_4.SEQ_MODE=4'b0000;
    defparam i1_3_lut_LC_17_18_4.LUT_INIT=16'b1100110001000100;
    LogicCell40 i1_3_lut_LC_17_18_4 (
            .in0(N__4056),
            .in1(N__3877),
            .in2(_gnd_net_),
            .in3(N__3678),
            .lcout(),
            .ltout(n12_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.state__i1_LC_17_18_5 .C_ON=1'b0;
    defparam \eeprom.state__i1_LC_17_18_5 .SEQ_MODE=4'b1000;
    defparam \eeprom.state__i1_LC_17_18_5 .LUT_INIT=16'b1100010011000000;
    LogicCell40 \eeprom.state__i1_LC_17_18_5  (
            .in0(N__3679),
            .in1(N__3431),
            .in2(N__3425),
            .in3(N__4006),
            .lcout(state_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3928),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.delay_counter_i0_i0_LC_17_19_0 .C_ON=1'b1;
    defparam \eeprom.delay_counter_i0_i0_LC_17_19_0 .SEQ_MODE=4'b1000;
    defparam \eeprom.delay_counter_i0_i0_LC_17_19_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.delay_counter_i0_i0_LC_17_19_0  (
            .in0(_gnd_net_),
            .in1(N__3560),
            .in2(N__3665),
            .in3(_gnd_net_),
            .lcout(\eeprom.delay_counter_0 ),
            .ltout(),
            .carryin(bfn_17_19_0_),
            .carryout(\eeprom.n2516 ),
            .clk(N__3932),
            .ce(N__3517),
            .sr(N__3503));
    defparam \eeprom.delay_counter_i0_i1_LC_17_19_1 .C_ON=1'b1;
    defparam \eeprom.delay_counter_i0_i1_LC_17_19_1 .SEQ_MODE=4'b1000;
    defparam \eeprom.delay_counter_i0_i1_LC_17_19_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.delay_counter_i0_i1_LC_17_19_1  (
            .in0(_gnd_net_),
            .in1(N__3791),
            .in2(N__3592),
            .in3(N__3422),
            .lcout(\eeprom.delay_counter_1 ),
            .ltout(),
            .carryin(\eeprom.n2516 ),
            .carryout(\eeprom.n2517 ),
            .clk(N__3932),
            .ce(N__3517),
            .sr(N__3503));
    defparam \eeprom.delay_counter_i0_i2_LC_17_19_2 .C_ON=1'b1;
    defparam \eeprom.delay_counter_i0_i2_LC_17_19_2 .SEQ_MODE=4'b1000;
    defparam \eeprom.delay_counter_i0_i2_LC_17_19_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.delay_counter_i0_i2_LC_17_19_2  (
            .in0(_gnd_net_),
            .in1(N__3564),
            .in2(N__3650),
            .in3(N__3419),
            .lcout(\eeprom.delay_counter_2 ),
            .ltout(),
            .carryin(\eeprom.n2517 ),
            .carryout(\eeprom.n2518 ),
            .clk(N__3932),
            .ce(N__3517),
            .sr(N__3503));
    defparam \eeprom.delay_counter_i0_i3_LC_17_19_3 .C_ON=1'b1;
    defparam \eeprom.delay_counter_i0_i3_LC_17_19_3 .SEQ_MODE=4'b1000;
    defparam \eeprom.delay_counter_i0_i3_LC_17_19_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.delay_counter_i0_i3_LC_17_19_3  (
            .in0(_gnd_net_),
            .in1(N__3764),
            .in2(N__3593),
            .in3(N__3416),
            .lcout(\eeprom.delay_counter_3 ),
            .ltout(),
            .carryin(\eeprom.n2518 ),
            .carryout(\eeprom.n2519 ),
            .clk(N__3932),
            .ce(N__3517),
            .sr(N__3503));
    defparam \eeprom.delay_counter_i0_i4_LC_17_19_4 .C_ON=1'b1;
    defparam \eeprom.delay_counter_i0_i4_LC_17_19_4 .SEQ_MODE=4'b1001;
    defparam \eeprom.delay_counter_i0_i4_LC_17_19_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.delay_counter_i0_i4_LC_17_19_4  (
            .in0(_gnd_net_),
            .in1(N__3568),
            .in2(N__3719),
            .in3(N__3413),
            .lcout(\eeprom.delay_counter_4 ),
            .ltout(),
            .carryin(\eeprom.n2519 ),
            .carryout(\eeprom.n2520 ),
            .clk(N__3932),
            .ce(N__3517),
            .sr(N__3503));
    defparam \eeprom.delay_counter_i0_i5_LC_17_19_5 .C_ON=1'b1;
    defparam \eeprom.delay_counter_i0_i5_LC_17_19_5 .SEQ_MODE=4'b1000;
    defparam \eeprom.delay_counter_i0_i5_LC_17_19_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.delay_counter_i0_i5_LC_17_19_5  (
            .in0(_gnd_net_),
            .in1(N__3632),
            .in2(N__3594),
            .in3(N__3410),
            .lcout(\eeprom.delay_counter_5 ),
            .ltout(),
            .carryin(\eeprom.n2520 ),
            .carryout(\eeprom.n2521 ),
            .clk(N__3932),
            .ce(N__3517),
            .sr(N__3503));
    defparam \eeprom.delay_counter_i0_i6_LC_17_19_6 .C_ON=1'b1;
    defparam \eeprom.delay_counter_i0_i6_LC_17_19_6 .SEQ_MODE=4'b1001;
    defparam \eeprom.delay_counter_i0_i6_LC_17_19_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.delay_counter_i0_i6_LC_17_19_6  (
            .in0(_gnd_net_),
            .in1(N__3488),
            .in2(N__3596),
            .in3(N__3407),
            .lcout(\eeprom.delay_counter_6 ),
            .ltout(),
            .carryin(\eeprom.n2521 ),
            .carryout(\eeprom.n2522 ),
            .clk(N__3932),
            .ce(N__3517),
            .sr(N__3503));
    defparam \eeprom.delay_counter_i0_i7_LC_17_19_7 .C_ON=1'b1;
    defparam \eeprom.delay_counter_i0_i7_LC_17_19_7 .SEQ_MODE=4'b1001;
    defparam \eeprom.delay_counter_i0_i7_LC_17_19_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.delay_counter_i0_i7_LC_17_19_7  (
            .in0(_gnd_net_),
            .in1(N__3779),
            .in2(N__3595),
            .in3(N__3404),
            .lcout(\eeprom.delay_counter_7 ),
            .ltout(),
            .carryin(\eeprom.n2522 ),
            .carryout(\eeprom.n2523 ),
            .clk(N__3932),
            .ce(N__3517),
            .sr(N__3503));
    defparam \eeprom.delay_counter_i0_i8_LC_17_20_0 .C_ON=1'b1;
    defparam \eeprom.delay_counter_i0_i8_LC_17_20_0 .SEQ_MODE=4'b1001;
    defparam \eeprom.delay_counter_i0_i8_LC_17_20_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.delay_counter_i0_i8_LC_17_20_0  (
            .in0(_gnd_net_),
            .in1(N__3578),
            .in2(N__3734),
            .in3(N__3455),
            .lcout(\eeprom.delay_counter_8 ),
            .ltout(),
            .carryin(bfn_17_20_0_),
            .carryout(\eeprom.n2524 ),
            .clk(N__3935),
            .ce(N__3518),
            .sr(N__3502));
    defparam \eeprom.delay_counter_i0_i9_LC_17_20_1 .C_ON=1'b1;
    defparam \eeprom.delay_counter_i0_i9_LC_17_20_1 .SEQ_MODE=4'b1001;
    defparam \eeprom.delay_counter_i0_i9_LC_17_20_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.delay_counter_i0_i9_LC_17_20_1  (
            .in0(_gnd_net_),
            .in1(N__3803),
            .in2(N__3597),
            .in3(N__3452),
            .lcout(\eeprom.delay_counter_9 ),
            .ltout(),
            .carryin(\eeprom.n2524 ),
            .carryout(\eeprom.n2525 ),
            .clk(N__3935),
            .ce(N__3518),
            .sr(N__3502));
    defparam \eeprom.delay_counter_i0_i10_LC_17_20_2 .C_ON=1'b1;
    defparam \eeprom.delay_counter_i0_i10_LC_17_20_2 .SEQ_MODE=4'b1001;
    defparam \eeprom.delay_counter_i0_i10_LC_17_20_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.delay_counter_i0_i10_LC_17_20_2  (
            .in0(_gnd_net_),
            .in1(N__3582),
            .in2(N__3620),
            .in3(N__3449),
            .lcout(\eeprom.delay_counter_10 ),
            .ltout(),
            .carryin(\eeprom.n2525 ),
            .carryout(\eeprom.n2526 ),
            .clk(N__3935),
            .ce(N__3518),
            .sr(N__3502));
    defparam \eeprom.delay_counter_i0_i11_LC_17_20_3 .C_ON=1'b1;
    defparam \eeprom.delay_counter_i0_i11_LC_17_20_3 .SEQ_MODE=4'b1000;
    defparam \eeprom.delay_counter_i0_i11_LC_17_20_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.delay_counter_i0_i11_LC_17_20_3  (
            .in0(_gnd_net_),
            .in1(N__3830),
            .in2(N__3598),
            .in3(N__3446),
            .lcout(\eeprom.delay_counter_11 ),
            .ltout(),
            .carryin(\eeprom.n2526 ),
            .carryout(\eeprom.n2527 ),
            .clk(N__3935),
            .ce(N__3518),
            .sr(N__3502));
    defparam \eeprom.delay_counter_i0_i12_LC_17_20_4 .C_ON=1'b1;
    defparam \eeprom.delay_counter_i0_i12_LC_17_20_4 .SEQ_MODE=4'b1000;
    defparam \eeprom.delay_counter_i0_i12_LC_17_20_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.delay_counter_i0_i12_LC_17_20_4  (
            .in0(_gnd_net_),
            .in1(N__3586),
            .in2(N__3476),
            .in3(N__3443),
            .lcout(\eeprom.delay_counter_12 ),
            .ltout(),
            .carryin(\eeprom.n2527 ),
            .carryout(\eeprom.n2528 ),
            .clk(N__3935),
            .ce(N__3518),
            .sr(N__3502));
    defparam \eeprom.delay_counter_i0_i13_LC_17_20_5 .C_ON=1'b1;
    defparam \eeprom.delay_counter_i0_i13_LC_17_20_5 .SEQ_MODE=4'b1000;
    defparam \eeprom.delay_counter_i0_i13_LC_17_20_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.delay_counter_i0_i13_LC_17_20_5  (
            .in0(_gnd_net_),
            .in1(N__3746),
            .in2(N__3599),
            .in3(N__3440),
            .lcout(\eeprom.delay_counter_13 ),
            .ltout(),
            .carryin(\eeprom.n2528 ),
            .carryout(\eeprom.n2529 ),
            .clk(N__3935),
            .ce(N__3518),
            .sr(N__3502));
    defparam \eeprom.delay_counter_i0_i14_LC_17_20_6 .C_ON=1'b1;
    defparam \eeprom.delay_counter_i0_i14_LC_17_20_6 .SEQ_MODE=4'b1000;
    defparam \eeprom.delay_counter_i0_i14_LC_17_20_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.delay_counter_i0_i14_LC_17_20_6  (
            .in0(_gnd_net_),
            .in1(N__3590),
            .in2(N__3845),
            .in3(N__3437),
            .lcout(\eeprom.delay_counter_14 ),
            .ltout(),
            .carryin(\eeprom.n2529 ),
            .carryout(\eeprom.n2530 ),
            .clk(N__3935),
            .ce(N__3518),
            .sr(N__3502));
    defparam \eeprom.delay_counter_i0_i15_LC_17_20_7 .C_ON=1'b0;
    defparam \eeprom.delay_counter_i0_i15_LC_17_20_7 .SEQ_MODE=4'b1000;
    defparam \eeprom.delay_counter_i0_i15_LC_17_20_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \eeprom.delay_counter_i0_i15_LC_17_20_7  (
            .in0(N__3591),
            .in1(N__3817),
            .in2(_gnd_net_),
            .in3(N__3434),
            .lcout(\eeprom.delay_counter_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3935),
            .ce(N__3518),
            .sr(N__3502));
    defparam \eeprom.i2_2_lut_adj_14_LC_18_18_0 .C_ON=1'b0;
    defparam \eeprom.i2_2_lut_adj_14_LC_18_18_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.i2_2_lut_adj_14_LC_18_18_0 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \eeprom.i2_2_lut_adj_14_LC_18_18_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__3962),
            .in3(N__5579),
            .lcout(),
            .ltout(n6_adj_397_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1779_4_lut_LC_18_18_1.C_ON=1'b0;
    defparam i1779_4_lut_LC_18_18_1.SEQ_MODE=4'b0000;
    defparam i1779_4_lut_LC_18_18_1.LUT_INIT=16'b1010101010101000;
    LogicCell40 i1779_4_lut_LC_18_18_1 (
            .in0(N__3998),
            .in1(N__4286),
            .in2(N__3686),
            .in3(N__5429),
            .lcout(),
            .ltout(n2662_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i1785_4_lut_4_lut_LC_18_18_2 .C_ON=1'b0;
    defparam \eeprom.i1785_4_lut_4_lut_LC_18_18_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.i1785_4_lut_4_lut_LC_18_18_2 .LUT_INIT=16'b1111111011110000;
    LogicCell40 \eeprom.i1785_4_lut_4_lut_LC_18_18_2  (
            .in0(N__4218),
            .in1(N__3999),
            .in2(N__3683),
            .in3(N__3873),
            .lcout(n2668),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i11_4_lut_LC_18_19_0 .C_ON=1'b0;
    defparam \eeprom.i11_4_lut_LC_18_19_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.i11_4_lut_LC_18_19_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \eeprom.i11_4_lut_LC_18_19_0  (
            .in0(N__3661),
            .in1(N__3461),
            .in2(N__3649),
            .in3(N__3752),
            .lcout(),
            .ltout(\eeprom.n24_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i12_4_lut_LC_18_19_1 .C_ON=1'b0;
    defparam \eeprom.i12_4_lut_LC_18_19_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.i12_4_lut_LC_18_19_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \eeprom.i12_4_lut_LC_18_19_1  (
            .in0(N__3631),
            .in1(N__3616),
            .in2(N__3605),
            .in3(N__3704),
            .lcout(\eeprom.n1338 ),
            .ltout(\eeprom.n1338_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i1902_2_lut_LC_18_19_2 .C_ON=1'b0;
    defparam \eeprom.i1902_2_lut_LC_18_19_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.i1902_2_lut_LC_18_19_2 .LUT_INIT=16'b0000000011110000;
    LogicCell40 \eeprom.i1902_2_lut_LC_18_19_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__3602),
            .in3(N__4219),
            .lcout(\eeprom.n575 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i1_3_lut_LC_18_19_3 .C_ON=1'b0;
    defparam \eeprom.i1_3_lut_LC_18_19_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.i1_3_lut_LC_18_19_3 .LUT_INIT=16'b0011001100100010;
    LogicCell40 \eeprom.i1_3_lut_LC_18_19_3  (
            .in0(N__4052),
            .in1(N__3874),
            .in2(_gnd_net_),
            .in3(N__4000),
            .lcout(\eeprom.n1435 ),
            .ltout(\eeprom.n1435_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i717_2_lut_LC_18_19_4 .C_ON=1'b0;
    defparam \eeprom.i717_2_lut_LC_18_19_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.i717_2_lut_LC_18_19_4 .LUT_INIT=16'b0101000001010000;
    LogicCell40 \eeprom.i717_2_lut_LC_18_19_4  (
            .in0(N__4001),
            .in1(_gnd_net_),
            .in2(N__3506),
            .in3(_gnd_net_),
            .lcout(\eeprom.n1503 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i3_2_lut_LC_18_19_5 .C_ON=1'b0;
    defparam \eeprom.i3_2_lut_LC_18_19_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.i3_2_lut_LC_18_19_5 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \eeprom.i3_2_lut_LC_18_19_5  (
            .in0(_gnd_net_),
            .in1(N__3487),
            .in2(_gnd_net_),
            .in3(N__3472),
            .lcout(\eeprom.n16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.mux_161_Mux_0_i1_4_lut_LC_18_19_6 .C_ON=1'b0;
    defparam \eeprom.mux_161_Mux_0_i1_4_lut_LC_18_19_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.mux_161_Mux_0_i1_4_lut_LC_18_19_6 .LUT_INIT=16'b0101000001110010;
    LogicCell40 \eeprom.mux_161_Mux_0_i1_4_lut_LC_18_19_6  (
            .in0(N__4002),
            .in1(N__4220),
            .in2(N__4058),
            .in3(N__3960),
            .lcout(),
            .ltout(n624_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rw_43_LC_18_19_7 .C_ON=1'b0;
    defparam \eeprom.rw_43_LC_18_19_7 .SEQ_MODE=4'b1000;
    defparam \eeprom.rw_43_LC_18_19_7 .LUT_INIT=16'b1011101010001010;
    LogicCell40 \eeprom.rw_43_LC_18_19_7  (
            .in0(N__4231),
            .in1(N__3875),
            .in2(N__3848),
            .in3(N__4003),
            .lcout(rw),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3936),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i3_4_lut_LC_18_20_1 .C_ON=1'b0;
    defparam \eeprom.i3_4_lut_LC_18_20_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.i3_4_lut_LC_18_20_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \eeprom.i3_4_lut_LC_18_20_1  (
            .in0(N__3841),
            .in1(N__3829),
            .in2(N__3818),
            .in3(N__3802),
            .lcout(),
            .ltout(\eeprom.n2685_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i9_4_lut_LC_18_20_2 .C_ON=1'b0;
    defparam \eeprom.i9_4_lut_LC_18_20_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.i9_4_lut_LC_18_20_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \eeprom.i9_4_lut_LC_18_20_2  (
            .in0(N__3790),
            .in1(N__3778),
            .in2(N__3767),
            .in3(N__3763),
            .lcout(\eeprom.n22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i7_3_lut_LC_18_20_5 .C_ON=1'b0;
    defparam \eeprom.i7_3_lut_LC_18_20_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.i7_3_lut_LC_18_20_5 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \eeprom.i7_3_lut_LC_18_20_5  (
            .in0(N__3745),
            .in1(N__3730),
            .in2(_gnd_net_),
            .in3(N__3715),
            .lcout(\eeprom.n20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i2c.enable_slow_121_LC_19_15_5 .C_ON=1'b0;
    defparam \eeprom.i2c.enable_slow_121_LC_19_15_5 .SEQ_MODE=4'b1001;
    defparam \eeprom.i2c.enable_slow_121_LC_19_15_5 .LUT_INIT=16'b0011001111111111;
    LogicCell40 \eeprom.i2c.enable_slow_121_LC_19_15_5  (
            .in0(_gnd_net_),
            .in1(N__4896),
            .in2(_gnd_net_),
            .in3(N__4075),
            .lcout(state_7_N_269_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3941),
            .ce(N__3692),
            .sr(N__4351));
    defparam \eeprom.i2c.i1_2_lut_LC_19_16_1 .C_ON=1'b0;
    defparam \eeprom.i2c.i1_2_lut_LC_19_16_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.i2c.i1_2_lut_LC_19_16_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \eeprom.i2c.i1_2_lut_LC_19_16_1  (
            .in0(_gnd_net_),
            .in1(N__4156),
            .in2(_gnd_net_),
            .in3(N__4093),
            .lcout(),
            .ltout(\eeprom.i2c.n6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i2c.i4_4_lut_LC_19_16_2 .C_ON=1'b0;
    defparam \eeprom.i2c.i4_4_lut_LC_19_16_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.i2c.i4_4_lut_LC_19_16_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \eeprom.i2c.i4_4_lut_LC_19_16_2  (
            .in0(N__4141),
            .in1(N__4126),
            .in2(N__3698),
            .in3(N__4111),
            .lcout(\eeprom.i2c.counter2_7__N_256 ),
            .ltout(\eeprom.i2c.counter2_7__N_256_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i2c.i1_2_lut_3_lut_LC_19_16_3 .C_ON=1'b0;
    defparam \eeprom.i2c.i1_2_lut_3_lut_LC_19_16_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.i2c.i1_2_lut_3_lut_LC_19_16_3 .LUT_INIT=16'b1111111110100000;
    LogicCell40 \eeprom.i2c.i1_2_lut_3_lut_LC_19_16_3  (
            .in0(N__4894),
            .in1(_gnd_net_),
            .in2(N__3695),
            .in3(N__4341),
            .lcout(\eeprom.i2c.n1384 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i2c.i2c_clk_122_LC_19_16_7 .C_ON=1'b0;
    defparam \eeprom.i2c.i2c_clk_122_LC_19_16_7 .SEQ_MODE=4'b1000;
    defparam \eeprom.i2c.i2c_clk_122_LC_19_16_7 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \eeprom.i2c.i2c_clk_122_LC_19_16_7  (
            .in0(N__4895),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4074),
            .lcout(\eeprom.i2c.i2c_clk ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3937),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i2c.counter2_333_334__i1_LC_19_17_0 .C_ON=1'b1;
    defparam \eeprom.i2c.counter2_333_334__i1_LC_19_17_0 .SEQ_MODE=4'b1000;
    defparam \eeprom.i2c.counter2_333_334__i1_LC_19_17_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.i2c.counter2_333_334__i1_LC_19_17_0  (
            .in0(_gnd_net_),
            .in1(N__4157),
            .in2(_gnd_net_),
            .in3(N__4145),
            .lcout(\eeprom.i2c.counter2_0 ),
            .ltout(),
            .carryin(bfn_19_17_0_),
            .carryout(\eeprom.i2c.n2531 ),
            .clk(N__3929),
            .ce(),
            .sr(N__4082));
    defparam \eeprom.i2c.counter2_333_334__i2_LC_19_17_1 .C_ON=1'b1;
    defparam \eeprom.i2c.counter2_333_334__i2_LC_19_17_1 .SEQ_MODE=4'b1000;
    defparam \eeprom.i2c.counter2_333_334__i2_LC_19_17_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.i2c.counter2_333_334__i2_LC_19_17_1  (
            .in0(_gnd_net_),
            .in1(N__4142),
            .in2(_gnd_net_),
            .in3(N__4130),
            .lcout(\eeprom.i2c.counter2_1 ),
            .ltout(),
            .carryin(\eeprom.i2c.n2531 ),
            .carryout(\eeprom.i2c.n2532 ),
            .clk(N__3929),
            .ce(),
            .sr(N__4082));
    defparam \eeprom.i2c.counter2_333_334__i3_LC_19_17_2 .C_ON=1'b1;
    defparam \eeprom.i2c.counter2_333_334__i3_LC_19_17_2 .SEQ_MODE=4'b1000;
    defparam \eeprom.i2c.counter2_333_334__i3_LC_19_17_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.i2c.counter2_333_334__i3_LC_19_17_2  (
            .in0(_gnd_net_),
            .in1(N__4127),
            .in2(_gnd_net_),
            .in3(N__4115),
            .lcout(\eeprom.i2c.counter2_2 ),
            .ltout(),
            .carryin(\eeprom.i2c.n2532 ),
            .carryout(\eeprom.i2c.n2533 ),
            .clk(N__3929),
            .ce(),
            .sr(N__4082));
    defparam \eeprom.i2c.counter2_333_334__i4_LC_19_17_3 .C_ON=1'b1;
    defparam \eeprom.i2c.counter2_333_334__i4_LC_19_17_3 .SEQ_MODE=4'b1000;
    defparam \eeprom.i2c.counter2_333_334__i4_LC_19_17_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.i2c.counter2_333_334__i4_LC_19_17_3  (
            .in0(_gnd_net_),
            .in1(N__4112),
            .in2(_gnd_net_),
            .in3(N__4100),
            .lcout(\eeprom.i2c.counter2_3 ),
            .ltout(),
            .carryin(\eeprom.i2c.n2533 ),
            .carryout(\eeprom.i2c.n2534 ),
            .clk(N__3929),
            .ce(),
            .sr(N__4082));
    defparam \eeprom.i2c.counter2_333_334__i5_LC_19_17_4 .C_ON=1'b0;
    defparam \eeprom.i2c.counter2_333_334__i5_LC_19_17_4 .SEQ_MODE=4'b1000;
    defparam \eeprom.i2c.counter2_333_334__i5_LC_19_17_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.i2c.counter2_333_334__i5_LC_19_17_4  (
            .in0(_gnd_net_),
            .in1(N__4094),
            .in2(_gnd_net_),
            .in3(N__4097),
            .lcout(\eeprom.i2c.counter2_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3929),
            .ce(),
            .sr(N__4082));
    defparam \eeprom.enable_39_LC_19_18_1 .C_ON=1'b0;
    defparam \eeprom.enable_39_LC_19_18_1 .SEQ_MODE=4'b1000;
    defparam \eeprom.enable_39_LC_19_18_1 .LUT_INIT=16'b0010001000101110;
    LogicCell40 \eeprom.enable_39_LC_19_18_1  (
            .in0(N__4051),
            .in1(N__4010),
            .in2(N__4217),
            .in3(N__3961),
            .lcout(\eeprom.enable ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3938),
            .ce(),
            .sr(N__3884));
    defparam \eeprom.i2c.i1878_2_lut_3_lut_LC_20_14_0 .C_ON=1'b0;
    defparam \eeprom.i2c.i1878_2_lut_3_lut_LC_20_14_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.i2c.i1878_2_lut_3_lut_LC_20_14_0 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \eeprom.i2c.i1878_2_lut_3_lut_LC_20_14_0  (
            .in0(N__4443),
            .in1(N__4820),
            .in2(_gnd_net_),
            .in3(N__4789),
            .lcout(),
            .ltout(\eeprom.i2c.n2740_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i2c.i1880_4_lut_LC_20_14_1 .C_ON=1'b0;
    defparam \eeprom.i2c.i1880_4_lut_LC_20_14_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.i2c.i1880_4_lut_LC_20_14_1 .LUT_INIT=16'b1011100000000000;
    LogicCell40 \eeprom.i2c.i1880_4_lut_LC_20_14_1  (
            .in0(N__4790),
            .in1(N__4596),
            .in2(N__4268),
            .in3(N__5266),
            .lcout(\eeprom.i2c.n2734 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i2c.i1_2_lut_3_lut_adj_11_LC_20_14_4 .C_ON=1'b0;
    defparam \eeprom.i2c.i1_2_lut_3_lut_adj_11_LC_20_14_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.i2c.i1_2_lut_3_lut_adj_11_LC_20_14_4 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \eeprom.i2c.i1_2_lut_3_lut_adj_11_LC_20_14_4  (
            .in0(N__5546),
            .in1(N__5131),
            .in2(_gnd_net_),
            .in3(N__5424),
            .lcout(\eeprom.i2c.n970 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i2c.i1881_2_lut_3_lut_LC_20_14_6 .C_ON=1'b0;
    defparam \eeprom.i2c.i1881_2_lut_3_lut_LC_20_14_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.i2c.i1881_2_lut_3_lut_LC_20_14_6 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \eeprom.i2c.i1881_2_lut_3_lut_LC_20_14_6  (
            .in0(N__4844),
            .in1(N__4821),
            .in2(_gnd_net_),
            .in3(N__4791),
            .lcout(),
            .ltout(\eeprom.i2c.n2747_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i2c.i17_4_lut_LC_20_14_7 .C_ON=1'b0;
    defparam \eeprom.i2c.i17_4_lut_LC_20_14_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.i2c.i17_4_lut_LC_20_14_7 .LUT_INIT=16'b0100000011101010;
    LogicCell40 \eeprom.i2c.i17_4_lut_LC_20_14_7  (
            .in0(N__4265),
            .in1(N__4295),
            .in2(N__4259),
            .in3(N__4253),
            .lcout(\eeprom.i2c.n1413 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i2c.equal_31_i11_2_lut_3_lut_4_lut_LC_20_15_0 .C_ON=1'b0;
    defparam \eeprom.i2c.equal_31_i11_2_lut_3_lut_4_lut_LC_20_15_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.i2c.equal_31_i11_2_lut_3_lut_4_lut_LC_20_15_0 .LUT_INIT=16'b1111111111101111;
    LogicCell40 \eeprom.i2c.equal_31_i11_2_lut_3_lut_4_lut_LC_20_15_0  (
            .in0(N__5129),
            .in1(N__5270),
            .in2(N__5428),
            .in3(N__5566),
            .lcout(),
            .ltout(\eeprom.i2c.n15_adj_381_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i2c.i1788_2_lut_3_lut_LC_20_15_1 .C_ON=1'b0;
    defparam \eeprom.i2c.i1788_2_lut_3_lut_LC_20_15_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.i2c.i1788_2_lut_3_lut_LC_20_15_1 .LUT_INIT=16'b1100000000000000;
    LogicCell40 \eeprom.i2c.i1788_2_lut_3_lut_LC_20_15_1  (
            .in0(_gnd_net_),
            .in1(N__5706),
            .in2(N__4256),
            .in3(N__5650),
            .lcout(\eeprom.i2c.n2671 ),
            .ltout(\eeprom.i2c.n2671_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i2c.i1787_2_lut_4_lut_LC_20_15_2 .C_ON=1'b0;
    defparam \eeprom.i2c.i1787_2_lut_4_lut_LC_20_15_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.i2c.i1787_2_lut_4_lut_LC_20_15_2 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \eeprom.i2c.i1787_2_lut_4_lut_LC_20_15_2  (
            .in0(N__5130),
            .in1(N__5420),
            .in2(N__4247),
            .in3(N__5568),
            .lcout(\eeprom.i2c.n1495 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i2c.saved_addr__i1_LC_20_15_4 .C_ON=1'b0;
    defparam \eeprom.i2c.saved_addr__i1_LC_20_15_4 .SEQ_MODE=4'b1000;
    defparam \eeprom.i2c.saved_addr__i1_LC_20_15_4 .LUT_INIT=16'b1111110100100000;
    LogicCell40 \eeprom.i2c.saved_addr__i1_LC_20_15_4  (
            .in0(N__4166),
            .in1(N__4184),
            .in2(N__4244),
            .in3(N__4444),
            .lcout(saved_addr_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4954),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i2c.i1844_2_lut_3_lut_4_lut_LC_20_15_5 .C_ON=1'b0;
    defparam \eeprom.i2c.i1844_2_lut_3_lut_4_lut_LC_20_15_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.i2c.i1844_2_lut_3_lut_4_lut_LC_20_15_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \eeprom.i2c.i1844_2_lut_3_lut_4_lut_LC_20_15_5  (
            .in0(N__5567),
            .in1(N__5419),
            .in2(N__5280),
            .in3(N__5128),
            .lcout(n15),
            .ltout(n15_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i2c.i2_2_lut_LC_20_15_6 .C_ON=1'b0;
    defparam \eeprom.i2c.i2_2_lut_LC_20_15_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.i2c.i2_2_lut_LC_20_15_6 .LUT_INIT=16'b0000101000001010;
    LogicCell40 \eeprom.i2c.i2_2_lut_LC_20_15_6  (
            .in0(N__4165),
            .in1(_gnd_net_),
            .in2(N__4298),
            .in3(_gnd_net_),
            .lcout(\eeprom.i2c.n2714 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i2c.i1_2_lut_adj_9_LC_20_15_7 .C_ON=1'b0;
    defparam \eeprom.i2c.i1_2_lut_adj_9_LC_20_15_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.i2c.i1_2_lut_adj_9_LC_20_15_7 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \eeprom.i2c.i1_2_lut_adj_9_LC_20_15_7  (
            .in0(_gnd_net_),
            .in1(N__5565),
            .in2(_gnd_net_),
            .in3(N__4535),
            .lcout(\eeprom.i2c.n37 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i2c.i375_2_lut_LC_20_16_2 .C_ON=1'b0;
    defparam \eeprom.i2c.i375_2_lut_LC_20_16_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.i2c.i375_2_lut_LC_20_16_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \eeprom.i2c.i375_2_lut_LC_20_16_2  (
            .in0(_gnd_net_),
            .in1(N__5705),
            .in2(_gnd_net_),
            .in3(N__5649),
            .lcout(state_7_N_285_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i2c.i1781_2_lut_LC_20_16_3 .C_ON=1'b0;
    defparam \eeprom.i2c.i1781_2_lut_LC_20_16_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.i2c.i1781_2_lut_LC_20_16_3 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \eeprom.i2c.i1781_2_lut_LC_20_16_3  (
            .in0(_gnd_net_),
            .in1(N__5573),
            .in2(_gnd_net_),
            .in3(N__5133),
            .lcout(\eeprom.i2c.n2664 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i2c.state_7__I_0_145_i11_2_lut_3_lut_4_lut_LC_20_16_5 .C_ON=1'b0;
    defparam \eeprom.i2c.state_7__I_0_145_i11_2_lut_3_lut_4_lut_LC_20_16_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.i2c.state_7__I_0_145_i11_2_lut_3_lut_4_lut_LC_20_16_5 .LUT_INIT=16'b1111101111111111;
    LogicCell40 \eeprom.i2c.state_7__I_0_145_i11_2_lut_3_lut_4_lut_LC_20_16_5  (
            .in0(N__5574),
            .in1(N__5423),
            .in2(N__5281),
            .in3(N__5134),
            .lcout(\eeprom.i2c.n11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i2_2_lut_LC_20_18_7 .C_ON=1'b0;
    defparam \eeprom.i2_2_lut_LC_20_18_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.i2_2_lut_LC_20_18_7 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \eeprom.i2_2_lut_LC_20_18_7  (
            .in0(_gnd_net_),
            .in1(N__5278),
            .in2(_gnd_net_),
            .in3(N__5135),
            .lcout(n7_adj_385),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam CONSTANT_ONE_LUT4_LC_21_13_7.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_21_13_7.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_21_13_7.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_21_13_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i2c.counter_i0_LC_21_14_0 .C_ON=1'b1;
    defparam \eeprom.i2c.counter_i0_LC_21_14_0 .SEQ_MODE=4'b1001;
    defparam \eeprom.i2c.counter_i0_LC_21_14_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.i2c.counter_i0_LC_21_14_0  (
            .in0(_gnd_net_),
            .in1(N__4795),
            .in2(_gnd_net_),
            .in3(N__4277),
            .lcout(\eeprom.i2c.counter_0 ),
            .ltout(),
            .carryin(bfn_21_14_0_),
            .carryout(\eeprom.i2c.n2509 ),
            .clk(N__4953),
            .ce(N__4379),
            .sr(N__4370));
    defparam \eeprom.i2c.counter_i1_LC_21_14_1 .C_ON=1'b1;
    defparam \eeprom.i2c.counter_i1_LC_21_14_1 .SEQ_MODE=4'b1001;
    defparam \eeprom.i2c.counter_i1_LC_21_14_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.i2c.counter_i1_LC_21_14_1  (
            .in0(_gnd_net_),
            .in1(N__4825),
            .in2(N__4413),
            .in3(N__4274),
            .lcout(\eeprom.i2c.counter_1 ),
            .ltout(),
            .carryin(\eeprom.i2c.n2509 ),
            .carryout(\eeprom.i2c.n2510 ),
            .clk(N__4953),
            .ce(N__4379),
            .sr(N__4370));
    defparam \eeprom.i2c.counter_i2_LC_21_14_2 .C_ON=1'b1;
    defparam \eeprom.i2c.counter_i2_LC_21_14_2 .SEQ_MODE=4'b1001;
    defparam \eeprom.i2c.counter_i2_LC_21_14_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.i2c.counter_i2_LC_21_14_2  (
            .in0(_gnd_net_),
            .in1(N__4403),
            .in2(N__4601),
            .in3(N__4271),
            .lcout(\eeprom.i2c.counter_2 ),
            .ltout(),
            .carryin(\eeprom.i2c.n2510 ),
            .carryout(\eeprom.i2c.n2511 ),
            .clk(N__4953),
            .ce(N__4379),
            .sr(N__4370));
    defparam \eeprom.i2c.counter_i3_LC_21_14_3 .C_ON=1'b1;
    defparam \eeprom.i2c.counter_i3_LC_21_14_3 .SEQ_MODE=4'b1000;
    defparam \eeprom.i2c.counter_i3_LC_21_14_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.i2c.counter_i3_LC_21_14_3  (
            .in0(_gnd_net_),
            .in1(N__4618),
            .in2(N__4414),
            .in3(N__4427),
            .lcout(\eeprom.i2c.counter_3 ),
            .ltout(),
            .carryin(\eeprom.i2c.n2511 ),
            .carryout(\eeprom.i2c.n2512 ),
            .clk(N__4953),
            .ce(N__4379),
            .sr(N__4370));
    defparam \eeprom.i2c.counter_i4_LC_21_14_4 .C_ON=1'b1;
    defparam \eeprom.i2c.counter_i4_LC_21_14_4 .SEQ_MODE=4'b1000;
    defparam \eeprom.i2c.counter_i4_LC_21_14_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.i2c.counter_i4_LC_21_14_4  (
            .in0(_gnd_net_),
            .in1(N__4407),
            .in2(N__4688),
            .in3(N__4424),
            .lcout(\eeprom.i2c.counter_4 ),
            .ltout(),
            .carryin(\eeprom.i2c.n2512 ),
            .carryout(\eeprom.i2c.n2513 ),
            .clk(N__4953),
            .ce(N__4379),
            .sr(N__4370));
    defparam \eeprom.i2c.counter_i5_LC_21_14_5 .C_ON=1'b1;
    defparam \eeprom.i2c.counter_i5_LC_21_14_5 .SEQ_MODE=4'b1000;
    defparam \eeprom.i2c.counter_i5_LC_21_14_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.i2c.counter_i5_LC_21_14_5  (
            .in0(_gnd_net_),
            .in1(N__4633),
            .in2(N__4415),
            .in3(N__4421),
            .lcout(\eeprom.i2c.counter_5 ),
            .ltout(),
            .carryin(\eeprom.i2c.n2513 ),
            .carryout(\eeprom.i2c.n2514 ),
            .clk(N__4953),
            .ce(N__4379),
            .sr(N__4370));
    defparam \eeprom.i2c.counter_i6_LC_21_14_6 .C_ON=1'b1;
    defparam \eeprom.i2c.counter_i6_LC_21_14_6 .SEQ_MODE=4'b1000;
    defparam \eeprom.i2c.counter_i6_LC_21_14_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.i2c.counter_i6_LC_21_14_6  (
            .in0(_gnd_net_),
            .in1(N__4411),
            .in2(N__4670),
            .in3(N__4418),
            .lcout(\eeprom.i2c.counter_6 ),
            .ltout(),
            .carryin(\eeprom.i2c.n2514 ),
            .carryout(\eeprom.i2c.n2515 ),
            .clk(N__4953),
            .ce(N__4379),
            .sr(N__4370));
    defparam \eeprom.i2c.counter_i7_LC_21_14_7 .C_ON=1'b0;
    defparam \eeprom.i2c.counter_i7_LC_21_14_7 .SEQ_MODE=4'b1000;
    defparam \eeprom.i2c.counter_i7_LC_21_14_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \eeprom.i2c.counter_i7_LC_21_14_7  (
            .in0(N__4412),
            .in1(N__4648),
            .in2(_gnd_net_),
            .in3(N__4382),
            .lcout(\eeprom.i2c.counter_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4953),
            .ce(N__4379),
            .sr(N__4370));
    defparam \eeprom.i2c.sda_out_133_LC_21_15_3 .C_ON=1'b0;
    defparam \eeprom.i2c.sda_out_133_LC_21_15_3 .SEQ_MODE=4'b1000;
    defparam \eeprom.i2c.sda_out_133_LC_21_15_3 .LUT_INIT=16'b0000000001011100;
    LogicCell40 \eeprom.i2c.sda_out_133_LC_21_15_3  (
            .in0(N__5421),
            .in1(N__4358),
            .in2(N__4718),
            .in3(N__5132),
            .lcout(\eeprom.i2c.sda_out ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVeeprom.i2c.sda_out_133C_net ),
            .ce(N__4544),
            .sr(_gnd_net_));
    defparam \eeprom.i2c.i1865_4_lut_LC_21_15_7 .C_ON=1'b0;
    defparam \eeprom.i2c.i1865_4_lut_LC_21_15_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.i2c.i1865_4_lut_LC_21_15_7 .LUT_INIT=16'b0111011100000011;
    LogicCell40 \eeprom.i2c.i1865_4_lut_LC_21_15_7  (
            .in0(N__5682),
            .in1(N__5747),
            .in2(N__4352),
            .in3(N__4479),
            .lcout(\eeprom.i2c.n2736 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i2c.write_enable_132_LC_21_16_0 .C_ON=1'b0;
    defparam \eeprom.i2c.write_enable_132_LC_21_16_0 .SEQ_MODE=4'b1001;
    defparam \eeprom.i2c.write_enable_132_LC_21_16_0 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \eeprom.i2c.write_enable_132_LC_21_16_0  (
            .in0(N__4714),
            .in1(N__5422),
            .in2(_gnd_net_),
            .in3(N__5119),
            .lcout(sda_enable),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVeeprom.i2c.write_enable_132C_net ),
            .ce(N__4568),
            .sr(N__4505));
    defparam \eeprom.i2c.state_i0_i3_LC_22_14_0 .C_ON=1'b0;
    defparam \eeprom.i2c.state_i0_i3_LC_22_14_0 .SEQ_MODE=4'b1001;
    defparam \eeprom.i2c.state_i0_i3_LC_22_14_0 .LUT_INIT=16'b1000100000001010;
    LogicCell40 \eeprom.i2c.state_i0_i3_LC_22_14_0  (
            .in0(N__5261),
            .in1(N__4319),
            .in2(N__4313),
            .in3(N__5399),
            .lcout(\eeprom.state_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4956),
            .ce(N__5631),
            .sr(N__4577));
    defparam \eeprom.i2c.i1_2_lut_4_lut_LC_22_15_0 .C_ON=1'b0;
    defparam \eeprom.i2c.i1_2_lut_4_lut_LC_22_15_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.i2c.i1_2_lut_4_lut_LC_22_15_0 .LUT_INIT=16'b0010111100100010;
    LogicCell40 \eeprom.i2c.i1_2_lut_4_lut_LC_22_15_0  (
            .in0(N__4530),
            .in1(N__5498),
            .in2(N__5236),
            .in3(N__4516),
            .lcout(),
            .ltout(\eeprom.i2c.n39_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i2c.i1897_4_lut_4_lut_LC_22_15_1 .C_ON=1'b0;
    defparam \eeprom.i2c.i1897_4_lut_4_lut_LC_22_15_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.i2c.i1897_4_lut_4_lut_LC_22_15_1 .LUT_INIT=16'b1111000010110000;
    LogicCell40 \eeprom.i2c.i1897_4_lut_4_lut_LC_22_15_1  (
            .in0(N__4713),
            .in1(N__5200),
            .in2(N__4571),
            .in3(N__5067),
            .lcout(\eeprom.i2c.n952 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i2c.i1_4_lut_4_lut_LC_22_15_2 .C_ON=1'b0;
    defparam \eeprom.i2c.i1_4_lut_4_lut_LC_22_15_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.i2c.i1_4_lut_4_lut_LC_22_15_2 .LUT_INIT=16'b1000100011001000;
    LogicCell40 \eeprom.i2c.i1_4_lut_4_lut_LC_22_15_2  (
            .in0(N__5066),
            .in1(N__5193),
            .in2(N__5401),
            .in3(N__5499),
            .lcout(\eeprom.i2c.n16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i2c.i56_3_lut_LC_22_15_3 .C_ON=1'b0;
    defparam \eeprom.i2c.i56_3_lut_LC_22_15_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.i2c.i56_3_lut_LC_22_15_3 .LUT_INIT=16'b0011000000111100;
    LogicCell40 \eeprom.i2c.i56_3_lut_LC_22_15_3  (
            .in0(_gnd_net_),
            .in1(N__5496),
            .in2(N__5400),
            .in3(N__5064),
            .lcout(\eeprom.i2c.n33 ),
            .ltout(\eeprom.i2c.n33_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i2c.i1_2_lut_adj_13_LC_22_15_4 .C_ON=1'b0;
    defparam \eeprom.i2c.i1_2_lut_adj_13_LC_22_15_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.i2c.i1_2_lut_adj_13_LC_22_15_4 .LUT_INIT=16'b0000000011110000;
    LogicCell40 \eeprom.i2c.i1_2_lut_adj_13_LC_22_15_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__4556),
            .in3(N__5194),
            .lcout(),
            .ltout(\eeprom.i2c.n34_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i2c.i1891_4_lut_LC_22_15_5 .C_ON=1'b0;
    defparam \eeprom.i2c.i1891_4_lut_LC_22_15_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.i2c.i1891_4_lut_LC_22_15_5 .LUT_INIT=16'b0011000100110000;
    LogicCell40 \eeprom.i2c.i1891_4_lut_LC_22_15_5  (
            .in0(N__5500),
            .in1(N__4553),
            .in2(N__4547),
            .in3(N__4531),
            .lcout(\eeprom.i2c.n2616 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i2c.i57_3_lut_3_lut_LC_22_15_6 .C_ON=1'b0;
    defparam \eeprom.i2c.i57_3_lut_3_lut_LC_22_15_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.i2c.i57_3_lut_3_lut_LC_22_15_6 .LUT_INIT=16'b0111011101100110;
    LogicCell40 \eeprom.i2c.i57_3_lut_3_lut_LC_22_15_6  (
            .in0(N__5065),
            .in1(N__5356),
            .in2(_gnd_net_),
            .in3(N__5192),
            .lcout(\eeprom.i2c.n36 ),
            .ltout(\eeprom.i2c.n36_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i2c.i1_3_lut_4_lut_LC_22_15_7 .C_ON=1'b0;
    defparam \eeprom.i2c.i1_3_lut_4_lut_LC_22_15_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.i2c.i1_3_lut_4_lut_LC_22_15_7 .LUT_INIT=16'b0000000010111010;
    LogicCell40 \eeprom.i2c.i1_3_lut_4_lut_LC_22_15_7  (
            .in0(N__4517),
            .in1(N__5497),
            .in2(N__4508),
            .in3(N__5199),
            .lcout(\eeprom.i2c.n1493 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i2c.state_i0_i1_LC_22_16_2 .C_ON=1'b0;
    defparam \eeprom.i2c.state_i0_i1_LC_22_16_2 .SEQ_MODE=4'b1001;
    defparam \eeprom.i2c.state_i0_i1_LC_22_16_2 .LUT_INIT=16'b0001111100001111;
    LogicCell40 \eeprom.i2c.state_i0_i1_LC_22_16_2  (
            .in0(N__4697),
            .in1(N__4486),
            .in2(N__4463),
            .in3(N__4451),
            .lcout(\eeprom.state_1_adj_383 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4955),
            .ce(N__5632),
            .sr(N__4754));
    defparam \eeprom.i2c.i22_3_lut_3_lut_LC_22_16_4 .C_ON=1'b0;
    defparam \eeprom.i2c.i22_3_lut_3_lut_LC_22_16_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.i2c.i22_3_lut_3_lut_LC_22_16_4 .LUT_INIT=16'b0011001101000100;
    LogicCell40 \eeprom.i2c.i22_3_lut_3_lut_LC_22_16_4  (
            .in0(N__5195),
            .in1(N__5535),
            .in2(_gnd_net_),
            .in3(N__5360),
            .lcout(\eeprom.i2c.n11_adj_377 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i2c.equal_25_i10_2_lut_LC_22_17_5 .C_ON=1'b0;
    defparam \eeprom.i2c.equal_25_i10_2_lut_LC_22_17_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.i2c.equal_25_i10_2_lut_LC_22_17_5 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \eeprom.i2c.equal_25_i10_2_lut_LC_22_17_5  (
            .in0(_gnd_net_),
            .in1(N__5086),
            .in2(_gnd_net_),
            .in3(N__5562),
            .lcout(\eeprom.i2c.n10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i2c.state_7__I_0_140_i11_2_lut_4_lut_LC_22_18_1 .C_ON=1'b0;
    defparam \eeprom.i2c.state_7__I_0_140_i11_2_lut_4_lut_LC_22_18_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.i2c.state_7__I_0_140_i11_2_lut_4_lut_LC_22_18_1 .LUT_INIT=16'b1111111111011111;
    LogicCell40 \eeprom.i2c.state_7__I_0_140_i11_2_lut_4_lut_LC_22_18_1  (
            .in0(N__5415),
            .in1(N__5578),
            .in2(N__5279),
            .in3(N__5127),
            .lcout(\eeprom.i2c.n11_adj_378 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i2c.i1221_2_lut_LC_23_14_0 .C_ON=1'b0;
    defparam \eeprom.i2c.i1221_2_lut_LC_23_14_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.i2c.i1221_2_lut_LC_23_14_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \eeprom.i2c.i1221_2_lut_LC_23_14_0  (
            .in0(_gnd_net_),
            .in1(N__5257),
            .in2(_gnd_net_),
            .in3(N__5364),
            .lcout(\eeprom.i2c.n2018 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i2c.i4_4_lut_adj_12_LC_23_14_1 .C_ON=1'b0;
    defparam \eeprom.i2c.i4_4_lut_adj_12_LC_23_14_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.i2c.i4_4_lut_adj_12_LC_23_14_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \eeprom.i2c.i4_4_lut_adj_12_LC_23_14_1  (
            .in0(N__4687),
            .in1(N__4669),
            .in2(N__4652),
            .in3(N__4634),
            .lcout(),
            .ltout(\eeprom.i2c.n10_adj_380_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i2c.i5_3_lut_LC_23_14_2 .C_ON=1'b0;
    defparam \eeprom.i2c.i5_3_lut_LC_23_14_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.i2c.i5_3_lut_LC_23_14_2 .LUT_INIT=16'b1111111111111010;
    LogicCell40 \eeprom.i2c.i5_3_lut_LC_23_14_2  (
            .in0(N__4619),
            .in1(_gnd_net_),
            .in2(N__4604),
            .in3(N__4600),
            .lcout(\eeprom.i2c.n2654 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i2c.i1_2_lut_3_lut_2_lut_LC_23_14_3 .C_ON=1'b0;
    defparam \eeprom.i2c.i1_2_lut_3_lut_2_lut_LC_23_14_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.i2c.i1_2_lut_3_lut_2_lut_LC_23_14_3 .LUT_INIT=16'b1010101001010101;
    LogicCell40 \eeprom.i2c.i1_2_lut_3_lut_2_lut_LC_23_14_3  (
            .in0(N__5365),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5260),
            .lcout(\eeprom.i2c.n2726 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i2c.i1900_3_lut_4_lut_LC_23_14_4 .C_ON=1'b0;
    defparam \eeprom.i2c.i1900_3_lut_4_lut_LC_23_14_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.i2c.i1900_3_lut_4_lut_LC_23_14_4 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \eeprom.i2c.i1900_3_lut_4_lut_LC_23_14_4  (
            .in0(N__5125),
            .in1(N__5258),
            .in2(N__5633),
            .in3(N__5531),
            .lcout(\eeprom.i2c.n2706 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i2c.i2_3_lut_4_lut_LC_23_14_5 .C_ON=1'b0;
    defparam \eeprom.i2c.i2_3_lut_4_lut_LC_23_14_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.i2c.i2_3_lut_4_lut_LC_23_14_5 .LUT_INIT=16'b1111111111011111;
    LogicCell40 \eeprom.i2c.i2_3_lut_4_lut_LC_23_14_5  (
            .in0(N__5366),
            .in1(N__5259),
            .in2(N__5563),
            .in3(N__5123),
            .lcout(\eeprom.i2c.n11_adj_376 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i2c.i1_4_lut_2_lut_4_lut_LC_23_14_6 .C_ON=1'b0;
    defparam \eeprom.i2c.i1_4_lut_2_lut_4_lut_LC_23_14_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.i2c.i1_4_lut_2_lut_4_lut_LC_23_14_6 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \eeprom.i2c.i1_4_lut_2_lut_4_lut_LC_23_14_6  (
            .in0(N__5124),
            .in1(N__5530),
            .in2(_gnd_net_),
            .in3(N__5367),
            .lcout(\eeprom.i2c.n21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i2c.i1904_4_lut_LC_23_15_0 .C_ON=1'b0;
    defparam \eeprom.i2c.i1904_4_lut_LC_23_15_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.i2c.i1904_4_lut_LC_23_15_0 .LUT_INIT=16'b0011011100000000;
    LogicCell40 \eeprom.i2c.i1904_4_lut_LC_23_15_0  (
            .in0(N__5746),
            .in1(N__4747),
            .in2(N__5588),
            .in3(N__5625),
            .lcout(\eeprom.i2c.n2008 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i2c.i1264_3_lut_4_lut_LC_23_15_1 .C_ON=1'b0;
    defparam \eeprom.i2c.i1264_3_lut_4_lut_LC_23_15_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.i2c.i1264_3_lut_4_lut_LC_23_15_1 .LUT_INIT=16'b1111111110101011;
    LogicCell40 \eeprom.i2c.i1264_3_lut_4_lut_LC_23_15_1  (
            .in0(N__5524),
            .in1(N__5068),
            .in2(N__5237),
            .in3(N__5395),
            .lcout(),
            .ltout(\eeprom.i2c.n2063_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i2c.i1_4_lut_LC_23_15_2 .C_ON=1'b0;
    defparam \eeprom.i2c.i1_4_lut_LC_23_15_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.i2c.i1_4_lut_LC_23_15_2 .LUT_INIT=16'b0000111100001110;
    LogicCell40 \eeprom.i2c.i1_4_lut_LC_23_15_2  (
            .in0(N__4840),
            .in1(N__4829),
            .in2(N__4802),
            .in3(N__4799),
            .lcout(),
            .ltout(\eeprom.i2c.n1358_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i2c.i1888_4_lut_LC_23_15_3 .C_ON=1'b0;
    defparam \eeprom.i2c.i1888_4_lut_LC_23_15_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.i2c.i1888_4_lut_LC_23_15_3 .LUT_INIT=16'b0000010100000111;
    LogicCell40 \eeprom.i2c.i1888_4_lut_LC_23_15_3  (
            .in0(N__5526),
            .in1(N__5070),
            .in2(N__4769),
            .in3(N__5731),
            .lcout(\eeprom.i2c.n876 ),
            .ltout(\eeprom.i2c.n876_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i2c.i1913_4_lut_LC_23_15_4 .C_ON=1'b0;
    defparam \eeprom.i2c.i1913_4_lut_LC_23_15_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.i2c.i1913_4_lut_LC_23_15_4 .LUT_INIT=16'b0001000011110000;
    LogicCell40 \eeprom.i2c.i1913_4_lut_LC_23_15_4  (
            .in0(N__4766),
            .in1(N__5683),
            .in2(N__4757),
            .in3(N__4748),
            .lcout(\eeprom.i2c.n2078 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i2c.i1874_4_lut_LC_23_15_5 .C_ON=1'b0;
    defparam \eeprom.i2c.i1874_4_lut_LC_23_15_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.i2c.i1874_4_lut_LC_23_15_5 .LUT_INIT=16'b1111111111011111;
    LogicCell40 \eeprom.i2c.i1874_4_lut_LC_23_15_5  (
            .in0(N__4746),
            .in1(N__4736),
            .in2(N__5009),
            .in3(N__4730),
            .lcout(),
            .ltout(\eeprom.i2c.n2741_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i2c.state_i0_i0_LC_23_15_6 .C_ON=1'b0;
    defparam \eeprom.i2c.state_i0_i0_LC_23_15_6 .SEQ_MODE=4'b1000;
    defparam \eeprom.i2c.state_i0_i0_LC_23_15_6 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \eeprom.i2c.state_i0_i0_LC_23_15_6  (
            .in0(N__5396),
            .in1(_gnd_net_),
            .in2(N__4721),
            .in3(N__5626),
            .lcout(state_0_adj_386),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4973),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i2c.state_7__I_0_141_i10_2_lut_LC_23_15_7 .C_ON=1'b0;
    defparam \eeprom.i2c.state_7__I_0_141_i10_2_lut_LC_23_15_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.i2c.state_7__I_0_141_i10_2_lut_LC_23_15_7 .LUT_INIT=16'b1011101110111011;
    LogicCell40 \eeprom.i2c.state_7__I_0_141_i10_2_lut_LC_23_15_7  (
            .in0(N__5525),
            .in1(N__5069),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\eeprom.i2c.n10_adj_379 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i2c.state_i0_i2_LC_23_16_0 .C_ON=1'b0;
    defparam \eeprom.i2c.state_i0_i2_LC_23_16_0 .SEQ_MODE=4'b1001;
    defparam \eeprom.i2c.state_i0_i2_LC_23_16_0 .LUT_INIT=16'b0000001000001010;
    LogicCell40 \eeprom.i2c.state_i0_i2_LC_23_16_0  (
            .in0(N__5732),
            .in1(N__5713),
            .in2(N__5684),
            .in3(N__5657),
            .lcout(\eeprom.state_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4976),
            .ce(N__5630),
            .sr(N__5597));
    defparam \eeprom.i2c.i2c_scl_enable_124_LC_23_17_6 .C_ON=1'b0;
    defparam \eeprom.i2c.i2c_scl_enable_124_LC_23_17_6 .SEQ_MODE=4'b1000;
    defparam \eeprom.i2c.i2c_scl_enable_124_LC_23_17_6 .LUT_INIT=16'b1111111111111000;
    LogicCell40 \eeprom.i2c.i2c_scl_enable_124_LC_23_17_6  (
            .in0(N__5569),
            .in1(N__5414),
            .in2(N__5262),
            .in3(N__5097),
            .lcout(scl_enable),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVeeprom.i2c.i2c_scl_enable_124C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i2c.state_7__I_0_139_i9_2_lut_LC_24_14_1 .C_ON=1'b0;
    defparam \eeprom.i2c.state_7__I_0_139_i9_2_lut_LC_24_14_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.i2c.state_7__I_0_139_i9_2_lut_LC_24_14_1 .LUT_INIT=16'b1100110011111111;
    LogicCell40 \eeprom.i2c.state_7__I_0_139_i9_2_lut_LC_24_14_1  (
            .in0(_gnd_net_),
            .in1(N__5397),
            .in2(_gnd_net_),
            .in3(N__5277),
            .lcout(\eeprom.i2c.n9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i2c.state_7__I_0_139_i11_2_lut_4_lut_LC_24_14_4 .C_ON=1'b0;
    defparam \eeprom.i2c.state_7__I_0_139_i11_2_lut_4_lut_LC_24_14_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.i2c.state_7__I_0_139_i11_2_lut_4_lut_LC_24_14_4 .LUT_INIT=16'b1111111111101111;
    LogicCell40 \eeprom.i2c.state_7__I_0_139_i11_2_lut_4_lut_LC_24_14_4  (
            .in0(N__5564),
            .in1(N__5398),
            .in2(N__5282),
            .in3(N__5126),
            .lcout(\eeprom.i2c.n11_adj_382 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i2c.i1198_2_lut_LC_26_17_2 .C_ON=1'b0;
    defparam \eeprom.i2c.i1198_2_lut_LC_26_17_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.i2c.i1198_2_lut_LC_26_17_2 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \eeprom.i2c.i1198_2_lut_LC_26_17_2  (
            .in0(N__4990),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4972),
            .lcout(scl_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
endmodule // TinyFPGA_B
