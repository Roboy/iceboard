-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2017.08.27940

-- Build Date:         Sep 12 2017 08:26:01

-- File Generated:     Jan 31 2020 00:08:55

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "TinyFPGA_B" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of TinyFPGA_B
entity TinyFPGA_B is
port (
    USBPU : out std_logic;
    TX : out std_logic;
    SDA : inout std_logic;
    SCL : inout std_logic;
    RX : in std_logic;
    NEOPXL : out std_logic;
    LED : out std_logic;
    INLC : out std_logic;
    INLB : out std_logic;
    INLA : out std_logic;
    INHC : out std_logic;
    INHB : out std_logic;
    INHA : out std_logic;
    HALL3 : in std_logic;
    HALL2 : in std_logic;
    HALL1 : in std_logic;
    FAULT_N : in std_logic;
    ENCODER1_B : in std_logic;
    ENCODER1_A : in std_logic;
    ENCODER0_B : in std_logic;
    ENCODER0_A : in std_logic;
    DE : out std_logic;
    CS_MISO : in std_logic;
    CS_CLK : out std_logic;
    CS : out std_logic;
    CLK : in std_logic);
end TinyFPGA_B;

-- Architecture of TinyFPGA_B
-- View name is \INTERFACE\
architecture \INTERFACE\ of TinyFPGA_B is

signal \N__6937\ : std_logic;
signal \N__6936\ : std_logic;
signal \N__6935\ : std_logic;
signal \N__6928\ : std_logic;
signal \N__6927\ : std_logic;
signal \N__6926\ : std_logic;
signal \N__6919\ : std_logic;
signal \N__6918\ : std_logic;
signal \N__6917\ : std_logic;
signal \N__6910\ : std_logic;
signal \N__6909\ : std_logic;
signal \N__6908\ : std_logic;
signal \N__6901\ : std_logic;
signal \N__6900\ : std_logic;
signal \N__6899\ : std_logic;
signal \N__6892\ : std_logic;
signal \N__6891\ : std_logic;
signal \N__6890\ : std_logic;
signal \N__6883\ : std_logic;
signal \N__6882\ : std_logic;
signal \N__6881\ : std_logic;
signal \N__6874\ : std_logic;
signal \N__6873\ : std_logic;
signal \N__6872\ : std_logic;
signal \N__6865\ : std_logic;
signal \N__6864\ : std_logic;
signal \N__6863\ : std_logic;
signal \N__6856\ : std_logic;
signal \N__6855\ : std_logic;
signal \N__6854\ : std_logic;
signal \N__6847\ : std_logic;
signal \N__6846\ : std_logic;
signal \N__6845\ : std_logic;
signal \N__6838\ : std_logic;
signal \N__6837\ : std_logic;
signal \N__6836\ : std_logic;
signal \N__6829\ : std_logic;
signal \N__6828\ : std_logic;
signal \N__6827\ : std_logic;
signal \N__6820\ : std_logic;
signal \N__6819\ : std_logic;
signal \N__6818\ : std_logic;
signal \N__6811\ : std_logic;
signal \N__6810\ : std_logic;
signal \N__6809\ : std_logic;
signal \N__6802\ : std_logic;
signal \N__6801\ : std_logic;
signal \N__6800\ : std_logic;
signal \N__6783\ : std_logic;
signal \N__6782\ : std_logic;
signal \N__6779\ : std_logic;
signal \N__6776\ : std_logic;
signal \N__6773\ : std_logic;
signal \N__6768\ : std_logic;
signal \N__6765\ : std_logic;
signal \N__6762\ : std_logic;
signal \N__6761\ : std_logic;
signal \N__6758\ : std_logic;
signal \N__6755\ : std_logic;
signal \N__6750\ : std_logic;
signal \N__6749\ : std_logic;
signal \N__6748\ : std_logic;
signal \N__6747\ : std_logic;
signal \N__6746\ : std_logic;
signal \N__6745\ : std_logic;
signal \N__6744\ : std_logic;
signal \N__6743\ : std_logic;
signal \N__6742\ : std_logic;
signal \N__6741\ : std_logic;
signal \N__6740\ : std_logic;
signal \N__6739\ : std_logic;
signal \N__6738\ : std_logic;
signal \N__6737\ : std_logic;
signal \N__6736\ : std_logic;
signal \N__6735\ : std_logic;
signal \N__6734\ : std_logic;
signal \N__6733\ : std_logic;
signal \N__6732\ : std_logic;
signal \N__6693\ : std_logic;
signal \N__6690\ : std_logic;
signal \N__6687\ : std_logic;
signal \N__6684\ : std_logic;
signal \N__6681\ : std_logic;
signal \N__6680\ : std_logic;
signal \N__6677\ : std_logic;
signal \N__6674\ : std_logic;
signal \N__6669\ : std_logic;
signal \N__6666\ : std_logic;
signal \N__6665\ : std_logic;
signal \N__6662\ : std_logic;
signal \N__6659\ : std_logic;
signal \N__6658\ : std_logic;
signal \N__6657\ : std_logic;
signal \N__6652\ : std_logic;
signal \N__6651\ : std_logic;
signal \N__6648\ : std_logic;
signal \N__6645\ : std_logic;
signal \N__6642\ : std_logic;
signal \N__6639\ : std_logic;
signal \N__6630\ : std_logic;
signal \N__6629\ : std_logic;
signal \N__6626\ : std_logic;
signal \N__6623\ : std_logic;
signal \N__6620\ : std_logic;
signal \N__6617\ : std_logic;
signal \N__6614\ : std_logic;
signal \N__6611\ : std_logic;
signal \N__6606\ : std_logic;
signal \N__6603\ : std_logic;
signal \N__6600\ : std_logic;
signal \N__6599\ : std_logic;
signal \N__6596\ : std_logic;
signal \N__6593\ : std_logic;
signal \N__6590\ : std_logic;
signal \N__6587\ : std_logic;
signal \N__6582\ : std_logic;
signal \N__6581\ : std_logic;
signal \N__6580\ : std_logic;
signal \N__6579\ : std_logic;
signal \N__6576\ : std_logic;
signal \N__6575\ : std_logic;
signal \N__6572\ : std_logic;
signal \N__6571\ : std_logic;
signal \N__6568\ : std_logic;
signal \N__6567\ : std_logic;
signal \N__6566\ : std_logic;
signal \N__6551\ : std_logic;
signal \N__6548\ : std_logic;
signal \N__6543\ : std_logic;
signal \N__6540\ : std_logic;
signal \N__6537\ : std_logic;
signal \N__6534\ : std_logic;
signal \N__6531\ : std_logic;
signal \N__6528\ : std_logic;
signal \N__6525\ : std_logic;
signal \N__6522\ : std_logic;
signal \N__6519\ : std_logic;
signal \N__6518\ : std_logic;
signal \N__6515\ : std_logic;
signal \N__6512\ : std_logic;
signal \N__6507\ : std_logic;
signal \N__6504\ : std_logic;
signal \N__6501\ : std_logic;
signal \N__6498\ : std_logic;
signal \N__6495\ : std_logic;
signal \N__6492\ : std_logic;
signal \N__6489\ : std_logic;
signal \N__6486\ : std_logic;
signal \N__6483\ : std_logic;
signal \N__6482\ : std_logic;
signal \N__6479\ : std_logic;
signal \N__6478\ : std_logic;
signal \N__6477\ : std_logic;
signal \N__6476\ : std_logic;
signal \N__6475\ : std_logic;
signal \N__6472\ : std_logic;
signal \N__6469\ : std_logic;
signal \N__6466\ : std_logic;
signal \N__6463\ : std_logic;
signal \N__6460\ : std_logic;
signal \N__6459\ : std_logic;
signal \N__6458\ : std_logic;
signal \N__6455\ : std_logic;
signal \N__6452\ : std_logic;
signal \N__6447\ : std_logic;
signal \N__6446\ : std_logic;
signal \N__6443\ : std_logic;
signal \N__6440\ : std_logic;
signal \N__6437\ : std_logic;
signal \N__6436\ : std_logic;
signal \N__6433\ : std_logic;
signal \N__6432\ : std_logic;
signal \N__6431\ : std_logic;
signal \N__6428\ : std_logic;
signal \N__6427\ : std_logic;
signal \N__6424\ : std_logic;
signal \N__6421\ : std_logic;
signal \N__6418\ : std_logic;
signal \N__6415\ : std_logic;
signal \N__6410\ : std_logic;
signal \N__6407\ : std_logic;
signal \N__6404\ : std_logic;
signal \N__6401\ : std_logic;
signal \N__6398\ : std_logic;
signal \N__6395\ : std_logic;
signal \N__6392\ : std_logic;
signal \N__6391\ : std_logic;
signal \N__6384\ : std_logic;
signal \N__6381\ : std_logic;
signal \N__6378\ : std_logic;
signal \N__6369\ : std_logic;
signal \N__6368\ : std_logic;
signal \N__6367\ : std_logic;
signal \N__6362\ : std_logic;
signal \N__6359\ : std_logic;
signal \N__6356\ : std_logic;
signal \N__6349\ : std_logic;
signal \N__6346\ : std_logic;
signal \N__6343\ : std_logic;
signal \N__6330\ : std_logic;
signal \N__6327\ : std_logic;
signal \N__6326\ : std_logic;
signal \N__6323\ : std_logic;
signal \N__6320\ : std_logic;
signal \N__6317\ : std_logic;
signal \N__6314\ : std_logic;
signal \N__6311\ : std_logic;
signal \N__6308\ : std_logic;
signal \N__6303\ : std_logic;
signal \N__6300\ : std_logic;
signal \N__6297\ : std_logic;
signal \N__6294\ : std_logic;
signal \N__6293\ : std_logic;
signal \N__6290\ : std_logic;
signal \N__6287\ : std_logic;
signal \N__6282\ : std_logic;
signal \N__6279\ : std_logic;
signal \N__6276\ : std_logic;
signal \N__6273\ : std_logic;
signal \N__6270\ : std_logic;
signal \N__6267\ : std_logic;
signal \N__6264\ : std_logic;
signal \N__6261\ : std_logic;
signal \N__6258\ : std_logic;
signal \N__6255\ : std_logic;
signal \N__6252\ : std_logic;
signal \N__6249\ : std_logic;
signal \N__6248\ : std_logic;
signal \N__6245\ : std_logic;
signal \N__6242\ : std_logic;
signal \N__6237\ : std_logic;
signal \N__6236\ : std_logic;
signal \N__6233\ : std_logic;
signal \N__6230\ : std_logic;
signal \N__6229\ : std_logic;
signal \N__6228\ : std_logic;
signal \N__6221\ : std_logic;
signal \N__6218\ : std_logic;
signal \N__6215\ : std_logic;
signal \N__6214\ : std_logic;
signal \N__6211\ : std_logic;
signal \N__6210\ : std_logic;
signal \N__6207\ : std_logic;
signal \N__6204\ : std_logic;
signal \N__6201\ : std_logic;
signal \N__6198\ : std_logic;
signal \N__6189\ : std_logic;
signal \N__6188\ : std_logic;
signal \N__6187\ : std_logic;
signal \N__6186\ : std_logic;
signal \N__6179\ : std_logic;
signal \N__6178\ : std_logic;
signal \N__6175\ : std_logic;
signal \N__6172\ : std_logic;
signal \N__6169\ : std_logic;
signal \N__6166\ : std_logic;
signal \N__6165\ : std_logic;
signal \N__6162\ : std_logic;
signal \N__6159\ : std_logic;
signal \N__6156\ : std_logic;
signal \N__6153\ : std_logic;
signal \N__6144\ : std_logic;
signal \N__6141\ : std_logic;
signal \N__6140\ : std_logic;
signal \N__6139\ : std_logic;
signal \N__6136\ : std_logic;
signal \N__6131\ : std_logic;
signal \N__6126\ : std_logic;
signal \N__6125\ : std_logic;
signal \N__6122\ : std_logic;
signal \N__6121\ : std_logic;
signal \N__6118\ : std_logic;
signal \N__6117\ : std_logic;
signal \N__6116\ : std_logic;
signal \N__6113\ : std_logic;
signal \N__6110\ : std_logic;
signal \N__6107\ : std_logic;
signal \N__6106\ : std_logic;
signal \N__6105\ : std_logic;
signal \N__6102\ : std_logic;
signal \N__6101\ : std_logic;
signal \N__6098\ : std_logic;
signal \N__6097\ : std_logic;
signal \N__6096\ : std_logic;
signal \N__6095\ : std_logic;
signal \N__6094\ : std_logic;
signal \N__6089\ : std_logic;
signal \N__6086\ : std_logic;
signal \N__6083\ : std_logic;
signal \N__6080\ : std_logic;
signal \N__6077\ : std_logic;
signal \N__6076\ : std_logic;
signal \N__6075\ : std_logic;
signal \N__6074\ : std_logic;
signal \N__6071\ : std_logic;
signal \N__6070\ : std_logic;
signal \N__6067\ : std_logic;
signal \N__6060\ : std_logic;
signal \N__6059\ : std_logic;
signal \N__6058\ : std_logic;
signal \N__6057\ : std_logic;
signal \N__6056\ : std_logic;
signal \N__6055\ : std_logic;
signal \N__6052\ : std_logic;
signal \N__6049\ : std_logic;
signal \N__6040\ : std_logic;
signal \N__6033\ : std_logic;
signal \N__6028\ : std_logic;
signal \N__6023\ : std_logic;
signal \N__6020\ : std_logic;
signal \N__6011\ : std_logic;
signal \N__5994\ : std_logic;
signal \N__5993\ : std_logic;
signal \N__5990\ : std_logic;
signal \N__5989\ : std_logic;
signal \N__5988\ : std_logic;
signal \N__5987\ : std_logic;
signal \N__5984\ : std_logic;
signal \N__5981\ : std_logic;
signal \N__5976\ : std_logic;
signal \N__5975\ : std_logic;
signal \N__5972\ : std_logic;
signal \N__5971\ : std_logic;
signal \N__5968\ : std_logic;
signal \N__5967\ : std_logic;
signal \N__5966\ : std_logic;
signal \N__5961\ : std_logic;
signal \N__5960\ : std_logic;
signal \N__5959\ : std_logic;
signal \N__5958\ : std_logic;
signal \N__5957\ : std_logic;
signal \N__5954\ : std_logic;
signal \N__5953\ : std_logic;
signal \N__5952\ : std_logic;
signal \N__5951\ : std_logic;
signal \N__5950\ : std_logic;
signal \N__5949\ : std_logic;
signal \N__5948\ : std_logic;
signal \N__5945\ : std_logic;
signal \N__5942\ : std_logic;
signal \N__5939\ : std_logic;
signal \N__5934\ : std_logic;
signal \N__5931\ : std_logic;
signal \N__5926\ : std_logic;
signal \N__5915\ : std_logic;
signal \N__5912\ : std_logic;
signal \N__5909\ : std_logic;
signal \N__5904\ : std_logic;
signal \N__5883\ : std_logic;
signal \N__5882\ : std_logic;
signal \N__5881\ : std_logic;
signal \N__5880\ : std_logic;
signal \N__5877\ : std_logic;
signal \N__5876\ : std_logic;
signal \N__5875\ : std_logic;
signal \N__5874\ : std_logic;
signal \N__5871\ : std_logic;
signal \N__5868\ : std_logic;
signal \N__5867\ : std_logic;
signal \N__5866\ : std_logic;
signal \N__5863\ : std_logic;
signal \N__5860\ : std_logic;
signal \N__5859\ : std_logic;
signal \N__5858\ : std_logic;
signal \N__5853\ : std_logic;
signal \N__5852\ : std_logic;
signal \N__5851\ : std_logic;
signal \N__5848\ : std_logic;
signal \N__5847\ : std_logic;
signal \N__5846\ : std_logic;
signal \N__5845\ : std_logic;
signal \N__5842\ : std_logic;
signal \N__5839\ : std_logic;
signal \N__5836\ : std_logic;
signal \N__5835\ : std_logic;
signal \N__5832\ : std_logic;
signal \N__5829\ : std_logic;
signal \N__5826\ : std_logic;
signal \N__5823\ : std_logic;
signal \N__5820\ : std_logic;
signal \N__5817\ : std_logic;
signal \N__5808\ : std_logic;
signal \N__5805\ : std_logic;
signal \N__5804\ : std_logic;
signal \N__5803\ : std_logic;
signal \N__5802\ : std_logic;
signal \N__5801\ : std_logic;
signal \N__5798\ : std_logic;
signal \N__5797\ : std_logic;
signal \N__5792\ : std_logic;
signal \N__5789\ : std_logic;
signal \N__5786\ : std_logic;
signal \N__5783\ : std_logic;
signal \N__5778\ : std_logic;
signal \N__5775\ : std_logic;
signal \N__5766\ : std_logic;
signal \N__5761\ : std_logic;
signal \N__5758\ : std_logic;
signal \N__5751\ : std_logic;
signal \N__5730\ : std_logic;
signal \N__5729\ : std_logic;
signal \N__5728\ : std_logic;
signal \N__5727\ : std_logic;
signal \N__5726\ : std_logic;
signal \N__5725\ : std_logic;
signal \N__5724\ : std_logic;
signal \N__5723\ : std_logic;
signal \N__5718\ : std_logic;
signal \N__5715\ : std_logic;
signal \N__5710\ : std_logic;
signal \N__5709\ : std_logic;
signal \N__5706\ : std_logic;
signal \N__5705\ : std_logic;
signal \N__5704\ : std_logic;
signal \N__5703\ : std_logic;
signal \N__5702\ : std_logic;
signal \N__5701\ : std_logic;
signal \N__5700\ : std_logic;
signal \N__5697\ : std_logic;
signal \N__5694\ : std_logic;
signal \N__5691\ : std_logic;
signal \N__5690\ : std_logic;
signal \N__5689\ : std_logic;
signal \N__5688\ : std_logic;
signal \N__5683\ : std_logic;
signal \N__5680\ : std_logic;
signal \N__5677\ : std_logic;
signal \N__5666\ : std_logic;
signal \N__5665\ : std_logic;
signal \N__5664\ : std_logic;
signal \N__5663\ : std_logic;
signal \N__5660\ : std_logic;
signal \N__5657\ : std_logic;
signal \N__5652\ : std_logic;
signal \N__5649\ : std_logic;
signal \N__5644\ : std_logic;
signal \N__5641\ : std_logic;
signal \N__5634\ : std_logic;
signal \N__5627\ : std_logic;
signal \N__5610\ : std_logic;
signal \N__5609\ : std_logic;
signal \N__5606\ : std_logic;
signal \N__5603\ : std_logic;
signal \N__5598\ : std_logic;
signal \N__5595\ : std_logic;
signal \N__5594\ : std_logic;
signal \N__5591\ : std_logic;
signal \N__5588\ : std_logic;
signal \N__5583\ : std_logic;
signal \N__5580\ : std_logic;
signal \N__5579\ : std_logic;
signal \N__5576\ : std_logic;
signal \N__5573\ : std_logic;
signal \N__5568\ : std_logic;
signal \N__5565\ : std_logic;
signal \N__5564\ : std_logic;
signal \N__5561\ : std_logic;
signal \N__5558\ : std_logic;
signal \N__5553\ : std_logic;
signal \N__5550\ : std_logic;
signal \N__5547\ : std_logic;
signal \N__5544\ : std_logic;
signal \N__5541\ : std_logic;
signal \N__5540\ : std_logic;
signal \N__5537\ : std_logic;
signal \N__5534\ : std_logic;
signal \N__5533\ : std_logic;
signal \N__5532\ : std_logic;
signal \N__5531\ : std_logic;
signal \N__5530\ : std_logic;
signal \N__5527\ : std_logic;
signal \N__5524\ : std_logic;
signal \N__5523\ : std_logic;
signal \N__5520\ : std_logic;
signal \N__5517\ : std_logic;
signal \N__5514\ : std_logic;
signal \N__5513\ : std_logic;
signal \N__5510\ : std_logic;
signal \N__5507\ : std_logic;
signal \N__5504\ : std_logic;
signal \N__5501\ : std_logic;
signal \N__5496\ : std_logic;
signal \N__5493\ : std_logic;
signal \N__5490\ : std_logic;
signal \N__5487\ : std_logic;
signal \N__5472\ : std_logic;
signal \N__5469\ : std_logic;
signal \N__5468\ : std_logic;
signal \N__5465\ : std_logic;
signal \N__5462\ : std_logic;
signal \N__5457\ : std_logic;
signal \N__5454\ : std_logic;
signal \N__5453\ : std_logic;
signal \N__5450\ : std_logic;
signal \N__5447\ : std_logic;
signal \N__5446\ : std_logic;
signal \N__5445\ : std_logic;
signal \N__5444\ : std_logic;
signal \N__5443\ : std_logic;
signal \N__5442\ : std_logic;
signal \N__5439\ : std_logic;
signal \N__5436\ : std_logic;
signal \N__5433\ : std_logic;
signal \N__5432\ : std_logic;
signal \N__5429\ : std_logic;
signal \N__5426\ : std_logic;
signal \N__5423\ : std_logic;
signal \N__5422\ : std_logic;
signal \N__5419\ : std_logic;
signal \N__5418\ : std_logic;
signal \N__5415\ : std_logic;
signal \N__5412\ : std_logic;
signal \N__5411\ : std_logic;
signal \N__5410\ : std_logic;
signal \N__5405\ : std_logic;
signal \N__5400\ : std_logic;
signal \N__5397\ : std_logic;
signal \N__5392\ : std_logic;
signal \N__5389\ : std_logic;
signal \N__5386\ : std_logic;
signal \N__5383\ : std_logic;
signal \N__5380\ : std_logic;
signal \N__5377\ : std_logic;
signal \N__5366\ : std_logic;
signal \N__5363\ : std_logic;
signal \N__5356\ : std_logic;
signal \N__5353\ : std_logic;
signal \N__5348\ : std_logic;
signal \N__5343\ : std_logic;
signal \N__5342\ : std_logic;
signal \N__5341\ : std_logic;
signal \N__5338\ : std_logic;
signal \N__5337\ : std_logic;
signal \N__5332\ : std_logic;
signal \N__5329\ : std_logic;
signal \N__5326\ : std_logic;
signal \N__5323\ : std_logic;
signal \N__5320\ : std_logic;
signal \N__5317\ : std_logic;
signal \N__5310\ : std_logic;
signal \N__5307\ : std_logic;
signal \N__5304\ : std_logic;
signal \N__5303\ : std_logic;
signal \N__5300\ : std_logic;
signal \N__5297\ : std_logic;
signal \N__5292\ : std_logic;
signal \N__5291\ : std_logic;
signal \N__5288\ : std_logic;
signal \N__5285\ : std_logic;
signal \N__5280\ : std_logic;
signal \N__5277\ : std_logic;
signal \N__5276\ : std_logic;
signal \N__5273\ : std_logic;
signal \N__5270\ : std_logic;
signal \N__5265\ : std_logic;
signal \N__5264\ : std_logic;
signal \N__5261\ : std_logic;
signal \N__5258\ : std_logic;
signal \N__5255\ : std_logic;
signal \N__5252\ : std_logic;
signal \N__5247\ : std_logic;
signal \N__5246\ : std_logic;
signal \N__5243\ : std_logic;
signal \N__5240\ : std_logic;
signal \N__5235\ : std_logic;
signal \N__5234\ : std_logic;
signal \N__5233\ : std_logic;
signal \N__5232\ : std_logic;
signal \N__5229\ : std_logic;
signal \N__5226\ : std_logic;
signal \N__5221\ : std_logic;
signal \N__5214\ : std_logic;
signal \N__5211\ : std_logic;
signal \N__5210\ : std_logic;
signal \N__5209\ : std_logic;
signal \N__5208\ : std_logic;
signal \N__5205\ : std_logic;
signal \N__5202\ : std_logic;
signal \N__5197\ : std_logic;
signal \N__5192\ : std_logic;
signal \N__5191\ : std_logic;
signal \N__5190\ : std_logic;
signal \N__5189\ : std_logic;
signal \N__5188\ : std_logic;
signal \N__5187\ : std_logic;
signal \N__5186\ : std_logic;
signal \N__5183\ : std_logic;
signal \N__5180\ : std_logic;
signal \N__5177\ : std_logic;
signal \N__5166\ : std_logic;
signal \N__5163\ : std_logic;
signal \N__5154\ : std_logic;
signal \N__5153\ : std_logic;
signal \N__5152\ : std_logic;
signal \N__5151\ : std_logic;
signal \N__5150\ : std_logic;
signal \N__5149\ : std_logic;
signal \N__5146\ : std_logic;
signal \N__5143\ : std_logic;
signal \N__5134\ : std_logic;
signal \N__5133\ : std_logic;
signal \N__5130\ : std_logic;
signal \N__5127\ : std_logic;
signal \N__5126\ : std_logic;
signal \N__5125\ : std_logic;
signal \N__5124\ : std_logic;
signal \N__5123\ : std_logic;
signal \N__5122\ : std_logic;
signal \N__5121\ : std_logic;
signal \N__5118\ : std_logic;
signal \N__5115\ : std_logic;
signal \N__5112\ : std_logic;
signal \N__5109\ : std_logic;
signal \N__5096\ : std_logic;
signal \N__5093\ : std_logic;
signal \N__5082\ : std_logic;
signal \N__5079\ : std_logic;
signal \N__5076\ : std_logic;
signal \N__5073\ : std_logic;
signal \N__5072\ : std_logic;
signal \N__5069\ : std_logic;
signal \N__5066\ : std_logic;
signal \N__5063\ : std_logic;
signal \N__5058\ : std_logic;
signal \N__5055\ : std_logic;
signal \N__5052\ : std_logic;
signal \N__5049\ : std_logic;
signal \N__5046\ : std_logic;
signal \N__5043\ : std_logic;
signal \N__5040\ : std_logic;
signal \N__5037\ : std_logic;
signal \N__5034\ : std_logic;
signal \N__5033\ : std_logic;
signal \N__5030\ : std_logic;
signal \N__5027\ : std_logic;
signal \N__5022\ : std_logic;
signal \N__5021\ : std_logic;
signal \N__5018\ : std_logic;
signal \N__5017\ : std_logic;
signal \N__5014\ : std_logic;
signal \N__5011\ : std_logic;
signal \N__5008\ : std_logic;
signal \N__5007\ : std_logic;
signal \N__5006\ : std_logic;
signal \N__5001\ : std_logic;
signal \N__4998\ : std_logic;
signal \N__4995\ : std_logic;
signal \N__4992\ : std_logic;
signal \N__4991\ : std_logic;
signal \N__4986\ : std_logic;
signal \N__4981\ : std_logic;
signal \N__4978\ : std_logic;
signal \N__4971\ : std_logic;
signal \N__4968\ : std_logic;
signal \N__4965\ : std_logic;
signal \N__4962\ : std_logic;
signal \N__4959\ : std_logic;
signal \N__4958\ : std_logic;
signal \N__4957\ : std_logic;
signal \N__4950\ : std_logic;
signal \N__4947\ : std_logic;
signal \N__4944\ : std_logic;
signal \N__4943\ : std_logic;
signal \N__4940\ : std_logic;
signal \N__4937\ : std_logic;
signal \N__4936\ : std_logic;
signal \N__4935\ : std_logic;
signal \N__4934\ : std_logic;
signal \N__4929\ : std_logic;
signal \N__4924\ : std_logic;
signal \N__4921\ : std_logic;
signal \N__4918\ : std_logic;
signal \N__4915\ : std_logic;
signal \N__4908\ : std_logic;
signal \N__4905\ : std_logic;
signal \N__4902\ : std_logic;
signal \N__4901\ : std_logic;
signal \N__4900\ : std_logic;
signal \N__4897\ : std_logic;
signal \N__4894\ : std_logic;
signal \N__4891\ : std_logic;
signal \N__4888\ : std_logic;
signal \N__4885\ : std_logic;
signal \N__4882\ : std_logic;
signal \N__4875\ : std_logic;
signal \N__4872\ : std_logic;
signal \N__4869\ : std_logic;
signal \N__4868\ : std_logic;
signal \N__4865\ : std_logic;
signal \N__4862\ : std_logic;
signal \N__4857\ : std_logic;
signal \N__4854\ : std_logic;
signal \N__4851\ : std_logic;
signal \N__4850\ : std_logic;
signal \N__4847\ : std_logic;
signal \N__4844\ : std_logic;
signal \N__4843\ : std_logic;
signal \N__4842\ : std_logic;
signal \N__4839\ : std_logic;
signal \N__4836\ : std_logic;
signal \N__4833\ : std_logic;
signal \N__4830\ : std_logic;
signal \N__4821\ : std_logic;
signal \N__4818\ : std_logic;
signal \N__4817\ : std_logic;
signal \N__4814\ : std_logic;
signal \N__4811\ : std_logic;
signal \N__4806\ : std_logic;
signal \N__4805\ : std_logic;
signal \N__4802\ : std_logic;
signal \N__4799\ : std_logic;
signal \N__4796\ : std_logic;
signal \N__4791\ : std_logic;
signal \N__4790\ : std_logic;
signal \N__4789\ : std_logic;
signal \N__4786\ : std_logic;
signal \N__4783\ : std_logic;
signal \N__4780\ : std_logic;
signal \N__4773\ : std_logic;
signal \N__4770\ : std_logic;
signal \N__4767\ : std_logic;
signal \N__4766\ : std_logic;
signal \N__4763\ : std_logic;
signal \N__4760\ : std_logic;
signal \N__4755\ : std_logic;
signal \N__4752\ : std_logic;
signal \N__4751\ : std_logic;
signal \N__4750\ : std_logic;
signal \N__4749\ : std_logic;
signal \N__4746\ : std_logic;
signal \N__4743\ : std_logic;
signal \N__4740\ : std_logic;
signal \N__4737\ : std_logic;
signal \N__4736\ : std_logic;
signal \N__4733\ : std_logic;
signal \N__4730\ : std_logic;
signal \N__4727\ : std_logic;
signal \N__4724\ : std_logic;
signal \N__4721\ : std_logic;
signal \N__4720\ : std_logic;
signal \N__4719\ : std_logic;
signal \N__4716\ : std_logic;
signal \N__4709\ : std_logic;
signal \N__4706\ : std_logic;
signal \N__4703\ : std_logic;
signal \N__4700\ : std_logic;
signal \N__4689\ : std_logic;
signal \N__4686\ : std_logic;
signal \N__4683\ : std_logic;
signal \N__4680\ : std_logic;
signal \N__4677\ : std_logic;
signal \N__4674\ : std_logic;
signal \N__4671\ : std_logic;
signal \N__4670\ : std_logic;
signal \N__4667\ : std_logic;
signal \N__4664\ : std_logic;
signal \N__4661\ : std_logic;
signal \N__4658\ : std_logic;
signal \N__4653\ : std_logic;
signal \N__4650\ : std_logic;
signal \N__4647\ : std_logic;
signal \N__4644\ : std_logic;
signal \N__4641\ : std_logic;
signal \N__4638\ : std_logic;
signal \N__4637\ : std_logic;
signal \N__4634\ : std_logic;
signal \N__4631\ : std_logic;
signal \N__4626\ : std_logic;
signal \N__4623\ : std_logic;
signal \N__4620\ : std_logic;
signal \N__4617\ : std_logic;
signal \N__4614\ : std_logic;
signal \N__4613\ : std_logic;
signal \N__4610\ : std_logic;
signal \N__4607\ : std_logic;
signal \N__4602\ : std_logic;
signal \N__4599\ : std_logic;
signal \N__4596\ : std_logic;
signal \N__4593\ : std_logic;
signal \N__4590\ : std_logic;
signal \N__4589\ : std_logic;
signal \N__4586\ : std_logic;
signal \N__4583\ : std_logic;
signal \N__4580\ : std_logic;
signal \N__4577\ : std_logic;
signal \N__4572\ : std_logic;
signal \N__4569\ : std_logic;
signal \N__4566\ : std_logic;
signal \N__4563\ : std_logic;
signal \N__4560\ : std_logic;
signal \N__4559\ : std_logic;
signal \N__4558\ : std_logic;
signal \N__4555\ : std_logic;
signal \N__4552\ : std_logic;
signal \N__4549\ : std_logic;
signal \N__4546\ : std_logic;
signal \N__4541\ : std_logic;
signal \N__4538\ : std_logic;
signal \N__4533\ : std_logic;
signal \N__4530\ : std_logic;
signal \N__4527\ : std_logic;
signal \N__4524\ : std_logic;
signal \N__4521\ : std_logic;
signal \N__4518\ : std_logic;
signal \N__4515\ : std_logic;
signal \N__4512\ : std_logic;
signal \N__4509\ : std_logic;
signal \N__4508\ : std_logic;
signal \N__4505\ : std_logic;
signal \N__4502\ : std_logic;
signal \N__4497\ : std_logic;
signal \N__4494\ : std_logic;
signal \N__4491\ : std_logic;
signal \N__4488\ : std_logic;
signal \N__4485\ : std_logic;
signal \N__4482\ : std_logic;
signal \N__4479\ : std_logic;
signal \N__4476\ : std_logic;
signal \N__4473\ : std_logic;
signal \N__4470\ : std_logic;
signal \N__4467\ : std_logic;
signal \N__4464\ : std_logic;
signal \N__4461\ : std_logic;
signal \N__4458\ : std_logic;
signal \N__4455\ : std_logic;
signal \N__4452\ : std_logic;
signal \N__4449\ : std_logic;
signal \N__4446\ : std_logic;
signal \N__4445\ : std_logic;
signal \N__4440\ : std_logic;
signal \N__4437\ : std_logic;
signal \N__4436\ : std_logic;
signal \N__4435\ : std_logic;
signal \N__4428\ : std_logic;
signal \N__4425\ : std_logic;
signal \N__4424\ : std_logic;
signal \N__4419\ : std_logic;
signal \N__4416\ : std_logic;
signal \N__4413\ : std_logic;
signal \N__4410\ : std_logic;
signal \N__4407\ : std_logic;
signal \N__4404\ : std_logic;
signal \N__4401\ : std_logic;
signal \N__4398\ : std_logic;
signal \N__4395\ : std_logic;
signal \N__4392\ : std_logic;
signal \N__4389\ : std_logic;
signal \N__4386\ : std_logic;
signal \N__4383\ : std_logic;
signal \N__4382\ : std_logic;
signal \N__4379\ : std_logic;
signal \N__4376\ : std_logic;
signal \N__4371\ : std_logic;
signal \N__4370\ : std_logic;
signal \N__4365\ : std_logic;
signal \N__4362\ : std_logic;
signal \N__4359\ : std_logic;
signal \N__4356\ : std_logic;
signal \N__4355\ : std_logic;
signal \N__4352\ : std_logic;
signal \N__4349\ : std_logic;
signal \N__4344\ : std_logic;
signal \N__4341\ : std_logic;
signal \N__4338\ : std_logic;
signal \N__4335\ : std_logic;
signal \N__4332\ : std_logic;
signal \N__4331\ : std_logic;
signal \N__4326\ : std_logic;
signal \N__4323\ : std_logic;
signal \N__4320\ : std_logic;
signal \N__4319\ : std_logic;
signal \N__4316\ : std_logic;
signal \N__4315\ : std_logic;
signal \N__4312\ : std_logic;
signal \N__4311\ : std_logic;
signal \N__4308\ : std_logic;
signal \N__4305\ : std_logic;
signal \N__4302\ : std_logic;
signal \N__4299\ : std_logic;
signal \N__4298\ : std_logic;
signal \N__4295\ : std_logic;
signal \N__4292\ : std_logic;
signal \N__4289\ : std_logic;
signal \N__4286\ : std_logic;
signal \N__4283\ : std_logic;
signal \N__4272\ : std_logic;
signal \N__4271\ : std_logic;
signal \N__4266\ : std_logic;
signal \N__4263\ : std_logic;
signal \N__4262\ : std_logic;
signal \N__4261\ : std_logic;
signal \N__4254\ : std_logic;
signal \N__4251\ : std_logic;
signal \N__4248\ : std_logic;
signal \N__4247\ : std_logic;
signal \N__4246\ : std_logic;
signal \N__4245\ : std_logic;
signal \N__4242\ : std_logic;
signal \N__4241\ : std_logic;
signal \N__4240\ : std_logic;
signal \N__4235\ : std_logic;
signal \N__4226\ : std_logic;
signal \N__4223\ : std_logic;
signal \N__4218\ : std_logic;
signal \N__4217\ : std_logic;
signal \N__4214\ : std_logic;
signal \N__4213\ : std_logic;
signal \N__4210\ : std_logic;
signal \N__4209\ : std_logic;
signal \N__4208\ : std_logic;
signal \N__4207\ : std_logic;
signal \N__4204\ : std_logic;
signal \N__4195\ : std_logic;
signal \N__4192\ : std_logic;
signal \N__4185\ : std_logic;
signal \N__4184\ : std_logic;
signal \N__4179\ : std_logic;
signal \N__4176\ : std_logic;
signal \N__4175\ : std_logic;
signal \N__4172\ : std_logic;
signal \N__4169\ : std_logic;
signal \N__4164\ : std_logic;
signal \N__4163\ : std_logic;
signal \N__4160\ : std_logic;
signal \N__4157\ : std_logic;
signal \N__4152\ : std_logic;
signal \N__4151\ : std_logic;
signal \N__4148\ : std_logic;
signal \N__4145\ : std_logic;
signal \N__4142\ : std_logic;
signal \N__4137\ : std_logic;
signal \N__4136\ : std_logic;
signal \N__4133\ : std_logic;
signal \N__4130\ : std_logic;
signal \N__4125\ : std_logic;
signal \N__4122\ : std_logic;
signal \N__4119\ : std_logic;
signal \N__4116\ : std_logic;
signal \N__4113\ : std_logic;
signal \N__4112\ : std_logic;
signal \N__4109\ : std_logic;
signal \N__4106\ : std_logic;
signal \N__4101\ : std_logic;
signal \N__4100\ : std_logic;
signal \N__4097\ : std_logic;
signal \N__4094\ : std_logic;
signal \N__4089\ : std_logic;
signal \N__4088\ : std_logic;
signal \N__4085\ : std_logic;
signal \N__4082\ : std_logic;
signal \N__4079\ : std_logic;
signal \N__4074\ : std_logic;
signal \N__4073\ : std_logic;
signal \N__4070\ : std_logic;
signal \N__4067\ : std_logic;
signal \N__4062\ : std_logic;
signal \N__4059\ : std_logic;
signal \N__4056\ : std_logic;
signal \N__4053\ : std_logic;
signal \N__4050\ : std_logic;
signal \N__4047\ : std_logic;
signal \N__4046\ : std_logic;
signal \N__4043\ : std_logic;
signal \N__4040\ : std_logic;
signal \N__4037\ : std_logic;
signal \N__4032\ : std_logic;
signal \N__4031\ : std_logic;
signal \N__4028\ : std_logic;
signal \N__4025\ : std_logic;
signal \N__4020\ : std_logic;
signal \N__4017\ : std_logic;
signal \N__4016\ : std_logic;
signal \N__4013\ : std_logic;
signal \N__4010\ : std_logic;
signal \N__4007\ : std_logic;
signal \N__4002\ : std_logic;
signal \N__4001\ : std_logic;
signal \N__3998\ : std_logic;
signal \N__3995\ : std_logic;
signal \N__3992\ : std_logic;
signal \N__3987\ : std_logic;
signal \N__3984\ : std_logic;
signal \N__3983\ : std_logic;
signal \N__3980\ : std_logic;
signal \N__3977\ : std_logic;
signal \N__3972\ : std_logic;
signal \N__3969\ : std_logic;
signal \N__3968\ : std_logic;
signal \N__3965\ : std_logic;
signal \N__3962\ : std_logic;
signal \N__3959\ : std_logic;
signal \N__3954\ : std_logic;
signal \N__3951\ : std_logic;
signal \N__3948\ : std_logic;
signal \N__3945\ : std_logic;
signal \N__3942\ : std_logic;
signal \N__3941\ : std_logic;
signal \N__3940\ : std_logic;
signal \N__3939\ : std_logic;
signal \N__3936\ : std_logic;
signal \N__3933\ : std_logic;
signal \N__3930\ : std_logic;
signal \N__3927\ : std_logic;
signal \N__3918\ : std_logic;
signal \N__3917\ : std_logic;
signal \N__3914\ : std_logic;
signal \N__3911\ : std_logic;
signal \N__3906\ : std_logic;
signal \N__3905\ : std_logic;
signal \N__3902\ : std_logic;
signal \N__3899\ : std_logic;
signal \N__3894\ : std_logic;
signal \N__3891\ : std_logic;
signal \N__3890\ : std_logic;
signal \N__3887\ : std_logic;
signal \N__3884\ : std_logic;
signal \N__3881\ : std_logic;
signal \N__3876\ : std_logic;
signal \N__3875\ : std_logic;
signal \N__3872\ : std_logic;
signal \N__3869\ : std_logic;
signal \N__3864\ : std_logic;
signal \N__3861\ : std_logic;
signal \N__3858\ : std_logic;
signal \N__3855\ : std_logic;
signal \N__3852\ : std_logic;
signal \N__3849\ : std_logic;
signal \N__3848\ : std_logic;
signal \N__3843\ : std_logic;
signal \N__3840\ : std_logic;
signal \N__3837\ : std_logic;
signal \N__3834\ : std_logic;
signal \N__3831\ : std_logic;
signal \N__3830\ : std_logic;
signal \N__3827\ : std_logic;
signal \N__3824\ : std_logic;
signal \N__3819\ : std_logic;
signal \N__3816\ : std_logic;
signal \N__3813\ : std_logic;
signal \N__3810\ : std_logic;
signal \N__3807\ : std_logic;
signal \N__3806\ : std_logic;
signal \N__3803\ : std_logic;
signal \N__3800\ : std_logic;
signal \N__3797\ : std_logic;
signal \N__3794\ : std_logic;
signal \N__3791\ : std_logic;
signal \N__3788\ : std_logic;
signal \N__3783\ : std_logic;
signal \N__3782\ : std_logic;
signal \N__3777\ : std_logic;
signal \N__3774\ : std_logic;
signal \N__3773\ : std_logic;
signal \N__3770\ : std_logic;
signal \N__3767\ : std_logic;
signal \N__3762\ : std_logic;
signal \N__3761\ : std_logic;
signal \N__3758\ : std_logic;
signal \N__3755\ : std_logic;
signal \N__3750\ : std_logic;
signal \N__3749\ : std_logic;
signal \N__3746\ : std_logic;
signal \N__3743\ : std_logic;
signal \N__3740\ : std_logic;
signal \N__3735\ : std_logic;
signal \N__3732\ : std_logic;
signal \N__3729\ : std_logic;
signal \N__3726\ : std_logic;
signal \N__3723\ : std_logic;
signal \N__3722\ : std_logic;
signal \N__3719\ : std_logic;
signal \N__3716\ : std_logic;
signal \N__3713\ : std_logic;
signal \N__3708\ : std_logic;
signal \N__3705\ : std_logic;
signal \N__3702\ : std_logic;
signal \N__3701\ : std_logic;
signal \N__3698\ : std_logic;
signal \N__3695\ : std_logic;
signal \N__3692\ : std_logic;
signal \N__3687\ : std_logic;
signal \N__3684\ : std_logic;
signal \N__3681\ : std_logic;
signal \N__3680\ : std_logic;
signal \N__3677\ : std_logic;
signal \N__3674\ : std_logic;
signal \N__3671\ : std_logic;
signal \N__3666\ : std_logic;
signal \N__3663\ : std_logic;
signal \N__3662\ : std_logic;
signal \N__3659\ : std_logic;
signal \N__3656\ : std_logic;
signal \N__3653\ : std_logic;
signal \N__3648\ : std_logic;
signal \N__3645\ : std_logic;
signal \N__3644\ : std_logic;
signal \N__3643\ : std_logic;
signal \N__3642\ : std_logic;
signal \N__3641\ : std_logic;
signal \N__3640\ : std_logic;
signal \N__3639\ : std_logic;
signal \N__3636\ : std_logic;
signal \N__3633\ : std_logic;
signal \N__3630\ : std_logic;
signal \N__3629\ : std_logic;
signal \N__3626\ : std_logic;
signal \N__3623\ : std_logic;
signal \N__3620\ : std_logic;
signal \N__3617\ : std_logic;
signal \N__3616\ : std_logic;
signal \N__3615\ : std_logic;
signal \N__3614\ : std_logic;
signal \N__3613\ : std_logic;
signal \N__3612\ : std_logic;
signal \N__3611\ : std_logic;
signal \N__3610\ : std_logic;
signal \N__3609\ : std_logic;
signal \N__3602\ : std_logic;
signal \N__3591\ : std_logic;
signal \N__3588\ : std_logic;
signal \N__3585\ : std_logic;
signal \N__3582\ : std_logic;
signal \N__3579\ : std_logic;
signal \N__3576\ : std_logic;
signal \N__3573\ : std_logic;
signal \N__3570\ : std_logic;
signal \N__3567\ : std_logic;
signal \N__3562\ : std_logic;
signal \N__3553\ : std_logic;
signal \N__3544\ : std_logic;
signal \N__3537\ : std_logic;
signal \N__3534\ : std_logic;
signal \N__3533\ : std_logic;
signal \N__3530\ : std_logic;
signal \N__3527\ : std_logic;
signal \N__3524\ : std_logic;
signal \N__3519\ : std_logic;
signal \N__3518\ : std_logic;
signal \N__3515\ : std_logic;
signal \N__3512\ : std_logic;
signal \N__3509\ : std_logic;
signal \N__3504\ : std_logic;
signal \N__3503\ : std_logic;
signal \N__3500\ : std_logic;
signal \N__3497\ : std_logic;
signal \N__3494\ : std_logic;
signal \N__3489\ : std_logic;
signal \N__3486\ : std_logic;
signal \N__3485\ : std_logic;
signal \N__3482\ : std_logic;
signal \N__3479\ : std_logic;
signal \N__3474\ : std_logic;
signal \N__3471\ : std_logic;
signal \N__3470\ : std_logic;
signal \N__3467\ : std_logic;
signal \N__3464\ : std_logic;
signal \N__3459\ : std_logic;
signal \N__3456\ : std_logic;
signal \N__3455\ : std_logic;
signal \N__3452\ : std_logic;
signal \N__3449\ : std_logic;
signal \N__3444\ : std_logic;
signal \N__3441\ : std_logic;
signal \N__3440\ : std_logic;
signal \N__3437\ : std_logic;
signal \N__3434\ : std_logic;
signal \N__3431\ : std_logic;
signal \N__3426\ : std_logic;
signal \N__3423\ : std_logic;
signal \N__3420\ : std_logic;
signal \N__3419\ : std_logic;
signal \N__3416\ : std_logic;
signal \N__3413\ : std_logic;
signal \N__3408\ : std_logic;
signal \N__3405\ : std_logic;
signal \N__3402\ : std_logic;
signal \N__3399\ : std_logic;
signal \N__3396\ : std_logic;
signal \N__3393\ : std_logic;
signal \N__3390\ : std_logic;
signal \N__3387\ : std_logic;
signal \N__3384\ : std_logic;
signal \N__3381\ : std_logic;
signal \N__3378\ : std_logic;
signal \N__3375\ : std_logic;
signal \N__3372\ : std_logic;
signal \N__3369\ : std_logic;
signal \N__3366\ : std_logic;
signal \N__3363\ : std_logic;
signal \N__3360\ : std_logic;
signal \N__3357\ : std_logic;
signal \N__3354\ : std_logic;
signal \N__3351\ : std_logic;
signal \N__3348\ : std_logic;
signal \N__3345\ : std_logic;
signal \N__3344\ : std_logic;
signal \N__3341\ : std_logic;
signal \N__3338\ : std_logic;
signal \N__3335\ : std_logic;
signal \N__3330\ : std_logic;
signal \N__3327\ : std_logic;
signal \N__3326\ : std_logic;
signal \N__3323\ : std_logic;
signal \N__3320\ : std_logic;
signal \N__3317\ : std_logic;
signal \N__3312\ : std_logic;
signal \N__3309\ : std_logic;
signal \N__3308\ : std_logic;
signal \N__3305\ : std_logic;
signal \N__3302\ : std_logic;
signal \N__3299\ : std_logic;
signal \N__3294\ : std_logic;
signal \N__3291\ : std_logic;
signal \N__3290\ : std_logic;
signal \N__3287\ : std_logic;
signal \N__3284\ : std_logic;
signal \N__3281\ : std_logic;
signal \N__3276\ : std_logic;
signal \N__3273\ : std_logic;
signal \N__3272\ : std_logic;
signal \N__3269\ : std_logic;
signal \N__3266\ : std_logic;
signal \N__3263\ : std_logic;
signal \N__3258\ : std_logic;
signal \N__3255\ : std_logic;
signal \N__3252\ : std_logic;
signal \N__3249\ : std_logic;
signal \N__3246\ : std_logic;
signal \N__3243\ : std_logic;
signal \N__3242\ : std_logic;
signal \N__3239\ : std_logic;
signal \N__3236\ : std_logic;
signal \N__3231\ : std_logic;
signal \N__3228\ : std_logic;
signal \N__3227\ : std_logic;
signal \N__3224\ : std_logic;
signal \N__3221\ : std_logic;
signal \N__3218\ : std_logic;
signal \N__3213\ : std_logic;
signal \N__3210\ : std_logic;
signal \N__3209\ : std_logic;
signal \N__3206\ : std_logic;
signal \N__3203\ : std_logic;
signal \N__3198\ : std_logic;
signal \N__3195\ : std_logic;
signal \N__3194\ : std_logic;
signal \N__3191\ : std_logic;
signal \N__3188\ : std_logic;
signal \N__3183\ : std_logic;
signal \N__3180\ : std_logic;
signal \N__3179\ : std_logic;
signal \N__3176\ : std_logic;
signal \N__3173\ : std_logic;
signal \N__3168\ : std_logic;
signal \N__3165\ : std_logic;
signal \N__3164\ : std_logic;
signal \N__3161\ : std_logic;
signal \N__3158\ : std_logic;
signal \N__3153\ : std_logic;
signal \N__3150\ : std_logic;
signal \N__3149\ : std_logic;
signal \N__3146\ : std_logic;
signal \N__3143\ : std_logic;
signal \N__3140\ : std_logic;
signal \N__3135\ : std_logic;
signal \N__3132\ : std_logic;
signal \N__3131\ : std_logic;
signal \N__3128\ : std_logic;
signal \N__3125\ : std_logic;
signal \N__3122\ : std_logic;
signal \N__3117\ : std_logic;
signal \N__3114\ : std_logic;
signal \N__3111\ : std_logic;
signal \N__3108\ : std_logic;
signal \N__3107\ : std_logic;
signal \N__3106\ : std_logic;
signal \N__3101\ : std_logic;
signal \N__3098\ : std_logic;
signal \N__3093\ : std_logic;
signal \N__3092\ : std_logic;
signal \N__3091\ : std_logic;
signal \N__3084\ : std_logic;
signal \N__3081\ : std_logic;
signal \N__3080\ : std_logic;
signal \N__3077\ : std_logic;
signal \N__3074\ : std_logic;
signal \N__3073\ : std_logic;
signal \N__3068\ : std_logic;
signal \N__3065\ : std_logic;
signal \N__3060\ : std_logic;
signal \N__3059\ : std_logic;
signal \N__3058\ : std_logic;
signal \N__3053\ : std_logic;
signal \N__3050\ : std_logic;
signal \N__3045\ : std_logic;
signal \N__3042\ : std_logic;
signal \N__3039\ : std_logic;
signal \N__3036\ : std_logic;
signal \N__3033\ : std_logic;
signal \N__3030\ : std_logic;
signal \N__3027\ : std_logic;
signal \N__3024\ : std_logic;
signal \N__3023\ : std_logic;
signal \N__3020\ : std_logic;
signal \N__3017\ : std_logic;
signal \N__3014\ : std_logic;
signal \N__3009\ : std_logic;
signal \N__3006\ : std_logic;
signal \N__3005\ : std_logic;
signal \N__3002\ : std_logic;
signal \N__2999\ : std_logic;
signal \N__2994\ : std_logic;
signal \N__2991\ : std_logic;
signal \N__2988\ : std_logic;
signal \N__2985\ : std_logic;
signal \N__2982\ : std_logic;
signal \N__2979\ : std_logic;
signal \N__2976\ : std_logic;
signal \N__2973\ : std_logic;
signal \N__2970\ : std_logic;
signal \N__2967\ : std_logic;
signal \N__2964\ : std_logic;
signal \N__2961\ : std_logic;
signal \N__2958\ : std_logic;
signal \N__2955\ : std_logic;
signal \N__2952\ : std_logic;
signal \N__2949\ : std_logic;
signal \N__2946\ : std_logic;
signal \N__2943\ : std_logic;
signal \N__2940\ : std_logic;
signal \N__2939\ : std_logic;
signal \N__2936\ : std_logic;
signal \N__2933\ : std_logic;
signal \N__2928\ : std_logic;
signal \N__2925\ : std_logic;
signal \N__2922\ : std_logic;
signal \N__2919\ : std_logic;
signal \N__2916\ : std_logic;
signal \N__2913\ : std_logic;
signal \N__2910\ : std_logic;
signal \N__2907\ : std_logic;
signal \N__2904\ : std_logic;
signal \N__2901\ : std_logic;
signal \N__2898\ : std_logic;
signal \N__2895\ : std_logic;
signal \N__2892\ : std_logic;
signal \N__2889\ : std_logic;
signal \N__2886\ : std_logic;
signal \N__2883\ : std_logic;
signal \N__2880\ : std_logic;
signal \N__2877\ : std_logic;
signal \N__2874\ : std_logic;
signal \N__2871\ : std_logic;
signal \N__2868\ : std_logic;
signal \N__2865\ : std_logic;
signal \N__2862\ : std_logic;
signal \N__2859\ : std_logic;
signal \N__2856\ : std_logic;
signal \N__2853\ : std_logic;
signal \N__2850\ : std_logic;
signal \N__2847\ : std_logic;
signal \N__2844\ : std_logic;
signal \N__2841\ : std_logic;
signal \N__2838\ : std_logic;
signal \N__2835\ : std_logic;
signal \N__2832\ : std_logic;
signal \N__2829\ : std_logic;
signal \N__2826\ : std_logic;
signal \N__2823\ : std_logic;
signal \N__2820\ : std_logic;
signal \N__2817\ : std_logic;
signal \N__2814\ : std_logic;
signal \N__2811\ : std_logic;
signal \N__2808\ : std_logic;
signal \N__2805\ : std_logic;
signal \N__2802\ : std_logic;
signal \N__2799\ : std_logic;
signal \N__2796\ : std_logic;
signal \N__2793\ : std_logic;
signal \N__2790\ : std_logic;
signal \N__2787\ : std_logic;
signal \N__2784\ : std_logic;
signal \N__2781\ : std_logic;
signal \N__2778\ : std_logic;
signal \N__2775\ : std_logic;
signal \N__2772\ : std_logic;
signal \N__2769\ : std_logic;
signal \N__2766\ : std_logic;
signal \N__2763\ : std_logic;
signal \N__2760\ : std_logic;
signal \N__2757\ : std_logic;
signal \N__2754\ : std_logic;
signal \N__2751\ : std_logic;
signal \N__2748\ : std_logic;
signal \N__2745\ : std_logic;
signal \N__2742\ : std_logic;
signal \CLK_pad_gb_input\ : std_logic;
signal \VCCG0\ : std_logic;
signal \GNDG0\ : std_logic;
signal \LED_c\ : std_logic;
signal n26 : std_logic;
signal \bfn_17_17_0_\ : std_logic;
signal n25_adj_402 : std_logic;
signal n2876 : std_logic;
signal n24_adj_401 : std_logic;
signal n2877 : std_logic;
signal n23_adj_400 : std_logic;
signal n2878 : std_logic;
signal n22_adj_399 : std_logic;
signal n2879 : std_logic;
signal n21 : std_logic;
signal n2880 : std_logic;
signal n20_adj_398 : std_logic;
signal n2881 : std_logic;
signal n19 : std_logic;
signal n2882 : std_logic;
signal n2883 : std_logic;
signal n18_adj_397 : std_logic;
signal \bfn_17_18_0_\ : std_logic;
signal n17 : std_logic;
signal n2884 : std_logic;
signal n16 : std_logic;
signal n2885 : std_logic;
signal n15_adj_396 : std_logic;
signal n2886 : std_logic;
signal n14_adj_395 : std_logic;
signal n2887 : std_logic;
signal n13_adj_394 : std_logic;
signal n2888 : std_logic;
signal n12_adj_393 : std_logic;
signal n2889 : std_logic;
signal n11 : std_logic;
signal n2890 : std_logic;
signal n2891 : std_logic;
signal n10 : std_logic;
signal \bfn_17_19_0_\ : std_logic;
signal n9 : std_logic;
signal n2892 : std_logic;
signal n8 : std_logic;
signal n2893 : std_logic;
signal n7 : std_logic;
signal n2894 : std_logic;
signal n6_adj_392 : std_logic;
signal n2895 : std_logic;
signal n2896 : std_logic;
signal n2897 : std_logic;
signal n2898 : std_logic;
signal n2899 : std_logic;
signal \bfn_17_20_0_\ : std_logic;
signal n2900 : std_logic;
signal blink_counter_25 : std_logic;
signal n3119 : std_logic;
signal blink_counter_21 : std_logic;
signal blink_counter_24 : std_logic;
signal blink_counter_23 : std_logic;
signal blink_counter_22 : std_logic;
signal n3120 : std_logic;
signal \n13_adj_391_cascade_\ : std_logic;
signal n14 : std_logic;
signal \n18_cascade_\ : std_logic;
signal \n3114_cascade_\ : std_logic;
signal delay_counter_0 : std_logic;
signal \bfn_20_17_0_\ : std_logic;
signal delay_counter_1 : std_logic;
signal n2818 : std_logic;
signal delay_counter_2 : std_logic;
signal n2819 : std_logic;
signal delay_counter_3 : std_logic;
signal n2820 : std_logic;
signal delay_counter_4 : std_logic;
signal n2821 : std_logic;
signal delay_counter_5 : std_logic;
signal n2822 : std_logic;
signal delay_counter_6 : std_logic;
signal n2823 : std_logic;
signal delay_counter_7 : std_logic;
signal n2824 : std_logic;
signal n2825 : std_logic;
signal delay_counter_8 : std_logic;
signal \bfn_20_18_0_\ : std_logic;
signal delay_counter_9 : std_logic;
signal n2826 : std_logic;
signal delay_counter_10 : std_logic;
signal n2827 : std_logic;
signal delay_counter_11 : std_logic;
signal n2828 : std_logic;
signal delay_counter_12 : std_logic;
signal n2829 : std_logic;
signal delay_counter_13 : std_logic;
signal n2830 : std_logic;
signal delay_counter_14 : std_logic;
signal n2831 : std_logic;
signal n2832 : std_logic;
signal n2833 : std_logic;
signal \bfn_20_19_0_\ : std_logic;
signal n2834 : std_logic;
signal n2835 : std_logic;
signal n2836 : std_logic;
signal n2837 : std_logic;
signal n2838 : std_logic;
signal n2839 : std_logic;
signal n2840 : std_logic;
signal n2841 : std_logic;
signal \bfn_20_20_0_\ : std_logic;
signal n2842 : std_logic;
signal n2843 : std_logic;
signal n2844 : std_logic;
signal n2845 : std_logic;
signal n2846 : std_logic;
signal n2847 : std_logic;
signal n2848 : std_logic;
signal \eeprom.n1704_cascade_\ : std_logic;
signal \eeprom.n25\ : std_logic;
signal \eeprom.n26_adj_385\ : std_logic;
signal \eeprom.n27\ : std_logic;
signal \eeprom.delay_counter_0\ : std_logic;
signal \bfn_21_13_0_\ : std_logic;
signal \eeprom.delay_counter_1\ : std_logic;
signal \eeprom.n2856\ : std_logic;
signal \eeprom.delay_counter_2\ : std_logic;
signal \eeprom.n2857\ : std_logic;
signal \eeprom.delay_counter_3\ : std_logic;
signal \eeprom.n2858\ : std_logic;
signal \eeprom.delay_counter_4\ : std_logic;
signal \eeprom.n2859\ : std_logic;
signal \eeprom.delay_counter_5\ : std_logic;
signal \eeprom.n2860\ : std_logic;
signal \eeprom.n2861\ : std_logic;
signal \eeprom.delay_counter_7\ : std_logic;
signal \eeprom.n2862\ : std_logic;
signal \eeprom.n2863\ : std_logic;
signal \bfn_21_14_0_\ : std_logic;
signal \eeprom.delay_counter_9\ : std_logic;
signal \eeprom.n2864\ : std_logic;
signal \eeprom.n2865\ : std_logic;
signal \eeprom.delay_counter_11\ : std_logic;
signal \eeprom.n2866\ : std_logic;
signal \eeprom.n2867\ : std_logic;
signal \eeprom.delay_counter_13\ : std_logic;
signal \eeprom.n2868\ : std_logic;
signal \eeprom.delay_counter_14\ : std_logic;
signal \eeprom.n2869\ : std_logic;
signal \eeprom.n730\ : std_logic;
signal \eeprom.n2870\ : std_logic;
signal \eeprom.delay_counter_15\ : std_logic;
signal \n805_cascade_\ : std_logic;
signal \eeprom.n1796\ : std_logic;
signal \eeprom.n1796_cascade_\ : std_logic;
signal \eeprom.n1929\ : std_logic;
signal data_ready : std_logic;
signal delay_counter_16 : std_logic;
signal delay_counter_17 : std_logic;
signal delay_counter_15 : std_logic;
signal n3069 : std_logic;
signal delay_counter_29 : std_logic;
signal delay_counter_18 : std_logic;
signal \n36_cascade_\ : std_logic;
signal delay_counter_24 : std_logic;
signal delay_counter_27 : std_logic;
signal \n22_cascade_\ : std_logic;
signal delay_counter_23 : std_logic;
signal delay_counter_31 : std_logic;
signal \n25_cascade_\ : std_logic;
signal \n104_cascade_\ : std_logic;
signal n1891 : std_logic;
signal delay_counter_21 : std_logic;
signal delay_counter_25 : std_logic;
signal delay_counter_20 : std_logic;
signal delay_counter_19 : std_logic;
signal n23 : std_logic;
signal n20 : std_logic;
signal \n20_cascade_\ : std_logic;
signal n6 : std_logic;
signal \n1836_cascade_\ : std_logic;
signal n1507 : std_logic;
signal n104 : std_logic;
signal n15 : std_logic;
signal \ID_READOUT_FSM_state_1\ : std_logic;
signal \ID_READOUT_FSM_state_0\ : std_logic;
signal n2414 : std_logic;
signal delay_counter_22 : std_logic;
signal delay_counter_30 : std_logic;
signal delay_counter_26 : std_logic;
signal delay_counter_28 : std_logic;
signal n24 : std_logic;
signal \eeprom.i2c.n10_adj_381_cascade_\ : std_logic;
signal \eeprom.delay_counter_12\ : std_logic;
signal \eeprom.delay_counter_10\ : std_logic;
signal \eeprom.delay_counter_8\ : std_logic;
signal \eeprom.delay_counter_6\ : std_logic;
signal \eeprom.n28\ : std_logic;
signal \eeprom.i2c.n2388\ : std_logic;
signal data_5 : std_logic;
signal data_0 : std_logic;
signal data_3 : std_logic;
signal n13 : std_logic;
signal n12 : std_logic;
signal data_4 : std_logic;
signal \n1718_cascade_\ : std_logic;
signal data_2 : std_logic;
signal n1718 : std_logic;
signal data_6 : std_logic;
signal \INVeeprom.i2c.write_enable_131C_net\ : std_logic;
signal \eeprom.i2c.n1928\ : std_logic;
signal \eeprom.i2c.n3130_cascade_\ : std_logic;
signal \eeprom.i2c.n1153\ : std_logic;
signal \eeprom.i2c.n37_cascade_\ : std_logic;
signal \eeprom.i2c.n33\ : std_logic;
signal \eeprom.i2c.n39\ : std_logic;
signal \eeprom.i2c.n39_cascade_\ : std_logic;
signal \eeprom.i2c.n3133\ : std_logic;
signal \eeprom.i2c.n7\ : std_logic;
signal \eeprom.i2c.n3082\ : std_logic;
signal \eeprom.i2c.n13\ : std_logic;
signal \eeprom.i2c.n15_cascade_\ : std_logic;
signal \eeprom.i2c.n10_adj_381\ : std_logic;
signal \eeprom.i2c.n11_adj_378_cascade_\ : std_logic;
signal \eeprom.i2c.n2352\ : std_logic;
signal \eeprom.i2c.n1734_cascade_\ : std_logic;
signal \eeprom.i2c.n2358\ : std_logic;
signal \eeprom.i2c.n1063_cascade_\ : std_logic;
signal \eeprom.i2c.n1923\ : std_logic;
signal \eeprom.enable\ : std_logic;
signal \eeprom.i2c.n1761\ : std_logic;
signal \eeprom.n1704\ : std_logic;
signal \eeprom.n26_cascade_\ : std_logic;
signal \eeprom.i2c.n3123\ : std_logic;
signal \INVeeprom.i2c.sda_out_132C_net\ : std_logic;
signal \eeprom.i2c.n2967\ : std_logic;
signal \eeprom.i2c.n11\ : std_logic;
signal rw : std_logic;
signal \state_7_N_270_0\ : std_logic;
signal \eeprom.i2c.n11_adj_374\ : std_logic;
signal \eeprom.i2c.n11_adj_378\ : std_logic;
signal saved_addr_0 : std_logic;
signal n4 : std_logic;
signal \eeprom.i2c.n1063\ : std_logic;
signal \eeprom.i2c.n9_adj_377_cascade_\ : std_logic;
signal \eeprom.i2c.n3050\ : std_logic;
signal n4_adj_389 : std_logic;
signal n2344 : std_logic;
signal \n2344_cascade_\ : std_logic;
signal data_7 : std_logic;
signal \enable_slow_N_373\ : std_logic;
signal \eeprom.n14_cascade_\ : std_logic;
signal n2382 : std_logic;
signal \n3051_cascade_\ : std_logic;
signal n2913 : std_logic;
signal \n1113_cascade_\ : std_logic;
signal read : std_logic;
signal n3109 : std_logic;
signal \eeprom.n9\ : std_logic;
signal state_1 : std_logic;
signal state_0 : std_logic;
signal \eeprom.n3142\ : std_logic;
signal \eeprom.i2c.n10_adj_380_cascade_\ : std_logic;
signal \eeprom.i2c.n15\ : std_logic;
signal \bfn_26_14_0_\ : std_logic;
signal \eeprom.i2c.n2849\ : std_logic;
signal \eeprom.i2c.n2850\ : std_logic;
signal \eeprom.i2c.n2851\ : std_logic;
signal \eeprom.i2c.n2852\ : std_logic;
signal \eeprom.i2c.n2853\ : std_logic;
signal \eeprom.i2c.n2854\ : std_logic;
signal \eeprom.i2c.n2855\ : std_logic;
signal \eeprom.n10\ : std_logic;
signal \eeprom.i2c.n9_adj_377\ : std_logic;
signal \eeprom.i2c.n3039_cascade_\ : std_logic;
signal \state_7_N_286_3\ : std_logic;
signal n1723 : std_logic;
signal data_1 : std_logic;
signal \eeprom.i2c.counter_6\ : std_logic;
signal \eeprom.i2c.counter_3\ : std_logic;
signal \eeprom.i2c.counter_5\ : std_logic;
signal \eeprom.i2c.counter_7\ : std_logic;
signal \eeprom.i2c.counter_4\ : std_logic;
signal \eeprom.i2c.n12_cascade_\ : std_logic;
signal \eeprom.i2c.n1056\ : std_logic;
signal \eeprom.i2c.n1172\ : std_logic;
signal \eeprom.i2c.n3039\ : std_logic;
signal \eeprom.i2c.n1056_cascade_\ : std_logic;
signal \eeprom.i2c.n37\ : std_logic;
signal \eeprom.i2c.counter_2\ : std_logic;
signal \eeprom.i2c.counter_1\ : std_logic;
signal n4_adj_390 : std_logic;
signal \eeprom.state_1_adj_386\ : std_logic;
signal \eeprom.state_3\ : std_logic;
signal \eeprom.state_0_adj_384\ : std_logic;
signal \eeprom.i2c.state_2\ : std_logic;
signal \INVeeprom.i2c.i2c_scl_enable_123C_net\ : std_logic;
signal \eeprom.i2c.counter2_0\ : std_logic;
signal \bfn_27_13_0_\ : std_logic;
signal \eeprom.i2c.counter2_1\ : std_logic;
signal \eeprom.i2c.n2871\ : std_logic;
signal \eeprom.i2c.counter2_2\ : std_logic;
signal \eeprom.i2c.n2872\ : std_logic;
signal \eeprom.i2c.counter2_3\ : std_logic;
signal \eeprom.i2c.n2873\ : std_logic;
signal \eeprom.i2c.counter2_4\ : std_logic;
signal \eeprom.i2c.n2874\ : std_logic;
signal \eeprom.i2c.n2875\ : std_logic;
signal \eeprom.i2c.counter2_5\ : std_logic;
signal \CLK_c\ : std_logic;
signal \eeprom.i2c.n1930\ : std_logic;
signal \eeprom.i2c.counter_0\ : std_logic;
signal \eeprom.i2c.n1757\ : std_logic;
signal \eeprom.i2c.n1924\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \eeprom.i2c.sda_out_adj_375\ : std_logic;
signal sda_enable : std_logic;
signal sda_out : std_logic;
signal \eeprom.i2c.i2c_clk\ : std_logic;
signal scl_enable : std_logic;
signal scl_c : std_logic;
signal \_gnd_net_\ : std_logic;

signal \CS_CLK_wire\ : std_logic;
signal \CS_wire\ : std_logic;
signal \DE_wire\ : std_logic;
signal \INHA_wire\ : std_logic;
signal \INHB_wire\ : std_logic;
signal \INHC_wire\ : std_logic;
signal \INLA_wire\ : std_logic;
signal \INLB_wire\ : std_logic;
signal \INLC_wire\ : std_logic;
signal \LED_wire\ : std_logic;
signal \NEOPXL_wire\ : std_logic;
signal \TX_wire\ : std_logic;
signal \USBPU_wire\ : std_logic;
signal \CLK_wire\ : std_logic;

begin
    CS_CLK <= \CS_CLK_wire\;
    CS <= \CS_wire\;
    DE <= \DE_wire\;
    INHA <= \INHA_wire\;
    INHB <= \INHB_wire\;
    INHC <= \INHC_wire\;
    INLA <= \INLA_wire\;
    INLB <= \INLB_wire\;
    INLC <= \INLC_wire\;
    LED <= \LED_wire\;
    NEOPXL <= \NEOPXL_wire\;
    TX <= \TX_wire\;
    USBPU <= \USBPU_wire\;
    \CLK_wire\ <= CLK;

    \CS_CLK_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6937\,
            DIN => \N__6936\,
            DOUT => \N__6935\,
            PACKAGEPIN => \CS_CLK_wire\
        );

    \CS_CLK_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__6937\,
            PADOUT => \N__6936\,
            PADIN => \N__6935\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \CS_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6928\,
            DIN => \N__6927\,
            DOUT => \N__6926\,
            PACKAGEPIN => \CS_wire\
        );

    \CS_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__6928\,
            PADOUT => \N__6927\,
            PADIN => \N__6926\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \DE_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6919\,
            DIN => \N__6918\,
            DOUT => \N__6917\,
            PACKAGEPIN => \DE_wire\
        );

    \DE_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__6919\,
            PADOUT => \N__6918\,
            PADIN => \N__6917\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \INHA_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6910\,
            DIN => \N__6909\,
            DOUT => \N__6908\,
            PACKAGEPIN => \INHA_wire\
        );

    \INHA_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__6910\,
            PADOUT => \N__6909\,
            PADIN => \N__6908\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \INHB_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6901\,
            DIN => \N__6900\,
            DOUT => \N__6899\,
            PACKAGEPIN => \INHB_wire\
        );

    \INHB_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__6901\,
            PADOUT => \N__6900\,
            PADIN => \N__6899\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \INHC_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6892\,
            DIN => \N__6891\,
            DOUT => \N__6890\,
            PACKAGEPIN => \INHC_wire\
        );

    \INHC_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__6892\,
            PADOUT => \N__6891\,
            PADIN => \N__6890\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \INLA_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6883\,
            DIN => \N__6882\,
            DOUT => \N__6881\,
            PACKAGEPIN => \INLA_wire\
        );

    \INLA_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__6883\,
            PADOUT => \N__6882\,
            PADIN => \N__6881\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \INLB_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6874\,
            DIN => \N__6873\,
            DOUT => \N__6872\,
            PACKAGEPIN => \INLB_wire\
        );

    \INLB_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__6874\,
            PADOUT => \N__6873\,
            PADIN => \N__6872\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \INLC_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6865\,
            DIN => \N__6864\,
            DOUT => \N__6863\,
            PACKAGEPIN => \INLC_wire\
        );

    \INLC_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__6865\,
            PADOUT => \N__6864\,
            PADIN => \N__6863\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \LED_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6856\,
            DIN => \N__6855\,
            DOUT => \N__6854\,
            PACKAGEPIN => \LED_wire\
        );

    \LED_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__6856\,
            PADOUT => \N__6855\,
            PADIN => \N__6854\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__2775\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \NEOPXL_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6847\,
            DIN => \N__6846\,
            DOUT => \N__6845\,
            PACKAGEPIN => \NEOPXL_wire\
        );

    \NEOPXL_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__6847\,
            PADOUT => \N__6846\,
            PADIN => \N__6845\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \TX_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6838\,
            DIN => \N__6837\,
            DOUT => \N__6836\,
            PACKAGEPIN => \TX_wire\
        );

    \TX_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__6838\,
            PADOUT => \N__6837\,
            PADIN => \N__6836\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \USBPU_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6829\,
            DIN => \N__6828\,
            DOUT => \N__6827\,
            PACKAGEPIN => \USBPU_wire\
        );

    \USBPU_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__6829\,
            PADOUT => \N__6828\,
            PADIN => \N__6827\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \scl_output_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__6820\,
            DIN => \N__6819\,
            DOUT => \N__6818\,
            PACKAGEPIN => SCL
        );

    \scl_output_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__6820\,
            PADOUT => \N__6819\,
            PADIN => \N__6818\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__6300\,
            DOUT1 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__6330\
        );

    \sda_output_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__6811\,
            DIN => \N__6810\,
            DOUT => \N__6809\,
            PACKAGEPIN => SDA
        );

    \sda_output_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__6811\,
            PADOUT => \N__6810\,
            PADIN => \N__6809\,
            CLOCKENABLE => 'H',
            DIN0 => \state_7_N_286_3\,
            DIN1 => OPEN,
            DOUT0 => \N__6498\,
            DOUT1 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__6525\
        );

    \CLK_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6802\,
            DIN => \N__6801\,
            DOUT => \N__6800\,
            PACKAGEPIN => \CLK_wire\
        );

    \CLK_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__6802\,
            PADOUT => \N__6801\,
            PADIN => \N__6800\,
            CLOCKENABLE => 'H',
            DIN0 => \CLK_pad_gb_input\,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \I__1582\ : CascadeMux
    port map (
            O => \N__6783\,
            I => \N__6779\
        );

    \I__1581\ : InMux
    port map (
            O => \N__6782\,
            I => \N__6776\
        );

    \I__1580\ : InMux
    port map (
            O => \N__6779\,
            I => \N__6773\
        );

    \I__1579\ : LocalMux
    port map (
            O => \N__6776\,
            I => \eeprom.i2c.counter2_4\
        );

    \I__1578\ : LocalMux
    port map (
            O => \N__6773\,
            I => \eeprom.i2c.counter2_4\
        );

    \I__1577\ : InMux
    port map (
            O => \N__6768\,
            I => \eeprom.i2c.n2874\
        );

    \I__1576\ : InMux
    port map (
            O => \N__6765\,
            I => \eeprom.i2c.n2875\
        );

    \I__1575\ : InMux
    port map (
            O => \N__6762\,
            I => \N__6758\
        );

    \I__1574\ : InMux
    port map (
            O => \N__6761\,
            I => \N__6755\
        );

    \I__1573\ : LocalMux
    port map (
            O => \N__6758\,
            I => \eeprom.i2c.counter2_5\
        );

    \I__1572\ : LocalMux
    port map (
            O => \N__6755\,
            I => \eeprom.i2c.counter2_5\
        );

    \I__1571\ : ClkMux
    port map (
            O => \N__6750\,
            I => \N__6693\
        );

    \I__1570\ : ClkMux
    port map (
            O => \N__6749\,
            I => \N__6693\
        );

    \I__1569\ : ClkMux
    port map (
            O => \N__6748\,
            I => \N__6693\
        );

    \I__1568\ : ClkMux
    port map (
            O => \N__6747\,
            I => \N__6693\
        );

    \I__1567\ : ClkMux
    port map (
            O => \N__6746\,
            I => \N__6693\
        );

    \I__1566\ : ClkMux
    port map (
            O => \N__6745\,
            I => \N__6693\
        );

    \I__1565\ : ClkMux
    port map (
            O => \N__6744\,
            I => \N__6693\
        );

    \I__1564\ : ClkMux
    port map (
            O => \N__6743\,
            I => \N__6693\
        );

    \I__1563\ : ClkMux
    port map (
            O => \N__6742\,
            I => \N__6693\
        );

    \I__1562\ : ClkMux
    port map (
            O => \N__6741\,
            I => \N__6693\
        );

    \I__1561\ : ClkMux
    port map (
            O => \N__6740\,
            I => \N__6693\
        );

    \I__1560\ : ClkMux
    port map (
            O => \N__6739\,
            I => \N__6693\
        );

    \I__1559\ : ClkMux
    port map (
            O => \N__6738\,
            I => \N__6693\
        );

    \I__1558\ : ClkMux
    port map (
            O => \N__6737\,
            I => \N__6693\
        );

    \I__1557\ : ClkMux
    port map (
            O => \N__6736\,
            I => \N__6693\
        );

    \I__1556\ : ClkMux
    port map (
            O => \N__6735\,
            I => \N__6693\
        );

    \I__1555\ : ClkMux
    port map (
            O => \N__6734\,
            I => \N__6693\
        );

    \I__1554\ : ClkMux
    port map (
            O => \N__6733\,
            I => \N__6693\
        );

    \I__1553\ : ClkMux
    port map (
            O => \N__6732\,
            I => \N__6693\
        );

    \I__1552\ : GlobalMux
    port map (
            O => \N__6693\,
            I => \N__6690\
        );

    \I__1551\ : gio2CtrlBuf
    port map (
            O => \N__6690\,
            I => \CLK_c\
        );

    \I__1550\ : SRMux
    port map (
            O => \N__6687\,
            I => \N__6684\
        );

    \I__1549\ : LocalMux
    port map (
            O => \N__6684\,
            I => \N__6681\
        );

    \I__1548\ : Span4Mux_v
    port map (
            O => \N__6681\,
            I => \N__6677\
        );

    \I__1547\ : InMux
    port map (
            O => \N__6680\,
            I => \N__6674\
        );

    \I__1546\ : Odrv4
    port map (
            O => \N__6677\,
            I => \eeprom.i2c.n1930\
        );

    \I__1545\ : LocalMux
    port map (
            O => \N__6674\,
            I => \eeprom.i2c.n1930\
        );

    \I__1544\ : InMux
    port map (
            O => \N__6669\,
            I => \N__6666\
        );

    \I__1543\ : LocalMux
    port map (
            O => \N__6666\,
            I => \N__6662\
        );

    \I__1542\ : InMux
    port map (
            O => \N__6665\,
            I => \N__6659\
        );

    \I__1541\ : Span4Mux_v
    port map (
            O => \N__6662\,
            I => \N__6652\
        );

    \I__1540\ : LocalMux
    port map (
            O => \N__6659\,
            I => \N__6652\
        );

    \I__1539\ : InMux
    port map (
            O => \N__6658\,
            I => \N__6648\
        );

    \I__1538\ : InMux
    port map (
            O => \N__6657\,
            I => \N__6645\
        );

    \I__1537\ : Span4Mux_h
    port map (
            O => \N__6652\,
            I => \N__6642\
        );

    \I__1536\ : InMux
    port map (
            O => \N__6651\,
            I => \N__6639\
        );

    \I__1535\ : LocalMux
    port map (
            O => \N__6648\,
            I => \eeprom.i2c.counter_0\
        );

    \I__1534\ : LocalMux
    port map (
            O => \N__6645\,
            I => \eeprom.i2c.counter_0\
        );

    \I__1533\ : Odrv4
    port map (
            O => \N__6642\,
            I => \eeprom.i2c.counter_0\
        );

    \I__1532\ : LocalMux
    port map (
            O => \N__6639\,
            I => \eeprom.i2c.counter_0\
        );

    \I__1531\ : CEMux
    port map (
            O => \N__6630\,
            I => \N__6626\
        );

    \I__1530\ : CEMux
    port map (
            O => \N__6629\,
            I => \N__6623\
        );

    \I__1529\ : LocalMux
    port map (
            O => \N__6626\,
            I => \N__6620\
        );

    \I__1528\ : LocalMux
    port map (
            O => \N__6623\,
            I => \N__6617\
        );

    \I__1527\ : Span4Mux_v
    port map (
            O => \N__6620\,
            I => \N__6614\
        );

    \I__1526\ : Span4Mux_h
    port map (
            O => \N__6617\,
            I => \N__6611\
        );

    \I__1525\ : Odrv4
    port map (
            O => \N__6614\,
            I => \eeprom.i2c.n1757\
        );

    \I__1524\ : Odrv4
    port map (
            O => \N__6611\,
            I => \eeprom.i2c.n1757\
        );

    \I__1523\ : SRMux
    port map (
            O => \N__6606\,
            I => \N__6603\
        );

    \I__1522\ : LocalMux
    port map (
            O => \N__6603\,
            I => \N__6600\
        );

    \I__1521\ : Span4Mux_v
    port map (
            O => \N__6600\,
            I => \N__6596\
        );

    \I__1520\ : SRMux
    port map (
            O => \N__6599\,
            I => \N__6593\
        );

    \I__1519\ : Span4Mux_h
    port map (
            O => \N__6596\,
            I => \N__6590\
        );

    \I__1518\ : LocalMux
    port map (
            O => \N__6593\,
            I => \N__6587\
        );

    \I__1517\ : Odrv4
    port map (
            O => \N__6590\,
            I => \eeprom.i2c.n1924\
        );

    \I__1516\ : Odrv12
    port map (
            O => \N__6587\,
            I => \eeprom.i2c.n1924\
        );

    \I__1515\ : CascadeMux
    port map (
            O => \N__6582\,
            I => \N__6576\
        );

    \I__1514\ : CascadeMux
    port map (
            O => \N__6581\,
            I => \N__6572\
        );

    \I__1513\ : CascadeMux
    port map (
            O => \N__6580\,
            I => \N__6568\
        );

    \I__1512\ : InMux
    port map (
            O => \N__6579\,
            I => \N__6551\
        );

    \I__1511\ : InMux
    port map (
            O => \N__6576\,
            I => \N__6551\
        );

    \I__1510\ : InMux
    port map (
            O => \N__6575\,
            I => \N__6551\
        );

    \I__1509\ : InMux
    port map (
            O => \N__6572\,
            I => \N__6551\
        );

    \I__1508\ : InMux
    port map (
            O => \N__6571\,
            I => \N__6551\
        );

    \I__1507\ : InMux
    port map (
            O => \N__6568\,
            I => \N__6551\
        );

    \I__1506\ : InMux
    port map (
            O => \N__6567\,
            I => \N__6551\
        );

    \I__1505\ : InMux
    port map (
            O => \N__6566\,
            I => \N__6548\
        );

    \I__1504\ : LocalMux
    port map (
            O => \N__6551\,
            I => \CONSTANT_ONE_NET\
        );

    \I__1503\ : LocalMux
    port map (
            O => \N__6548\,
            I => \CONSTANT_ONE_NET\
        );

    \I__1502\ : InMux
    port map (
            O => \N__6543\,
            I => \N__6540\
        );

    \I__1501\ : LocalMux
    port map (
            O => \N__6540\,
            I => \N__6537\
        );

    \I__1500\ : Span4Mux_v
    port map (
            O => \N__6537\,
            I => \N__6534\
        );

    \I__1499\ : Span4Mux_v
    port map (
            O => \N__6534\,
            I => \N__6531\
        );

    \I__1498\ : Span4Mux_h
    port map (
            O => \N__6531\,
            I => \N__6528\
        );

    \I__1497\ : Odrv4
    port map (
            O => \N__6528\,
            I => \eeprom.i2c.sda_out_adj_375\
        );

    \I__1496\ : IoInMux
    port map (
            O => \N__6525\,
            I => \N__6522\
        );

    \I__1495\ : LocalMux
    port map (
            O => \N__6522\,
            I => \N__6519\
        );

    \I__1494\ : IoSpan4Mux
    port map (
            O => \N__6519\,
            I => \N__6515\
        );

    \I__1493\ : InMux
    port map (
            O => \N__6518\,
            I => \N__6512\
        );

    \I__1492\ : Span4Mux_s1_h
    port map (
            O => \N__6515\,
            I => \N__6507\
        );

    \I__1491\ : LocalMux
    port map (
            O => \N__6512\,
            I => \N__6507\
        );

    \I__1490\ : Span4Mux_h
    port map (
            O => \N__6507\,
            I => \N__6504\
        );

    \I__1489\ : Span4Mux_v
    port map (
            O => \N__6504\,
            I => \N__6501\
        );

    \I__1488\ : Odrv4
    port map (
            O => \N__6501\,
            I => sda_enable
        );

    \I__1487\ : IoInMux
    port map (
            O => \N__6498\,
            I => \N__6495\
        );

    \I__1486\ : LocalMux
    port map (
            O => \N__6495\,
            I => \N__6492\
        );

    \I__1485\ : Span4Mux_s2_h
    port map (
            O => \N__6492\,
            I => \N__6489\
        );

    \I__1484\ : Odrv4
    port map (
            O => \N__6489\,
            I => sda_out
        );

    \I__1483\ : ClkMux
    port map (
            O => \N__6486\,
            I => \N__6483\
        );

    \I__1482\ : LocalMux
    port map (
            O => \N__6483\,
            I => \N__6479\
        );

    \I__1481\ : ClkMux
    port map (
            O => \N__6482\,
            I => \N__6472\
        );

    \I__1480\ : Span4Mux_v
    port map (
            O => \N__6479\,
            I => \N__6469\
        );

    \I__1479\ : ClkMux
    port map (
            O => \N__6478\,
            I => \N__6466\
        );

    \I__1478\ : InMux
    port map (
            O => \N__6477\,
            I => \N__6463\
        );

    \I__1477\ : ClkMux
    port map (
            O => \N__6476\,
            I => \N__6460\
        );

    \I__1476\ : ClkMux
    port map (
            O => \N__6475\,
            I => \N__6455\
        );

    \I__1475\ : LocalMux
    port map (
            O => \N__6472\,
            I => \N__6452\
        );

    \I__1474\ : Span4Mux_h
    port map (
            O => \N__6469\,
            I => \N__6447\
        );

    \I__1473\ : LocalMux
    port map (
            O => \N__6466\,
            I => \N__6447\
        );

    \I__1472\ : LocalMux
    port map (
            O => \N__6463\,
            I => \N__6443\
        );

    \I__1471\ : LocalMux
    port map (
            O => \N__6460\,
            I => \N__6440\
        );

    \I__1470\ : ClkMux
    port map (
            O => \N__6459\,
            I => \N__6437\
        );

    \I__1469\ : ClkMux
    port map (
            O => \N__6458\,
            I => \N__6433\
        );

    \I__1468\ : LocalMux
    port map (
            O => \N__6455\,
            I => \N__6428\
        );

    \I__1467\ : Span4Mux_v
    port map (
            O => \N__6452\,
            I => \N__6424\
        );

    \I__1466\ : Span4Mux_v
    port map (
            O => \N__6447\,
            I => \N__6421\
        );

    \I__1465\ : ClkMux
    port map (
            O => \N__6446\,
            I => \N__6418\
        );

    \I__1464\ : Span4Mux_v
    port map (
            O => \N__6443\,
            I => \N__6415\
        );

    \I__1463\ : Span4Mux_v
    port map (
            O => \N__6440\,
            I => \N__6410\
        );

    \I__1462\ : LocalMux
    port map (
            O => \N__6437\,
            I => \N__6410\
        );

    \I__1461\ : ClkMux
    port map (
            O => \N__6436\,
            I => \N__6407\
        );

    \I__1460\ : LocalMux
    port map (
            O => \N__6433\,
            I => \N__6404\
        );

    \I__1459\ : ClkMux
    port map (
            O => \N__6432\,
            I => \N__6401\
        );

    \I__1458\ : ClkMux
    port map (
            O => \N__6431\,
            I => \N__6398\
        );

    \I__1457\ : Span4Mux_v
    port map (
            O => \N__6428\,
            I => \N__6395\
        );

    \I__1456\ : ClkMux
    port map (
            O => \N__6427\,
            I => \N__6392\
        );

    \I__1455\ : Span4Mux_h
    port map (
            O => \N__6424\,
            I => \N__6384\
        );

    \I__1454\ : Span4Mux_h
    port map (
            O => \N__6421\,
            I => \N__6384\
        );

    \I__1453\ : LocalMux
    port map (
            O => \N__6418\,
            I => \N__6384\
        );

    \I__1452\ : Span4Mux_h
    port map (
            O => \N__6415\,
            I => \N__6381\
        );

    \I__1451\ : Span4Mux_v
    port map (
            O => \N__6410\,
            I => \N__6378\
        );

    \I__1450\ : LocalMux
    port map (
            O => \N__6407\,
            I => \N__6369\
        );

    \I__1449\ : Span4Mux_v
    port map (
            O => \N__6404\,
            I => \N__6369\
        );

    \I__1448\ : LocalMux
    port map (
            O => \N__6401\,
            I => \N__6369\
        );

    \I__1447\ : LocalMux
    port map (
            O => \N__6398\,
            I => \N__6369\
        );

    \I__1446\ : Sp12to4
    port map (
            O => \N__6395\,
            I => \N__6362\
        );

    \I__1445\ : LocalMux
    port map (
            O => \N__6392\,
            I => \N__6362\
        );

    \I__1444\ : ClkMux
    port map (
            O => \N__6391\,
            I => \N__6359\
        );

    \I__1443\ : Span4Mux_v
    port map (
            O => \N__6384\,
            I => \N__6356\
        );

    \I__1442\ : Span4Mux_v
    port map (
            O => \N__6381\,
            I => \N__6349\
        );

    \I__1441\ : Span4Mux_v
    port map (
            O => \N__6378\,
            I => \N__6349\
        );

    \I__1440\ : Span4Mux_v
    port map (
            O => \N__6369\,
            I => \N__6349\
        );

    \I__1439\ : ClkMux
    port map (
            O => \N__6368\,
            I => \N__6346\
        );

    \I__1438\ : InMux
    port map (
            O => \N__6367\,
            I => \N__6343\
        );

    \I__1437\ : Odrv12
    port map (
            O => \N__6362\,
            I => \eeprom.i2c.i2c_clk\
        );

    \I__1436\ : LocalMux
    port map (
            O => \N__6359\,
            I => \eeprom.i2c.i2c_clk\
        );

    \I__1435\ : Odrv4
    port map (
            O => \N__6356\,
            I => \eeprom.i2c.i2c_clk\
        );

    \I__1434\ : Odrv4
    port map (
            O => \N__6349\,
            I => \eeprom.i2c.i2c_clk\
        );

    \I__1433\ : LocalMux
    port map (
            O => \N__6346\,
            I => \eeprom.i2c.i2c_clk\
        );

    \I__1432\ : LocalMux
    port map (
            O => \N__6343\,
            I => \eeprom.i2c.i2c_clk\
        );

    \I__1431\ : IoInMux
    port map (
            O => \N__6330\,
            I => \N__6327\
        );

    \I__1430\ : LocalMux
    port map (
            O => \N__6327\,
            I => \N__6323\
        );

    \I__1429\ : InMux
    port map (
            O => \N__6326\,
            I => \N__6320\
        );

    \I__1428\ : IoSpan4Mux
    port map (
            O => \N__6323\,
            I => \N__6317\
        );

    \I__1427\ : LocalMux
    port map (
            O => \N__6320\,
            I => \N__6314\
        );

    \I__1426\ : Span4Mux_s3_h
    port map (
            O => \N__6317\,
            I => \N__6311\
        );

    \I__1425\ : Span4Mux_s3_h
    port map (
            O => \N__6314\,
            I => \N__6308\
        );

    \I__1424\ : Span4Mux_v
    port map (
            O => \N__6311\,
            I => \N__6303\
        );

    \I__1423\ : Span4Mux_v
    port map (
            O => \N__6308\,
            I => \N__6303\
        );

    \I__1422\ : Odrv4
    port map (
            O => \N__6303\,
            I => scl_enable
        );

    \I__1421\ : IoInMux
    port map (
            O => \N__6300\,
            I => \N__6297\
        );

    \I__1420\ : LocalMux
    port map (
            O => \N__6297\,
            I => scl_c
        );

    \I__1419\ : InMux
    port map (
            O => \N__6294\,
            I => \N__6290\
        );

    \I__1418\ : InMux
    port map (
            O => \N__6293\,
            I => \N__6287\
        );

    \I__1417\ : LocalMux
    port map (
            O => \N__6290\,
            I => \eeprom.i2c.counter_4\
        );

    \I__1416\ : LocalMux
    port map (
            O => \N__6287\,
            I => \eeprom.i2c.counter_4\
        );

    \I__1415\ : CascadeMux
    port map (
            O => \N__6282\,
            I => \eeprom.i2c.n12_cascade_\
        );

    \I__1414\ : InMux
    port map (
            O => \N__6279\,
            I => \N__6276\
        );

    \I__1413\ : LocalMux
    port map (
            O => \N__6276\,
            I => \N__6273\
        );

    \I__1412\ : Odrv4
    port map (
            O => \N__6273\,
            I => \eeprom.i2c.n1056\
        );

    \I__1411\ : InMux
    port map (
            O => \N__6270\,
            I => \N__6267\
        );

    \I__1410\ : LocalMux
    port map (
            O => \N__6267\,
            I => \eeprom.i2c.n1172\
        );

    \I__1409\ : InMux
    port map (
            O => \N__6264\,
            I => \N__6261\
        );

    \I__1408\ : LocalMux
    port map (
            O => \N__6261\,
            I => \eeprom.i2c.n3039\
        );

    \I__1407\ : CascadeMux
    port map (
            O => \N__6258\,
            I => \eeprom.i2c.n1056_cascade_\
        );

    \I__1406\ : InMux
    port map (
            O => \N__6255\,
            I => \N__6252\
        );

    \I__1405\ : LocalMux
    port map (
            O => \N__6252\,
            I => \N__6249\
        );

    \I__1404\ : Span4Mux_v
    port map (
            O => \N__6249\,
            I => \N__6245\
        );

    \I__1403\ : InMux
    port map (
            O => \N__6248\,
            I => \N__6242\
        );

    \I__1402\ : Odrv4
    port map (
            O => \N__6245\,
            I => \eeprom.i2c.n37\
        );

    \I__1401\ : LocalMux
    port map (
            O => \N__6242\,
            I => \eeprom.i2c.n37\
        );

    \I__1400\ : CascadeMux
    port map (
            O => \N__6237\,
            I => \N__6233\
        );

    \I__1399\ : CascadeMux
    port map (
            O => \N__6236\,
            I => \N__6230\
        );

    \I__1398\ : InMux
    port map (
            O => \N__6233\,
            I => \N__6221\
        );

    \I__1397\ : InMux
    port map (
            O => \N__6230\,
            I => \N__6221\
        );

    \I__1396\ : InMux
    port map (
            O => \N__6229\,
            I => \N__6221\
        );

    \I__1395\ : InMux
    port map (
            O => \N__6228\,
            I => \N__6218\
        );

    \I__1394\ : LocalMux
    port map (
            O => \N__6221\,
            I => \N__6215\
        );

    \I__1393\ : LocalMux
    port map (
            O => \N__6218\,
            I => \N__6211\
        );

    \I__1392\ : Span4Mux_h
    port map (
            O => \N__6215\,
            I => \N__6207\
        );

    \I__1391\ : InMux
    port map (
            O => \N__6214\,
            I => \N__6204\
        );

    \I__1390\ : Span4Mux_v
    port map (
            O => \N__6211\,
            I => \N__6201\
        );

    \I__1389\ : InMux
    port map (
            O => \N__6210\,
            I => \N__6198\
        );

    \I__1388\ : Odrv4
    port map (
            O => \N__6207\,
            I => \eeprom.i2c.counter_2\
        );

    \I__1387\ : LocalMux
    port map (
            O => \N__6204\,
            I => \eeprom.i2c.counter_2\
        );

    \I__1386\ : Odrv4
    port map (
            O => \N__6201\,
            I => \eeprom.i2c.counter_2\
        );

    \I__1385\ : LocalMux
    port map (
            O => \N__6198\,
            I => \eeprom.i2c.counter_2\
        );

    \I__1384\ : InMux
    port map (
            O => \N__6189\,
            I => \N__6179\
        );

    \I__1383\ : InMux
    port map (
            O => \N__6188\,
            I => \N__6179\
        );

    \I__1382\ : InMux
    port map (
            O => \N__6187\,
            I => \N__6179\
        );

    \I__1381\ : InMux
    port map (
            O => \N__6186\,
            I => \N__6175\
        );

    \I__1380\ : LocalMux
    port map (
            O => \N__6179\,
            I => \N__6172\
        );

    \I__1379\ : CascadeMux
    port map (
            O => \N__6178\,
            I => \N__6169\
        );

    \I__1378\ : LocalMux
    port map (
            O => \N__6175\,
            I => \N__6166\
        );

    \I__1377\ : Span4Mux_h
    port map (
            O => \N__6172\,
            I => \N__6162\
        );

    \I__1376\ : InMux
    port map (
            O => \N__6169\,
            I => \N__6159\
        );

    \I__1375\ : Span4Mux_h
    port map (
            O => \N__6166\,
            I => \N__6156\
        );

    \I__1374\ : InMux
    port map (
            O => \N__6165\,
            I => \N__6153\
        );

    \I__1373\ : Odrv4
    port map (
            O => \N__6162\,
            I => \eeprom.i2c.counter_1\
        );

    \I__1372\ : LocalMux
    port map (
            O => \N__6159\,
            I => \eeprom.i2c.counter_1\
        );

    \I__1371\ : Odrv4
    port map (
            O => \N__6156\,
            I => \eeprom.i2c.counter_1\
        );

    \I__1370\ : LocalMux
    port map (
            O => \N__6153\,
            I => \eeprom.i2c.counter_1\
        );

    \I__1369\ : InMux
    port map (
            O => \N__6144\,
            I => \N__6141\
        );

    \I__1368\ : LocalMux
    port map (
            O => \N__6141\,
            I => \N__6136\
        );

    \I__1367\ : InMux
    port map (
            O => \N__6140\,
            I => \N__6131\
        );

    \I__1366\ : InMux
    port map (
            O => \N__6139\,
            I => \N__6131\
        );

    \I__1365\ : Odrv12
    port map (
            O => \N__6136\,
            I => n4_adj_390
        );

    \I__1364\ : LocalMux
    port map (
            O => \N__6131\,
            I => n4_adj_390
        );

    \I__1363\ : InMux
    port map (
            O => \N__6126\,
            I => \N__6122\
        );

    \I__1362\ : CascadeMux
    port map (
            O => \N__6125\,
            I => \N__6118\
        );

    \I__1361\ : LocalMux
    port map (
            O => \N__6122\,
            I => \N__6113\
        );

    \I__1360\ : InMux
    port map (
            O => \N__6121\,
            I => \N__6110\
        );

    \I__1359\ : InMux
    port map (
            O => \N__6118\,
            I => \N__6107\
        );

    \I__1358\ : InMux
    port map (
            O => \N__6117\,
            I => \N__6102\
        );

    \I__1357\ : InMux
    port map (
            O => \N__6116\,
            I => \N__6098\
        );

    \I__1356\ : Span4Mux_v
    port map (
            O => \N__6113\,
            I => \N__6089\
        );

    \I__1355\ : LocalMux
    port map (
            O => \N__6110\,
            I => \N__6089\
        );

    \I__1354\ : LocalMux
    port map (
            O => \N__6107\,
            I => \N__6086\
        );

    \I__1353\ : InMux
    port map (
            O => \N__6106\,
            I => \N__6083\
        );

    \I__1352\ : InMux
    port map (
            O => \N__6105\,
            I => \N__6080\
        );

    \I__1351\ : LocalMux
    port map (
            O => \N__6102\,
            I => \N__6077\
        );

    \I__1350\ : CascadeMux
    port map (
            O => \N__6101\,
            I => \N__6071\
        );

    \I__1349\ : LocalMux
    port map (
            O => \N__6098\,
            I => \N__6067\
        );

    \I__1348\ : InMux
    port map (
            O => \N__6097\,
            I => \N__6060\
        );

    \I__1347\ : InMux
    port map (
            O => \N__6096\,
            I => \N__6060\
        );

    \I__1346\ : InMux
    port map (
            O => \N__6095\,
            I => \N__6060\
        );

    \I__1345\ : InMux
    port map (
            O => \N__6094\,
            I => \N__6052\
        );

    \I__1344\ : Span4Mux_h
    port map (
            O => \N__6089\,
            I => \N__6049\
        );

    \I__1343\ : Span4Mux_h
    port map (
            O => \N__6086\,
            I => \N__6040\
        );

    \I__1342\ : LocalMux
    port map (
            O => \N__6083\,
            I => \N__6040\
        );

    \I__1341\ : LocalMux
    port map (
            O => \N__6080\,
            I => \N__6040\
        );

    \I__1340\ : Span4Mux_h
    port map (
            O => \N__6077\,
            I => \N__6040\
        );

    \I__1339\ : InMux
    port map (
            O => \N__6076\,
            I => \N__6033\
        );

    \I__1338\ : InMux
    port map (
            O => \N__6075\,
            I => \N__6033\
        );

    \I__1337\ : InMux
    port map (
            O => \N__6074\,
            I => \N__6033\
        );

    \I__1336\ : InMux
    port map (
            O => \N__6071\,
            I => \N__6028\
        );

    \I__1335\ : InMux
    port map (
            O => \N__6070\,
            I => \N__6028\
        );

    \I__1334\ : Span4Mux_h
    port map (
            O => \N__6067\,
            I => \N__6023\
        );

    \I__1333\ : LocalMux
    port map (
            O => \N__6060\,
            I => \N__6023\
        );

    \I__1332\ : InMux
    port map (
            O => \N__6059\,
            I => \N__6020\
        );

    \I__1331\ : InMux
    port map (
            O => \N__6058\,
            I => \N__6011\
        );

    \I__1330\ : InMux
    port map (
            O => \N__6057\,
            I => \N__6011\
        );

    \I__1329\ : InMux
    port map (
            O => \N__6056\,
            I => \N__6011\
        );

    \I__1328\ : InMux
    port map (
            O => \N__6055\,
            I => \N__6011\
        );

    \I__1327\ : LocalMux
    port map (
            O => \N__6052\,
            I => \eeprom.state_1_adj_386\
        );

    \I__1326\ : Odrv4
    port map (
            O => \N__6049\,
            I => \eeprom.state_1_adj_386\
        );

    \I__1325\ : Odrv4
    port map (
            O => \N__6040\,
            I => \eeprom.state_1_adj_386\
        );

    \I__1324\ : LocalMux
    port map (
            O => \N__6033\,
            I => \eeprom.state_1_adj_386\
        );

    \I__1323\ : LocalMux
    port map (
            O => \N__6028\,
            I => \eeprom.state_1_adj_386\
        );

    \I__1322\ : Odrv4
    port map (
            O => \N__6023\,
            I => \eeprom.state_1_adj_386\
        );

    \I__1321\ : LocalMux
    port map (
            O => \N__6020\,
            I => \eeprom.state_1_adj_386\
        );

    \I__1320\ : LocalMux
    port map (
            O => \N__6011\,
            I => \eeprom.state_1_adj_386\
        );

    \I__1319\ : InMux
    port map (
            O => \N__5994\,
            I => \N__5990\
        );

    \I__1318\ : InMux
    port map (
            O => \N__5993\,
            I => \N__5984\
        );

    \I__1317\ : LocalMux
    port map (
            O => \N__5990\,
            I => \N__5981\
        );

    \I__1316\ : InMux
    port map (
            O => \N__5989\,
            I => \N__5976\
        );

    \I__1315\ : InMux
    port map (
            O => \N__5988\,
            I => \N__5976\
        );

    \I__1314\ : InMux
    port map (
            O => \N__5987\,
            I => \N__5972\
        );

    \I__1313\ : LocalMux
    port map (
            O => \N__5984\,
            I => \N__5968\
        );

    \I__1312\ : Span4Mux_v
    port map (
            O => \N__5981\,
            I => \N__5961\
        );

    \I__1311\ : LocalMux
    port map (
            O => \N__5976\,
            I => \N__5961\
        );

    \I__1310\ : CascadeMux
    port map (
            O => \N__5975\,
            I => \N__5954\
        );

    \I__1309\ : LocalMux
    port map (
            O => \N__5972\,
            I => \N__5945\
        );

    \I__1308\ : InMux
    port map (
            O => \N__5971\,
            I => \N__5942\
        );

    \I__1307\ : Span4Mux_h
    port map (
            O => \N__5968\,
            I => \N__5939\
        );

    \I__1306\ : InMux
    port map (
            O => \N__5967\,
            I => \N__5934\
        );

    \I__1305\ : InMux
    port map (
            O => \N__5966\,
            I => \N__5934\
        );

    \I__1304\ : Span4Mux_h
    port map (
            O => \N__5961\,
            I => \N__5931\
        );

    \I__1303\ : InMux
    port map (
            O => \N__5960\,
            I => \N__5926\
        );

    \I__1302\ : InMux
    port map (
            O => \N__5959\,
            I => \N__5926\
        );

    \I__1301\ : InMux
    port map (
            O => \N__5958\,
            I => \N__5915\
        );

    \I__1300\ : InMux
    port map (
            O => \N__5957\,
            I => \N__5915\
        );

    \I__1299\ : InMux
    port map (
            O => \N__5954\,
            I => \N__5915\
        );

    \I__1298\ : InMux
    port map (
            O => \N__5953\,
            I => \N__5915\
        );

    \I__1297\ : InMux
    port map (
            O => \N__5952\,
            I => \N__5915\
        );

    \I__1296\ : InMux
    port map (
            O => \N__5951\,
            I => \N__5912\
        );

    \I__1295\ : InMux
    port map (
            O => \N__5950\,
            I => \N__5909\
        );

    \I__1294\ : InMux
    port map (
            O => \N__5949\,
            I => \N__5904\
        );

    \I__1293\ : InMux
    port map (
            O => \N__5948\,
            I => \N__5904\
        );

    \I__1292\ : Odrv12
    port map (
            O => \N__5945\,
            I => \eeprom.state_3\
        );

    \I__1291\ : LocalMux
    port map (
            O => \N__5942\,
            I => \eeprom.state_3\
        );

    \I__1290\ : Odrv4
    port map (
            O => \N__5939\,
            I => \eeprom.state_3\
        );

    \I__1289\ : LocalMux
    port map (
            O => \N__5934\,
            I => \eeprom.state_3\
        );

    \I__1288\ : Odrv4
    port map (
            O => \N__5931\,
            I => \eeprom.state_3\
        );

    \I__1287\ : LocalMux
    port map (
            O => \N__5926\,
            I => \eeprom.state_3\
        );

    \I__1286\ : LocalMux
    port map (
            O => \N__5915\,
            I => \eeprom.state_3\
        );

    \I__1285\ : LocalMux
    port map (
            O => \N__5912\,
            I => \eeprom.state_3\
        );

    \I__1284\ : LocalMux
    port map (
            O => \N__5909\,
            I => \eeprom.state_3\
        );

    \I__1283\ : LocalMux
    port map (
            O => \N__5904\,
            I => \eeprom.state_3\
        );

    \I__1282\ : CascadeMux
    port map (
            O => \N__5883\,
            I => \N__5877\
        );

    \I__1281\ : InMux
    port map (
            O => \N__5882\,
            I => \N__5871\
        );

    \I__1280\ : InMux
    port map (
            O => \N__5881\,
            I => \N__5868\
        );

    \I__1279\ : InMux
    port map (
            O => \N__5880\,
            I => \N__5863\
        );

    \I__1278\ : InMux
    port map (
            O => \N__5877\,
            I => \N__5860\
        );

    \I__1277\ : InMux
    port map (
            O => \N__5876\,
            I => \N__5853\
        );

    \I__1276\ : InMux
    port map (
            O => \N__5875\,
            I => \N__5853\
        );

    \I__1275\ : CascadeMux
    port map (
            O => \N__5874\,
            I => \N__5848\
        );

    \I__1274\ : LocalMux
    port map (
            O => \N__5871\,
            I => \N__5842\
        );

    \I__1273\ : LocalMux
    port map (
            O => \N__5868\,
            I => \N__5839\
        );

    \I__1272\ : InMux
    port map (
            O => \N__5867\,
            I => \N__5836\
        );

    \I__1271\ : CascadeMux
    port map (
            O => \N__5866\,
            I => \N__5832\
        );

    \I__1270\ : LocalMux
    port map (
            O => \N__5863\,
            I => \N__5829\
        );

    \I__1269\ : LocalMux
    port map (
            O => \N__5860\,
            I => \N__5826\
        );

    \I__1268\ : InMux
    port map (
            O => \N__5859\,
            I => \N__5823\
        );

    \I__1267\ : InMux
    port map (
            O => \N__5858\,
            I => \N__5820\
        );

    \I__1266\ : LocalMux
    port map (
            O => \N__5853\,
            I => \N__5817\
        );

    \I__1265\ : InMux
    port map (
            O => \N__5852\,
            I => \N__5808\
        );

    \I__1264\ : InMux
    port map (
            O => \N__5851\,
            I => \N__5808\
        );

    \I__1263\ : InMux
    port map (
            O => \N__5848\,
            I => \N__5808\
        );

    \I__1262\ : InMux
    port map (
            O => \N__5847\,
            I => \N__5808\
        );

    \I__1261\ : InMux
    port map (
            O => \N__5846\,
            I => \N__5805\
        );

    \I__1260\ : CascadeMux
    port map (
            O => \N__5845\,
            I => \N__5798\
        );

    \I__1259\ : Span4Mux_v
    port map (
            O => \N__5842\,
            I => \N__5792\
        );

    \I__1258\ : Span4Mux_v
    port map (
            O => \N__5839\,
            I => \N__5792\
        );

    \I__1257\ : LocalMux
    port map (
            O => \N__5836\,
            I => \N__5789\
        );

    \I__1256\ : InMux
    port map (
            O => \N__5835\,
            I => \N__5786\
        );

    \I__1255\ : InMux
    port map (
            O => \N__5832\,
            I => \N__5783\
        );

    \I__1254\ : Span4Mux_v
    port map (
            O => \N__5829\,
            I => \N__5778\
        );

    \I__1253\ : Span4Mux_v
    port map (
            O => \N__5826\,
            I => \N__5778\
        );

    \I__1252\ : LocalMux
    port map (
            O => \N__5823\,
            I => \N__5775\
        );

    \I__1251\ : LocalMux
    port map (
            O => \N__5820\,
            I => \N__5766\
        );

    \I__1250\ : Span4Mux_h
    port map (
            O => \N__5817\,
            I => \N__5766\
        );

    \I__1249\ : LocalMux
    port map (
            O => \N__5808\,
            I => \N__5766\
        );

    \I__1248\ : LocalMux
    port map (
            O => \N__5805\,
            I => \N__5766\
        );

    \I__1247\ : InMux
    port map (
            O => \N__5804\,
            I => \N__5761\
        );

    \I__1246\ : InMux
    port map (
            O => \N__5803\,
            I => \N__5761\
        );

    \I__1245\ : InMux
    port map (
            O => \N__5802\,
            I => \N__5758\
        );

    \I__1244\ : InMux
    port map (
            O => \N__5801\,
            I => \N__5751\
        );

    \I__1243\ : InMux
    port map (
            O => \N__5798\,
            I => \N__5751\
        );

    \I__1242\ : InMux
    port map (
            O => \N__5797\,
            I => \N__5751\
        );

    \I__1241\ : Odrv4
    port map (
            O => \N__5792\,
            I => \eeprom.state_0_adj_384\
        );

    \I__1240\ : Odrv12
    port map (
            O => \N__5789\,
            I => \eeprom.state_0_adj_384\
        );

    \I__1239\ : LocalMux
    port map (
            O => \N__5786\,
            I => \eeprom.state_0_adj_384\
        );

    \I__1238\ : LocalMux
    port map (
            O => \N__5783\,
            I => \eeprom.state_0_adj_384\
        );

    \I__1237\ : Odrv4
    port map (
            O => \N__5778\,
            I => \eeprom.state_0_adj_384\
        );

    \I__1236\ : Odrv4
    port map (
            O => \N__5775\,
            I => \eeprom.state_0_adj_384\
        );

    \I__1235\ : Odrv4
    port map (
            O => \N__5766\,
            I => \eeprom.state_0_adj_384\
        );

    \I__1234\ : LocalMux
    port map (
            O => \N__5761\,
            I => \eeprom.state_0_adj_384\
        );

    \I__1233\ : LocalMux
    port map (
            O => \N__5758\,
            I => \eeprom.state_0_adj_384\
        );

    \I__1232\ : LocalMux
    port map (
            O => \N__5751\,
            I => \eeprom.state_0_adj_384\
        );

    \I__1231\ : InMux
    port map (
            O => \N__5730\,
            I => \N__5718\
        );

    \I__1230\ : InMux
    port map (
            O => \N__5729\,
            I => \N__5718\
        );

    \I__1229\ : InMux
    port map (
            O => \N__5728\,
            I => \N__5715\
        );

    \I__1228\ : InMux
    port map (
            O => \N__5727\,
            I => \N__5710\
        );

    \I__1227\ : InMux
    port map (
            O => \N__5726\,
            I => \N__5710\
        );

    \I__1226\ : InMux
    port map (
            O => \N__5725\,
            I => \N__5706\
        );

    \I__1225\ : InMux
    port map (
            O => \N__5724\,
            I => \N__5697\
        );

    \I__1224\ : InMux
    port map (
            O => \N__5723\,
            I => \N__5694\
        );

    \I__1223\ : LocalMux
    port map (
            O => \N__5718\,
            I => \N__5691\
        );

    \I__1222\ : LocalMux
    port map (
            O => \N__5715\,
            I => \N__5683\
        );

    \I__1221\ : LocalMux
    port map (
            O => \N__5710\,
            I => \N__5683\
        );

    \I__1220\ : InMux
    port map (
            O => \N__5709\,
            I => \N__5680\
        );

    \I__1219\ : LocalMux
    port map (
            O => \N__5706\,
            I => \N__5677\
        );

    \I__1218\ : InMux
    port map (
            O => \N__5705\,
            I => \N__5666\
        );

    \I__1217\ : InMux
    port map (
            O => \N__5704\,
            I => \N__5666\
        );

    \I__1216\ : InMux
    port map (
            O => \N__5703\,
            I => \N__5666\
        );

    \I__1215\ : InMux
    port map (
            O => \N__5702\,
            I => \N__5666\
        );

    \I__1214\ : InMux
    port map (
            O => \N__5701\,
            I => \N__5666\
        );

    \I__1213\ : InMux
    port map (
            O => \N__5700\,
            I => \N__5660\
        );

    \I__1212\ : LocalMux
    port map (
            O => \N__5697\,
            I => \N__5657\
        );

    \I__1211\ : LocalMux
    port map (
            O => \N__5694\,
            I => \N__5652\
        );

    \I__1210\ : Span4Mux_h
    port map (
            O => \N__5691\,
            I => \N__5652\
        );

    \I__1209\ : InMux
    port map (
            O => \N__5690\,
            I => \N__5649\
        );

    \I__1208\ : InMux
    port map (
            O => \N__5689\,
            I => \N__5644\
        );

    \I__1207\ : InMux
    port map (
            O => \N__5688\,
            I => \N__5644\
        );

    \I__1206\ : Span4Mux_v
    port map (
            O => \N__5683\,
            I => \N__5641\
        );

    \I__1205\ : LocalMux
    port map (
            O => \N__5680\,
            I => \N__5634\
        );

    \I__1204\ : Span4Mux_h
    port map (
            O => \N__5677\,
            I => \N__5634\
        );

    \I__1203\ : LocalMux
    port map (
            O => \N__5666\,
            I => \N__5634\
        );

    \I__1202\ : InMux
    port map (
            O => \N__5665\,
            I => \N__5627\
        );

    \I__1201\ : InMux
    port map (
            O => \N__5664\,
            I => \N__5627\
        );

    \I__1200\ : InMux
    port map (
            O => \N__5663\,
            I => \N__5627\
        );

    \I__1199\ : LocalMux
    port map (
            O => \N__5660\,
            I => \eeprom.i2c.state_2\
        );

    \I__1198\ : Odrv4
    port map (
            O => \N__5657\,
            I => \eeprom.i2c.state_2\
        );

    \I__1197\ : Odrv4
    port map (
            O => \N__5652\,
            I => \eeprom.i2c.state_2\
        );

    \I__1196\ : LocalMux
    port map (
            O => \N__5649\,
            I => \eeprom.i2c.state_2\
        );

    \I__1195\ : LocalMux
    port map (
            O => \N__5644\,
            I => \eeprom.i2c.state_2\
        );

    \I__1194\ : Odrv4
    port map (
            O => \N__5641\,
            I => \eeprom.i2c.state_2\
        );

    \I__1193\ : Odrv4
    port map (
            O => \N__5634\,
            I => \eeprom.i2c.state_2\
        );

    \I__1192\ : LocalMux
    port map (
            O => \N__5627\,
            I => \eeprom.i2c.state_2\
        );

    \I__1191\ : InMux
    port map (
            O => \N__5610\,
            I => \N__5606\
        );

    \I__1190\ : InMux
    port map (
            O => \N__5609\,
            I => \N__5603\
        );

    \I__1189\ : LocalMux
    port map (
            O => \N__5606\,
            I => \eeprom.i2c.counter2_0\
        );

    \I__1188\ : LocalMux
    port map (
            O => \N__5603\,
            I => \eeprom.i2c.counter2_0\
        );

    \I__1187\ : InMux
    port map (
            O => \N__5598\,
            I => \bfn_27_13_0_\
        );

    \I__1186\ : InMux
    port map (
            O => \N__5595\,
            I => \N__5591\
        );

    \I__1185\ : InMux
    port map (
            O => \N__5594\,
            I => \N__5588\
        );

    \I__1184\ : LocalMux
    port map (
            O => \N__5591\,
            I => \eeprom.i2c.counter2_1\
        );

    \I__1183\ : LocalMux
    port map (
            O => \N__5588\,
            I => \eeprom.i2c.counter2_1\
        );

    \I__1182\ : InMux
    port map (
            O => \N__5583\,
            I => \eeprom.i2c.n2871\
        );

    \I__1181\ : InMux
    port map (
            O => \N__5580\,
            I => \N__5576\
        );

    \I__1180\ : InMux
    port map (
            O => \N__5579\,
            I => \N__5573\
        );

    \I__1179\ : LocalMux
    port map (
            O => \N__5576\,
            I => \eeprom.i2c.counter2_2\
        );

    \I__1178\ : LocalMux
    port map (
            O => \N__5573\,
            I => \eeprom.i2c.counter2_2\
        );

    \I__1177\ : InMux
    port map (
            O => \N__5568\,
            I => \eeprom.i2c.n2872\
        );

    \I__1176\ : InMux
    port map (
            O => \N__5565\,
            I => \N__5561\
        );

    \I__1175\ : InMux
    port map (
            O => \N__5564\,
            I => \N__5558\
        );

    \I__1174\ : LocalMux
    port map (
            O => \N__5561\,
            I => \eeprom.i2c.counter2_3\
        );

    \I__1173\ : LocalMux
    port map (
            O => \N__5558\,
            I => \eeprom.i2c.counter2_3\
        );

    \I__1172\ : InMux
    port map (
            O => \N__5553\,
            I => \eeprom.i2c.n2873\
        );

    \I__1171\ : InMux
    port map (
            O => \N__5550\,
            I => \eeprom.i2c.n2853\
        );

    \I__1170\ : InMux
    port map (
            O => \N__5547\,
            I => \eeprom.i2c.n2854\
        );

    \I__1169\ : InMux
    port map (
            O => \N__5544\,
            I => \eeprom.i2c.n2855\
        );

    \I__1168\ : InMux
    port map (
            O => \N__5541\,
            I => \N__5537\
        );

    \I__1167\ : CascadeMux
    port map (
            O => \N__5540\,
            I => \N__5534\
        );

    \I__1166\ : LocalMux
    port map (
            O => \N__5537\,
            I => \N__5527\
        );

    \I__1165\ : InMux
    port map (
            O => \N__5534\,
            I => \N__5524\
        );

    \I__1164\ : CascadeMux
    port map (
            O => \N__5533\,
            I => \N__5520\
        );

    \I__1163\ : CascadeMux
    port map (
            O => \N__5532\,
            I => \N__5517\
        );

    \I__1162\ : CascadeMux
    port map (
            O => \N__5531\,
            I => \N__5514\
        );

    \I__1161\ : InMux
    port map (
            O => \N__5530\,
            I => \N__5510\
        );

    \I__1160\ : Span4Mux_v
    port map (
            O => \N__5527\,
            I => \N__5507\
        );

    \I__1159\ : LocalMux
    port map (
            O => \N__5524\,
            I => \N__5504\
        );

    \I__1158\ : InMux
    port map (
            O => \N__5523\,
            I => \N__5501\
        );

    \I__1157\ : InMux
    port map (
            O => \N__5520\,
            I => \N__5496\
        );

    \I__1156\ : InMux
    port map (
            O => \N__5517\,
            I => \N__5496\
        );

    \I__1155\ : InMux
    port map (
            O => \N__5514\,
            I => \N__5493\
        );

    \I__1154\ : InMux
    port map (
            O => \N__5513\,
            I => \N__5490\
        );

    \I__1153\ : LocalMux
    port map (
            O => \N__5510\,
            I => \N__5487\
        );

    \I__1152\ : Odrv4
    port map (
            O => \N__5507\,
            I => \eeprom.n10\
        );

    \I__1151\ : Odrv4
    port map (
            O => \N__5504\,
            I => \eeprom.n10\
        );

    \I__1150\ : LocalMux
    port map (
            O => \N__5501\,
            I => \eeprom.n10\
        );

    \I__1149\ : LocalMux
    port map (
            O => \N__5496\,
            I => \eeprom.n10\
        );

    \I__1148\ : LocalMux
    port map (
            O => \N__5493\,
            I => \eeprom.n10\
        );

    \I__1147\ : LocalMux
    port map (
            O => \N__5490\,
            I => \eeprom.n10\
        );

    \I__1146\ : Odrv12
    port map (
            O => \N__5487\,
            I => \eeprom.n10\
        );

    \I__1145\ : InMux
    port map (
            O => \N__5472\,
            I => \N__5469\
        );

    \I__1144\ : LocalMux
    port map (
            O => \N__5469\,
            I => \N__5465\
        );

    \I__1143\ : InMux
    port map (
            O => \N__5468\,
            I => \N__5462\
        );

    \I__1142\ : Odrv4
    port map (
            O => \N__5465\,
            I => \eeprom.i2c.n9_adj_377\
        );

    \I__1141\ : LocalMux
    port map (
            O => \N__5462\,
            I => \eeprom.i2c.n9_adj_377\
        );

    \I__1140\ : CascadeMux
    port map (
            O => \N__5457\,
            I => \eeprom.i2c.n3039_cascade_\
        );

    \I__1139\ : InMux
    port map (
            O => \N__5454\,
            I => \N__5450\
        );

    \I__1138\ : CascadeMux
    port map (
            O => \N__5453\,
            I => \N__5447\
        );

    \I__1137\ : LocalMux
    port map (
            O => \N__5450\,
            I => \N__5439\
        );

    \I__1136\ : InMux
    port map (
            O => \N__5447\,
            I => \N__5436\
        );

    \I__1135\ : CascadeMux
    port map (
            O => \N__5446\,
            I => \N__5433\
        );

    \I__1134\ : CascadeMux
    port map (
            O => \N__5445\,
            I => \N__5429\
        );

    \I__1133\ : CascadeMux
    port map (
            O => \N__5444\,
            I => \N__5426\
        );

    \I__1132\ : CascadeMux
    port map (
            O => \N__5443\,
            I => \N__5423\
        );

    \I__1131\ : CascadeMux
    port map (
            O => \N__5442\,
            I => \N__5419\
        );

    \I__1130\ : Span4Mux_v
    port map (
            O => \N__5439\,
            I => \N__5415\
        );

    \I__1129\ : LocalMux
    port map (
            O => \N__5436\,
            I => \N__5412\
        );

    \I__1128\ : InMux
    port map (
            O => \N__5433\,
            I => \N__5405\
        );

    \I__1127\ : InMux
    port map (
            O => \N__5432\,
            I => \N__5405\
        );

    \I__1126\ : InMux
    port map (
            O => \N__5429\,
            I => \N__5400\
        );

    \I__1125\ : InMux
    port map (
            O => \N__5426\,
            I => \N__5400\
        );

    \I__1124\ : InMux
    port map (
            O => \N__5423\,
            I => \N__5397\
        );

    \I__1123\ : InMux
    port map (
            O => \N__5422\,
            I => \N__5392\
        );

    \I__1122\ : InMux
    port map (
            O => \N__5419\,
            I => \N__5392\
        );

    \I__1121\ : InMux
    port map (
            O => \N__5418\,
            I => \N__5389\
        );

    \I__1120\ : Span4Mux_v
    port map (
            O => \N__5415\,
            I => \N__5386\
        );

    \I__1119\ : Span4Mux_h
    port map (
            O => \N__5412\,
            I => \N__5383\
        );

    \I__1118\ : InMux
    port map (
            O => \N__5411\,
            I => \N__5380\
        );

    \I__1117\ : InMux
    port map (
            O => \N__5410\,
            I => \N__5377\
        );

    \I__1116\ : LocalMux
    port map (
            O => \N__5405\,
            I => \N__5366\
        );

    \I__1115\ : LocalMux
    port map (
            O => \N__5400\,
            I => \N__5366\
        );

    \I__1114\ : LocalMux
    port map (
            O => \N__5397\,
            I => \N__5366\
        );

    \I__1113\ : LocalMux
    port map (
            O => \N__5392\,
            I => \N__5366\
        );

    \I__1112\ : LocalMux
    port map (
            O => \N__5389\,
            I => \N__5366\
        );

    \I__1111\ : Span4Mux_v
    port map (
            O => \N__5386\,
            I => \N__5363\
        );

    \I__1110\ : Sp12to4
    port map (
            O => \N__5383\,
            I => \N__5356\
        );

    \I__1109\ : LocalMux
    port map (
            O => \N__5380\,
            I => \N__5356\
        );

    \I__1108\ : LocalMux
    port map (
            O => \N__5377\,
            I => \N__5356\
        );

    \I__1107\ : Span12Mux_v
    port map (
            O => \N__5366\,
            I => \N__5353\
        );

    \I__1106\ : Sp12to4
    port map (
            O => \N__5363\,
            I => \N__5348\
        );

    \I__1105\ : Span12Mux_v
    port map (
            O => \N__5356\,
            I => \N__5348\
        );

    \I__1104\ : Odrv12
    port map (
            O => \N__5353\,
            I => \state_7_N_286_3\
        );

    \I__1103\ : Odrv12
    port map (
            O => \N__5348\,
            I => \state_7_N_286_3\
        );

    \I__1102\ : InMux
    port map (
            O => \N__5343\,
            I => \N__5338\
        );

    \I__1101\ : InMux
    port map (
            O => \N__5342\,
            I => \N__5332\
        );

    \I__1100\ : InMux
    port map (
            O => \N__5341\,
            I => \N__5332\
        );

    \I__1099\ : LocalMux
    port map (
            O => \N__5338\,
            I => \N__5329\
        );

    \I__1098\ : CascadeMux
    port map (
            O => \N__5337\,
            I => \N__5326\
        );

    \I__1097\ : LocalMux
    port map (
            O => \N__5332\,
            I => \N__5323\
        );

    \I__1096\ : Span4Mux_h
    port map (
            O => \N__5329\,
            I => \N__5320\
        );

    \I__1095\ : InMux
    port map (
            O => \N__5326\,
            I => \N__5317\
        );

    \I__1094\ : Odrv12
    port map (
            O => \N__5323\,
            I => n1723
        );

    \I__1093\ : Odrv4
    port map (
            O => \N__5320\,
            I => n1723
        );

    \I__1092\ : LocalMux
    port map (
            O => \N__5317\,
            I => n1723
        );

    \I__1091\ : InMux
    port map (
            O => \N__5310\,
            I => \N__5307\
        );

    \I__1090\ : LocalMux
    port map (
            O => \N__5307\,
            I => \N__5304\
        );

    \I__1089\ : Span4Mux_h
    port map (
            O => \N__5304\,
            I => \N__5300\
        );

    \I__1088\ : InMux
    port map (
            O => \N__5303\,
            I => \N__5297\
        );

    \I__1087\ : Odrv4
    port map (
            O => \N__5300\,
            I => data_1
        );

    \I__1086\ : LocalMux
    port map (
            O => \N__5297\,
            I => data_1
        );

    \I__1085\ : InMux
    port map (
            O => \N__5292\,
            I => \N__5288\
        );

    \I__1084\ : InMux
    port map (
            O => \N__5291\,
            I => \N__5285\
        );

    \I__1083\ : LocalMux
    port map (
            O => \N__5288\,
            I => \eeprom.i2c.counter_6\
        );

    \I__1082\ : LocalMux
    port map (
            O => \N__5285\,
            I => \eeprom.i2c.counter_6\
        );

    \I__1081\ : CascadeMux
    port map (
            O => \N__5280\,
            I => \N__5277\
        );

    \I__1080\ : InMux
    port map (
            O => \N__5277\,
            I => \N__5273\
        );

    \I__1079\ : InMux
    port map (
            O => \N__5276\,
            I => \N__5270\
        );

    \I__1078\ : LocalMux
    port map (
            O => \N__5273\,
            I => \eeprom.i2c.counter_3\
        );

    \I__1077\ : LocalMux
    port map (
            O => \N__5270\,
            I => \eeprom.i2c.counter_3\
        );

    \I__1076\ : CascadeMux
    port map (
            O => \N__5265\,
            I => \N__5261\
        );

    \I__1075\ : CascadeMux
    port map (
            O => \N__5264\,
            I => \N__5258\
        );

    \I__1074\ : InMux
    port map (
            O => \N__5261\,
            I => \N__5255\
        );

    \I__1073\ : InMux
    port map (
            O => \N__5258\,
            I => \N__5252\
        );

    \I__1072\ : LocalMux
    port map (
            O => \N__5255\,
            I => \eeprom.i2c.counter_5\
        );

    \I__1071\ : LocalMux
    port map (
            O => \N__5252\,
            I => \eeprom.i2c.counter_5\
        );

    \I__1070\ : InMux
    port map (
            O => \N__5247\,
            I => \N__5243\
        );

    \I__1069\ : InMux
    port map (
            O => \N__5246\,
            I => \N__5240\
        );

    \I__1068\ : LocalMux
    port map (
            O => \N__5243\,
            I => \eeprom.i2c.counter_7\
        );

    \I__1067\ : LocalMux
    port map (
            O => \N__5240\,
            I => \eeprom.i2c.counter_7\
        );

    \I__1066\ : InMux
    port map (
            O => \N__5235\,
            I => \N__5229\
        );

    \I__1065\ : InMux
    port map (
            O => \N__5234\,
            I => \N__5226\
        );

    \I__1064\ : InMux
    port map (
            O => \N__5233\,
            I => \N__5221\
        );

    \I__1063\ : InMux
    port map (
            O => \N__5232\,
            I => \N__5221\
        );

    \I__1062\ : LocalMux
    port map (
            O => \N__5229\,
            I => \eeprom.n9\
        );

    \I__1061\ : LocalMux
    port map (
            O => \N__5226\,
            I => \eeprom.n9\
        );

    \I__1060\ : LocalMux
    port map (
            O => \N__5221\,
            I => \eeprom.n9\
        );

    \I__1059\ : SRMux
    port map (
            O => \N__5214\,
            I => \N__5211\
        );

    \I__1058\ : LocalMux
    port map (
            O => \N__5211\,
            I => \N__5205\
        );

    \I__1057\ : InMux
    port map (
            O => \N__5210\,
            I => \N__5202\
        );

    \I__1056\ : InMux
    port map (
            O => \N__5209\,
            I => \N__5197\
        );

    \I__1055\ : InMux
    port map (
            O => \N__5208\,
            I => \N__5197\
        );

    \I__1054\ : Span4Mux_h
    port map (
            O => \N__5205\,
            I => \N__5192\
        );

    \I__1053\ : LocalMux
    port map (
            O => \N__5202\,
            I => \N__5192\
        );

    \I__1052\ : LocalMux
    port map (
            O => \N__5197\,
            I => \N__5183\
        );

    \I__1051\ : Span4Mux_v
    port map (
            O => \N__5192\,
            I => \N__5180\
        );

    \I__1050\ : InMux
    port map (
            O => \N__5191\,
            I => \N__5177\
        );

    \I__1049\ : InMux
    port map (
            O => \N__5190\,
            I => \N__5166\
        );

    \I__1048\ : InMux
    port map (
            O => \N__5189\,
            I => \N__5166\
        );

    \I__1047\ : InMux
    port map (
            O => \N__5188\,
            I => \N__5166\
        );

    \I__1046\ : InMux
    port map (
            O => \N__5187\,
            I => \N__5166\
        );

    \I__1045\ : InMux
    port map (
            O => \N__5186\,
            I => \N__5166\
        );

    \I__1044\ : Span4Mux_h
    port map (
            O => \N__5183\,
            I => \N__5163\
        );

    \I__1043\ : Odrv4
    port map (
            O => \N__5180\,
            I => state_1
        );

    \I__1042\ : LocalMux
    port map (
            O => \N__5177\,
            I => state_1
        );

    \I__1041\ : LocalMux
    port map (
            O => \N__5166\,
            I => state_1
        );

    \I__1040\ : Odrv4
    port map (
            O => \N__5163\,
            I => state_1
        );

    \I__1039\ : CascadeMux
    port map (
            O => \N__5154\,
            I => \N__5146\
        );

    \I__1038\ : InMux
    port map (
            O => \N__5153\,
            I => \N__5143\
        );

    \I__1037\ : InMux
    port map (
            O => \N__5152\,
            I => \N__5134\
        );

    \I__1036\ : InMux
    port map (
            O => \N__5151\,
            I => \N__5134\
        );

    \I__1035\ : InMux
    port map (
            O => \N__5150\,
            I => \N__5134\
        );

    \I__1034\ : InMux
    port map (
            O => \N__5149\,
            I => \N__5134\
        );

    \I__1033\ : InMux
    port map (
            O => \N__5146\,
            I => \N__5130\
        );

    \I__1032\ : LocalMux
    port map (
            O => \N__5143\,
            I => \N__5127\
        );

    \I__1031\ : LocalMux
    port map (
            O => \N__5134\,
            I => \N__5118\
        );

    \I__1030\ : InMux
    port map (
            O => \N__5133\,
            I => \N__5115\
        );

    \I__1029\ : LocalMux
    port map (
            O => \N__5130\,
            I => \N__5112\
        );

    \I__1028\ : Span4Mux_h
    port map (
            O => \N__5127\,
            I => \N__5109\
        );

    \I__1027\ : InMux
    port map (
            O => \N__5126\,
            I => \N__5096\
        );

    \I__1026\ : InMux
    port map (
            O => \N__5125\,
            I => \N__5096\
        );

    \I__1025\ : InMux
    port map (
            O => \N__5124\,
            I => \N__5096\
        );

    \I__1024\ : InMux
    port map (
            O => \N__5123\,
            I => \N__5096\
        );

    \I__1023\ : InMux
    port map (
            O => \N__5122\,
            I => \N__5096\
        );

    \I__1022\ : InMux
    port map (
            O => \N__5121\,
            I => \N__5096\
        );

    \I__1021\ : Span4Mux_h
    port map (
            O => \N__5118\,
            I => \N__5093\
        );

    \I__1020\ : LocalMux
    port map (
            O => \N__5115\,
            I => state_0
        );

    \I__1019\ : Odrv4
    port map (
            O => \N__5112\,
            I => state_0
        );

    \I__1018\ : Odrv4
    port map (
            O => \N__5109\,
            I => state_0
        );

    \I__1017\ : LocalMux
    port map (
            O => \N__5096\,
            I => state_0
        );

    \I__1016\ : Odrv4
    port map (
            O => \N__5093\,
            I => state_0
        );

    \I__1015\ : CEMux
    port map (
            O => \N__5082\,
            I => \N__5079\
        );

    \I__1014\ : LocalMux
    port map (
            O => \N__5079\,
            I => \eeprom.n3142\
        );

    \I__1013\ : CascadeMux
    port map (
            O => \N__5076\,
            I => \eeprom.i2c.n10_adj_380_cascade_\
        );

    \I__1012\ : InMux
    port map (
            O => \N__5073\,
            I => \N__5069\
        );

    \I__1011\ : InMux
    port map (
            O => \N__5072\,
            I => \N__5066\
        );

    \I__1010\ : LocalMux
    port map (
            O => \N__5069\,
            I => \N__5063\
        );

    \I__1009\ : LocalMux
    port map (
            O => \N__5066\,
            I => \N__5058\
        );

    \I__1008\ : Span4Mux_v
    port map (
            O => \N__5063\,
            I => \N__5058\
        );

    \I__1007\ : Odrv4
    port map (
            O => \N__5058\,
            I => \eeprom.i2c.n15\
        );

    \I__1006\ : InMux
    port map (
            O => \N__5055\,
            I => \eeprom.i2c.n2849\
        );

    \I__1005\ : InMux
    port map (
            O => \N__5052\,
            I => \eeprom.i2c.n2850\
        );

    \I__1004\ : InMux
    port map (
            O => \N__5049\,
            I => \eeprom.i2c.n2851\
        );

    \I__1003\ : InMux
    port map (
            O => \N__5046\,
            I => \eeprom.i2c.n2852\
        );

    \I__1002\ : CascadeMux
    port map (
            O => \N__5043\,
            I => \N__5040\
        );

    \I__1001\ : InMux
    port map (
            O => \N__5040\,
            I => \N__5037\
        );

    \I__1000\ : LocalMux
    port map (
            O => \N__5037\,
            I => \N__5034\
        );

    \I__999\ : Span4Mux_h
    port map (
            O => \N__5034\,
            I => \N__5030\
        );

    \I__998\ : InMux
    port map (
            O => \N__5033\,
            I => \N__5027\
        );

    \I__997\ : Odrv4
    port map (
            O => \N__5030\,
            I => data_7
        );

    \I__996\ : LocalMux
    port map (
            O => \N__5027\,
            I => data_7
        );

    \I__995\ : CascadeMux
    port map (
            O => \N__5022\,
            I => \N__5018\
        );

    \I__994\ : InMux
    port map (
            O => \N__5021\,
            I => \N__5014\
        );

    \I__993\ : InMux
    port map (
            O => \N__5018\,
            I => \N__5011\
        );

    \I__992\ : CascadeMux
    port map (
            O => \N__5017\,
            I => \N__5008\
        );

    \I__991\ : LocalMux
    port map (
            O => \N__5014\,
            I => \N__5001\
        );

    \I__990\ : LocalMux
    port map (
            O => \N__5011\,
            I => \N__5001\
        );

    \I__989\ : InMux
    port map (
            O => \N__5008\,
            I => \N__4998\
        );

    \I__988\ : InMux
    port map (
            O => \N__5007\,
            I => \N__4995\
        );

    \I__987\ : InMux
    port map (
            O => \N__5006\,
            I => \N__4992\
        );

    \I__986\ : Span4Mux_v
    port map (
            O => \N__5001\,
            I => \N__4986\
        );

    \I__985\ : LocalMux
    port map (
            O => \N__4998\,
            I => \N__4986\
        );

    \I__984\ : LocalMux
    port map (
            O => \N__4995\,
            I => \N__4981\
        );

    \I__983\ : LocalMux
    port map (
            O => \N__4992\,
            I => \N__4981\
        );

    \I__982\ : InMux
    port map (
            O => \N__4991\,
            I => \N__4978\
        );

    \I__981\ : Odrv4
    port map (
            O => \N__4986\,
            I => \enable_slow_N_373\
        );

    \I__980\ : Odrv4
    port map (
            O => \N__4981\,
            I => \enable_slow_N_373\
        );

    \I__979\ : LocalMux
    port map (
            O => \N__4978\,
            I => \enable_slow_N_373\
        );

    \I__978\ : CascadeMux
    port map (
            O => \N__4971\,
            I => \eeprom.n14_cascade_\
        );

    \I__977\ : InMux
    port map (
            O => \N__4968\,
            I => \N__4965\
        );

    \I__976\ : LocalMux
    port map (
            O => \N__4965\,
            I => n2382
        );

    \I__975\ : CascadeMux
    port map (
            O => \N__4962\,
            I => \n3051_cascade_\
        );

    \I__974\ : InMux
    port map (
            O => \N__4959\,
            I => \N__4950\
        );

    \I__973\ : InMux
    port map (
            O => \N__4958\,
            I => \N__4950\
        );

    \I__972\ : InMux
    port map (
            O => \N__4957\,
            I => \N__4950\
        );

    \I__971\ : LocalMux
    port map (
            O => \N__4950\,
            I => n2913
        );

    \I__970\ : CascadeMux
    port map (
            O => \N__4947\,
            I => \n1113_cascade_\
        );

    \I__969\ : InMux
    port map (
            O => \N__4944\,
            I => \N__4940\
        );

    \I__968\ : InMux
    port map (
            O => \N__4943\,
            I => \N__4937\
        );

    \I__967\ : LocalMux
    port map (
            O => \N__4940\,
            I => \N__4929\
        );

    \I__966\ : LocalMux
    port map (
            O => \N__4937\,
            I => \N__4929\
        );

    \I__965\ : InMux
    port map (
            O => \N__4936\,
            I => \N__4924\
        );

    \I__964\ : InMux
    port map (
            O => \N__4935\,
            I => \N__4924\
        );

    \I__963\ : InMux
    port map (
            O => \N__4934\,
            I => \N__4921\
        );

    \I__962\ : Span4Mux_h
    port map (
            O => \N__4929\,
            I => \N__4918\
        );

    \I__961\ : LocalMux
    port map (
            O => \N__4924\,
            I => \N__4915\
        );

    \I__960\ : LocalMux
    port map (
            O => \N__4921\,
            I => read
        );

    \I__959\ : Odrv4
    port map (
            O => \N__4918\,
            I => read
        );

    \I__958\ : Odrv4
    port map (
            O => \N__4915\,
            I => read
        );

    \I__957\ : InMux
    port map (
            O => \N__4908\,
            I => \N__4905\
        );

    \I__956\ : LocalMux
    port map (
            O => \N__4905\,
            I => n3109
        );

    \I__955\ : CascadeMux
    port map (
            O => \N__4902\,
            I => \N__4897\
        );

    \I__954\ : InMux
    port map (
            O => \N__4901\,
            I => \N__4894\
        );

    \I__953\ : CascadeMux
    port map (
            O => \N__4900\,
            I => \N__4891\
        );

    \I__952\ : InMux
    port map (
            O => \N__4897\,
            I => \N__4888\
        );

    \I__951\ : LocalMux
    port map (
            O => \N__4894\,
            I => \N__4885\
        );

    \I__950\ : InMux
    port map (
            O => \N__4891\,
            I => \N__4882\
        );

    \I__949\ : LocalMux
    port map (
            O => \N__4888\,
            I => \eeprom.i2c.n11\
        );

    \I__948\ : Odrv4
    port map (
            O => \N__4885\,
            I => \eeprom.i2c.n11\
        );

    \I__947\ : LocalMux
    port map (
            O => \N__4882\,
            I => \eeprom.i2c.n11\
        );

    \I__946\ : InMux
    port map (
            O => \N__4875\,
            I => \N__4872\
        );

    \I__945\ : LocalMux
    port map (
            O => \N__4872\,
            I => \N__4869\
        );

    \I__944\ : Span4Mux_v
    port map (
            O => \N__4869\,
            I => \N__4865\
        );

    \I__943\ : InMux
    port map (
            O => \N__4868\,
            I => \N__4862\
        );

    \I__942\ : Odrv4
    port map (
            O => \N__4865\,
            I => rw
        );

    \I__941\ : LocalMux
    port map (
            O => \N__4862\,
            I => rw
        );

    \I__940\ : CascadeMux
    port map (
            O => \N__4857\,
            I => \N__4854\
        );

    \I__939\ : InMux
    port map (
            O => \N__4854\,
            I => \N__4851\
        );

    \I__938\ : LocalMux
    port map (
            O => \N__4851\,
            I => \N__4847\
        );

    \I__937\ : InMux
    port map (
            O => \N__4850\,
            I => \N__4844\
        );

    \I__936\ : Span4Mux_v
    port map (
            O => \N__4847\,
            I => \N__4839\
        );

    \I__935\ : LocalMux
    port map (
            O => \N__4844\,
            I => \N__4836\
        );

    \I__934\ : InMux
    port map (
            O => \N__4843\,
            I => \N__4833\
        );

    \I__933\ : InMux
    port map (
            O => \N__4842\,
            I => \N__4830\
        );

    \I__932\ : Odrv4
    port map (
            O => \N__4839\,
            I => \state_7_N_270_0\
        );

    \I__931\ : Odrv4
    port map (
            O => \N__4836\,
            I => \state_7_N_270_0\
        );

    \I__930\ : LocalMux
    port map (
            O => \N__4833\,
            I => \state_7_N_270_0\
        );

    \I__929\ : LocalMux
    port map (
            O => \N__4830\,
            I => \state_7_N_270_0\
        );

    \I__928\ : InMux
    port map (
            O => \N__4821\,
            I => \N__4818\
        );

    \I__927\ : LocalMux
    port map (
            O => \N__4818\,
            I => \N__4814\
        );

    \I__926\ : InMux
    port map (
            O => \N__4817\,
            I => \N__4811\
        );

    \I__925\ : Odrv12
    port map (
            O => \N__4814\,
            I => \eeprom.i2c.n11_adj_374\
        );

    \I__924\ : LocalMux
    port map (
            O => \N__4811\,
            I => \eeprom.i2c.n11_adj_374\
        );

    \I__923\ : InMux
    port map (
            O => \N__4806\,
            I => \N__4802\
        );

    \I__922\ : InMux
    port map (
            O => \N__4805\,
            I => \N__4799\
        );

    \I__921\ : LocalMux
    port map (
            O => \N__4802\,
            I => \N__4796\
        );

    \I__920\ : LocalMux
    port map (
            O => \N__4799\,
            I => \eeprom.i2c.n11_adj_378\
        );

    \I__919\ : Odrv4
    port map (
            O => \N__4796\,
            I => \eeprom.i2c.n11_adj_378\
        );

    \I__918\ : InMux
    port map (
            O => \N__4791\,
            I => \N__4786\
        );

    \I__917\ : InMux
    port map (
            O => \N__4790\,
            I => \N__4783\
        );

    \I__916\ : InMux
    port map (
            O => \N__4789\,
            I => \N__4780\
        );

    \I__915\ : LocalMux
    port map (
            O => \N__4786\,
            I => saved_addr_0
        );

    \I__914\ : LocalMux
    port map (
            O => \N__4783\,
            I => saved_addr_0
        );

    \I__913\ : LocalMux
    port map (
            O => \N__4780\,
            I => saved_addr_0
        );

    \I__912\ : InMux
    port map (
            O => \N__4773\,
            I => \N__4770\
        );

    \I__911\ : LocalMux
    port map (
            O => \N__4770\,
            I => \N__4767\
        );

    \I__910\ : Span4Mux_v
    port map (
            O => \N__4767\,
            I => \N__4763\
        );

    \I__909\ : InMux
    port map (
            O => \N__4766\,
            I => \N__4760\
        );

    \I__908\ : Sp12to4
    port map (
            O => \N__4763\,
            I => \N__4755\
        );

    \I__907\ : LocalMux
    port map (
            O => \N__4760\,
            I => \N__4755\
        );

    \I__906\ : Odrv12
    port map (
            O => \N__4755\,
            I => n4
        );

    \I__905\ : CEMux
    port map (
            O => \N__4752\,
            I => \N__4746\
        );

    \I__904\ : CEMux
    port map (
            O => \N__4751\,
            I => \N__4743\
        );

    \I__903\ : CEMux
    port map (
            O => \N__4750\,
            I => \N__4740\
        );

    \I__902\ : CEMux
    port map (
            O => \N__4749\,
            I => \N__4737\
        );

    \I__901\ : LocalMux
    port map (
            O => \N__4746\,
            I => \N__4733\
        );

    \I__900\ : LocalMux
    port map (
            O => \N__4743\,
            I => \N__4730\
        );

    \I__899\ : LocalMux
    port map (
            O => \N__4740\,
            I => \N__4727\
        );

    \I__898\ : LocalMux
    port map (
            O => \N__4737\,
            I => \N__4724\
        );

    \I__897\ : CascadeMux
    port map (
            O => \N__4736\,
            I => \N__4721\
        );

    \I__896\ : Span4Mux_h
    port map (
            O => \N__4733\,
            I => \N__4716\
        );

    \I__895\ : Span4Mux_h
    port map (
            O => \N__4730\,
            I => \N__4709\
        );

    \I__894\ : Span4Mux_v
    port map (
            O => \N__4727\,
            I => \N__4709\
        );

    \I__893\ : Span4Mux_h
    port map (
            O => \N__4724\,
            I => \N__4709\
        );

    \I__892\ : InMux
    port map (
            O => \N__4721\,
            I => \N__4706\
        );

    \I__891\ : InMux
    port map (
            O => \N__4720\,
            I => \N__4703\
        );

    \I__890\ : InMux
    port map (
            O => \N__4719\,
            I => \N__4700\
        );

    \I__889\ : Odrv4
    port map (
            O => \N__4716\,
            I => \eeprom.i2c.n1063\
        );

    \I__888\ : Odrv4
    port map (
            O => \N__4709\,
            I => \eeprom.i2c.n1063\
        );

    \I__887\ : LocalMux
    port map (
            O => \N__4706\,
            I => \eeprom.i2c.n1063\
        );

    \I__886\ : LocalMux
    port map (
            O => \N__4703\,
            I => \eeprom.i2c.n1063\
        );

    \I__885\ : LocalMux
    port map (
            O => \N__4700\,
            I => \eeprom.i2c.n1063\
        );

    \I__884\ : CascadeMux
    port map (
            O => \N__4689\,
            I => \eeprom.i2c.n9_adj_377_cascade_\
        );

    \I__883\ : SRMux
    port map (
            O => \N__4686\,
            I => \N__4683\
        );

    \I__882\ : LocalMux
    port map (
            O => \N__4683\,
            I => \N__4680\
        );

    \I__881\ : Span4Mux_h
    port map (
            O => \N__4680\,
            I => \N__4677\
        );

    \I__880\ : Odrv4
    port map (
            O => \N__4677\,
            I => \eeprom.i2c.n3050\
        );

    \I__879\ : InMux
    port map (
            O => \N__4674\,
            I => \N__4671\
        );

    \I__878\ : LocalMux
    port map (
            O => \N__4671\,
            I => \N__4667\
        );

    \I__877\ : InMux
    port map (
            O => \N__4670\,
            I => \N__4664\
        );

    \I__876\ : Span4Mux_h
    port map (
            O => \N__4667\,
            I => \N__4661\
        );

    \I__875\ : LocalMux
    port map (
            O => \N__4664\,
            I => \N__4658\
        );

    \I__874\ : Odrv4
    port map (
            O => \N__4661\,
            I => n4_adj_389
        );

    \I__873\ : Odrv4
    port map (
            O => \N__4658\,
            I => n4_adj_389
        );

    \I__872\ : InMux
    port map (
            O => \N__4653\,
            I => \N__4650\
        );

    \I__871\ : LocalMux
    port map (
            O => \N__4650\,
            I => \N__4647\
        );

    \I__870\ : Odrv12
    port map (
            O => \N__4647\,
            I => n2344
        );

    \I__869\ : CascadeMux
    port map (
            O => \N__4644\,
            I => \n2344_cascade_\
        );

    \I__868\ : CascadeMux
    port map (
            O => \N__4641\,
            I => \N__4638\
        );

    \I__867\ : InMux
    port map (
            O => \N__4638\,
            I => \N__4634\
        );

    \I__866\ : InMux
    port map (
            O => \N__4637\,
            I => \N__4631\
        );

    \I__865\ : LocalMux
    port map (
            O => \N__4634\,
            I => \eeprom.i2c.n10_adj_381\
        );

    \I__864\ : LocalMux
    port map (
            O => \N__4631\,
            I => \eeprom.i2c.n10_adj_381\
        );

    \I__863\ : CascadeMux
    port map (
            O => \N__4626\,
            I => \eeprom.i2c.n11_adj_378_cascade_\
        );

    \I__862\ : InMux
    port map (
            O => \N__4623\,
            I => \N__4620\
        );

    \I__861\ : LocalMux
    port map (
            O => \N__4620\,
            I => \eeprom.i2c.n2352\
        );

    \I__860\ : CascadeMux
    port map (
            O => \N__4617\,
            I => \eeprom.i2c.n1734_cascade_\
        );

    \I__859\ : InMux
    port map (
            O => \N__4614\,
            I => \N__4610\
        );

    \I__858\ : InMux
    port map (
            O => \N__4613\,
            I => \N__4607\
        );

    \I__857\ : LocalMux
    port map (
            O => \N__4610\,
            I => \eeprom.i2c.n2358\
        );

    \I__856\ : LocalMux
    port map (
            O => \N__4607\,
            I => \eeprom.i2c.n2358\
        );

    \I__855\ : CascadeMux
    port map (
            O => \N__4602\,
            I => \eeprom.i2c.n1063_cascade_\
        );

    \I__854\ : SRMux
    port map (
            O => \N__4599\,
            I => \N__4596\
        );

    \I__853\ : LocalMux
    port map (
            O => \N__4596\,
            I => \N__4593\
        );

    \I__852\ : Odrv4
    port map (
            O => \N__4593\,
            I => \eeprom.i2c.n1923\
        );

    \I__851\ : InMux
    port map (
            O => \N__4590\,
            I => \N__4586\
        );

    \I__850\ : InMux
    port map (
            O => \N__4589\,
            I => \N__4583\
        );

    \I__849\ : LocalMux
    port map (
            O => \N__4586\,
            I => \N__4580\
        );

    \I__848\ : LocalMux
    port map (
            O => \N__4583\,
            I => \N__4577\
        );

    \I__847\ : Odrv4
    port map (
            O => \N__4580\,
            I => \eeprom.enable\
        );

    \I__846\ : Odrv4
    port map (
            O => \N__4577\,
            I => \eeprom.enable\
        );

    \I__845\ : CEMux
    port map (
            O => \N__4572\,
            I => \N__4569\
        );

    \I__844\ : LocalMux
    port map (
            O => \N__4569\,
            I => \N__4566\
        );

    \I__843\ : Span4Mux_h
    port map (
            O => \N__4566\,
            I => \N__4563\
        );

    \I__842\ : Odrv4
    port map (
            O => \N__4563\,
            I => \eeprom.i2c.n1761\
        );

    \I__841\ : InMux
    port map (
            O => \N__4560\,
            I => \N__4555\
        );

    \I__840\ : InMux
    port map (
            O => \N__4559\,
            I => \N__4552\
        );

    \I__839\ : InMux
    port map (
            O => \N__4558\,
            I => \N__4549\
        );

    \I__838\ : LocalMux
    port map (
            O => \N__4555\,
            I => \N__4546\
        );

    \I__837\ : LocalMux
    port map (
            O => \N__4552\,
            I => \N__4541\
        );

    \I__836\ : LocalMux
    port map (
            O => \N__4549\,
            I => \N__4541\
        );

    \I__835\ : Span4Mux_v
    port map (
            O => \N__4546\,
            I => \N__4538\
        );

    \I__834\ : Odrv12
    port map (
            O => \N__4541\,
            I => \eeprom.n1704\
        );

    \I__833\ : Odrv4
    port map (
            O => \N__4538\,
            I => \eeprom.n1704\
        );

    \I__832\ : CascadeMux
    port map (
            O => \N__4533\,
            I => \eeprom.n26_cascade_\
        );

    \I__831\ : InMux
    port map (
            O => \N__4530\,
            I => \N__4527\
        );

    \I__830\ : LocalMux
    port map (
            O => \N__4527\,
            I => \eeprom.i2c.n3123\
        );

    \I__829\ : CEMux
    port map (
            O => \N__4524\,
            I => \N__4521\
        );

    \I__828\ : LocalMux
    port map (
            O => \N__4521\,
            I => \N__4518\
        );

    \I__827\ : Span4Mux_h
    port map (
            O => \N__4518\,
            I => \N__4515\
        );

    \I__826\ : Odrv4
    port map (
            O => \N__4515\,
            I => \eeprom.i2c.n2967\
        );

    \I__825\ : CascadeMux
    port map (
            O => \N__4512\,
            I => \eeprom.i2c.n37_cascade_\
        );

    \I__824\ : InMux
    port map (
            O => \N__4509\,
            I => \N__4505\
        );

    \I__823\ : InMux
    port map (
            O => \N__4508\,
            I => \N__4502\
        );

    \I__822\ : LocalMux
    port map (
            O => \N__4505\,
            I => \eeprom.i2c.n33\
        );

    \I__821\ : LocalMux
    port map (
            O => \N__4502\,
            I => \eeprom.i2c.n33\
        );

    \I__820\ : InMux
    port map (
            O => \N__4497\,
            I => \N__4494\
        );

    \I__819\ : LocalMux
    port map (
            O => \N__4494\,
            I => \eeprom.i2c.n39\
        );

    \I__818\ : CascadeMux
    port map (
            O => \N__4491\,
            I => \eeprom.i2c.n39_cascade_\
        );

    \I__817\ : InMux
    port map (
            O => \N__4488\,
            I => \N__4485\
        );

    \I__816\ : LocalMux
    port map (
            O => \N__4485\,
            I => \eeprom.i2c.n3133\
        );

    \I__815\ : CascadeMux
    port map (
            O => \N__4482\,
            I => \N__4479\
        );

    \I__814\ : InMux
    port map (
            O => \N__4479\,
            I => \N__4476\
        );

    \I__813\ : LocalMux
    port map (
            O => \N__4476\,
            I => \N__4473\
        );

    \I__812\ : Span4Mux_h
    port map (
            O => \N__4473\,
            I => \N__4470\
        );

    \I__811\ : Odrv4
    port map (
            O => \N__4470\,
            I => \eeprom.i2c.n7\
        );

    \I__810\ : SRMux
    port map (
            O => \N__4467\,
            I => \N__4464\
        );

    \I__809\ : LocalMux
    port map (
            O => \N__4464\,
            I => \N__4461\
        );

    \I__808\ : Odrv4
    port map (
            O => \N__4461\,
            I => \eeprom.i2c.n3082\
        );

    \I__807\ : InMux
    port map (
            O => \N__4458\,
            I => \N__4455\
        );

    \I__806\ : LocalMux
    port map (
            O => \N__4455\,
            I => \eeprom.i2c.n13\
        );

    \I__805\ : CascadeMux
    port map (
            O => \N__4452\,
            I => \eeprom.i2c.n15_cascade_\
        );

    \I__804\ : CascadeMux
    port map (
            O => \N__4449\,
            I => \n1718_cascade_\
        );

    \I__803\ : InMux
    port map (
            O => \N__4446\,
            I => \N__4440\
        );

    \I__802\ : InMux
    port map (
            O => \N__4445\,
            I => \N__4440\
        );

    \I__801\ : LocalMux
    port map (
            O => \N__4440\,
            I => data_2
        );

    \I__800\ : InMux
    port map (
            O => \N__4437\,
            I => \N__4428\
        );

    \I__799\ : InMux
    port map (
            O => \N__4436\,
            I => \N__4428\
        );

    \I__798\ : InMux
    port map (
            O => \N__4435\,
            I => \N__4428\
        );

    \I__797\ : LocalMux
    port map (
            O => \N__4428\,
            I => n1718
        );

    \I__796\ : InMux
    port map (
            O => \N__4425\,
            I => \N__4419\
        );

    \I__795\ : InMux
    port map (
            O => \N__4424\,
            I => \N__4419\
        );

    \I__794\ : LocalMux
    port map (
            O => \N__4419\,
            I => data_6
        );

    \I__793\ : SRMux
    port map (
            O => \N__4416\,
            I => \N__4413\
        );

    \I__792\ : LocalMux
    port map (
            O => \N__4413\,
            I => \N__4410\
        );

    \I__791\ : Odrv4
    port map (
            O => \N__4410\,
            I => \eeprom.i2c.n1928\
        );

    \I__790\ : CascadeMux
    port map (
            O => \N__4407\,
            I => \eeprom.i2c.n3130_cascade_\
        );

    \I__789\ : CEMux
    port map (
            O => \N__4404\,
            I => \N__4401\
        );

    \I__788\ : LocalMux
    port map (
            O => \N__4401\,
            I => \N__4398\
        );

    \I__787\ : Odrv4
    port map (
            O => \N__4398\,
            I => \eeprom.i2c.n1153\
        );

    \I__786\ : SRMux
    port map (
            O => \N__4395\,
            I => \N__4392\
        );

    \I__785\ : LocalMux
    port map (
            O => \N__4392\,
            I => \N__4389\
        );

    \I__784\ : Span4Mux_h
    port map (
            O => \N__4389\,
            I => \N__4386\
        );

    \I__783\ : Odrv4
    port map (
            O => \N__4386\,
            I => \eeprom.i2c.n2388\
        );

    \I__782\ : InMux
    port map (
            O => \N__4383\,
            I => \N__4379\
        );

    \I__781\ : InMux
    port map (
            O => \N__4382\,
            I => \N__4376\
        );

    \I__780\ : LocalMux
    port map (
            O => \N__4379\,
            I => data_5
        );

    \I__779\ : LocalMux
    port map (
            O => \N__4376\,
            I => data_5
        );

    \I__778\ : InMux
    port map (
            O => \N__4371\,
            I => \N__4365\
        );

    \I__777\ : InMux
    port map (
            O => \N__4370\,
            I => \N__4365\
        );

    \I__776\ : LocalMux
    port map (
            O => \N__4365\,
            I => data_0
        );

    \I__775\ : CascadeMux
    port map (
            O => \N__4362\,
            I => \N__4359\
        );

    \I__774\ : InMux
    port map (
            O => \N__4359\,
            I => \N__4356\
        );

    \I__773\ : LocalMux
    port map (
            O => \N__4356\,
            I => \N__4352\
        );

    \I__772\ : InMux
    port map (
            O => \N__4355\,
            I => \N__4349\
        );

    \I__771\ : Odrv4
    port map (
            O => \N__4352\,
            I => data_3
        );

    \I__770\ : LocalMux
    port map (
            O => \N__4349\,
            I => data_3
        );

    \I__769\ : InMux
    port map (
            O => \N__4344\,
            I => \N__4341\
        );

    \I__768\ : LocalMux
    port map (
            O => \N__4341\,
            I => n13
        );

    \I__767\ : InMux
    port map (
            O => \N__4338\,
            I => \N__4335\
        );

    \I__766\ : LocalMux
    port map (
            O => \N__4335\,
            I => n12
        );

    \I__765\ : InMux
    port map (
            O => \N__4332\,
            I => \N__4326\
        );

    \I__764\ : InMux
    port map (
            O => \N__4331\,
            I => \N__4326\
        );

    \I__763\ : LocalMux
    port map (
            O => \N__4326\,
            I => data_4
        );

    \I__762\ : CascadeMux
    port map (
            O => \N__4323\,
            I => \n1836_cascade_\
        );

    \I__761\ : CEMux
    port map (
            O => \N__4320\,
            I => \N__4316\
        );

    \I__760\ : CEMux
    port map (
            O => \N__4319\,
            I => \N__4312\
        );

    \I__759\ : LocalMux
    port map (
            O => \N__4316\,
            I => \N__4308\
        );

    \I__758\ : CEMux
    port map (
            O => \N__4315\,
            I => \N__4305\
        );

    \I__757\ : LocalMux
    port map (
            O => \N__4312\,
            I => \N__4302\
        );

    \I__756\ : CEMux
    port map (
            O => \N__4311\,
            I => \N__4299\
        );

    \I__755\ : Span4Mux_h
    port map (
            O => \N__4308\,
            I => \N__4295\
        );

    \I__754\ : LocalMux
    port map (
            O => \N__4305\,
            I => \N__4292\
        );

    \I__753\ : Span4Mux_h
    port map (
            O => \N__4302\,
            I => \N__4289\
        );

    \I__752\ : LocalMux
    port map (
            O => \N__4299\,
            I => \N__4286\
        );

    \I__751\ : InMux
    port map (
            O => \N__4298\,
            I => \N__4283\
        );

    \I__750\ : Odrv4
    port map (
            O => \N__4295\,
            I => n1507
        );

    \I__749\ : Odrv4
    port map (
            O => \N__4292\,
            I => n1507
        );

    \I__748\ : Odrv4
    port map (
            O => \N__4289\,
            I => n1507
        );

    \I__747\ : Odrv12
    port map (
            O => \N__4286\,
            I => n1507
        );

    \I__746\ : LocalMux
    port map (
            O => \N__4283\,
            I => n1507
        );

    \I__745\ : InMux
    port map (
            O => \N__4272\,
            I => \N__4266\
        );

    \I__744\ : InMux
    port map (
            O => \N__4271\,
            I => \N__4266\
        );

    \I__743\ : LocalMux
    port map (
            O => \N__4266\,
            I => n104
        );

    \I__742\ : InMux
    port map (
            O => \N__4263\,
            I => \N__4254\
        );

    \I__741\ : InMux
    port map (
            O => \N__4262\,
            I => \N__4254\
        );

    \I__740\ : InMux
    port map (
            O => \N__4261\,
            I => \N__4254\
        );

    \I__739\ : LocalMux
    port map (
            O => \N__4254\,
            I => \N__4251\
        );

    \I__738\ : Odrv12
    port map (
            O => \N__4251\,
            I => n15
        );

    \I__737\ : CascadeMux
    port map (
            O => \N__4248\,
            I => \N__4242\
        );

    \I__736\ : InMux
    port map (
            O => \N__4247\,
            I => \N__4235\
        );

    \I__735\ : InMux
    port map (
            O => \N__4246\,
            I => \N__4235\
        );

    \I__734\ : InMux
    port map (
            O => \N__4245\,
            I => \N__4226\
        );

    \I__733\ : InMux
    port map (
            O => \N__4242\,
            I => \N__4226\
        );

    \I__732\ : InMux
    port map (
            O => \N__4241\,
            I => \N__4226\
        );

    \I__731\ : InMux
    port map (
            O => \N__4240\,
            I => \N__4226\
        );

    \I__730\ : LocalMux
    port map (
            O => \N__4235\,
            I => \N__4223\
        );

    \I__729\ : LocalMux
    port map (
            O => \N__4226\,
            I => \ID_READOUT_FSM_state_1\
        );

    \I__728\ : Odrv4
    port map (
            O => \N__4223\,
            I => \ID_READOUT_FSM_state_1\
        );

    \I__727\ : InMux
    port map (
            O => \N__4218\,
            I => \N__4214\
        );

    \I__726\ : CascadeMux
    port map (
            O => \N__4217\,
            I => \N__4210\
        );

    \I__725\ : LocalMux
    port map (
            O => \N__4214\,
            I => \N__4204\
        );

    \I__724\ : InMux
    port map (
            O => \N__4213\,
            I => \N__4195\
        );

    \I__723\ : InMux
    port map (
            O => \N__4210\,
            I => \N__4195\
        );

    \I__722\ : InMux
    port map (
            O => \N__4209\,
            I => \N__4195\
        );

    \I__721\ : InMux
    port map (
            O => \N__4208\,
            I => \N__4195\
        );

    \I__720\ : InMux
    port map (
            O => \N__4207\,
            I => \N__4192\
        );

    \I__719\ : Odrv4
    port map (
            O => \N__4204\,
            I => \ID_READOUT_FSM_state_0\
        );

    \I__718\ : LocalMux
    port map (
            O => \N__4195\,
            I => \ID_READOUT_FSM_state_0\
        );

    \I__717\ : LocalMux
    port map (
            O => \N__4192\,
            I => \ID_READOUT_FSM_state_0\
        );

    \I__716\ : InMux
    port map (
            O => \N__4185\,
            I => \N__4179\
        );

    \I__715\ : InMux
    port map (
            O => \N__4184\,
            I => \N__4179\
        );

    \I__714\ : LocalMux
    port map (
            O => \N__4179\,
            I => n2414
        );

    \I__713\ : InMux
    port map (
            O => \N__4176\,
            I => \N__4172\
        );

    \I__712\ : InMux
    port map (
            O => \N__4175\,
            I => \N__4169\
        );

    \I__711\ : LocalMux
    port map (
            O => \N__4172\,
            I => delay_counter_22
        );

    \I__710\ : LocalMux
    port map (
            O => \N__4169\,
            I => delay_counter_22
        );

    \I__709\ : InMux
    port map (
            O => \N__4164\,
            I => \N__4160\
        );

    \I__708\ : InMux
    port map (
            O => \N__4163\,
            I => \N__4157\
        );

    \I__707\ : LocalMux
    port map (
            O => \N__4160\,
            I => delay_counter_30
        );

    \I__706\ : LocalMux
    port map (
            O => \N__4157\,
            I => delay_counter_30
        );

    \I__705\ : CascadeMux
    port map (
            O => \N__4152\,
            I => \N__4148\
        );

    \I__704\ : InMux
    port map (
            O => \N__4151\,
            I => \N__4145\
        );

    \I__703\ : InMux
    port map (
            O => \N__4148\,
            I => \N__4142\
        );

    \I__702\ : LocalMux
    port map (
            O => \N__4145\,
            I => delay_counter_26
        );

    \I__701\ : LocalMux
    port map (
            O => \N__4142\,
            I => delay_counter_26
        );

    \I__700\ : InMux
    port map (
            O => \N__4137\,
            I => \N__4133\
        );

    \I__699\ : InMux
    port map (
            O => \N__4136\,
            I => \N__4130\
        );

    \I__698\ : LocalMux
    port map (
            O => \N__4133\,
            I => delay_counter_28
        );

    \I__697\ : LocalMux
    port map (
            O => \N__4130\,
            I => delay_counter_28
        );

    \I__696\ : InMux
    port map (
            O => \N__4125\,
            I => \N__4122\
        );

    \I__695\ : LocalMux
    port map (
            O => \N__4122\,
            I => \N__4119\
        );

    \I__694\ : Odrv4
    port map (
            O => \N__4119\,
            I => n24
        );

    \I__693\ : CascadeMux
    port map (
            O => \N__4116\,
            I => \eeprom.i2c.n10_adj_381_cascade_\
        );

    \I__692\ : InMux
    port map (
            O => \N__4113\,
            I => \N__4109\
        );

    \I__691\ : InMux
    port map (
            O => \N__4112\,
            I => \N__4106\
        );

    \I__690\ : LocalMux
    port map (
            O => \N__4109\,
            I => \eeprom.delay_counter_12\
        );

    \I__689\ : LocalMux
    port map (
            O => \N__4106\,
            I => \eeprom.delay_counter_12\
        );

    \I__688\ : InMux
    port map (
            O => \N__4101\,
            I => \N__4097\
        );

    \I__687\ : InMux
    port map (
            O => \N__4100\,
            I => \N__4094\
        );

    \I__686\ : LocalMux
    port map (
            O => \N__4097\,
            I => \eeprom.delay_counter_10\
        );

    \I__685\ : LocalMux
    port map (
            O => \N__4094\,
            I => \eeprom.delay_counter_10\
        );

    \I__684\ : CascadeMux
    port map (
            O => \N__4089\,
            I => \N__4085\
        );

    \I__683\ : InMux
    port map (
            O => \N__4088\,
            I => \N__4082\
        );

    \I__682\ : InMux
    port map (
            O => \N__4085\,
            I => \N__4079\
        );

    \I__681\ : LocalMux
    port map (
            O => \N__4082\,
            I => \eeprom.delay_counter_8\
        );

    \I__680\ : LocalMux
    port map (
            O => \N__4079\,
            I => \eeprom.delay_counter_8\
        );

    \I__679\ : InMux
    port map (
            O => \N__4074\,
            I => \N__4070\
        );

    \I__678\ : InMux
    port map (
            O => \N__4073\,
            I => \N__4067\
        );

    \I__677\ : LocalMux
    port map (
            O => \N__4070\,
            I => \eeprom.delay_counter_6\
        );

    \I__676\ : LocalMux
    port map (
            O => \N__4067\,
            I => \eeprom.delay_counter_6\
        );

    \I__675\ : CascadeMux
    port map (
            O => \N__4062\,
            I => \N__4059\
        );

    \I__674\ : InMux
    port map (
            O => \N__4059\,
            I => \N__4056\
        );

    \I__673\ : LocalMux
    port map (
            O => \N__4056\,
            I => \N__4053\
        );

    \I__672\ : Span4Mux_v
    port map (
            O => \N__4053\,
            I => \N__4050\
        );

    \I__671\ : Odrv4
    port map (
            O => \N__4050\,
            I => \eeprom.n28\
        );

    \I__670\ : InMux
    port map (
            O => \N__4047\,
            I => \N__4043\
        );

    \I__669\ : InMux
    port map (
            O => \N__4046\,
            I => \N__4040\
        );

    \I__668\ : LocalMux
    port map (
            O => \N__4043\,
            I => \N__4037\
        );

    \I__667\ : LocalMux
    port map (
            O => \N__4040\,
            I => delay_counter_29
        );

    \I__666\ : Odrv4
    port map (
            O => \N__4037\,
            I => delay_counter_29
        );

    \I__665\ : InMux
    port map (
            O => \N__4032\,
            I => \N__4028\
        );

    \I__664\ : InMux
    port map (
            O => \N__4031\,
            I => \N__4025\
        );

    \I__663\ : LocalMux
    port map (
            O => \N__4028\,
            I => delay_counter_18
        );

    \I__662\ : LocalMux
    port map (
            O => \N__4025\,
            I => delay_counter_18
        );

    \I__661\ : CascadeMux
    port map (
            O => \N__4020\,
            I => \n36_cascade_\
        );

    \I__660\ : InMux
    port map (
            O => \N__4017\,
            I => \N__4013\
        );

    \I__659\ : InMux
    port map (
            O => \N__4016\,
            I => \N__4010\
        );

    \I__658\ : LocalMux
    port map (
            O => \N__4013\,
            I => \N__4007\
        );

    \I__657\ : LocalMux
    port map (
            O => \N__4010\,
            I => delay_counter_24
        );

    \I__656\ : Odrv4
    port map (
            O => \N__4007\,
            I => delay_counter_24
        );

    \I__655\ : InMux
    port map (
            O => \N__4002\,
            I => \N__3998\
        );

    \I__654\ : InMux
    port map (
            O => \N__4001\,
            I => \N__3995\
        );

    \I__653\ : LocalMux
    port map (
            O => \N__3998\,
            I => \N__3992\
        );

    \I__652\ : LocalMux
    port map (
            O => \N__3995\,
            I => delay_counter_27
        );

    \I__651\ : Odrv4
    port map (
            O => \N__3992\,
            I => delay_counter_27
        );

    \I__650\ : CascadeMux
    port map (
            O => \N__3987\,
            I => \n22_cascade_\
        );

    \I__649\ : InMux
    port map (
            O => \N__3984\,
            I => \N__3980\
        );

    \I__648\ : InMux
    port map (
            O => \N__3983\,
            I => \N__3977\
        );

    \I__647\ : LocalMux
    port map (
            O => \N__3980\,
            I => delay_counter_23
        );

    \I__646\ : LocalMux
    port map (
            O => \N__3977\,
            I => delay_counter_23
        );

    \I__645\ : InMux
    port map (
            O => \N__3972\,
            I => \N__3969\
        );

    \I__644\ : LocalMux
    port map (
            O => \N__3969\,
            I => \N__3965\
        );

    \I__643\ : InMux
    port map (
            O => \N__3968\,
            I => \N__3962\
        );

    \I__642\ : Span4Mux_h
    port map (
            O => \N__3965\,
            I => \N__3959\
        );

    \I__641\ : LocalMux
    port map (
            O => \N__3962\,
            I => delay_counter_31
        );

    \I__640\ : Odrv4
    port map (
            O => \N__3959\,
            I => delay_counter_31
        );

    \I__639\ : CascadeMux
    port map (
            O => \N__3954\,
            I => \n25_cascade_\
        );

    \I__638\ : CascadeMux
    port map (
            O => \N__3951\,
            I => \n104_cascade_\
        );

    \I__637\ : SRMux
    port map (
            O => \N__3948\,
            I => \N__3945\
        );

    \I__636\ : LocalMux
    port map (
            O => \N__3945\,
            I => \N__3942\
        );

    \I__635\ : Span4Mux_h
    port map (
            O => \N__3942\,
            I => \N__3936\
        );

    \I__634\ : SRMux
    port map (
            O => \N__3941\,
            I => \N__3933\
        );

    \I__633\ : SRMux
    port map (
            O => \N__3940\,
            I => \N__3930\
        );

    \I__632\ : SRMux
    port map (
            O => \N__3939\,
            I => \N__3927\
        );

    \I__631\ : Odrv4
    port map (
            O => \N__3936\,
            I => n1891
        );

    \I__630\ : LocalMux
    port map (
            O => \N__3933\,
            I => n1891
        );

    \I__629\ : LocalMux
    port map (
            O => \N__3930\,
            I => n1891
        );

    \I__628\ : LocalMux
    port map (
            O => \N__3927\,
            I => n1891
        );

    \I__627\ : InMux
    port map (
            O => \N__3918\,
            I => \N__3914\
        );

    \I__626\ : InMux
    port map (
            O => \N__3917\,
            I => \N__3911\
        );

    \I__625\ : LocalMux
    port map (
            O => \N__3914\,
            I => delay_counter_21
        );

    \I__624\ : LocalMux
    port map (
            O => \N__3911\,
            I => delay_counter_21
        );

    \I__623\ : InMux
    port map (
            O => \N__3906\,
            I => \N__3902\
        );

    \I__622\ : InMux
    port map (
            O => \N__3905\,
            I => \N__3899\
        );

    \I__621\ : LocalMux
    port map (
            O => \N__3902\,
            I => delay_counter_25
        );

    \I__620\ : LocalMux
    port map (
            O => \N__3899\,
            I => delay_counter_25
        );

    \I__619\ : CascadeMux
    port map (
            O => \N__3894\,
            I => \N__3891\
        );

    \I__618\ : InMux
    port map (
            O => \N__3891\,
            I => \N__3887\
        );

    \I__617\ : InMux
    port map (
            O => \N__3890\,
            I => \N__3884\
        );

    \I__616\ : LocalMux
    port map (
            O => \N__3887\,
            I => \N__3881\
        );

    \I__615\ : LocalMux
    port map (
            O => \N__3884\,
            I => delay_counter_20
        );

    \I__614\ : Odrv4
    port map (
            O => \N__3881\,
            I => delay_counter_20
        );

    \I__613\ : InMux
    port map (
            O => \N__3876\,
            I => \N__3872\
        );

    \I__612\ : InMux
    port map (
            O => \N__3875\,
            I => \N__3869\
        );

    \I__611\ : LocalMux
    port map (
            O => \N__3872\,
            I => delay_counter_19
        );

    \I__610\ : LocalMux
    port map (
            O => \N__3869\,
            I => delay_counter_19
        );

    \I__609\ : InMux
    port map (
            O => \N__3864\,
            I => \N__3861\
        );

    \I__608\ : LocalMux
    port map (
            O => \N__3861\,
            I => n23
        );

    \I__607\ : InMux
    port map (
            O => \N__3858\,
            I => \N__3855\
        );

    \I__606\ : LocalMux
    port map (
            O => \N__3855\,
            I => n20
        );

    \I__605\ : CascadeMux
    port map (
            O => \N__3852\,
            I => \n20_cascade_\
        );

    \I__604\ : InMux
    port map (
            O => \N__3849\,
            I => \N__3843\
        );

    \I__603\ : InMux
    port map (
            O => \N__3848\,
            I => \N__3843\
        );

    \I__602\ : LocalMux
    port map (
            O => \N__3843\,
            I => \N__3840\
        );

    \I__601\ : Odrv4
    port map (
            O => \N__3840\,
            I => n6
        );

    \I__600\ : CascadeMux
    port map (
            O => \N__3837\,
            I => \n805_cascade_\
        );

    \I__599\ : CEMux
    port map (
            O => \N__3834\,
            I => \N__3831\
        );

    \I__598\ : LocalMux
    port map (
            O => \N__3831\,
            I => \N__3827\
        );

    \I__597\ : CEMux
    port map (
            O => \N__3830\,
            I => \N__3824\
        );

    \I__596\ : Span4Mux_v
    port map (
            O => \N__3827\,
            I => \N__3819\
        );

    \I__595\ : LocalMux
    port map (
            O => \N__3824\,
            I => \N__3819\
        );

    \I__594\ : Span4Mux_v
    port map (
            O => \N__3819\,
            I => \N__3816\
        );

    \I__593\ : Span4Mux_v
    port map (
            O => \N__3816\,
            I => \N__3813\
        );

    \I__592\ : Odrv4
    port map (
            O => \N__3813\,
            I => \eeprom.n1796\
        );

    \I__591\ : CascadeMux
    port map (
            O => \N__3810\,
            I => \eeprom.n1796_cascade_\
        );

    \I__590\ : SRMux
    port map (
            O => \N__3807\,
            I => \N__3803\
        );

    \I__589\ : SRMux
    port map (
            O => \N__3806\,
            I => \N__3800\
        );

    \I__588\ : LocalMux
    port map (
            O => \N__3803\,
            I => \N__3797\
        );

    \I__587\ : LocalMux
    port map (
            O => \N__3800\,
            I => \N__3794\
        );

    \I__586\ : Span4Mux_h
    port map (
            O => \N__3797\,
            I => \N__3791\
        );

    \I__585\ : Sp12to4
    port map (
            O => \N__3794\,
            I => \N__3788\
        );

    \I__584\ : Odrv4
    port map (
            O => \N__3791\,
            I => \eeprom.n1929\
        );

    \I__583\ : Odrv12
    port map (
            O => \N__3788\,
            I => \eeprom.n1929\
        );

    \I__582\ : InMux
    port map (
            O => \N__3783\,
            I => \N__3777\
        );

    \I__581\ : InMux
    port map (
            O => \N__3782\,
            I => \N__3777\
        );

    \I__580\ : LocalMux
    port map (
            O => \N__3777\,
            I => data_ready
        );

    \I__579\ : InMux
    port map (
            O => \N__3774\,
            I => \N__3770\
        );

    \I__578\ : InMux
    port map (
            O => \N__3773\,
            I => \N__3767\
        );

    \I__577\ : LocalMux
    port map (
            O => \N__3770\,
            I => delay_counter_16
        );

    \I__576\ : LocalMux
    port map (
            O => \N__3767\,
            I => delay_counter_16
        );

    \I__575\ : InMux
    port map (
            O => \N__3762\,
            I => \N__3758\
        );

    \I__574\ : InMux
    port map (
            O => \N__3761\,
            I => \N__3755\
        );

    \I__573\ : LocalMux
    port map (
            O => \N__3758\,
            I => delay_counter_17
        );

    \I__572\ : LocalMux
    port map (
            O => \N__3755\,
            I => delay_counter_17
        );

    \I__571\ : CascadeMux
    port map (
            O => \N__3750\,
            I => \N__3746\
        );

    \I__570\ : InMux
    port map (
            O => \N__3749\,
            I => \N__3743\
        );

    \I__569\ : InMux
    port map (
            O => \N__3746\,
            I => \N__3740\
        );

    \I__568\ : LocalMux
    port map (
            O => \N__3743\,
            I => delay_counter_15
        );

    \I__567\ : LocalMux
    port map (
            O => \N__3740\,
            I => delay_counter_15
        );

    \I__566\ : InMux
    port map (
            O => \N__3735\,
            I => \N__3732\
        );

    \I__565\ : LocalMux
    port map (
            O => \N__3732\,
            I => \N__3729\
        );

    \I__564\ : Odrv4
    port map (
            O => \N__3729\,
            I => n3069
        );

    \I__563\ : InMux
    port map (
            O => \N__3726\,
            I => \bfn_21_14_0_\
        );

    \I__562\ : InMux
    port map (
            O => \N__3723\,
            I => \N__3719\
        );

    \I__561\ : InMux
    port map (
            O => \N__3722\,
            I => \N__3716\
        );

    \I__560\ : LocalMux
    port map (
            O => \N__3719\,
            I => \N__3713\
        );

    \I__559\ : LocalMux
    port map (
            O => \N__3716\,
            I => \eeprom.delay_counter_9\
        );

    \I__558\ : Odrv4
    port map (
            O => \N__3713\,
            I => \eeprom.delay_counter_9\
        );

    \I__557\ : InMux
    port map (
            O => \N__3708\,
            I => \eeprom.n2864\
        );

    \I__556\ : InMux
    port map (
            O => \N__3705\,
            I => \eeprom.n2865\
        );

    \I__555\ : InMux
    port map (
            O => \N__3702\,
            I => \N__3698\
        );

    \I__554\ : InMux
    port map (
            O => \N__3701\,
            I => \N__3695\
        );

    \I__553\ : LocalMux
    port map (
            O => \N__3698\,
            I => \N__3692\
        );

    \I__552\ : LocalMux
    port map (
            O => \N__3695\,
            I => \eeprom.delay_counter_11\
        );

    \I__551\ : Odrv4
    port map (
            O => \N__3692\,
            I => \eeprom.delay_counter_11\
        );

    \I__550\ : InMux
    port map (
            O => \N__3687\,
            I => \eeprom.n2866\
        );

    \I__549\ : InMux
    port map (
            O => \N__3684\,
            I => \eeprom.n2867\
        );

    \I__548\ : InMux
    port map (
            O => \N__3681\,
            I => \N__3677\
        );

    \I__547\ : InMux
    port map (
            O => \N__3680\,
            I => \N__3674\
        );

    \I__546\ : LocalMux
    port map (
            O => \N__3677\,
            I => \N__3671\
        );

    \I__545\ : LocalMux
    port map (
            O => \N__3674\,
            I => \eeprom.delay_counter_13\
        );

    \I__544\ : Odrv4
    port map (
            O => \N__3671\,
            I => \eeprom.delay_counter_13\
        );

    \I__543\ : InMux
    port map (
            O => \N__3666\,
            I => \eeprom.n2868\
        );

    \I__542\ : InMux
    port map (
            O => \N__3663\,
            I => \N__3659\
        );

    \I__541\ : InMux
    port map (
            O => \N__3662\,
            I => \N__3656\
        );

    \I__540\ : LocalMux
    port map (
            O => \N__3659\,
            I => \N__3653\
        );

    \I__539\ : LocalMux
    port map (
            O => \N__3656\,
            I => \eeprom.delay_counter_14\
        );

    \I__538\ : Odrv4
    port map (
            O => \N__3653\,
            I => \eeprom.delay_counter_14\
        );

    \I__537\ : InMux
    port map (
            O => \N__3648\,
            I => \eeprom.n2869\
        );

    \I__536\ : CascadeMux
    port map (
            O => \N__3645\,
            I => \N__3636\
        );

    \I__535\ : CascadeMux
    port map (
            O => \N__3644\,
            I => \N__3633\
        );

    \I__534\ : CascadeMux
    port map (
            O => \N__3643\,
            I => \N__3630\
        );

    \I__533\ : CascadeMux
    port map (
            O => \N__3642\,
            I => \N__3626\
        );

    \I__532\ : CascadeMux
    port map (
            O => \N__3641\,
            I => \N__3623\
        );

    \I__531\ : CascadeMux
    port map (
            O => \N__3640\,
            I => \N__3620\
        );

    \I__530\ : CascadeMux
    port map (
            O => \N__3639\,
            I => \N__3617\
        );

    \I__529\ : InMux
    port map (
            O => \N__3636\,
            I => \N__3602\
        );

    \I__528\ : InMux
    port map (
            O => \N__3633\,
            I => \N__3602\
        );

    \I__527\ : InMux
    port map (
            O => \N__3630\,
            I => \N__3602\
        );

    \I__526\ : InMux
    port map (
            O => \N__3629\,
            I => \N__3591\
        );

    \I__525\ : InMux
    port map (
            O => \N__3626\,
            I => \N__3591\
        );

    \I__524\ : InMux
    port map (
            O => \N__3623\,
            I => \N__3591\
        );

    \I__523\ : InMux
    port map (
            O => \N__3620\,
            I => \N__3591\
        );

    \I__522\ : InMux
    port map (
            O => \N__3617\,
            I => \N__3591\
        );

    \I__521\ : CascadeMux
    port map (
            O => \N__3616\,
            I => \N__3588\
        );

    \I__520\ : CascadeMux
    port map (
            O => \N__3615\,
            I => \N__3585\
        );

    \I__519\ : CascadeMux
    port map (
            O => \N__3614\,
            I => \N__3582\
        );

    \I__518\ : CascadeMux
    port map (
            O => \N__3613\,
            I => \N__3579\
        );

    \I__517\ : CascadeMux
    port map (
            O => \N__3612\,
            I => \N__3576\
        );

    \I__516\ : CascadeMux
    port map (
            O => \N__3611\,
            I => \N__3573\
        );

    \I__515\ : CascadeMux
    port map (
            O => \N__3610\,
            I => \N__3570\
        );

    \I__514\ : CascadeMux
    port map (
            O => \N__3609\,
            I => \N__3567\
        );

    \I__513\ : LocalMux
    port map (
            O => \N__3602\,
            I => \N__3562\
        );

    \I__512\ : LocalMux
    port map (
            O => \N__3591\,
            I => \N__3562\
        );

    \I__511\ : InMux
    port map (
            O => \N__3588\,
            I => \N__3553\
        );

    \I__510\ : InMux
    port map (
            O => \N__3585\,
            I => \N__3553\
        );

    \I__509\ : InMux
    port map (
            O => \N__3582\,
            I => \N__3553\
        );

    \I__508\ : InMux
    port map (
            O => \N__3579\,
            I => \N__3553\
        );

    \I__507\ : InMux
    port map (
            O => \N__3576\,
            I => \N__3544\
        );

    \I__506\ : InMux
    port map (
            O => \N__3573\,
            I => \N__3544\
        );

    \I__505\ : InMux
    port map (
            O => \N__3570\,
            I => \N__3544\
        );

    \I__504\ : InMux
    port map (
            O => \N__3567\,
            I => \N__3544\
        );

    \I__503\ : Odrv12
    port map (
            O => \N__3562\,
            I => \eeprom.n730\
        );

    \I__502\ : LocalMux
    port map (
            O => \N__3553\,
            I => \eeprom.n730\
        );

    \I__501\ : LocalMux
    port map (
            O => \N__3544\,
            I => \eeprom.n730\
        );

    \I__500\ : InMux
    port map (
            O => \N__3537\,
            I => \eeprom.n2870\
        );

    \I__499\ : InMux
    port map (
            O => \N__3534\,
            I => \N__3530\
        );

    \I__498\ : InMux
    port map (
            O => \N__3533\,
            I => \N__3527\
        );

    \I__497\ : LocalMux
    port map (
            O => \N__3530\,
            I => \N__3524\
        );

    \I__496\ : LocalMux
    port map (
            O => \N__3527\,
            I => \eeprom.delay_counter_15\
        );

    \I__495\ : Odrv4
    port map (
            O => \N__3524\,
            I => \eeprom.delay_counter_15\
        );

    \I__494\ : CascadeMux
    port map (
            O => \N__3519\,
            I => \N__3515\
        );

    \I__493\ : InMux
    port map (
            O => \N__3518\,
            I => \N__3512\
        );

    \I__492\ : InMux
    port map (
            O => \N__3515\,
            I => \N__3509\
        );

    \I__491\ : LocalMux
    port map (
            O => \N__3512\,
            I => \eeprom.delay_counter_0\
        );

    \I__490\ : LocalMux
    port map (
            O => \N__3509\,
            I => \eeprom.delay_counter_0\
        );

    \I__489\ : CascadeMux
    port map (
            O => \N__3504\,
            I => \N__3500\
        );

    \I__488\ : InMux
    port map (
            O => \N__3503\,
            I => \N__3497\
        );

    \I__487\ : InMux
    port map (
            O => \N__3500\,
            I => \N__3494\
        );

    \I__486\ : LocalMux
    port map (
            O => \N__3497\,
            I => \eeprom.delay_counter_1\
        );

    \I__485\ : LocalMux
    port map (
            O => \N__3494\,
            I => \eeprom.delay_counter_1\
        );

    \I__484\ : InMux
    port map (
            O => \N__3489\,
            I => \eeprom.n2856\
        );

    \I__483\ : InMux
    port map (
            O => \N__3486\,
            I => \N__3482\
        );

    \I__482\ : InMux
    port map (
            O => \N__3485\,
            I => \N__3479\
        );

    \I__481\ : LocalMux
    port map (
            O => \N__3482\,
            I => \eeprom.delay_counter_2\
        );

    \I__480\ : LocalMux
    port map (
            O => \N__3479\,
            I => \eeprom.delay_counter_2\
        );

    \I__479\ : InMux
    port map (
            O => \N__3474\,
            I => \eeprom.n2857\
        );

    \I__478\ : InMux
    port map (
            O => \N__3471\,
            I => \N__3467\
        );

    \I__477\ : InMux
    port map (
            O => \N__3470\,
            I => \N__3464\
        );

    \I__476\ : LocalMux
    port map (
            O => \N__3467\,
            I => \eeprom.delay_counter_3\
        );

    \I__475\ : LocalMux
    port map (
            O => \N__3464\,
            I => \eeprom.delay_counter_3\
        );

    \I__474\ : InMux
    port map (
            O => \N__3459\,
            I => \eeprom.n2858\
        );

    \I__473\ : InMux
    port map (
            O => \N__3456\,
            I => \N__3452\
        );

    \I__472\ : InMux
    port map (
            O => \N__3455\,
            I => \N__3449\
        );

    \I__471\ : LocalMux
    port map (
            O => \N__3452\,
            I => \eeprom.delay_counter_4\
        );

    \I__470\ : LocalMux
    port map (
            O => \N__3449\,
            I => \eeprom.delay_counter_4\
        );

    \I__469\ : InMux
    port map (
            O => \N__3444\,
            I => \eeprom.n2859\
        );

    \I__468\ : CascadeMux
    port map (
            O => \N__3441\,
            I => \N__3437\
        );

    \I__467\ : InMux
    port map (
            O => \N__3440\,
            I => \N__3434\
        );

    \I__466\ : InMux
    port map (
            O => \N__3437\,
            I => \N__3431\
        );

    \I__465\ : LocalMux
    port map (
            O => \N__3434\,
            I => \eeprom.delay_counter_5\
        );

    \I__464\ : LocalMux
    port map (
            O => \N__3431\,
            I => \eeprom.delay_counter_5\
        );

    \I__463\ : InMux
    port map (
            O => \N__3426\,
            I => \eeprom.n2860\
        );

    \I__462\ : InMux
    port map (
            O => \N__3423\,
            I => \eeprom.n2861\
        );

    \I__461\ : InMux
    port map (
            O => \N__3420\,
            I => \N__3416\
        );

    \I__460\ : InMux
    port map (
            O => \N__3419\,
            I => \N__3413\
        );

    \I__459\ : LocalMux
    port map (
            O => \N__3416\,
            I => \eeprom.delay_counter_7\
        );

    \I__458\ : LocalMux
    port map (
            O => \N__3413\,
            I => \eeprom.delay_counter_7\
        );

    \I__457\ : InMux
    port map (
            O => \N__3408\,
            I => \eeprom.n2862\
        );

    \I__456\ : InMux
    port map (
            O => \N__3405\,
            I => n2845
        );

    \I__455\ : InMux
    port map (
            O => \N__3402\,
            I => n2846
        );

    \I__454\ : InMux
    port map (
            O => \N__3399\,
            I => n2847
        );

    \I__453\ : InMux
    port map (
            O => \N__3396\,
            I => n2848
        );

    \I__452\ : CascadeMux
    port map (
            O => \N__3393\,
            I => \eeprom.n1704_cascade_\
        );

    \I__451\ : InMux
    port map (
            O => \N__3390\,
            I => \N__3387\
        );

    \I__450\ : LocalMux
    port map (
            O => \N__3387\,
            I => \eeprom.n25\
        );

    \I__449\ : InMux
    port map (
            O => \N__3384\,
            I => \N__3381\
        );

    \I__448\ : LocalMux
    port map (
            O => \N__3381\,
            I => \eeprom.n26_adj_385\
        );

    \I__447\ : InMux
    port map (
            O => \N__3378\,
            I => \N__3375\
        );

    \I__446\ : LocalMux
    port map (
            O => \N__3375\,
            I => \eeprom.n27\
        );

    \I__445\ : InMux
    port map (
            O => \N__3372\,
            I => n2836
        );

    \I__444\ : InMux
    port map (
            O => \N__3369\,
            I => n2837
        );

    \I__443\ : InMux
    port map (
            O => \N__3366\,
            I => n2838
        );

    \I__442\ : InMux
    port map (
            O => \N__3363\,
            I => n2839
        );

    \I__441\ : InMux
    port map (
            O => \N__3360\,
            I => n2840
        );

    \I__440\ : InMux
    port map (
            O => \N__3357\,
            I => \bfn_20_20_0_\
        );

    \I__439\ : InMux
    port map (
            O => \N__3354\,
            I => n2842
        );

    \I__438\ : InMux
    port map (
            O => \N__3351\,
            I => n2843
        );

    \I__437\ : InMux
    port map (
            O => \N__3348\,
            I => n2844
        );

    \I__436\ : InMux
    port map (
            O => \N__3345\,
            I => \N__3341\
        );

    \I__435\ : InMux
    port map (
            O => \N__3344\,
            I => \N__3338\
        );

    \I__434\ : LocalMux
    port map (
            O => \N__3341\,
            I => \N__3335\
        );

    \I__433\ : LocalMux
    port map (
            O => \N__3338\,
            I => delay_counter_10
        );

    \I__432\ : Odrv4
    port map (
            O => \N__3335\,
            I => delay_counter_10
        );

    \I__431\ : InMux
    port map (
            O => \N__3330\,
            I => n2827
        );

    \I__430\ : InMux
    port map (
            O => \N__3327\,
            I => \N__3323\
        );

    \I__429\ : InMux
    port map (
            O => \N__3326\,
            I => \N__3320\
        );

    \I__428\ : LocalMux
    port map (
            O => \N__3323\,
            I => \N__3317\
        );

    \I__427\ : LocalMux
    port map (
            O => \N__3320\,
            I => delay_counter_11
        );

    \I__426\ : Odrv4
    port map (
            O => \N__3317\,
            I => delay_counter_11
        );

    \I__425\ : InMux
    port map (
            O => \N__3312\,
            I => n2828
        );

    \I__424\ : InMux
    port map (
            O => \N__3309\,
            I => \N__3305\
        );

    \I__423\ : InMux
    port map (
            O => \N__3308\,
            I => \N__3302\
        );

    \I__422\ : LocalMux
    port map (
            O => \N__3305\,
            I => \N__3299\
        );

    \I__421\ : LocalMux
    port map (
            O => \N__3302\,
            I => delay_counter_12
        );

    \I__420\ : Odrv4
    port map (
            O => \N__3299\,
            I => delay_counter_12
        );

    \I__419\ : InMux
    port map (
            O => \N__3294\,
            I => n2829
        );

    \I__418\ : InMux
    port map (
            O => \N__3291\,
            I => \N__3287\
        );

    \I__417\ : InMux
    port map (
            O => \N__3290\,
            I => \N__3284\
        );

    \I__416\ : LocalMux
    port map (
            O => \N__3287\,
            I => \N__3281\
        );

    \I__415\ : LocalMux
    port map (
            O => \N__3284\,
            I => delay_counter_13
        );

    \I__414\ : Odrv4
    port map (
            O => \N__3281\,
            I => delay_counter_13
        );

    \I__413\ : InMux
    port map (
            O => \N__3276\,
            I => n2830
        );

    \I__412\ : InMux
    port map (
            O => \N__3273\,
            I => \N__3269\
        );

    \I__411\ : InMux
    port map (
            O => \N__3272\,
            I => \N__3266\
        );

    \I__410\ : LocalMux
    port map (
            O => \N__3269\,
            I => \N__3263\
        );

    \I__409\ : LocalMux
    port map (
            O => \N__3266\,
            I => delay_counter_14
        );

    \I__408\ : Odrv4
    port map (
            O => \N__3263\,
            I => delay_counter_14
        );

    \I__407\ : InMux
    port map (
            O => \N__3258\,
            I => n2831
        );

    \I__406\ : InMux
    port map (
            O => \N__3255\,
            I => n2832
        );

    \I__405\ : InMux
    port map (
            O => \N__3252\,
            I => \bfn_20_19_0_\
        );

    \I__404\ : InMux
    port map (
            O => \N__3249\,
            I => n2834
        );

    \I__403\ : InMux
    port map (
            O => \N__3246\,
            I => n2835
        );

    \I__402\ : InMux
    port map (
            O => \N__3243\,
            I => \N__3239\
        );

    \I__401\ : InMux
    port map (
            O => \N__3242\,
            I => \N__3236\
        );

    \I__400\ : LocalMux
    port map (
            O => \N__3239\,
            I => delay_counter_2
        );

    \I__399\ : LocalMux
    port map (
            O => \N__3236\,
            I => delay_counter_2
        );

    \I__398\ : InMux
    port map (
            O => \N__3231\,
            I => n2819
        );

    \I__397\ : CascadeMux
    port map (
            O => \N__3228\,
            I => \N__3224\
        );

    \I__396\ : InMux
    port map (
            O => \N__3227\,
            I => \N__3221\
        );

    \I__395\ : InMux
    port map (
            O => \N__3224\,
            I => \N__3218\
        );

    \I__394\ : LocalMux
    port map (
            O => \N__3221\,
            I => delay_counter_3
        );

    \I__393\ : LocalMux
    port map (
            O => \N__3218\,
            I => delay_counter_3
        );

    \I__392\ : InMux
    port map (
            O => \N__3213\,
            I => n2820
        );

    \I__391\ : InMux
    port map (
            O => \N__3210\,
            I => \N__3206\
        );

    \I__390\ : InMux
    port map (
            O => \N__3209\,
            I => \N__3203\
        );

    \I__389\ : LocalMux
    port map (
            O => \N__3206\,
            I => delay_counter_4
        );

    \I__388\ : LocalMux
    port map (
            O => \N__3203\,
            I => delay_counter_4
        );

    \I__387\ : InMux
    port map (
            O => \N__3198\,
            I => n2821
        );

    \I__386\ : InMux
    port map (
            O => \N__3195\,
            I => \N__3191\
        );

    \I__385\ : InMux
    port map (
            O => \N__3194\,
            I => \N__3188\
        );

    \I__384\ : LocalMux
    port map (
            O => \N__3191\,
            I => delay_counter_5
        );

    \I__383\ : LocalMux
    port map (
            O => \N__3188\,
            I => delay_counter_5
        );

    \I__382\ : InMux
    port map (
            O => \N__3183\,
            I => n2822
        );

    \I__381\ : InMux
    port map (
            O => \N__3180\,
            I => \N__3176\
        );

    \I__380\ : InMux
    port map (
            O => \N__3179\,
            I => \N__3173\
        );

    \I__379\ : LocalMux
    port map (
            O => \N__3176\,
            I => delay_counter_6
        );

    \I__378\ : LocalMux
    port map (
            O => \N__3173\,
            I => delay_counter_6
        );

    \I__377\ : InMux
    port map (
            O => \N__3168\,
            I => n2823
        );

    \I__376\ : InMux
    port map (
            O => \N__3165\,
            I => \N__3161\
        );

    \I__375\ : InMux
    port map (
            O => \N__3164\,
            I => \N__3158\
        );

    \I__374\ : LocalMux
    port map (
            O => \N__3161\,
            I => delay_counter_7
        );

    \I__373\ : LocalMux
    port map (
            O => \N__3158\,
            I => delay_counter_7
        );

    \I__372\ : InMux
    port map (
            O => \N__3153\,
            I => n2824
        );

    \I__371\ : InMux
    port map (
            O => \N__3150\,
            I => \N__3146\
        );

    \I__370\ : InMux
    port map (
            O => \N__3149\,
            I => \N__3143\
        );

    \I__369\ : LocalMux
    port map (
            O => \N__3146\,
            I => \N__3140\
        );

    \I__368\ : LocalMux
    port map (
            O => \N__3143\,
            I => delay_counter_8
        );

    \I__367\ : Odrv4
    port map (
            O => \N__3140\,
            I => delay_counter_8
        );

    \I__366\ : InMux
    port map (
            O => \N__3135\,
            I => \bfn_20_18_0_\
        );

    \I__365\ : InMux
    port map (
            O => \N__3132\,
            I => \N__3128\
        );

    \I__364\ : InMux
    port map (
            O => \N__3131\,
            I => \N__3125\
        );

    \I__363\ : LocalMux
    port map (
            O => \N__3128\,
            I => \N__3122\
        );

    \I__362\ : LocalMux
    port map (
            O => \N__3125\,
            I => delay_counter_9
        );

    \I__361\ : Odrv4
    port map (
            O => \N__3122\,
            I => delay_counter_9
        );

    \I__360\ : InMux
    port map (
            O => \N__3117\,
            I => n2826
        );

    \I__359\ : InMux
    port map (
            O => \N__3114\,
            I => \N__3111\
        );

    \I__358\ : LocalMux
    port map (
            O => \N__3111\,
            I => n3119
        );

    \I__357\ : InMux
    port map (
            O => \N__3108\,
            I => \N__3101\
        );

    \I__356\ : InMux
    port map (
            O => \N__3107\,
            I => \N__3101\
        );

    \I__355\ : InMux
    port map (
            O => \N__3106\,
            I => \N__3098\
        );

    \I__354\ : LocalMux
    port map (
            O => \N__3101\,
            I => blink_counter_21
        );

    \I__353\ : LocalMux
    port map (
            O => \N__3098\,
            I => blink_counter_21
        );

    \I__352\ : InMux
    port map (
            O => \N__3093\,
            I => \N__3084\
        );

    \I__351\ : InMux
    port map (
            O => \N__3092\,
            I => \N__3084\
        );

    \I__350\ : InMux
    port map (
            O => \N__3091\,
            I => \N__3084\
        );

    \I__349\ : LocalMux
    port map (
            O => \N__3084\,
            I => blink_counter_24
        );

    \I__348\ : CascadeMux
    port map (
            O => \N__3081\,
            I => \N__3077\
        );

    \I__347\ : CascadeMux
    port map (
            O => \N__3080\,
            I => \N__3074\
        );

    \I__346\ : InMux
    port map (
            O => \N__3077\,
            I => \N__3068\
        );

    \I__345\ : InMux
    port map (
            O => \N__3074\,
            I => \N__3068\
        );

    \I__344\ : InMux
    port map (
            O => \N__3073\,
            I => \N__3065\
        );

    \I__343\ : LocalMux
    port map (
            O => \N__3068\,
            I => blink_counter_23
        );

    \I__342\ : LocalMux
    port map (
            O => \N__3065\,
            I => blink_counter_23
        );

    \I__341\ : InMux
    port map (
            O => \N__3060\,
            I => \N__3053\
        );

    \I__340\ : InMux
    port map (
            O => \N__3059\,
            I => \N__3053\
        );

    \I__339\ : InMux
    port map (
            O => \N__3058\,
            I => \N__3050\
        );

    \I__338\ : LocalMux
    port map (
            O => \N__3053\,
            I => blink_counter_22
        );

    \I__337\ : LocalMux
    port map (
            O => \N__3050\,
            I => blink_counter_22
        );

    \I__336\ : InMux
    port map (
            O => \N__3045\,
            I => \N__3042\
        );

    \I__335\ : LocalMux
    port map (
            O => \N__3042\,
            I => n3120
        );

    \I__334\ : CascadeMux
    port map (
            O => \N__3039\,
            I => \n13_adj_391_cascade_\
        );

    \I__333\ : InMux
    port map (
            O => \N__3036\,
            I => \N__3033\
        );

    \I__332\ : LocalMux
    port map (
            O => \N__3033\,
            I => n14
        );

    \I__331\ : CascadeMux
    port map (
            O => \N__3030\,
            I => \n18_cascade_\
        );

    \I__330\ : CascadeMux
    port map (
            O => \N__3027\,
            I => \n3114_cascade_\
        );

    \I__329\ : CascadeMux
    port map (
            O => \N__3024\,
            I => \N__3020\
        );

    \I__328\ : InMux
    port map (
            O => \N__3023\,
            I => \N__3017\
        );

    \I__327\ : InMux
    port map (
            O => \N__3020\,
            I => \N__3014\
        );

    \I__326\ : LocalMux
    port map (
            O => \N__3017\,
            I => delay_counter_0
        );

    \I__325\ : LocalMux
    port map (
            O => \N__3014\,
            I => delay_counter_0
        );

    \I__324\ : InMux
    port map (
            O => \N__3009\,
            I => \bfn_20_17_0_\
        );

    \I__323\ : InMux
    port map (
            O => \N__3006\,
            I => \N__3002\
        );

    \I__322\ : InMux
    port map (
            O => \N__3005\,
            I => \N__2999\
        );

    \I__321\ : LocalMux
    port map (
            O => \N__3002\,
            I => delay_counter_1
        );

    \I__320\ : LocalMux
    port map (
            O => \N__2999\,
            I => delay_counter_1
        );

    \I__319\ : InMux
    port map (
            O => \N__2994\,
            I => n2818
        );

    \I__318\ : InMux
    port map (
            O => \N__2991\,
            I => \N__2988\
        );

    \I__317\ : LocalMux
    port map (
            O => \N__2988\,
            I => n9
        );

    \I__316\ : InMux
    port map (
            O => \N__2985\,
            I => n2892
        );

    \I__315\ : InMux
    port map (
            O => \N__2982\,
            I => \N__2979\
        );

    \I__314\ : LocalMux
    port map (
            O => \N__2979\,
            I => n8
        );

    \I__313\ : InMux
    port map (
            O => \N__2976\,
            I => n2893
        );

    \I__312\ : InMux
    port map (
            O => \N__2973\,
            I => \N__2970\
        );

    \I__311\ : LocalMux
    port map (
            O => \N__2970\,
            I => n7
        );

    \I__310\ : InMux
    port map (
            O => \N__2967\,
            I => n2894
        );

    \I__309\ : InMux
    port map (
            O => \N__2964\,
            I => \N__2961\
        );

    \I__308\ : LocalMux
    port map (
            O => \N__2961\,
            I => n6_adj_392
        );

    \I__307\ : InMux
    port map (
            O => \N__2958\,
            I => n2895
        );

    \I__306\ : InMux
    port map (
            O => \N__2955\,
            I => n2896
        );

    \I__305\ : InMux
    port map (
            O => \N__2952\,
            I => n2897
        );

    \I__304\ : InMux
    port map (
            O => \N__2949\,
            I => n2898
        );

    \I__303\ : InMux
    port map (
            O => \N__2946\,
            I => \bfn_17_20_0_\
        );

    \I__302\ : InMux
    port map (
            O => \N__2943\,
            I => n2900
        );

    \I__301\ : InMux
    port map (
            O => \N__2940\,
            I => \N__2936\
        );

    \I__300\ : InMux
    port map (
            O => \N__2939\,
            I => \N__2933\
        );

    \I__299\ : LocalMux
    port map (
            O => \N__2936\,
            I => blink_counter_25
        );

    \I__298\ : LocalMux
    port map (
            O => \N__2933\,
            I => blink_counter_25
        );

    \I__297\ : InMux
    port map (
            O => \N__2928\,
            I => \N__2925\
        );

    \I__296\ : LocalMux
    port map (
            O => \N__2925\,
            I => n17
        );

    \I__295\ : InMux
    port map (
            O => \N__2922\,
            I => n2884
        );

    \I__294\ : InMux
    port map (
            O => \N__2919\,
            I => \N__2916\
        );

    \I__293\ : LocalMux
    port map (
            O => \N__2916\,
            I => n16
        );

    \I__292\ : InMux
    port map (
            O => \N__2913\,
            I => n2885
        );

    \I__291\ : InMux
    port map (
            O => \N__2910\,
            I => \N__2907\
        );

    \I__290\ : LocalMux
    port map (
            O => \N__2907\,
            I => n15_adj_396
        );

    \I__289\ : InMux
    port map (
            O => \N__2904\,
            I => n2886
        );

    \I__288\ : InMux
    port map (
            O => \N__2901\,
            I => \N__2898\
        );

    \I__287\ : LocalMux
    port map (
            O => \N__2898\,
            I => n14_adj_395
        );

    \I__286\ : InMux
    port map (
            O => \N__2895\,
            I => n2887
        );

    \I__285\ : InMux
    port map (
            O => \N__2892\,
            I => \N__2889\
        );

    \I__284\ : LocalMux
    port map (
            O => \N__2889\,
            I => n13_adj_394
        );

    \I__283\ : InMux
    port map (
            O => \N__2886\,
            I => n2888
        );

    \I__282\ : InMux
    port map (
            O => \N__2883\,
            I => \N__2880\
        );

    \I__281\ : LocalMux
    port map (
            O => \N__2880\,
            I => n12_adj_393
        );

    \I__280\ : InMux
    port map (
            O => \N__2877\,
            I => n2889
        );

    \I__279\ : InMux
    port map (
            O => \N__2874\,
            I => \N__2871\
        );

    \I__278\ : LocalMux
    port map (
            O => \N__2871\,
            I => n11
        );

    \I__277\ : InMux
    port map (
            O => \N__2868\,
            I => n2890
        );

    \I__276\ : InMux
    port map (
            O => \N__2865\,
            I => \N__2862\
        );

    \I__275\ : LocalMux
    port map (
            O => \N__2862\,
            I => n10
        );

    \I__274\ : InMux
    port map (
            O => \N__2859\,
            I => \bfn_17_19_0_\
        );

    \I__273\ : InMux
    port map (
            O => \N__2856\,
            I => \N__2853\
        );

    \I__272\ : LocalMux
    port map (
            O => \N__2853\,
            I => n26
        );

    \I__271\ : InMux
    port map (
            O => \N__2850\,
            I => \bfn_17_17_0_\
        );

    \I__270\ : InMux
    port map (
            O => \N__2847\,
            I => \N__2844\
        );

    \I__269\ : LocalMux
    port map (
            O => \N__2844\,
            I => n25_adj_402
        );

    \I__268\ : InMux
    port map (
            O => \N__2841\,
            I => n2876
        );

    \I__267\ : InMux
    port map (
            O => \N__2838\,
            I => \N__2835\
        );

    \I__266\ : LocalMux
    port map (
            O => \N__2835\,
            I => n24_adj_401
        );

    \I__265\ : InMux
    port map (
            O => \N__2832\,
            I => n2877
        );

    \I__264\ : InMux
    port map (
            O => \N__2829\,
            I => \N__2826\
        );

    \I__263\ : LocalMux
    port map (
            O => \N__2826\,
            I => n23_adj_400
        );

    \I__262\ : InMux
    port map (
            O => \N__2823\,
            I => n2878
        );

    \I__261\ : InMux
    port map (
            O => \N__2820\,
            I => \N__2817\
        );

    \I__260\ : LocalMux
    port map (
            O => \N__2817\,
            I => n22_adj_399
        );

    \I__259\ : InMux
    port map (
            O => \N__2814\,
            I => n2879
        );

    \I__258\ : InMux
    port map (
            O => \N__2811\,
            I => \N__2808\
        );

    \I__257\ : LocalMux
    port map (
            O => \N__2808\,
            I => n21
        );

    \I__256\ : InMux
    port map (
            O => \N__2805\,
            I => n2880
        );

    \I__255\ : InMux
    port map (
            O => \N__2802\,
            I => \N__2799\
        );

    \I__254\ : LocalMux
    port map (
            O => \N__2799\,
            I => n20_adj_398
        );

    \I__253\ : InMux
    port map (
            O => \N__2796\,
            I => n2881
        );

    \I__252\ : InMux
    port map (
            O => \N__2793\,
            I => \N__2790\
        );

    \I__251\ : LocalMux
    port map (
            O => \N__2790\,
            I => n19
        );

    \I__250\ : InMux
    port map (
            O => \N__2787\,
            I => n2882
        );

    \I__249\ : InMux
    port map (
            O => \N__2784\,
            I => \N__2781\
        );

    \I__248\ : LocalMux
    port map (
            O => \N__2781\,
            I => n18_adj_397
        );

    \I__247\ : InMux
    port map (
            O => \N__2778\,
            I => \bfn_17_18_0_\
        );

    \I__246\ : IoInMux
    port map (
            O => \N__2775\,
            I => \N__2772\
        );

    \I__245\ : LocalMux
    port map (
            O => \N__2772\,
            I => \N__2769\
        );

    \I__244\ : IoSpan4Mux
    port map (
            O => \N__2769\,
            I => \N__2766\
        );

    \I__243\ : Sp12to4
    port map (
            O => \N__2766\,
            I => \N__2763\
        );

    \I__242\ : Span12Mux_v
    port map (
            O => \N__2763\,
            I => \N__2760\
        );

    \I__241\ : Odrv12
    port map (
            O => \N__2760\,
            I => \LED_c\
        );

    \I__240\ : IoInMux
    port map (
            O => \N__2757\,
            I => \N__2754\
        );

    \I__239\ : LocalMux
    port map (
            O => \N__2754\,
            I => \N__2751\
        );

    \I__238\ : IoSpan4Mux
    port map (
            O => \N__2751\,
            I => \N__2748\
        );

    \I__237\ : IoSpan4Mux
    port map (
            O => \N__2748\,
            I => \N__2745\
        );

    \I__236\ : IoSpan4Mux
    port map (
            O => \N__2745\,
            I => \N__2742\
        );

    \I__235\ : Odrv4
    port map (
            O => \N__2742\,
            I => \CLK_pad_gb_input\
        );

    \INVeeprom.i2c.i2c_scl_enable_123C\ : INV
    port map (
            O => \INVeeprom.i2c.i2c_scl_enable_123C_net\,
            I => \N__6478\
        );

    \INVeeprom.i2c.sda_out_132C\ : INV
    port map (
            O => \INVeeprom.i2c.sda_out_132C_net\,
            I => \N__6459\
        );

    \INVeeprom.i2c.write_enable_131C\ : INV
    port map (
            O => \INVeeprom.i2c.write_enable_131C_net\,
            I => \N__6436\
        );

    \IN_MUX_bfv_26_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_26_14_0_\
        );

    \IN_MUX_bfv_27_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_27_13_0_\
        );

    \IN_MUX_bfv_21_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_21_13_0_\
        );

    \IN_MUX_bfv_21_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \eeprom.n2863\,
            carryinitout => \bfn_21_14_0_\
        );

    \IN_MUX_bfv_17_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_17_17_0_\
        );

    \IN_MUX_bfv_17_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n2883,
            carryinitout => \bfn_17_18_0_\
        );

    \IN_MUX_bfv_17_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n2891,
            carryinitout => \bfn_17_19_0_\
        );

    \IN_MUX_bfv_17_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n2899,
            carryinitout => \bfn_17_20_0_\
        );

    \IN_MUX_bfv_20_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_20_17_0_\
        );

    \IN_MUX_bfv_20_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n2825,
            carryinitout => \bfn_20_18_0_\
        );

    \IN_MUX_bfv_20_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n2833,
            carryinitout => \bfn_20_19_0_\
        );

    \IN_MUX_bfv_20_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n2841,
            carryinitout => \bfn_20_20_0_\
        );

    \CLK_pad_gb\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__2757\,
            GLOBALBUFFEROUTPUT => \CLK_c\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \i2105_3_lut_LC_16_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000110111011"
        )
    port map (
            in0 => \N__2940\,
            in1 => \N__3114\,
            in2 => \_gnd_net_\,
            in3 => \N__3045\,
            lcout => \LED_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_410__i0_LC_17_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2856\,
            in2 => \_gnd_net_\,
            in3 => \N__2850\,
            lcout => n26,
            ltout => OPEN,
            carryin => \bfn_17_17_0_\,
            carryout => n2876,
            clk => \N__6732\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_410__i1_LC_17_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2847\,
            in2 => \_gnd_net_\,
            in3 => \N__2841\,
            lcout => n25_adj_402,
            ltout => OPEN,
            carryin => n2876,
            carryout => n2877,
            clk => \N__6732\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_410__i2_LC_17_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2838\,
            in2 => \_gnd_net_\,
            in3 => \N__2832\,
            lcout => n24_adj_401,
            ltout => OPEN,
            carryin => n2877,
            carryout => n2878,
            clk => \N__6732\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_410__i3_LC_17_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2829\,
            in2 => \_gnd_net_\,
            in3 => \N__2823\,
            lcout => n23_adj_400,
            ltout => OPEN,
            carryin => n2878,
            carryout => n2879,
            clk => \N__6732\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_410__i4_LC_17_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2820\,
            in2 => \_gnd_net_\,
            in3 => \N__2814\,
            lcout => n22_adj_399,
            ltout => OPEN,
            carryin => n2879,
            carryout => n2880,
            clk => \N__6732\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_410__i5_LC_17_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2811\,
            in2 => \_gnd_net_\,
            in3 => \N__2805\,
            lcout => n21,
            ltout => OPEN,
            carryin => n2880,
            carryout => n2881,
            clk => \N__6732\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_410__i6_LC_17_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2802\,
            in2 => \_gnd_net_\,
            in3 => \N__2796\,
            lcout => n20_adj_398,
            ltout => OPEN,
            carryin => n2881,
            carryout => n2882,
            clk => \N__6732\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_410__i7_LC_17_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2793\,
            in2 => \_gnd_net_\,
            in3 => \N__2787\,
            lcout => n19,
            ltout => OPEN,
            carryin => n2882,
            carryout => n2883,
            clk => \N__6732\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_410__i8_LC_17_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2784\,
            in2 => \_gnd_net_\,
            in3 => \N__2778\,
            lcout => n18_adj_397,
            ltout => OPEN,
            carryin => \bfn_17_18_0_\,
            carryout => n2884,
            clk => \N__6733\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_410__i9_LC_17_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2928\,
            in2 => \_gnd_net_\,
            in3 => \N__2922\,
            lcout => n17,
            ltout => OPEN,
            carryin => n2884,
            carryout => n2885,
            clk => \N__6733\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_410__i10_LC_17_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2919\,
            in2 => \_gnd_net_\,
            in3 => \N__2913\,
            lcout => n16,
            ltout => OPEN,
            carryin => n2885,
            carryout => n2886,
            clk => \N__6733\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_410__i11_LC_17_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2910\,
            in2 => \_gnd_net_\,
            in3 => \N__2904\,
            lcout => n15_adj_396,
            ltout => OPEN,
            carryin => n2886,
            carryout => n2887,
            clk => \N__6733\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_410__i12_LC_17_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2901\,
            in2 => \_gnd_net_\,
            in3 => \N__2895\,
            lcout => n14_adj_395,
            ltout => OPEN,
            carryin => n2887,
            carryout => n2888,
            clk => \N__6733\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_410__i13_LC_17_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2892\,
            in2 => \_gnd_net_\,
            in3 => \N__2886\,
            lcout => n13_adj_394,
            ltout => OPEN,
            carryin => n2888,
            carryout => n2889,
            clk => \N__6733\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_410__i14_LC_17_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2883\,
            in2 => \_gnd_net_\,
            in3 => \N__2877\,
            lcout => n12_adj_393,
            ltout => OPEN,
            carryin => n2889,
            carryout => n2890,
            clk => \N__6733\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_410__i15_LC_17_18_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2874\,
            in2 => \_gnd_net_\,
            in3 => \N__2868\,
            lcout => n11,
            ltout => OPEN,
            carryin => n2890,
            carryout => n2891,
            clk => \N__6733\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_410__i16_LC_17_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2865\,
            in2 => \_gnd_net_\,
            in3 => \N__2859\,
            lcout => n10,
            ltout => OPEN,
            carryin => \bfn_17_19_0_\,
            carryout => n2892,
            clk => \N__6734\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_410__i17_LC_17_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2991\,
            in2 => \_gnd_net_\,
            in3 => \N__2985\,
            lcout => n9,
            ltout => OPEN,
            carryin => n2892,
            carryout => n2893,
            clk => \N__6734\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_410__i18_LC_17_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2982\,
            in2 => \_gnd_net_\,
            in3 => \N__2976\,
            lcout => n8,
            ltout => OPEN,
            carryin => n2893,
            carryout => n2894,
            clk => \N__6734\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_410__i19_LC_17_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2973\,
            in2 => \_gnd_net_\,
            in3 => \N__2967\,
            lcout => n7,
            ltout => OPEN,
            carryin => n2894,
            carryout => n2895,
            clk => \N__6734\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_410__i20_LC_17_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2964\,
            in2 => \_gnd_net_\,
            in3 => \N__2958\,
            lcout => n6_adj_392,
            ltout => OPEN,
            carryin => n2895,
            carryout => n2896,
            clk => \N__6734\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_410__i21_LC_17_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3106\,
            in2 => \_gnd_net_\,
            in3 => \N__2955\,
            lcout => blink_counter_21,
            ltout => OPEN,
            carryin => n2896,
            carryout => n2897,
            clk => \N__6734\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_410__i22_LC_17_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3058\,
            in2 => \_gnd_net_\,
            in3 => \N__2952\,
            lcout => blink_counter_22,
            ltout => OPEN,
            carryin => n2897,
            carryout => n2898,
            clk => \N__6734\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_410__i23_LC_17_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3073\,
            in2 => \_gnd_net_\,
            in3 => \N__2949\,
            lcout => blink_counter_23,
            ltout => OPEN,
            carryin => n2898,
            carryout => n2899,
            clk => \N__6734\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_410__i24_LC_17_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3091\,
            in2 => \_gnd_net_\,
            in3 => \N__2946\,
            lcout => blink_counter_24,
            ltout => OPEN,
            carryin => \bfn_17_20_0_\,
            carryout => n2900,
            clk => \N__6736\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_410__i25_LC_17_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2939\,
            in2 => \_gnd_net_\,
            in3 => \N__2943\,
            lcout => blink_counter_25,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6736\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2103_4_lut_LC_17_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101000100010"
        )
    port map (
            in0 => \N__3107\,
            in1 => \N__3092\,
            in2 => \N__3080\,
            in3 => \N__3059\,
            lcout => n3119,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2104_4_lut_LC_17_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101011111000"
        )
    port map (
            in0 => \N__3108\,
            in1 => \N__3093\,
            in2 => \N__3081\,
            in3 => \N__3060\,
            lcout => n3120,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i6_4_lut_LC_20_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__3209\,
            in1 => \N__3179\,
            in2 => \N__3228\,
            in3 => \N__3164\,
            lcout => n14,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i5_4_lut_LC_20_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__3005\,
            in1 => \N__3242\,
            in2 => \N__3024\,
            in3 => \N__3194\,
            lcout => OPEN,
            ltout => \n13_adj_391_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i530_3_lut_LC_20_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3150\,
            in2 => \N__3039\,
            in3 => \N__3036\,
            lcout => OPEN,
            ltout => \n18_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i3_4_lut_LC_20_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__3345\,
            in1 => \N__3327\,
            in2 => \N__3030\,
            in3 => \N__3132\,
            lcout => OPEN,
            ltout => \n3114_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i3_4_lut_adj_9_LC_20_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__3291\,
            in1 => \N__3273\,
            in2 => \N__3027\,
            in3 => \N__3309\,
            lcout => n3069,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_counter_i0_LC_20_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3023\,
            in2 => \_gnd_net_\,
            in3 => \N__3009\,
            lcout => delay_counter_0,
            ltout => OPEN,
            carryin => \bfn_20_17_0_\,
            carryout => n2818,
            clk => \N__6735\,
            ce => \N__4320\,
            sr => \N__3940\
        );

    \delay_counter_i1_LC_20_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3006\,
            in2 => \_gnd_net_\,
            in3 => \N__2994\,
            lcout => delay_counter_1,
            ltout => OPEN,
            carryin => n2818,
            carryout => n2819,
            clk => \N__6735\,
            ce => \N__4320\,
            sr => \N__3940\
        );

    \delay_counter_i2_LC_20_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3243\,
            in2 => \_gnd_net_\,
            in3 => \N__3231\,
            lcout => delay_counter_2,
            ltout => OPEN,
            carryin => n2819,
            carryout => n2820,
            clk => \N__6735\,
            ce => \N__4320\,
            sr => \N__3940\
        );

    \delay_counter_i3_LC_20_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3227\,
            in2 => \_gnd_net_\,
            in3 => \N__3213\,
            lcout => delay_counter_3,
            ltout => OPEN,
            carryin => n2820,
            carryout => n2821,
            clk => \N__6735\,
            ce => \N__4320\,
            sr => \N__3940\
        );

    \delay_counter_i4_LC_20_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3210\,
            in2 => \_gnd_net_\,
            in3 => \N__3198\,
            lcout => delay_counter_4,
            ltout => OPEN,
            carryin => n2821,
            carryout => n2822,
            clk => \N__6735\,
            ce => \N__4320\,
            sr => \N__3940\
        );

    \delay_counter_i5_LC_20_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3195\,
            in2 => \_gnd_net_\,
            in3 => \N__3183\,
            lcout => delay_counter_5,
            ltout => OPEN,
            carryin => n2822,
            carryout => n2823,
            clk => \N__6735\,
            ce => \N__4320\,
            sr => \N__3940\
        );

    \delay_counter_i6_LC_20_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3180\,
            in2 => \_gnd_net_\,
            in3 => \N__3168\,
            lcout => delay_counter_6,
            ltout => OPEN,
            carryin => n2823,
            carryout => n2824,
            clk => \N__6735\,
            ce => \N__4320\,
            sr => \N__3940\
        );

    \delay_counter_i7_LC_20_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3165\,
            in2 => \_gnd_net_\,
            in3 => \N__3153\,
            lcout => delay_counter_7,
            ltout => OPEN,
            carryin => n2824,
            carryout => n2825,
            clk => \N__6735\,
            ce => \N__4320\,
            sr => \N__3940\
        );

    \delay_counter_i8_LC_20_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3149\,
            in2 => \_gnd_net_\,
            in3 => \N__3135\,
            lcout => delay_counter_8,
            ltout => OPEN,
            carryin => \bfn_20_18_0_\,
            carryout => n2826,
            clk => \N__6738\,
            ce => \N__4319\,
            sr => \N__3939\
        );

    \delay_counter_i9_LC_20_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3131\,
            in2 => \_gnd_net_\,
            in3 => \N__3117\,
            lcout => delay_counter_9,
            ltout => OPEN,
            carryin => n2826,
            carryout => n2827,
            clk => \N__6738\,
            ce => \N__4319\,
            sr => \N__3939\
        );

    \delay_counter_i10_LC_20_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3344\,
            in2 => \_gnd_net_\,
            in3 => \N__3330\,
            lcout => delay_counter_10,
            ltout => OPEN,
            carryin => n2827,
            carryout => n2828,
            clk => \N__6738\,
            ce => \N__4319\,
            sr => \N__3939\
        );

    \delay_counter_i11_LC_20_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3326\,
            in2 => \_gnd_net_\,
            in3 => \N__3312\,
            lcout => delay_counter_11,
            ltout => OPEN,
            carryin => n2828,
            carryout => n2829,
            clk => \N__6738\,
            ce => \N__4319\,
            sr => \N__3939\
        );

    \delay_counter_i12_LC_20_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3308\,
            in2 => \_gnd_net_\,
            in3 => \N__3294\,
            lcout => delay_counter_12,
            ltout => OPEN,
            carryin => n2829,
            carryout => n2830,
            clk => \N__6738\,
            ce => \N__4319\,
            sr => \N__3939\
        );

    \delay_counter_i13_LC_20_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3290\,
            in2 => \_gnd_net_\,
            in3 => \N__3276\,
            lcout => delay_counter_13,
            ltout => OPEN,
            carryin => n2830,
            carryout => n2831,
            clk => \N__6738\,
            ce => \N__4319\,
            sr => \N__3939\
        );

    \delay_counter_i14_LC_20_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3272\,
            in2 => \_gnd_net_\,
            in3 => \N__3258\,
            lcout => delay_counter_14,
            ltout => OPEN,
            carryin => n2831,
            carryout => n2832,
            clk => \N__6738\,
            ce => \N__4319\,
            sr => \N__3939\
        );

    \delay_counter_i15_LC_20_18_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3749\,
            in2 => \_gnd_net_\,
            in3 => \N__3255\,
            lcout => delay_counter_15,
            ltout => OPEN,
            carryin => n2832,
            carryout => n2833,
            clk => \N__6738\,
            ce => \N__4319\,
            sr => \N__3939\
        );

    \delay_counter_i16_LC_20_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3774\,
            in2 => \_gnd_net_\,
            in3 => \N__3252\,
            lcout => delay_counter_16,
            ltout => OPEN,
            carryin => \bfn_20_19_0_\,
            carryout => n2834,
            clk => \N__6739\,
            ce => \N__4311\,
            sr => \N__3941\
        );

    \delay_counter_i17_LC_20_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3762\,
            in2 => \_gnd_net_\,
            in3 => \N__3249\,
            lcout => delay_counter_17,
            ltout => OPEN,
            carryin => n2834,
            carryout => n2835,
            clk => \N__6739\,
            ce => \N__4311\,
            sr => \N__3941\
        );

    \delay_counter_i18_LC_20_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4032\,
            in2 => \_gnd_net_\,
            in3 => \N__3246\,
            lcout => delay_counter_18,
            ltout => OPEN,
            carryin => n2835,
            carryout => n2836,
            clk => \N__6739\,
            ce => \N__4311\,
            sr => \N__3941\
        );

    \delay_counter_i19_LC_20_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3876\,
            in2 => \_gnd_net_\,
            in3 => \N__3372\,
            lcout => delay_counter_19,
            ltout => OPEN,
            carryin => n2836,
            carryout => n2837,
            clk => \N__6739\,
            ce => \N__4311\,
            sr => \N__3941\
        );

    \delay_counter_i20_LC_20_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3890\,
            in2 => \_gnd_net_\,
            in3 => \N__3369\,
            lcout => delay_counter_20,
            ltout => OPEN,
            carryin => n2837,
            carryout => n2838,
            clk => \N__6739\,
            ce => \N__4311\,
            sr => \N__3941\
        );

    \delay_counter_i21_LC_20_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3918\,
            in2 => \_gnd_net_\,
            in3 => \N__3366\,
            lcout => delay_counter_21,
            ltout => OPEN,
            carryin => n2838,
            carryout => n2839,
            clk => \N__6739\,
            ce => \N__4311\,
            sr => \N__3941\
        );

    \delay_counter_i22_LC_20_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4176\,
            in2 => \_gnd_net_\,
            in3 => \N__3363\,
            lcout => delay_counter_22,
            ltout => OPEN,
            carryin => n2839,
            carryout => n2840,
            clk => \N__6739\,
            ce => \N__4311\,
            sr => \N__3941\
        );

    \delay_counter_i23_LC_20_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3984\,
            in2 => \_gnd_net_\,
            in3 => \N__3360\,
            lcout => delay_counter_23,
            ltout => OPEN,
            carryin => n2840,
            carryout => n2841,
            clk => \N__6739\,
            ce => \N__4311\,
            sr => \N__3941\
        );

    \delay_counter_i24_LC_20_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4016\,
            in2 => \_gnd_net_\,
            in3 => \N__3357\,
            lcout => delay_counter_24,
            ltout => OPEN,
            carryin => \bfn_20_20_0_\,
            carryout => n2842,
            clk => \N__6741\,
            ce => \N__4315\,
            sr => \N__3948\
        );

    \delay_counter_i25_LC_20_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3906\,
            in2 => \_gnd_net_\,
            in3 => \N__3354\,
            lcout => delay_counter_25,
            ltout => OPEN,
            carryin => n2842,
            carryout => n2843,
            clk => \N__6741\,
            ce => \N__4315\,
            sr => \N__3948\
        );

    \delay_counter_i26_LC_20_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4151\,
            in2 => \_gnd_net_\,
            in3 => \N__3351\,
            lcout => delay_counter_26,
            ltout => OPEN,
            carryin => n2843,
            carryout => n2844,
            clk => \N__6741\,
            ce => \N__4315\,
            sr => \N__3948\
        );

    \delay_counter_i27_LC_20_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4001\,
            in2 => \_gnd_net_\,
            in3 => \N__3348\,
            lcout => delay_counter_27,
            ltout => OPEN,
            carryin => n2844,
            carryout => n2845,
            clk => \N__6741\,
            ce => \N__4315\,
            sr => \N__3948\
        );

    \delay_counter_i28_LC_20_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4137\,
            in2 => \_gnd_net_\,
            in3 => \N__3405\,
            lcout => delay_counter_28,
            ltout => OPEN,
            carryin => n2845,
            carryout => n2846,
            clk => \N__6741\,
            ce => \N__4315\,
            sr => \N__3948\
        );

    \delay_counter_i29_LC_20_20_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4046\,
            in2 => \_gnd_net_\,
            in3 => \N__3402\,
            lcout => delay_counter_29,
            ltout => OPEN,
            carryin => n2846,
            carryout => n2847,
            clk => \N__6741\,
            ce => \N__4315\,
            sr => \N__3948\
        );

    \delay_counter_i30_LC_20_20_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4164\,
            in2 => \_gnd_net_\,
            in3 => \N__3399\,
            lcout => delay_counter_30,
            ltout => OPEN,
            carryin => n2847,
            carryout => n2848,
            clk => \N__6741\,
            ce => \N__4315\,
            sr => \N__3948\
        );

    \delay_counter_i31_LC_20_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3968\,
            in2 => \_gnd_net_\,
            in3 => \N__3396\,
            lcout => delay_counter_31,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6741\,
            ce => \N__4315\,
            sr => \N__3948\
        );

    \eeprom.i15_4_lut_LC_21_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__3384\,
            in1 => \N__3378\,
            in2 => \N__4062\,
            in3 => \N__3390\,
            lcout => \eeprom.n1704\,
            ltout => \eeprom.n1704_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2156_2_lut_3_lut_4_lut_LC_21_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__6126\,
            in1 => \N__5541\,
            in2 => \N__3393\,
            in3 => \N__5881\,
            lcout => \eeprom.n730\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i9_4_lut_LC_21_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__3681\,
            in1 => \N__3723\,
            in2 => \N__3519\,
            in3 => \N__3455\,
            lcout => \eeprom.n25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i10_4_lut_LC_21_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__3485\,
            in1 => \N__3419\,
            in2 => \N__3441\,
            in3 => \N__3702\,
            lcout => \eeprom.n26_adj_385\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i11_4_lut_LC_21_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__3663\,
            in1 => \N__3470\,
            in2 => \N__3504\,
            in3 => \N__3534\,
            lcout => \eeprom.n27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.i1_2_lut_LC_21_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010001000100"
        )
    port map (
            in0 => \N__5700\,
            in1 => \N__5993\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \eeprom.i2c.n7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.delay_counter_i0_i0_LC_21_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3518\,
            in2 => \N__3609\,
            in3 => \_gnd_net_\,
            lcout => \eeprom.delay_counter_0\,
            ltout => OPEN,
            carryin => \bfn_21_13_0_\,
            carryout => \eeprom.n2856\,
            clk => \N__6747\,
            ce => \N__3834\,
            sr => \N__3807\
        );

    \eeprom.delay_counter_i0_i1_LC_21_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3503\,
            in2 => \N__3613\,
            in3 => \N__3489\,
            lcout => \eeprom.delay_counter_1\,
            ltout => OPEN,
            carryin => \eeprom.n2856\,
            carryout => \eeprom.n2857\,
            clk => \N__6747\,
            ce => \N__3834\,
            sr => \N__3807\
        );

    \eeprom.delay_counter_i0_i2_LC_21_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3486\,
            in2 => \N__3610\,
            in3 => \N__3474\,
            lcout => \eeprom.delay_counter_2\,
            ltout => OPEN,
            carryin => \eeprom.n2857\,
            carryout => \eeprom.n2858\,
            clk => \N__6747\,
            ce => \N__3834\,
            sr => \N__3807\
        );

    \eeprom.delay_counter_i0_i3_LC_21_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3471\,
            in2 => \N__3614\,
            in3 => \N__3459\,
            lcout => \eeprom.delay_counter_3\,
            ltout => OPEN,
            carryin => \eeprom.n2858\,
            carryout => \eeprom.n2859\,
            clk => \N__6747\,
            ce => \N__3834\,
            sr => \N__3807\
        );

    \eeprom.delay_counter_i0_i4_LC_21_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1001",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3456\,
            in2 => \N__3611\,
            in3 => \N__3444\,
            lcout => \eeprom.delay_counter_4\,
            ltout => OPEN,
            carryin => \eeprom.n2859\,
            carryout => \eeprom.n2860\,
            clk => \N__6747\,
            ce => \N__3834\,
            sr => \N__3807\
        );

    \eeprom.delay_counter_i0_i5_LC_21_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3440\,
            in2 => \N__3615\,
            in3 => \N__3426\,
            lcout => \eeprom.delay_counter_5\,
            ltout => OPEN,
            carryin => \eeprom.n2860\,
            carryout => \eeprom.n2861\,
            clk => \N__6747\,
            ce => \N__3834\,
            sr => \N__3807\
        );

    \eeprom.delay_counter_i0_i6_LC_21_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1001",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4074\,
            in2 => \N__3612\,
            in3 => \N__3423\,
            lcout => \eeprom.delay_counter_6\,
            ltout => OPEN,
            carryin => \eeprom.n2861\,
            carryout => \eeprom.n2862\,
            clk => \N__6747\,
            ce => \N__3834\,
            sr => \N__3807\
        );

    \eeprom.delay_counter_i0_i7_LC_21_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1001",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3420\,
            in2 => \N__3616\,
            in3 => \N__3408\,
            lcout => \eeprom.delay_counter_7\,
            ltout => OPEN,
            carryin => \eeprom.n2862\,
            carryout => \eeprom.n2863\,
            clk => \N__6747\,
            ce => \N__3834\,
            sr => \N__3807\
        );

    \eeprom.delay_counter_i0_i8_LC_21_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1001",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4088\,
            in2 => \N__3639\,
            in3 => \N__3726\,
            lcout => \eeprom.delay_counter_8\,
            ltout => OPEN,
            carryin => \bfn_21_14_0_\,
            carryout => \eeprom.n2864\,
            clk => \N__6746\,
            ce => \N__3830\,
            sr => \N__3806\
        );

    \eeprom.delay_counter_i0_i9_LC_21_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1001",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3722\,
            in2 => \N__3643\,
            in3 => \N__3708\,
            lcout => \eeprom.delay_counter_9\,
            ltout => OPEN,
            carryin => \eeprom.n2864\,
            carryout => \eeprom.n2865\,
            clk => \N__6746\,
            ce => \N__3830\,
            sr => \N__3806\
        );

    \eeprom.delay_counter_i0_i10_LC_21_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1001",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4101\,
            in2 => \N__3640\,
            in3 => \N__3705\,
            lcout => \eeprom.delay_counter_10\,
            ltout => OPEN,
            carryin => \eeprom.n2865\,
            carryout => \eeprom.n2866\,
            clk => \N__6746\,
            ce => \N__3830\,
            sr => \N__3806\
        );

    \eeprom.delay_counter_i0_i11_LC_21_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3701\,
            in2 => \N__3644\,
            in3 => \N__3687\,
            lcout => \eeprom.delay_counter_11\,
            ltout => OPEN,
            carryin => \eeprom.n2866\,
            carryout => \eeprom.n2867\,
            clk => \N__6746\,
            ce => \N__3830\,
            sr => \N__3806\
        );

    \eeprom.delay_counter_i0_i12_LC_21_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4113\,
            in2 => \N__3641\,
            in3 => \N__3684\,
            lcout => \eeprom.delay_counter_12\,
            ltout => OPEN,
            carryin => \eeprom.n2867\,
            carryout => \eeprom.n2868\,
            clk => \N__6746\,
            ce => \N__3830\,
            sr => \N__3806\
        );

    \eeprom.delay_counter_i0_i13_LC_21_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3680\,
            in2 => \N__3645\,
            in3 => \N__3666\,
            lcout => \eeprom.delay_counter_13\,
            ltout => OPEN,
            carryin => \eeprom.n2868\,
            carryout => \eeprom.n2869\,
            clk => \N__6746\,
            ce => \N__3830\,
            sr => \N__3806\
        );

    \eeprom.delay_counter_i0_i14_LC_21_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3662\,
            in2 => \N__3642\,
            in3 => \N__3648\,
            lcout => \eeprom.delay_counter_14\,
            ltout => OPEN,
            carryin => \eeprom.n2869\,
            carryout => \eeprom.n2870\,
            clk => \N__6746\,
            ce => \N__3830\,
            sr => \N__3806\
        );

    \eeprom.delay_counter_i0_i15_LC_21_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__3533\,
            in1 => \N__3629\,
            in2 => \_gnd_net_\,
            in3 => \N__3537\,
            lcout => \eeprom.delay_counter_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6746\,
            ce => \N__3830\,
            sr => \N__3806\
        );

    \i7_4_lut_LC_21_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101111"
        )
    port map (
            in0 => \N__4383\,
            in1 => \N__4344\,
            in2 => \N__5043\,
            in3 => \N__4338\,
            lcout => n15,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.mux_217_Mux_0_i1_4_lut_LC_21_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010001001110"
        )
    port map (
            in0 => \N__5151\,
            in1 => \N__4936\,
            in2 => \N__5017\,
            in3 => \N__4558\,
            lcout => OPEN,
            ltout => \n805_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rw_43_LC_21_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110010001100"
        )
    port map (
            in0 => \N__5209\,
            in1 => \N__4868\,
            in2 => \N__3837\,
            in3 => \N__5152\,
            lcout => rw,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6742\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i1_3_lut_LC_21_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100100010"
        )
    port map (
            in0 => \N__5149\,
            in1 => \N__5208\,
            in2 => \_gnd_net_\,
            in3 => \N__4935\,
            lcout => \eeprom.n1796\,
            ltout => \eeprom.n1796_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i1002_2_lut_LC_21_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__3810\,
            in3 => \N__5150\,
            lcout => \eeprom.n1929\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.enable_39_LC_21_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010001001110"
        )
    port map (
            in0 => \N__5153\,
            in1 => \N__4934\,
            in2 => \N__5022\,
            in3 => \N__4559\,
            lcout => \eeprom.enable\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6740\,
            ce => 'H',
            sr => \N__5214\
        );

    \eeprom.data_ready_42_LC_21_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101110100000"
        )
    port map (
            in0 => \N__3783\,
            in1 => \N__5021\,
            in2 => \N__5154\,
            in3 => \N__5210\,
            lcout => data_ready,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6737\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_LC_21_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4246\,
            in2 => \_gnd_net_\,
            in3 => \N__3782\,
            lcout => n6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \read_26_LC_21_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4218\,
            in2 => \_gnd_net_\,
            in3 => \N__4247\,
            lcout => read,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6737\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i526_4_lut_LC_21_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011001000"
        )
    port map (
            in0 => \N__3773\,
            in1 => \N__3761\,
            in2 => \N__3750\,
            in3 => \N__3735\,
            lcout => OPEN,
            ltout => \n36_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i8_4_lut_LC_21_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__4047\,
            in1 => \N__4031\,
            in2 => \N__4020\,
            in3 => \N__4017\,
            lcout => OPEN,
            ltout => \n22_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i11_3_lut_LC_21_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111010"
        )
    port map (
            in0 => \N__4002\,
            in1 => \_gnd_net_\,
            in2 => \N__3987\,
            in3 => \N__3983\,
            lcout => OPEN,
            ltout => \n25_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1422_4_lut_LC_21_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010100"
        )
    port map (
            in0 => \N__3972\,
            in1 => \N__4125\,
            in2 => \N__3954\,
            in3 => \N__3864\,
            lcout => n104,
            ltout => \n104_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i995_2_lut_LC_21_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__4298\,
            in1 => \_gnd_net_\,
            in2 => \N__3951\,
            in3 => \_gnd_net_\,
            lcout => n1891,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ID_READOUT_FSM_state__i0_LC_21_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000001011100"
        )
    port map (
            in0 => \N__3849\,
            in1 => \N__4185\,
            in2 => \N__4217\,
            in3 => \N__3858\,
            lcout => \ID_READOUT_FSM_state_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6743\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i9_4_lut_LC_21_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__3917\,
            in1 => \N__3905\,
            in2 => \N__3894\,
            in3 => \N__3875\,
            lcout => n23,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2007_2_lut_3_lut_LC_21_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010011001100"
        )
    port map (
            in0 => \N__4262\,
            in1 => \N__4240\,
            in2 => \_gnd_net_\,
            in3 => \N__4271\,
            lcout => n20,
            ltout => \n20_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i24_3_lut_LC_21_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4209\,
            in2 => \N__3852\,
            in3 => \N__3848\,
            lcout => OPEN,
            ltout => \n1836_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ID_READOUT_FSM_state__i1_LC_21_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010110000001100"
        )
    port map (
            in0 => \N__4213\,
            in1 => \N__4245\,
            in2 => \N__4323\,
            in3 => \N__4184\,
            lcout => \ID_READOUT_FSM_state_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6743\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i625_2_lut_3_lut_LC_21_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__4263\,
            in1 => \N__4207\,
            in2 => \_gnd_net_\,
            in3 => \N__4241\,
            lcout => n1507,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1484_2_lut_3_lut_4_lut_LC_21_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101111111"
        )
    port map (
            in0 => \N__4272\,
            in1 => \N__4261\,
            in2 => \N__4248\,
            in3 => \N__4208\,
            lcout => n2414,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i10_4_lut_LC_21_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__4175\,
            in1 => \N__4163\,
            in2 => \N__4152\,
            in3 => \N__4136\,
            lcout => n24,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.state_i0_i2_LC_22_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__5418\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4817\,
            lcout => \eeprom.i2c.state_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6427\,
            ce => \N__4752\,
            sr => \N__4395\
        );

    \eeprom.i2c.state_7__I_0_142_i10_2_lut_LC_22_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5959\,
            in2 => \_gnd_net_\,
            in3 => \N__5688\,
            lcout => \eeprom.i2c.n10_adj_381\,
            ltout => \eeprom.i2c.n10_adj_381_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.i2132_4_lut_LC_22_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110111001101"
        )
    port map (
            in0 => \N__4590\,
            in1 => \N__5422\,
            in2 => \N__4116\,
            in3 => \N__5513\,
            lcout => \eeprom.i2c.n3133\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i12_4_lut_LC_22_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__4112\,
            in1 => \N__4100\,
            in2 => \N__4089\,
            in3 => \N__4073\,
            lcout => \eeprom.n28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.i2178_2_lut_LC_22_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4613\,
            in2 => \_gnd_net_\,
            in3 => \N__4719\,
            lcout => \eeprom.i2c.n2388\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.state_7__I_0_139_i11_2_lut_4_lut_LC_22_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111011111"
        )
    port map (
            in0 => \N__6121\,
            in1 => \N__5960\,
            in2 => \N__5866\,
            in3 => \N__5689\,
            lcout => \eeprom.i2c.n11_adj_374\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.data_out_i0_i3_LC_22_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010111000"
        )
    port map (
            in0 => \N__4355\,
            in1 => \N__4773\,
            in2 => \N__5442\,
            in3 => \N__5341\,
            lcout => data_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6486\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.data_out_i0_i5_LC_22_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011011000"
        )
    port map (
            in0 => \N__5342\,
            in1 => \N__4382\,
            in2 => \N__5443\,
            in3 => \N__4674\,
            lcout => data_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6486\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.i2176_3_lut_4_lut_LC_22_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__5971\,
            in1 => \N__6116\,
            in2 => \N__4736\,
            in3 => \N__5723\,
            lcout => \eeprom.i2c.n3082\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.data_out_i0_i0_LC_22_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011011000"
        )
    port map (
            in0 => \N__4435\,
            in1 => \N__4370\,
            in2 => \N__5444\,
            in3 => \N__6144\,
            lcout => data_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6482\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i5_4_lut_adj_10_LC_22_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__4371\,
            in1 => \N__4446\,
            in2 => \N__4362\,
            in3 => \N__5310\,
            lcout => n13,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i4_2_lut_LC_22_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4425\,
            in2 => \_gnd_net_\,
            in3 => \N__4332\,
            lcout => n12,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.data_out_i0_i4_LC_22_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010111000"
        )
    port map (
            in0 => \N__4331\,
            in1 => \N__4670\,
            in2 => \N__5446\,
            in3 => \N__4436\,
            lcout => data_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6482\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.i1_2_lut_adj_7_LC_22_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__6669\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5072\,
            lcout => n1718,
            ltout => \n1718_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.data_out_i0_i2_LC_22_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001010"
        )
    port map (
            in0 => \N__5432\,
            in1 => \N__4445\,
            in2 => \N__4449\,
            in3 => \N__4766\,
            lcout => data_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6482\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.data_out_i0_i6_LC_22_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100011001100"
        )
    port map (
            in0 => \N__4437\,
            in1 => \N__4424\,
            in2 => \N__5445\,
            in3 => \N__4653\,
            lcout => data_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6482\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.enable_slow_120_LC_22_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000111111111"
        )
    port map (
            in0 => \N__5880\,
            in1 => \N__5523\,
            in2 => \N__6125\,
            in3 => \N__4843\,
            lcout => \state_7_N_270_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6744\,
            ce => \N__4572\,
            sr => \_gnd_net_\
        );

    \eeprom.i2c.write_enable_131_LC_23_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__4901\,
            in1 => \N__5859\,
            in2 => \_gnd_net_\,
            in3 => \N__5724\,
            lcout => sda_enable,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVeeprom.i2c.write_enable_131C_net\,
            ce => \N__4404\,
            sr => \N__4416\
        );

    \eeprom.i2c.i1_3_lut_adj_4_LC_23_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100100010"
        )
    port map (
            in0 => \N__6248\,
            in1 => \N__6095\,
            in2 => \_gnd_net_\,
            in3 => \N__4509\,
            lcout => \eeprom.i2c.n1928\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.i2129_2_lut_LC_23_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4789\,
            in2 => \_gnd_net_\,
            in3 => \N__6186\,
            lcout => OPEN,
            ltout => \eeprom.i2c.n3130_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.i2128_4_lut_LC_23_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100000000000"
        )
    port map (
            in0 => \N__6228\,
            in1 => \N__6665\,
            in2 => \N__4407\,
            in3 => \N__6097\,
            lcout => \eeprom.i2c.n3123\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.i2152_4_lut_4_lut_LC_23_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011000100"
        )
    port map (
            in0 => \N__6096\,
            in1 => \N__4497\,
            in2 => \N__4900\,
            in3 => \N__5690\,
            lcout => \eeprom.i2c.n1153\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.state_i0_i0_LC_23_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0011001100110111"
        )
    port map (
            in0 => \N__5801\,
            in1 => \N__4806\,
            in2 => \N__4641\,
            in3 => \N__6058\,
            lcout => \eeprom.state_0_adj_384\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6432\,
            ce => \N__4750\,
            sr => \N__4599\
        );

    \eeprom.i2c.i56_3_lut_3_lut_LC_23_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010001100110"
        )
    port map (
            in0 => \N__5948\,
            in1 => \N__5797\,
            in2 => \_gnd_net_\,
            in3 => \N__5663\,
            lcout => \eeprom.i2c.n33\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.i1_4_lut_4_lut_LC_23_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001100010010"
        )
    port map (
            in0 => \N__5664\,
            in1 => \N__5949\,
            in2 => \N__5845\,
            in3 => \N__6055\,
            lcout => \eeprom.i2c.n37\,
            ltout => \eeprom.i2c.n37_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.i1_3_lut_LC_23_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010111110000"
        )
    port map (
            in0 => \N__6056\,
            in1 => \_gnd_net_\,
            in2 => \N__4512\,
            in3 => \N__4508\,
            lcout => \eeprom.i2c.n39\,
            ltout => \eeprom.i2c.n39_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.i2148_4_lut_LC_23_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000011110000"
        )
    port map (
            in0 => \N__5665\,
            in1 => \N__4458\,
            in2 => \N__4491\,
            in3 => \N__6057\,
            lcout => \eeprom.i2c.n2967\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.state_i0_i3_LC_23_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1101100000000000"
        )
    port map (
            in0 => \N__5804\,
            in1 => \N__4488\,
            in2 => \N__4482\,
            in3 => \N__6094\,
            lcout => \eeprom.state_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6458\,
            ce => \N__4749\,
            sr => \N__4467\
        );

    \eeprom.i2c.i1_3_lut_3_lut_LC_23_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5803\,
            in2 => \_gnd_net_\,
            in3 => \N__5951\,
            lcout => \eeprom.i2c.n13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.state_7__I_0_143_i11_2_lut_3_lut_4_lut_LC_23_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110111111111"
        )
    port map (
            in0 => \N__5703\,
            in1 => \N__5851\,
            in2 => \N__5975\,
            in3 => \N__6076\,
            lcout => \eeprom.i2c.n15\,
            ltout => \eeprom.i2c.n15_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.i1433_4_lut_LC_23_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010110000"
        )
    port map (
            in0 => \N__5468\,
            in1 => \N__5958\,
            in2 => \N__4452\,
            in3 => \N__5705\,
            lcout => \eeprom.i2c.n2358\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.i1427_2_lut_LC_23_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5847\,
            in2 => \_gnd_net_\,
            in3 => \N__6074\,
            lcout => \eeprom.i2c.n2352\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.state_7__I_0_138_i11_2_lut_3_lut_4_lut_LC_23_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111101"
        )
    port map (
            in0 => \N__6075\,
            in1 => \N__5953\,
            in2 => \N__5874\,
            in3 => \N__5702\,
            lcout => \eeprom.i2c.n11_adj_378\,
            ltout => \eeprom.i2c.n11_adj_378_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.i1_4_lut_LC_23_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110001001100"
        )
    port map (
            in0 => \N__4637\,
            in1 => \N__6279\,
            in2 => \N__4626\,
            in3 => \N__5852\,
            lcout => OPEN,
            ltout => \eeprom.i2c.n1734_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.i2162_4_lut_LC_23_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001100000111"
        )
    port map (
            in0 => \N__4623\,
            in1 => \N__5957\,
            in2 => \N__4617\,
            in3 => \N__5704\,
            lcout => \eeprom.i2c.n1063\,
            ltout => \eeprom.i2c.n1063_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.i996_4_lut_LC_23_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000010110000"
        )
    port map (
            in0 => \N__4850\,
            in1 => \N__4614\,
            in2 => \N__4602\,
            in3 => \N__4991\,
            lcout => \eeprom.i2c.n1923\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.equal_40_i10_2_lut_LC_23_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5952\,
            in2 => \_gnd_net_\,
            in3 => \N__5701\,
            lcout => \eeprom.n10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.i1_2_lut_3_lut_4_lut_LC_23_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001000"
        )
    port map (
            in0 => \N__5234\,
            in1 => \N__4842\,
            in2 => \N__5531\,
            in3 => \N__4589\,
            lcout => \eeprom.i2c.n1761\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.i1_2_lut_adj_3_LC_23_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6106\,
            in2 => \_gnd_net_\,
            in3 => \N__5709\,
            lcout => OPEN,
            ltout => \eeprom.n26_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i3_4_lut_LC_23_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__4560\,
            in1 => \N__5867\,
            in2 => \N__4533\,
            in3 => \N__5987\,
            lcout => n2913,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.sda_out_132_LC_24_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000111010"
        )
    port map (
            in0 => \N__4530\,
            in1 => \N__5835\,
            in2 => \N__4902\,
            in3 => \N__5725\,
            lcout => \eeprom.i2c.sda_out_adj_375\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVeeprom.i2c.sda_out_132C_net\,
            ce => \N__4524\,
            sr => \_gnd_net_\
        );

    \eeprom.i2c.i22_3_lut_3_lut_LC_24_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000110101010"
        )
    port map (
            in0 => \N__5802\,
            in1 => \N__6059\,
            in2 => \_gnd_net_\,
            in3 => \N__5950\,
            lcout => \eeprom.i2c.n11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.saved_addr__i1_LC_24_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111100100000"
        )
    port map (
            in0 => \N__4875\,
            in1 => \N__5006\,
            in2 => \N__4857\,
            in3 => \N__4790\,
            lcout => saved_addr_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6431\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.state_i0_i1_LC_24_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0011011100110011"
        )
    port map (
            in0 => \N__4821\,
            in1 => \N__4805\,
            in2 => \N__5453\,
            in3 => \N__4791\,
            lcout => \eeprom.state_1_adj_386\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6476\,
            ce => \N__4751\,
            sr => \N__4686\
        );

    \eeprom.i2c.equal_58_i4_2_lut_LC_24_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__6236\,
            in3 => \N__6187\,
            lcout => n4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.equal_42_i9_2_lut_LC_24_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6070\,
            in2 => \_gnd_net_\,
            in3 => \N__5846\,
            lcout => \eeprom.i2c.n9_adj_377\,
            ltout => \eeprom.i2c.n9_adj_377_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.i2181_4_lut_LC_24_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000001100"
        )
    port map (
            in0 => \N__5967\,
            in1 => \N__4720\,
            in2 => \N__4689\,
            in3 => \N__5730\,
            lcout => \eeprom.i2c.n3050\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.equal_56_i4_2_lut_LC_24_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110111011"
        )
    port map (
            in0 => \N__6189\,
            in1 => \N__6229\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => n4_adj_389,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.i1419_2_lut_LC_24_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__6237\,
            in3 => \N__6188\,
            lcout => n2344,
            ltout => \n2344_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.data_out_i0_i7_LC_24_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101100"
        )
    port map (
            in0 => \N__5454\,
            in1 => \N__5033\,
            in2 => \N__4644\,
            in3 => \N__5343\,
            lcout => data_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6475\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.equal_40_i11_2_lut_4_lut_LC_24_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__5966\,
            in1 => \N__5858\,
            in2 => \N__6101\,
            in3 => \N__5729\,
            lcout => \enable_slow_N_373\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i1492_2_lut_3_lut_4_lut_LC_24_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111011"
        )
    port map (
            in0 => \N__5123\,
            in1 => \N__5187\,
            in2 => \N__5532\,
            in3 => \N__5232\,
            lcout => n2382,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.i1400_2_lut_LC_24_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__6105\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5882\,
            lcout => \eeprom.n9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i28_3_lut_LC_24_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010011101110"
        )
    port map (
            in0 => \N__5121\,
            in1 => \N__4943\,
            in2 => \_gnd_net_\,
            in3 => \N__4957\,
            lcout => OPEN,
            ltout => \eeprom.n14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2126_4_lut_LC_24_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000001110010"
        )
    port map (
            in0 => \N__5189\,
            in1 => \N__5007\,
            in2 => \N__4971\,
            in3 => \N__5125\,
            lcout => \eeprom.n3142\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2_3_lut_4_lut_LC_24_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__5126\,
            in1 => \N__5188\,
            in2 => \_gnd_net_\,
            in3 => \N__4959\,
            lcout => OPEN,
            ltout => \n3051_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.state__i1_LC_24_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100100011000000"
        )
    port map (
            in0 => \N__5190\,
            in1 => \N__4968\,
            in2 => \N__4962\,
            in3 => \N__4908\,
            lcout => state_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6748\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i546_3_lut_3_lut_4_lut_LC_24_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011001000"
        )
    port map (
            in0 => \N__5122\,
            in1 => \N__5186\,
            in2 => \N__5533\,
            in3 => \N__5233\,
            lcout => OPEN,
            ltout => \n1113_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2_4_lut_LC_24_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100011111111"
        )
    port map (
            in0 => \N__4958\,
            in1 => \N__5124\,
            in2 => \N__4947\,
            in3 => \N__4944\,
            lcout => n3109,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.state__i0_LC_24_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001000110011"
        )
    port map (
            in0 => \N__5235\,
            in1 => \N__5133\,
            in2 => \N__5540\,
            in3 => \N__5191\,
            lcout => state_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6745\,
            ce => \N__5082\,
            sr => \_gnd_net_\
        );

    \eeprom.i2c.i2c_clk_121_LC_26_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6367\,
            in2 => \_gnd_net_\,
            in3 => \N__6680\,
            lcout => \eeprom.i2c.i2c_clk\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6749\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.i4_4_lut_LC_26_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__5579\,
            in1 => \N__6761\,
            in2 => \N__6783\,
            in3 => \N__5564\,
            lcout => OPEN,
            ltout => \eeprom.i2c.n10_adj_380_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.i5_3_lut_LC_26_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5595\,
            in2 => \N__5076\,
            in3 => \N__5610\,
            lcout => \eeprom.i2c.n1930\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.i1_2_lut_adj_8_LC_26_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6657\,
            in2 => \_gnd_net_\,
            in3 => \N__5073\,
            lcout => n1723,
            ltout => OPEN,
            carryin => \bfn_26_14_0_\,
            carryout => \eeprom.i2c.n2849\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.counter_i1_LC_26_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1001",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6567\,
            in2 => \N__6178\,
            in3 => \N__5055\,
            lcout => \eeprom.i2c.counter_1\,
            ltout => OPEN,
            carryin => \eeprom.i2c.n2849\,
            carryout => \eeprom.i2c.n2850\,
            clk => \N__6368\,
            ce => \N__6629\,
            sr => \N__6599\
        );

    \eeprom.i2c.counter_i2_LC_26_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1001",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6214\,
            in2 => \N__6580\,
            in3 => \N__5052\,
            lcout => \eeprom.i2c.counter_2\,
            ltout => OPEN,
            carryin => \eeprom.i2c.n2850\,
            carryout => \eeprom.i2c.n2851\,
            clk => \N__6368\,
            ce => \N__6629\,
            sr => \N__6599\
        );

    \eeprom.i2c.counter_i3_LC_26_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6571\,
            in2 => \N__5280\,
            in3 => \N__5049\,
            lcout => \eeprom.i2c.counter_3\,
            ltout => OPEN,
            carryin => \eeprom.i2c.n2851\,
            carryout => \eeprom.i2c.n2852\,
            clk => \N__6368\,
            ce => \N__6629\,
            sr => \N__6599\
        );

    \eeprom.i2c.counter_i4_LC_26_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6294\,
            in2 => \N__6581\,
            in3 => \N__5046\,
            lcout => \eeprom.i2c.counter_4\,
            ltout => OPEN,
            carryin => \eeprom.i2c.n2852\,
            carryout => \eeprom.i2c.n2853\,
            clk => \N__6368\,
            ce => \N__6629\,
            sr => \N__6599\
        );

    \eeprom.i2c.counter_i5_LC_26_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6575\,
            in2 => \N__5265\,
            in3 => \N__5550\,
            lcout => \eeprom.i2c.counter_5\,
            ltout => OPEN,
            carryin => \eeprom.i2c.n2853\,
            carryout => \eeprom.i2c.n2854\,
            clk => \N__6368\,
            ce => \N__6629\,
            sr => \N__6599\
        );

    \eeprom.i2c.counter_i6_LC_26_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5292\,
            in2 => \N__6582\,
            in3 => \N__5547\,
            lcout => \eeprom.i2c.counter_6\,
            ltout => OPEN,
            carryin => \eeprom.i2c.n2854\,
            carryout => \eeprom.i2c.n2855\,
            clk => \N__6368\,
            ce => \N__6629\,
            sr => \N__6599\
        );

    \eeprom.i2c.counter_i7_LC_26_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__5247\,
            in1 => \N__6579\,
            in2 => \_gnd_net_\,
            in3 => \N__5544\,
            lcout => \eeprom.i2c.counter_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6368\,
            ce => \N__6629\,
            sr => \N__6599\
        );

    \eeprom.i2c.i2024_2_lut_3_lut_LC_26_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010001000"
        )
    port map (
            in0 => \N__5411\,
            in1 => \N__5530\,
            in2 => \_gnd_net_\,
            in3 => \N__5472\,
            lcout => \eeprom.i2c.n3039\,
            ltout => \eeprom.i2c.n3039_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.i2008_2_lut_4_lut_LC_26_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__5876\,
            in1 => \N__5989\,
            in2 => \N__5457\,
            in3 => \N__5727\,
            lcout => \eeprom.i2c.n1924\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.data_out_i0_i1_LC_26_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000000100"
        )
    port map (
            in0 => \N__6140\,
            in1 => \N__5410\,
            in2 => \N__5337\,
            in3 => \N__5303\,
            lcout => data_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6446\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.i1_2_lut_3_lut_LC_26_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__5875\,
            in1 => \N__5988\,
            in2 => \_gnd_net_\,
            in3 => \N__5726\,
            lcout => \eeprom.i2c.n1172\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.i5_4_lut_LC_26_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__5291\,
            in1 => \N__5276\,
            in2 => \N__5264\,
            in3 => \N__6651\,
            lcout => OPEN,
            ltout => \eeprom.i2c.n12_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.i6_4_lut_LC_26_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__5246\,
            in1 => \N__6293\,
            in2 => \N__6282\,
            in3 => \N__6139\,
            lcout => \eeprom.i2c.n1056\,
            ltout => \eeprom.i2c.n1056_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.i17_4_lut_LC_26_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111001000100010"
        )
    port map (
            in0 => \N__6270\,
            in1 => \N__6264\,
            in2 => \N__6258\,
            in3 => \N__6255\,
            lcout => \eeprom.i2c.n1757\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.equal_59_i4_2_lut_LC_26_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6210\,
            in2 => \_gnd_net_\,
            in3 => \N__6165\,
            lcout => n4_adj_390,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.i2c_scl_enable_123_LC_26_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111101010"
        )
    port map (
            in0 => \N__6117\,
            in1 => \N__5994\,
            in2 => \N__5883\,
            in3 => \N__5728\,
            lcout => scl_enable,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVeeprom.i2c.i2c_scl_enable_123C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.counter2_411_412__i1_LC_27_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5609\,
            in2 => \_gnd_net_\,
            in3 => \N__5598\,
            lcout => \eeprom.i2c.counter2_0\,
            ltout => OPEN,
            carryin => \bfn_27_13_0_\,
            carryout => \eeprom.i2c.n2871\,
            clk => \N__6750\,
            ce => 'H',
            sr => \N__6687\
        );

    \eeprom.i2c.counter2_411_412__i2_LC_27_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5594\,
            in2 => \_gnd_net_\,
            in3 => \N__5583\,
            lcout => \eeprom.i2c.counter2_1\,
            ltout => OPEN,
            carryin => \eeprom.i2c.n2871\,
            carryout => \eeprom.i2c.n2872\,
            clk => \N__6750\,
            ce => 'H',
            sr => \N__6687\
        );

    \eeprom.i2c.counter2_411_412__i3_LC_27_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5580\,
            in2 => \_gnd_net_\,
            in3 => \N__5568\,
            lcout => \eeprom.i2c.counter2_2\,
            ltout => OPEN,
            carryin => \eeprom.i2c.n2872\,
            carryout => \eeprom.i2c.n2873\,
            clk => \N__6750\,
            ce => 'H',
            sr => \N__6687\
        );

    \eeprom.i2c.counter2_411_412__i4_LC_27_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5565\,
            in2 => \_gnd_net_\,
            in3 => \N__5553\,
            lcout => \eeprom.i2c.counter2_3\,
            ltout => OPEN,
            carryin => \eeprom.i2c.n2873\,
            carryout => \eeprom.i2c.n2874\,
            clk => \N__6750\,
            ce => 'H',
            sr => \N__6687\
        );

    \eeprom.i2c.counter2_411_412__i5_LC_27_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6782\,
            in2 => \_gnd_net_\,
            in3 => \N__6768\,
            lcout => \eeprom.i2c.counter2_4\,
            ltout => OPEN,
            carryin => \eeprom.i2c.n2874\,
            carryout => \eeprom.i2c.n2875\,
            clk => \N__6750\,
            ce => 'H',
            sr => \N__6687\
        );

    \eeprom.i2c.counter2_411_412__i6_LC_27_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6762\,
            in2 => \_gnd_net_\,
            in3 => \N__6765\,
            lcout => \eeprom.i2c.counter2_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6750\,
            ce => 'H',
            sr => \N__6687\
        );

    \eeprom.i2c.counter_i0_LC_27_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__6566\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6658\,
            lcout => \eeprom.i2c.counter_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6391\,
            ce => \N__6630\,
            sr => \N__6606\
        );

    \CONSTANT_ONE_LUT4_LC_27_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.i471_2_lut_LC_30_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6543\,
            in2 => \_gnd_net_\,
            in3 => \N__6518\,
            lcout => sda_out,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.i1404_2_lut_LC_32_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6477\,
            in2 => \_gnd_net_\,
            in3 => \N__6326\,
            lcout => scl_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;
