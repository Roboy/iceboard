// ******************************************************************************

// iCEcube Netlister

// Version:            2017.08.27940

// Build Date:         Sep 12 2017 08:25:46

// File Generated:     Jan 29 2020 12:28:03

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "TinyFPGA_B" view "INTERFACE"

module TinyFPGA_B (
    USBPU,
    TX,
    SDA,
    SCL,
    RX,
    NEOPXL,
    LED,
    INLC,
    INLB,
    INLA,
    INHC,
    INHB,
    INHA,
    HALL3,
    HALL2,
    HALL1,
    FAULT_N,
    ENCODER1_B,
    ENCODER1_A,
    ENCODER0_B,
    ENCODER0_A,
    DE,
    CS_MISO,
    CS_CLK,
    CS,
    CLK);

    output USBPU;
    output TX;
    inout SDA;
    inout SCL;
    input RX;
    output NEOPXL;
    output LED;
    output INLC;
    output INLB;
    output INLA;
    output INHC;
    output INHB;
    output INHA;
    input HALL3;
    input HALL2;
    input HALL1;
    input FAULT_N;
    input ENCODER1_B;
    input ENCODER1_A;
    input ENCODER0_B;
    input ENCODER0_A;
    output DE;
    input CS_MISO;
    output CS_CLK;
    output CS;
    input CLK;

    wire N__28245;
    wire N__28244;
    wire N__28243;
    wire N__28236;
    wire N__28235;
    wire N__28234;
    wire N__28227;
    wire N__28226;
    wire N__28225;
    wire N__28218;
    wire N__28217;
    wire N__28216;
    wire N__28209;
    wire N__28208;
    wire N__28207;
    wire N__28200;
    wire N__28199;
    wire N__28198;
    wire N__28191;
    wire N__28190;
    wire N__28189;
    wire N__28182;
    wire N__28181;
    wire N__28180;
    wire N__28173;
    wire N__28172;
    wire N__28171;
    wire N__28164;
    wire N__28163;
    wire N__28162;
    wire N__28155;
    wire N__28154;
    wire N__28153;
    wire N__28146;
    wire N__28145;
    wire N__28144;
    wire N__28137;
    wire N__28136;
    wire N__28135;
    wire N__28128;
    wire N__28127;
    wire N__28126;
    wire N__28119;
    wire N__28118;
    wire N__28117;
    wire N__28110;
    wire N__28109;
    wire N__28108;
    wire N__28091;
    wire N__28088;
    wire N__28085;
    wire N__28082;
    wire N__28079;
    wire N__28076;
    wire N__28073;
    wire N__28072;
    wire N__28069;
    wire N__28066;
    wire N__28063;
    wire N__28062;
    wire N__28057;
    wire N__28054;
    wire N__28049;
    wire N__28046;
    wire N__28043;
    wire N__28040;
    wire N__28037;
    wire N__28034;
    wire N__28031;
    wire N__28030;
    wire N__28027;
    wire N__28026;
    wire N__28023;
    wire N__28020;
    wire N__28015;
    wire N__28010;
    wire N__28007;
    wire N__28004;
    wire N__28001;
    wire N__27998;
    wire N__27995;
    wire N__27994;
    wire N__27991;
    wire N__27988;
    wire N__27987;
    wire N__27984;
    wire N__27981;
    wire N__27978;
    wire N__27975;
    wire N__27970;
    wire N__27965;
    wire N__27962;
    wire N__27959;
    wire N__27956;
    wire N__27953;
    wire N__27950;
    wire N__27947;
    wire N__27944;
    wire N__27943;
    wire N__27940;
    wire N__27937;
    wire N__27934;
    wire N__27931;
    wire N__27928;
    wire N__27925;
    wire N__27920;
    wire N__27919;
    wire N__27916;
    wire N__27915;
    wire N__27912;
    wire N__27911;
    wire N__27910;
    wire N__27909;
    wire N__27908;
    wire N__27907;
    wire N__27904;
    wire N__27903;
    wire N__27902;
    wire N__27899;
    wire N__27894;
    wire N__27891;
    wire N__27890;
    wire N__27889;
    wire N__27888;
    wire N__27887;
    wire N__27886;
    wire N__27883;
    wire N__27882;
    wire N__27881;
    wire N__27878;
    wire N__27875;
    wire N__27874;
    wire N__27871;
    wire N__27864;
    wire N__27861;
    wire N__27856;
    wire N__27851;
    wire N__27848;
    wire N__27839;
    wire N__27832;
    wire N__27829;
    wire N__27824;
    wire N__27809;
    wire N__27806;
    wire N__27805;
    wire N__27802;
    wire N__27799;
    wire N__27794;
    wire N__27791;
    wire N__27788;
    wire N__27787;
    wire N__27786;
    wire N__27785;
    wire N__27784;
    wire N__27783;
    wire N__27782;
    wire N__27781;
    wire N__27780;
    wire N__27779;
    wire N__27778;
    wire N__27777;
    wire N__27776;
    wire N__27775;
    wire N__27774;
    wire N__27773;
    wire N__27770;
    wire N__27769;
    wire N__27768;
    wire N__27767;
    wire N__27766;
    wire N__27765;
    wire N__27762;
    wire N__27761;
    wire N__27760;
    wire N__27757;
    wire N__27756;
    wire N__27755;
    wire N__27754;
    wire N__27753;
    wire N__27752;
    wire N__27751;
    wire N__27750;
    wire N__27749;
    wire N__27748;
    wire N__27747;
    wire N__27746;
    wire N__27745;
    wire N__27744;
    wire N__27743;
    wire N__27742;
    wire N__27739;
    wire N__27736;
    wire N__27733;
    wire N__27732;
    wire N__27731;
    wire N__27730;
    wire N__27729;
    wire N__27728;
    wire N__27727;
    wire N__27726;
    wire N__27725;
    wire N__27724;
    wire N__27723;
    wire N__27722;
    wire N__27721;
    wire N__27716;
    wire N__27715;
    wire N__27714;
    wire N__27713;
    wire N__27712;
    wire N__27711;
    wire N__27710;
    wire N__27709;
    wire N__27708;
    wire N__27707;
    wire N__27706;
    wire N__27701;
    wire N__27694;
    wire N__27683;
    wire N__27680;
    wire N__27677;
    wire N__27674;
    wire N__27671;
    wire N__27670;
    wire N__27659;
    wire N__27654;
    wire N__27653;
    wire N__27650;
    wire N__27649;
    wire N__27648;
    wire N__27647;
    wire N__27644;
    wire N__27643;
    wire N__27642;
    wire N__27641;
    wire N__27638;
    wire N__27635;
    wire N__27630;
    wire N__27629;
    wire N__27628;
    wire N__27627;
    wire N__27624;
    wire N__27621;
    wire N__27620;
    wire N__27617;
    wire N__27614;
    wire N__27613;
    wire N__27612;
    wire N__27611;
    wire N__27608;
    wire N__27607;
    wire N__27606;
    wire N__27605;
    wire N__27604;
    wire N__27599;
    wire N__27596;
    wire N__27591;
    wire N__27590;
    wire N__27589;
    wire N__27588;
    wire N__27587;
    wire N__27586;
    wire N__27583;
    wire N__27582;
    wire N__27581;
    wire N__27578;
    wire N__27575;
    wire N__27570;
    wire N__27569;
    wire N__27566;
    wire N__27565;
    wire N__27564;
    wire N__27561;
    wire N__27560;
    wire N__27557;
    wire N__27556;
    wire N__27553;
    wire N__27550;
    wire N__27547;
    wire N__27546;
    wire N__27545;
    wire N__27544;
    wire N__27543;
    wire N__27542;
    wire N__27541;
    wire N__27538;
    wire N__27529;
    wire N__27520;
    wire N__27519;
    wire N__27518;
    wire N__27515;
    wire N__27514;
    wire N__27513;
    wire N__27510;
    wire N__27509;
    wire N__27504;
    wire N__27501;
    wire N__27490;
    wire N__27485;
    wire N__27476;
    wire N__27467;
    wire N__27460;
    wire N__27459;
    wire N__27456;
    wire N__27453;
    wire N__27448;
    wire N__27443;
    wire N__27436;
    wire N__27431;
    wire N__27428;
    wire N__27423;
    wire N__27422;
    wire N__27421;
    wire N__27418;
    wire N__27415;
    wire N__27412;
    wire N__27411;
    wire N__27410;
    wire N__27407;
    wire N__27402;
    wire N__27397;
    wire N__27394;
    wire N__27393;
    wire N__27390;
    wire N__27387;
    wire N__27386;
    wire N__27385;
    wire N__27384;
    wire N__27383;
    wire N__27382;
    wire N__27381;
    wire N__27378;
    wire N__27375;
    wire N__27372;
    wire N__27371;
    wire N__27368;
    wire N__27365;
    wire N__27362;
    wire N__27357;
    wire N__27348;
    wire N__27345;
    wire N__27342;
    wire N__27335;
    wire N__27334;
    wire N__27333;
    wire N__27332;
    wire N__27331;
    wire N__27330;
    wire N__27327;
    wire N__27326;
    wire N__27325;
    wire N__27322;
    wire N__27319;
    wire N__27318;
    wire N__27315;
    wire N__27312;
    wire N__27311;
    wire N__27310;
    wire N__27307;
    wire N__27306;
    wire N__27305;
    wire N__27304;
    wire N__27303;
    wire N__27302;
    wire N__27295;
    wire N__27290;
    wire N__27279;
    wire N__27272;
    wire N__27263;
    wire N__27260;
    wire N__27255;
    wire N__27252;
    wire N__27247;
    wire N__27240;
    wire N__27235;
    wire N__27226;
    wire N__27223;
    wire N__27218;
    wire N__27215;
    wire N__27206;
    wire N__27205;
    wire N__27202;
    wire N__27199;
    wire N__27196;
    wire N__27195;
    wire N__27194;
    wire N__27193;
    wire N__27192;
    wire N__27191;
    wire N__27190;
    wire N__27189;
    wire N__27188;
    wire N__27187;
    wire N__27186;
    wire N__27185;
    wire N__27182;
    wire N__27181;
    wire N__27180;
    wire N__27179;
    wire N__27176;
    wire N__27175;
    wire N__27174;
    wire N__27171;
    wire N__27166;
    wire N__27163;
    wire N__27160;
    wire N__27155;
    wire N__27142;
    wire N__27139;
    wire N__27136;
    wire N__27133;
    wire N__27130;
    wire N__27127;
    wire N__27126;
    wire N__27123;
    wire N__27118;
    wire N__27109;
    wire N__27106;
    wire N__27103;
    wire N__27098;
    wire N__27095;
    wire N__27092;
    wire N__27091;
    wire N__27088;
    wire N__27085;
    wire N__27084;
    wire N__27081;
    wire N__27080;
    wire N__27079;
    wire N__27078;
    wire N__27077;
    wire N__27076;
    wire N__27075;
    wire N__27074;
    wire N__27073;
    wire N__27066;
    wire N__27059;
    wire N__27048;
    wire N__27043;
    wire N__27036;
    wire N__27031;
    wire N__27026;
    wire N__27025;
    wire N__27024;
    wire N__27021;
    wire N__27018;
    wire N__27017;
    wire N__27016;
    wire N__27013;
    wire N__27010;
    wire N__27009;
    wire N__27008;
    wire N__27005;
    wire N__27002;
    wire N__26999;
    wire N__26998;
    wire N__26995;
    wire N__26992;
    wire N__26989;
    wire N__26988;
    wire N__26987;
    wire N__26984;
    wire N__26981;
    wire N__26978;
    wire N__26973;
    wire N__26964;
    wire N__26957;
    wire N__26952;
    wire N__26947;
    wire N__26938;
    wire N__26937;
    wire N__26936;
    wire N__26933;
    wire N__26922;
    wire N__26919;
    wire N__26904;
    wire N__26901;
    wire N__26898;
    wire N__26895;
    wire N__26892;
    wire N__26889;
    wire N__26886;
    wire N__26885;
    wire N__26882;
    wire N__26881;
    wire N__26880;
    wire N__26877;
    wire N__26870;
    wire N__26863;
    wire N__26858;
    wire N__26849;
    wire N__26840;
    wire N__26833;
    wire N__26822;
    wire N__26817;
    wire N__26800;
    wire N__26795;
    wire N__26786;
    wire N__26779;
    wire N__26768;
    wire N__26765;
    wire N__26764;
    wire N__26761;
    wire N__26756;
    wire N__26753;
    wire N__26740;
    wire N__26735;
    wire N__26728;
    wire N__26725;
    wire N__26720;
    wire N__26705;
    wire N__26704;
    wire N__26703;
    wire N__26700;
    wire N__26697;
    wire N__26694;
    wire N__26691;
    wire N__26684;
    wire N__26681;
    wire N__26678;
    wire N__26675;
    wire N__26672;
    wire N__26671;
    wire N__26668;
    wire N__26667;
    wire N__26664;
    wire N__26661;
    wire N__26658;
    wire N__26651;
    wire N__26648;
    wire N__26645;
    wire N__26642;
    wire N__26639;
    wire N__26636;
    wire N__26635;
    wire N__26634;
    wire N__26631;
    wire N__26628;
    wire N__26625;
    wire N__26620;
    wire N__26617;
    wire N__26614;
    wire N__26611;
    wire N__26606;
    wire N__26603;
    wire N__26600;
    wire N__26597;
    wire N__26594;
    wire N__26593;
    wire N__26590;
    wire N__26587;
    wire N__26586;
    wire N__26583;
    wire N__26580;
    wire N__26577;
    wire N__26574;
    wire N__26571;
    wire N__26568;
    wire N__26561;
    wire N__26558;
    wire N__26555;
    wire N__26552;
    wire N__26549;
    wire N__26546;
    wire N__26543;
    wire N__26540;
    wire N__26539;
    wire N__26538;
    wire N__26535;
    wire N__26532;
    wire N__26529;
    wire N__26522;
    wire N__26519;
    wire N__26516;
    wire N__26513;
    wire N__26512;
    wire N__26511;
    wire N__26508;
    wire N__26505;
    wire N__26502;
    wire N__26499;
    wire N__26496;
    wire N__26493;
    wire N__26490;
    wire N__26483;
    wire N__26480;
    wire N__26477;
    wire N__26474;
    wire N__26471;
    wire N__26468;
    wire N__26467;
    wire N__26464;
    wire N__26461;
    wire N__26460;
    wire N__26457;
    wire N__26454;
    wire N__26451;
    wire N__26444;
    wire N__26441;
    wire N__26438;
    wire N__26435;
    wire N__26432;
    wire N__26429;
    wire N__26426;
    wire N__26423;
    wire N__26420;
    wire N__26419;
    wire N__26418;
    wire N__26415;
    wire N__26410;
    wire N__26407;
    wire N__26404;
    wire N__26399;
    wire N__26396;
    wire N__26393;
    wire N__26390;
    wire N__26387;
    wire N__26386;
    wire N__26385;
    wire N__26382;
    wire N__26379;
    wire N__26376;
    wire N__26369;
    wire N__26366;
    wire N__26363;
    wire N__26360;
    wire N__26357;
    wire N__26354;
    wire N__26351;
    wire N__26348;
    wire N__26345;
    wire N__26342;
    wire N__26339;
    wire N__26336;
    wire N__26335;
    wire N__26332;
    wire N__26331;
    wire N__26328;
    wire N__26325;
    wire N__26322;
    wire N__26319;
    wire N__26312;
    wire N__26309;
    wire N__26306;
    wire N__26303;
    wire N__26300;
    wire N__26297;
    wire N__26294;
    wire N__26293;
    wire N__26290;
    wire N__26287;
    wire N__26284;
    wire N__26283;
    wire N__26278;
    wire N__26275;
    wire N__26272;
    wire N__26267;
    wire N__26264;
    wire N__26261;
    wire N__26258;
    wire N__26255;
    wire N__26252;
    wire N__26249;
    wire N__26246;
    wire N__26245;
    wire N__26244;
    wire N__26241;
    wire N__26238;
    wire N__26235;
    wire N__26232;
    wire N__26229;
    wire N__26224;
    wire N__26221;
    wire N__26218;
    wire N__26213;
    wire N__26210;
    wire N__26207;
    wire N__26204;
    wire N__26201;
    wire N__26198;
    wire N__26195;
    wire N__26192;
    wire N__26191;
    wire N__26188;
    wire N__26185;
    wire N__26184;
    wire N__26181;
    wire N__26178;
    wire N__26175;
    wire N__26172;
    wire N__26165;
    wire N__26162;
    wire N__26159;
    wire N__26156;
    wire N__26153;
    wire N__26150;
    wire N__26147;
    wire N__26146;
    wire N__26145;
    wire N__26142;
    wire N__26139;
    wire N__26136;
    wire N__26133;
    wire N__26130;
    wire N__26125;
    wire N__26120;
    wire N__26117;
    wire N__26114;
    wire N__26111;
    wire N__26108;
    wire N__26105;
    wire N__26102;
    wire N__26099;
    wire N__26096;
    wire N__26093;
    wire N__26092;
    wire N__26089;
    wire N__26088;
    wire N__26085;
    wire N__26082;
    wire N__26077;
    wire N__26074;
    wire N__26069;
    wire N__26066;
    wire N__26063;
    wire N__26060;
    wire N__26057;
    wire N__26056;
    wire N__26055;
    wire N__26052;
    wire N__26049;
    wire N__26046;
    wire N__26043;
    wire N__26040;
    wire N__26033;
    wire N__26030;
    wire N__26027;
    wire N__26024;
    wire N__26021;
    wire N__26018;
    wire N__26015;
    wire N__26014;
    wire N__26011;
    wire N__26008;
    wire N__26003;
    wire N__26000;
    wire N__25997;
    wire N__25994;
    wire N__25993;
    wire N__25990;
    wire N__25987;
    wire N__25984;
    wire N__25981;
    wire N__25980;
    wire N__25975;
    wire N__25972;
    wire N__25967;
    wire N__25964;
    wire N__25961;
    wire N__25958;
    wire N__25955;
    wire N__25952;
    wire N__25949;
    wire N__25948;
    wire N__25945;
    wire N__25942;
    wire N__25939;
    wire N__25934;
    wire N__25931;
    wire N__25928;
    wire N__25925;
    wire N__25922;
    wire N__25919;
    wire N__25916;
    wire N__25913;
    wire N__25912;
    wire N__25909;
    wire N__25906;
    wire N__25901;
    wire N__25898;
    wire N__25895;
    wire N__25892;
    wire N__25889;
    wire N__25886;
    wire N__25883;
    wire N__25880;
    wire N__25877;
    wire N__25876;
    wire N__25875;
    wire N__25872;
    wire N__25869;
    wire N__25866;
    wire N__25863;
    wire N__25860;
    wire N__25857;
    wire N__25852;
    wire N__25849;
    wire N__25846;
    wire N__25843;
    wire N__25840;
    wire N__25835;
    wire N__25834;
    wire N__25833;
    wire N__25832;
    wire N__25829;
    wire N__25826;
    wire N__25825;
    wire N__25824;
    wire N__25821;
    wire N__25818;
    wire N__25817;
    wire N__25816;
    wire N__25807;
    wire N__25804;
    wire N__25799;
    wire N__25796;
    wire N__25793;
    wire N__25784;
    wire N__25781;
    wire N__25778;
    wire N__25775;
    wire N__25772;
    wire N__25769;
    wire N__25766;
    wire N__25763;
    wire N__25762;
    wire N__25759;
    wire N__25756;
    wire N__25753;
    wire N__25750;
    wire N__25747;
    wire N__25744;
    wire N__25739;
    wire N__25736;
    wire N__25733;
    wire N__25730;
    wire N__25727;
    wire N__25724;
    wire N__25723;
    wire N__25720;
    wire N__25717;
    wire N__25714;
    wire N__25711;
    wire N__25706;
    wire N__25705;
    wire N__25704;
    wire N__25703;
    wire N__25700;
    wire N__25697;
    wire N__25696;
    wire N__25693;
    wire N__25690;
    wire N__25689;
    wire N__25686;
    wire N__25685;
    wire N__25684;
    wire N__25683;
    wire N__25682;
    wire N__25681;
    wire N__25680;
    wire N__25679;
    wire N__25678;
    wire N__25673;
    wire N__25672;
    wire N__25665;
    wire N__25664;
    wire N__25663;
    wire N__25662;
    wire N__25661;
    wire N__25660;
    wire N__25659;
    wire N__25656;
    wire N__25649;
    wire N__25642;
    wire N__25637;
    wire N__25634;
    wire N__25633;
    wire N__25632;
    wire N__25629;
    wire N__25628;
    wire N__25625;
    wire N__25616;
    wire N__25613;
    wire N__25610;
    wire N__25599;
    wire N__25590;
    wire N__25587;
    wire N__25574;
    wire N__25571;
    wire N__25568;
    wire N__25565;
    wire N__25562;
    wire N__25559;
    wire N__25558;
    wire N__25555;
    wire N__25552;
    wire N__25549;
    wire N__25544;
    wire N__25541;
    wire N__25538;
    wire N__25535;
    wire N__25532;
    wire N__25529;
    wire N__25526;
    wire N__25525;
    wire N__25522;
    wire N__25519;
    wire N__25514;
    wire N__25511;
    wire N__25508;
    wire N__25505;
    wire N__25502;
    wire N__25501;
    wire N__25498;
    wire N__25495;
    wire N__25494;
    wire N__25491;
    wire N__25488;
    wire N__25485;
    wire N__25478;
    wire N__25475;
    wire N__25472;
    wire N__25469;
    wire N__25466;
    wire N__25463;
    wire N__25462;
    wire N__25459;
    wire N__25456;
    wire N__25453;
    wire N__25450;
    wire N__25445;
    wire N__25442;
    wire N__25439;
    wire N__25436;
    wire N__25433;
    wire N__25430;
    wire N__25429;
    wire N__25426;
    wire N__25425;
    wire N__25422;
    wire N__25419;
    wire N__25416;
    wire N__25409;
    wire N__25406;
    wire N__25403;
    wire N__25400;
    wire N__25397;
    wire N__25394;
    wire N__25393;
    wire N__25390;
    wire N__25389;
    wire N__25386;
    wire N__25383;
    wire N__25380;
    wire N__25377;
    wire N__25374;
    wire N__25371;
    wire N__25368;
    wire N__25361;
    wire N__25358;
    wire N__25355;
    wire N__25352;
    wire N__25349;
    wire N__25348;
    wire N__25345;
    wire N__25342;
    wire N__25341;
    wire N__25336;
    wire N__25333;
    wire N__25328;
    wire N__25325;
    wire N__25322;
    wire N__25319;
    wire N__25316;
    wire N__25313;
    wire N__25312;
    wire N__25309;
    wire N__25308;
    wire N__25305;
    wire N__25302;
    wire N__25299;
    wire N__25292;
    wire N__25289;
    wire N__25286;
    wire N__25283;
    wire N__25280;
    wire N__25277;
    wire N__25276;
    wire N__25273;
    wire N__25270;
    wire N__25267;
    wire N__25264;
    wire N__25261;
    wire N__25256;
    wire N__25253;
    wire N__25250;
    wire N__25247;
    wire N__25244;
    wire N__25241;
    wire N__25240;
    wire N__25239;
    wire N__25236;
    wire N__25233;
    wire N__25230;
    wire N__25227;
    wire N__25224;
    wire N__25217;
    wire N__25214;
    wire N__25211;
    wire N__25208;
    wire N__25205;
    wire N__25202;
    wire N__25199;
    wire N__25198;
    wire N__25195;
    wire N__25192;
    wire N__25187;
    wire N__25186;
    wire N__25183;
    wire N__25180;
    wire N__25175;
    wire N__25174;
    wire N__25171;
    wire N__25168;
    wire N__25165;
    wire N__25162;
    wire N__25161;
    wire N__25158;
    wire N__25155;
    wire N__25152;
    wire N__25149;
    wire N__25144;
    wire N__25139;
    wire N__25136;
    wire N__25133;
    wire N__25130;
    wire N__25127;
    wire N__25124;
    wire N__25123;
    wire N__25120;
    wire N__25117;
    wire N__25114;
    wire N__25113;
    wire N__25110;
    wire N__25107;
    wire N__25104;
    wire N__25097;
    wire N__25094;
    wire N__25091;
    wire N__25088;
    wire N__25085;
    wire N__25082;
    wire N__25079;
    wire N__25076;
    wire N__25073;
    wire N__25072;
    wire N__25071;
    wire N__25068;
    wire N__25065;
    wire N__25062;
    wire N__25059;
    wire N__25052;
    wire N__25049;
    wire N__25046;
    wire N__25043;
    wire N__25040;
    wire N__25037;
    wire N__25034;
    wire N__25033;
    wire N__25030;
    wire N__25027;
    wire N__25026;
    wire N__25023;
    wire N__25018;
    wire N__25013;
    wire N__25010;
    wire N__25007;
    wire N__25004;
    wire N__25001;
    wire N__24998;
    wire N__24995;
    wire N__24994;
    wire N__24991;
    wire N__24988;
    wire N__24985;
    wire N__24984;
    wire N__24981;
    wire N__24978;
    wire N__24975;
    wire N__24968;
    wire N__24965;
    wire N__24962;
    wire N__24959;
    wire N__24956;
    wire N__24953;
    wire N__24950;
    wire N__24947;
    wire N__24946;
    wire N__24943;
    wire N__24940;
    wire N__24935;
    wire N__24932;
    wire N__24929;
    wire N__24926;
    wire N__24923;
    wire N__24922;
    wire N__24919;
    wire N__24918;
    wire N__24915;
    wire N__24912;
    wire N__24907;
    wire N__24902;
    wire N__24899;
    wire N__24896;
    wire N__24893;
    wire N__24890;
    wire N__24887;
    wire N__24884;
    wire N__24883;
    wire N__24880;
    wire N__24877;
    wire N__24874;
    wire N__24871;
    wire N__24870;
    wire N__24865;
    wire N__24862;
    wire N__24857;
    wire N__24854;
    wire N__24851;
    wire N__24848;
    wire N__24845;
    wire N__24842;
    wire N__24839;
    wire N__24836;
    wire N__24833;
    wire N__24832;
    wire N__24829;
    wire N__24826;
    wire N__24825;
    wire N__24822;
    wire N__24819;
    wire N__24816;
    wire N__24811;
    wire N__24808;
    wire N__24803;
    wire N__24800;
    wire N__24797;
    wire N__24796;
    wire N__24793;
    wire N__24790;
    wire N__24787;
    wire N__24784;
    wire N__24781;
    wire N__24776;
    wire N__24773;
    wire N__24770;
    wire N__24767;
    wire N__24764;
    wire N__24763;
    wire N__24762;
    wire N__24761;
    wire N__24760;
    wire N__24759;
    wire N__24758;
    wire N__24757;
    wire N__24754;
    wire N__24753;
    wire N__24750;
    wire N__24747;
    wire N__24742;
    wire N__24741;
    wire N__24738;
    wire N__24737;
    wire N__24736;
    wire N__24735;
    wire N__24732;
    wire N__24729;
    wire N__24728;
    wire N__24727;
    wire N__24722;
    wire N__24719;
    wire N__24714;
    wire N__24707;
    wire N__24706;
    wire N__24705;
    wire N__24702;
    wire N__24701;
    wire N__24698;
    wire N__24689;
    wire N__24680;
    wire N__24671;
    wire N__24668;
    wire N__24659;
    wire N__24658;
    wire N__24655;
    wire N__24654;
    wire N__24651;
    wire N__24648;
    wire N__24645;
    wire N__24642;
    wire N__24639;
    wire N__24636;
    wire N__24633;
    wire N__24630;
    wire N__24625;
    wire N__24620;
    wire N__24617;
    wire N__24614;
    wire N__24611;
    wire N__24608;
    wire N__24605;
    wire N__24604;
    wire N__24601;
    wire N__24600;
    wire N__24597;
    wire N__24594;
    wire N__24591;
    wire N__24584;
    wire N__24581;
    wire N__24578;
    wire N__24575;
    wire N__24574;
    wire N__24571;
    wire N__24568;
    wire N__24565;
    wire N__24560;
    wire N__24557;
    wire N__24554;
    wire N__24551;
    wire N__24550;
    wire N__24547;
    wire N__24544;
    wire N__24543;
    wire N__24540;
    wire N__24537;
    wire N__24534;
    wire N__24527;
    wire N__24524;
    wire N__24521;
    wire N__24518;
    wire N__24517;
    wire N__24514;
    wire N__24511;
    wire N__24508;
    wire N__24503;
    wire N__24500;
    wire N__24497;
    wire N__24494;
    wire N__24491;
    wire N__24488;
    wire N__24487;
    wire N__24484;
    wire N__24483;
    wire N__24480;
    wire N__24477;
    wire N__24474;
    wire N__24471;
    wire N__24466;
    wire N__24461;
    wire N__24458;
    wire N__24455;
    wire N__24452;
    wire N__24449;
    wire N__24446;
    wire N__24443;
    wire N__24440;
    wire N__24437;
    wire N__24434;
    wire N__24431;
    wire N__24428;
    wire N__24425;
    wire N__24422;
    wire N__24419;
    wire N__24416;
    wire N__24413;
    wire N__24410;
    wire N__24407;
    wire N__24404;
    wire N__24401;
    wire N__24398;
    wire N__24395;
    wire N__24392;
    wire N__24389;
    wire N__24386;
    wire N__24383;
    wire N__24380;
    wire N__24377;
    wire N__24374;
    wire N__24371;
    wire N__24368;
    wire N__24365;
    wire N__24362;
    wire N__24359;
    wire N__24356;
    wire N__24353;
    wire N__24350;
    wire N__24349;
    wire N__24348;
    wire N__24347;
    wire N__24346;
    wire N__24345;
    wire N__24344;
    wire N__24343;
    wire N__24342;
    wire N__24323;
    wire N__24320;
    wire N__24317;
    wire N__24314;
    wire N__24311;
    wire N__24308;
    wire N__24305;
    wire N__24302;
    wire N__24299;
    wire N__24296;
    wire N__24293;
    wire N__24290;
    wire N__24287;
    wire N__24284;
    wire N__24283;
    wire N__24280;
    wire N__24277;
    wire N__24274;
    wire N__24273;
    wire N__24270;
    wire N__24267;
    wire N__24264;
    wire N__24261;
    wire N__24258;
    wire N__24255;
    wire N__24248;
    wire N__24245;
    wire N__24244;
    wire N__24241;
    wire N__24238;
    wire N__24235;
    wire N__24232;
    wire N__24231;
    wire N__24228;
    wire N__24225;
    wire N__24222;
    wire N__24215;
    wire N__24212;
    wire N__24209;
    wire N__24208;
    wire N__24205;
    wire N__24202;
    wire N__24201;
    wire N__24198;
    wire N__24195;
    wire N__24192;
    wire N__24185;
    wire N__24182;
    wire N__24179;
    wire N__24178;
    wire N__24175;
    wire N__24172;
    wire N__24171;
    wire N__24168;
    wire N__24165;
    wire N__24162;
    wire N__24155;
    wire N__24152;
    wire N__24149;
    wire N__24146;
    wire N__24143;
    wire N__24140;
    wire N__24137;
    wire N__24134;
    wire N__24131;
    wire N__24128;
    wire N__24125;
    wire N__24122;
    wire N__24119;
    wire N__24116;
    wire N__24113;
    wire N__24110;
    wire N__24107;
    wire N__24104;
    wire N__24101;
    wire N__24098;
    wire N__24095;
    wire N__24092;
    wire N__24091;
    wire N__24088;
    wire N__24085;
    wire N__24080;
    wire N__24077;
    wire N__24076;
    wire N__24075;
    wire N__24074;
    wire N__24071;
    wire N__24070;
    wire N__24067;
    wire N__24066;
    wire N__24063;
    wire N__24062;
    wire N__24061;
    wire N__24060;
    wire N__24059;
    wire N__24044;
    wire N__24043;
    wire N__24042;
    wire N__24041;
    wire N__24038;
    wire N__24037;
    wire N__24034;
    wire N__24033;
    wire N__24030;
    wire N__24027;
    wire N__24024;
    wire N__24011;
    wire N__24008;
    wire N__24005;
    wire N__24004;
    wire N__23999;
    wire N__23996;
    wire N__23993;
    wire N__23990;
    wire N__23987;
    wire N__23984;
    wire N__23981;
    wire N__23978;
    wire N__23969;
    wire N__23966;
    wire N__23963;
    wire N__23960;
    wire N__23959;
    wire N__23956;
    wire N__23951;
    wire N__23948;
    wire N__23945;
    wire N__23942;
    wire N__23939;
    wire N__23936;
    wire N__23933;
    wire N__23930;
    wire N__23927;
    wire N__23924;
    wire N__23921;
    wire N__23918;
    wire N__23915;
    wire N__23912;
    wire N__23909;
    wire N__23908;
    wire N__23905;
    wire N__23902;
    wire N__23901;
    wire N__23898;
    wire N__23895;
    wire N__23892;
    wire N__23891;
    wire N__23886;
    wire N__23883;
    wire N__23880;
    wire N__23877;
    wire N__23874;
    wire N__23867;
    wire N__23864;
    wire N__23861;
    wire N__23858;
    wire N__23855;
    wire N__23852;
    wire N__23849;
    wire N__23846;
    wire N__23845;
    wire N__23842;
    wire N__23839;
    wire N__23838;
    wire N__23835;
    wire N__23832;
    wire N__23829;
    wire N__23828;
    wire N__23823;
    wire N__23820;
    wire N__23817;
    wire N__23814;
    wire N__23811;
    wire N__23804;
    wire N__23801;
    wire N__23798;
    wire N__23795;
    wire N__23792;
    wire N__23789;
    wire N__23788;
    wire N__23785;
    wire N__23782;
    wire N__23779;
    wire N__23776;
    wire N__23773;
    wire N__23772;
    wire N__23769;
    wire N__23768;
    wire N__23765;
    wire N__23762;
    wire N__23759;
    wire N__23756;
    wire N__23747;
    wire N__23744;
    wire N__23741;
    wire N__23738;
    wire N__23735;
    wire N__23732;
    wire N__23729;
    wire N__23726;
    wire N__23723;
    wire N__23722;
    wire N__23719;
    wire N__23716;
    wire N__23711;
    wire N__23710;
    wire N__23707;
    wire N__23704;
    wire N__23703;
    wire N__23698;
    wire N__23695;
    wire N__23692;
    wire N__23687;
    wire N__23684;
    wire N__23681;
    wire N__23678;
    wire N__23675;
    wire N__23672;
    wire N__23669;
    wire N__23666;
    wire N__23665;
    wire N__23662;
    wire N__23659;
    wire N__23658;
    wire N__23653;
    wire N__23650;
    wire N__23649;
    wire N__23646;
    wire N__23643;
    wire N__23640;
    wire N__23635;
    wire N__23630;
    wire N__23627;
    wire N__23624;
    wire N__23621;
    wire N__23618;
    wire N__23615;
    wire N__23612;
    wire N__23611;
    wire N__23608;
    wire N__23605;
    wire N__23600;
    wire N__23599;
    wire N__23596;
    wire N__23595;
    wire N__23592;
    wire N__23589;
    wire N__23586;
    wire N__23579;
    wire N__23576;
    wire N__23573;
    wire N__23570;
    wire N__23567;
    wire N__23564;
    wire N__23561;
    wire N__23558;
    wire N__23555;
    wire N__23552;
    wire N__23549;
    wire N__23546;
    wire N__23543;
    wire N__23540;
    wire N__23537;
    wire N__23534;
    wire N__23531;
    wire N__23528;
    wire N__23525;
    wire N__23522;
    wire N__23519;
    wire N__23516;
    wire N__23513;
    wire N__23510;
    wire N__23507;
    wire N__23504;
    wire N__23501;
    wire N__23498;
    wire N__23495;
    wire N__23492;
    wire N__23489;
    wire N__23488;
    wire N__23485;
    wire N__23482;
    wire N__23481;
    wire N__23476;
    wire N__23475;
    wire N__23472;
    wire N__23469;
    wire N__23466;
    wire N__23459;
    wire N__23456;
    wire N__23453;
    wire N__23450;
    wire N__23447;
    wire N__23444;
    wire N__23441;
    wire N__23438;
    wire N__23435;
    wire N__23432;
    wire N__23429;
    wire N__23426;
    wire N__23425;
    wire N__23422;
    wire N__23421;
    wire N__23418;
    wire N__23415;
    wire N__23412;
    wire N__23409;
    wire N__23406;
    wire N__23403;
    wire N__23400;
    wire N__23397;
    wire N__23392;
    wire N__23387;
    wire N__23384;
    wire N__23381;
    wire N__23378;
    wire N__23375;
    wire N__23374;
    wire N__23373;
    wire N__23372;
    wire N__23371;
    wire N__23370;
    wire N__23369;
    wire N__23366;
    wire N__23365;
    wire N__23364;
    wire N__23363;
    wire N__23362;
    wire N__23361;
    wire N__23354;
    wire N__23353;
    wire N__23352;
    wire N__23349;
    wire N__23348;
    wire N__23347;
    wire N__23346;
    wire N__23345;
    wire N__23342;
    wire N__23341;
    wire N__23338;
    wire N__23333;
    wire N__23332;
    wire N__23331;
    wire N__23328;
    wire N__23325;
    wire N__23324;
    wire N__23319;
    wire N__23316;
    wire N__23313;
    wire N__23306;
    wire N__23299;
    wire N__23294;
    wire N__23291;
    wire N__23288;
    wire N__23277;
    wire N__23272;
    wire N__23255;
    wire N__23254;
    wire N__23251;
    wire N__23248;
    wire N__23245;
    wire N__23244;
    wire N__23239;
    wire N__23236;
    wire N__23231;
    wire N__23228;
    wire N__23225;
    wire N__23222;
    wire N__23221;
    wire N__23220;
    wire N__23217;
    wire N__23214;
    wire N__23211;
    wire N__23208;
    wire N__23205;
    wire N__23202;
    wire N__23199;
    wire N__23194;
    wire N__23189;
    wire N__23188;
    wire N__23185;
    wire N__23182;
    wire N__23179;
    wire N__23178;
    wire N__23175;
    wire N__23172;
    wire N__23169;
    wire N__23166;
    wire N__23159;
    wire N__23156;
    wire N__23153;
    wire N__23150;
    wire N__23147;
    wire N__23144;
    wire N__23141;
    wire N__23140;
    wire N__23139;
    wire N__23136;
    wire N__23131;
    wire N__23126;
    wire N__23123;
    wire N__23120;
    wire N__23117;
    wire N__23114;
    wire N__23113;
    wire N__23110;
    wire N__23107;
    wire N__23106;
    wire N__23103;
    wire N__23100;
    wire N__23097;
    wire N__23092;
    wire N__23087;
    wire N__23084;
    wire N__23081;
    wire N__23078;
    wire N__23077;
    wire N__23074;
    wire N__23073;
    wire N__23070;
    wire N__23067;
    wire N__23064;
    wire N__23059;
    wire N__23054;
    wire N__23051;
    wire N__23048;
    wire N__23045;
    wire N__23042;
    wire N__23039;
    wire N__23036;
    wire N__23035;
    wire N__23032;
    wire N__23031;
    wire N__23028;
    wire N__23025;
    wire N__23022;
    wire N__23017;
    wire N__23012;
    wire N__23009;
    wire N__23006;
    wire N__23003;
    wire N__23000;
    wire N__22997;
    wire N__22994;
    wire N__22991;
    wire N__22990;
    wire N__22987;
    wire N__22984;
    wire N__22983;
    wire N__22980;
    wire N__22979;
    wire N__22978;
    wire N__22977;
    wire N__22974;
    wire N__22971;
    wire N__22970;
    wire N__22969;
    wire N__22966;
    wire N__22963;
    wire N__22960;
    wire N__22959;
    wire N__22958;
    wire N__22957;
    wire N__22956;
    wire N__22955;
    wire N__22954;
    wire N__22951;
    wire N__22950;
    wire N__22949;
    wire N__22944;
    wire N__22943;
    wire N__22942;
    wire N__22939;
    wire N__22938;
    wire N__22935;
    wire N__22930;
    wire N__22927;
    wire N__22924;
    wire N__22923;
    wire N__22922;
    wire N__22921;
    wire N__22920;
    wire N__22917;
    wire N__22912;
    wire N__22907;
    wire N__22906;
    wire N__22903;
    wire N__22898;
    wire N__22895;
    wire N__22892;
    wire N__22889;
    wire N__22888;
    wire N__22885;
    wire N__22882;
    wire N__22879;
    wire N__22874;
    wire N__22871;
    wire N__22862;
    wire N__22855;
    wire N__22854;
    wire N__22853;
    wire N__22852;
    wire N__22851;
    wire N__22850;
    wire N__22849;
    wire N__22848;
    wire N__22847;
    wire N__22846;
    wire N__22845;
    wire N__22842;
    wire N__22831;
    wire N__22828;
    wire N__22819;
    wire N__22812;
    wire N__22803;
    wire N__22794;
    wire N__22789;
    wire N__22772;
    wire N__22769;
    wire N__22766;
    wire N__22763;
    wire N__22760;
    wire N__22757;
    wire N__22754;
    wire N__22751;
    wire N__22748;
    wire N__22745;
    wire N__22742;
    wire N__22739;
    wire N__22736;
    wire N__22733;
    wire N__22732;
    wire N__22729;
    wire N__22726;
    wire N__22723;
    wire N__22720;
    wire N__22715;
    wire N__22712;
    wire N__22709;
    wire N__22706;
    wire N__22703;
    wire N__22700;
    wire N__22697;
    wire N__22694;
    wire N__22691;
    wire N__22688;
    wire N__22685;
    wire N__22684;
    wire N__22681;
    wire N__22678;
    wire N__22675;
    wire N__22674;
    wire N__22669;
    wire N__22666;
    wire N__22661;
    wire N__22658;
    wire N__22655;
    wire N__22652;
    wire N__22649;
    wire N__22646;
    wire N__22645;
    wire N__22642;
    wire N__22639;
    wire N__22636;
    wire N__22635;
    wire N__22630;
    wire N__22627;
    wire N__22622;
    wire N__22619;
    wire N__22616;
    wire N__22613;
    wire N__22610;
    wire N__22607;
    wire N__22606;
    wire N__22605;
    wire N__22602;
    wire N__22597;
    wire N__22592;
    wire N__22589;
    wire N__22586;
    wire N__22583;
    wire N__22580;
    wire N__22577;
    wire N__22574;
    wire N__22571;
    wire N__22570;
    wire N__22567;
    wire N__22564;
    wire N__22563;
    wire N__22560;
    wire N__22555;
    wire N__22552;
    wire N__22549;
    wire N__22544;
    wire N__22541;
    wire N__22538;
    wire N__22535;
    wire N__22532;
    wire N__22529;
    wire N__22528;
    wire N__22525;
    wire N__22524;
    wire N__22521;
    wire N__22518;
    wire N__22515;
    wire N__22510;
    wire N__22507;
    wire N__22502;
    wire N__22499;
    wire N__22496;
    wire N__22493;
    wire N__22490;
    wire N__22489;
    wire N__22486;
    wire N__22483;
    wire N__22480;
    wire N__22479;
    wire N__22476;
    wire N__22473;
    wire N__22470;
    wire N__22463;
    wire N__22460;
    wire N__22457;
    wire N__22454;
    wire N__22451;
    wire N__22448;
    wire N__22445;
    wire N__22444;
    wire N__22443;
    wire N__22440;
    wire N__22437;
    wire N__22434;
    wire N__22431;
    wire N__22428;
    wire N__22425;
    wire N__22418;
    wire N__22415;
    wire N__22412;
    wire N__22409;
    wire N__22406;
    wire N__22405;
    wire N__22402;
    wire N__22399;
    wire N__22396;
    wire N__22393;
    wire N__22388;
    wire N__22385;
    wire N__22382;
    wire N__22379;
    wire N__22376;
    wire N__22373;
    wire N__22370;
    wire N__22369;
    wire N__22366;
    wire N__22363;
    wire N__22360;
    wire N__22355;
    wire N__22352;
    wire N__22349;
    wire N__22346;
    wire N__22343;
    wire N__22340;
    wire N__22339;
    wire N__22338;
    wire N__22335;
    wire N__22332;
    wire N__22329;
    wire N__22326;
    wire N__22319;
    wire N__22316;
    wire N__22313;
    wire N__22310;
    wire N__22307;
    wire N__22304;
    wire N__22301;
    wire N__22298;
    wire N__22297;
    wire N__22294;
    wire N__22291;
    wire N__22286;
    wire N__22283;
    wire N__22280;
    wire N__22277;
    wire N__22274;
    wire N__22271;
    wire N__22270;
    wire N__22269;
    wire N__22266;
    wire N__22261;
    wire N__22258;
    wire N__22253;
    wire N__22250;
    wire N__22247;
    wire N__22244;
    wire N__22241;
    wire N__22240;
    wire N__22237;
    wire N__22234;
    wire N__22231;
    wire N__22230;
    wire N__22227;
    wire N__22224;
    wire N__22221;
    wire N__22214;
    wire N__22211;
    wire N__22208;
    wire N__22205;
    wire N__22202;
    wire N__22199;
    wire N__22198;
    wire N__22195;
    wire N__22192;
    wire N__22189;
    wire N__22186;
    wire N__22183;
    wire N__22178;
    wire N__22175;
    wire N__22172;
    wire N__22169;
    wire N__22166;
    wire N__22165;
    wire N__22162;
    wire N__22159;
    wire N__22156;
    wire N__22155;
    wire N__22150;
    wire N__22147;
    wire N__22142;
    wire N__22139;
    wire N__22136;
    wire N__22133;
    wire N__22130;
    wire N__22127;
    wire N__22126;
    wire N__22125;
    wire N__22122;
    wire N__22119;
    wire N__22116;
    wire N__22113;
    wire N__22110;
    wire N__22107;
    wire N__22100;
    wire N__22097;
    wire N__22094;
    wire N__22091;
    wire N__22088;
    wire N__22085;
    wire N__22082;
    wire N__22081;
    wire N__22080;
    wire N__22077;
    wire N__22074;
    wire N__22071;
    wire N__22068;
    wire N__22065;
    wire N__22062;
    wire N__22055;
    wire N__22052;
    wire N__22049;
    wire N__22046;
    wire N__22043;
    wire N__22042;
    wire N__22039;
    wire N__22038;
    wire N__22035;
    wire N__22030;
    wire N__22025;
    wire N__22022;
    wire N__22019;
    wire N__22016;
    wire N__22013;
    wire N__22012;
    wire N__22009;
    wire N__22006;
    wire N__22003;
    wire N__22002;
    wire N__21999;
    wire N__21996;
    wire N__21993;
    wire N__21986;
    wire N__21983;
    wire N__21980;
    wire N__21977;
    wire N__21976;
    wire N__21973;
    wire N__21970;
    wire N__21967;
    wire N__21962;
    wire N__21959;
    wire N__21956;
    wire N__21953;
    wire N__21952;
    wire N__21951;
    wire N__21948;
    wire N__21945;
    wire N__21942;
    wire N__21937;
    wire N__21932;
    wire N__21929;
    wire N__21926;
    wire N__21925;
    wire N__21922;
    wire N__21919;
    wire N__21916;
    wire N__21913;
    wire N__21912;
    wire N__21909;
    wire N__21906;
    wire N__21903;
    wire N__21896;
    wire N__21893;
    wire N__21890;
    wire N__21889;
    wire N__21886;
    wire N__21883;
    wire N__21880;
    wire N__21877;
    wire N__21876;
    wire N__21873;
    wire N__21870;
    wire N__21867;
    wire N__21860;
    wire N__21857;
    wire N__21854;
    wire N__21851;
    wire N__21848;
    wire N__21845;
    wire N__21844;
    wire N__21841;
    wire N__21838;
    wire N__21835;
    wire N__21832;
    wire N__21831;
    wire N__21826;
    wire N__21823;
    wire N__21818;
    wire N__21817;
    wire N__21814;
    wire N__21811;
    wire N__21808;
    wire N__21803;
    wire N__21800;
    wire N__21797;
    wire N__21794;
    wire N__21793;
    wire N__21792;
    wire N__21791;
    wire N__21790;
    wire N__21789;
    wire N__21788;
    wire N__21785;
    wire N__21784;
    wire N__21781;
    wire N__21778;
    wire N__21777;
    wire N__21776;
    wire N__21773;
    wire N__21772;
    wire N__21771;
    wire N__21766;
    wire N__21765;
    wire N__21764;
    wire N__21763;
    wire N__21762;
    wire N__21761;
    wire N__21758;
    wire N__21753;
    wire N__21750;
    wire N__21747;
    wire N__21746;
    wire N__21743;
    wire N__21742;
    wire N__21741;
    wire N__21738;
    wire N__21731;
    wire N__21728;
    wire N__21721;
    wire N__21716;
    wire N__21711;
    wire N__21706;
    wire N__21697;
    wire N__21680;
    wire N__21677;
    wire N__21676;
    wire N__21673;
    wire N__21670;
    wire N__21667;
    wire N__21664;
    wire N__21661;
    wire N__21658;
    wire N__21653;
    wire N__21650;
    wire N__21647;
    wire N__21644;
    wire N__21643;
    wire N__21640;
    wire N__21637;
    wire N__21632;
    wire N__21629;
    wire N__21626;
    wire N__21623;
    wire N__21620;
    wire N__21617;
    wire N__21616;
    wire N__21615;
    wire N__21612;
    wire N__21609;
    wire N__21606;
    wire N__21603;
    wire N__21598;
    wire N__21593;
    wire N__21590;
    wire N__21587;
    wire N__21584;
    wire N__21581;
    wire N__21580;
    wire N__21577;
    wire N__21574;
    wire N__21571;
    wire N__21568;
    wire N__21563;
    wire N__21560;
    wire N__21559;
    wire N__21556;
    wire N__21553;
    wire N__21552;
    wire N__21549;
    wire N__21546;
    wire N__21543;
    wire N__21536;
    wire N__21533;
    wire N__21530;
    wire N__21527;
    wire N__21524;
    wire N__21521;
    wire N__21518;
    wire N__21517;
    wire N__21514;
    wire N__21511;
    wire N__21510;
    wire N__21507;
    wire N__21504;
    wire N__21501;
    wire N__21494;
    wire N__21493;
    wire N__21490;
    wire N__21487;
    wire N__21482;
    wire N__21481;
    wire N__21478;
    wire N__21475;
    wire N__21470;
    wire N__21467;
    wire N__21464;
    wire N__21461;
    wire N__21458;
    wire N__21455;
    wire N__21454;
    wire N__21453;
    wire N__21450;
    wire N__21447;
    wire N__21444;
    wire N__21441;
    wire N__21438;
    wire N__21435;
    wire N__21428;
    wire N__21427;
    wire N__21424;
    wire N__21421;
    wire N__21416;
    wire N__21413;
    wire N__21410;
    wire N__21407;
    wire N__21404;
    wire N__21401;
    wire N__21398;
    wire N__21395;
    wire N__21392;
    wire N__21391;
    wire N__21390;
    wire N__21387;
    wire N__21384;
    wire N__21381;
    wire N__21378;
    wire N__21371;
    wire N__21370;
    wire N__21367;
    wire N__21364;
    wire N__21361;
    wire N__21356;
    wire N__21353;
    wire N__21350;
    wire N__21347;
    wire N__21344;
    wire N__21341;
    wire N__21340;
    wire N__21337;
    wire N__21334;
    wire N__21331;
    wire N__21326;
    wire N__21323;
    wire N__21320;
    wire N__21317;
    wire N__21314;
    wire N__21311;
    wire N__21310;
    wire N__21307;
    wire N__21306;
    wire N__21303;
    wire N__21300;
    wire N__21297;
    wire N__21294;
    wire N__21291;
    wire N__21288;
    wire N__21285;
    wire N__21278;
    wire N__21275;
    wire N__21272;
    wire N__21269;
    wire N__21266;
    wire N__21265;
    wire N__21264;
    wire N__21261;
    wire N__21258;
    wire N__21255;
    wire N__21252;
    wire N__21249;
    wire N__21246;
    wire N__21241;
    wire N__21238;
    wire N__21233;
    wire N__21230;
    wire N__21227;
    wire N__21224;
    wire N__21221;
    wire N__21218;
    wire N__21215;
    wire N__21212;
    wire N__21209;
    wire N__21206;
    wire N__21203;
    wire N__21200;
    wire N__21197;
    wire N__21194;
    wire N__21191;
    wire N__21188;
    wire N__21185;
    wire N__21182;
    wire N__21179;
    wire N__21176;
    wire N__21173;
    wire N__21170;
    wire N__21167;
    wire N__21164;
    wire N__21161;
    wire N__21158;
    wire N__21155;
    wire N__21152;
    wire N__21149;
    wire N__21146;
    wire N__21143;
    wire N__21140;
    wire N__21137;
    wire N__21134;
    wire N__21131;
    wire N__21128;
    wire N__21125;
    wire N__21122;
    wire N__21119;
    wire N__21116;
    wire N__21113;
    wire N__21110;
    wire N__21107;
    wire N__21106;
    wire N__21103;
    wire N__21100;
    wire N__21095;
    wire N__21092;
    wire N__21089;
    wire N__21086;
    wire N__21083;
    wire N__21080;
    wire N__21077;
    wire N__21076;
    wire N__21073;
    wire N__21072;
    wire N__21069;
    wire N__21066;
    wire N__21063;
    wire N__21056;
    wire N__21053;
    wire N__21050;
    wire N__21047;
    wire N__21044;
    wire N__21041;
    wire N__21038;
    wire N__21035;
    wire N__21032;
    wire N__21029;
    wire N__21026;
    wire N__21023;
    wire N__21020;
    wire N__21017;
    wire N__21014;
    wire N__21011;
    wire N__21008;
    wire N__21005;
    wire N__21002;
    wire N__20999;
    wire N__20996;
    wire N__20993;
    wire N__20990;
    wire N__20987;
    wire N__20984;
    wire N__20981;
    wire N__20978;
    wire N__20975;
    wire N__20974;
    wire N__20971;
    wire N__20968;
    wire N__20965;
    wire N__20960;
    wire N__20957;
    wire N__20954;
    wire N__20951;
    wire N__20948;
    wire N__20945;
    wire N__20942;
    wire N__20939;
    wire N__20936;
    wire N__20933;
    wire N__20930;
    wire N__20927;
    wire N__20924;
    wire N__20921;
    wire N__20918;
    wire N__20917;
    wire N__20914;
    wire N__20911;
    wire N__20906;
    wire N__20903;
    wire N__20900;
    wire N__20897;
    wire N__20894;
    wire N__20891;
    wire N__20888;
    wire N__20885;
    wire N__20882;
    wire N__20879;
    wire N__20876;
    wire N__20873;
    wire N__20870;
    wire N__20867;
    wire N__20864;
    wire N__20861;
    wire N__20858;
    wire N__20855;
    wire N__20852;
    wire N__20849;
    wire N__20846;
    wire N__20843;
    wire N__20840;
    wire N__20837;
    wire N__20834;
    wire N__20831;
    wire N__20830;
    wire N__20829;
    wire N__20826;
    wire N__20823;
    wire N__20820;
    wire N__20817;
    wire N__20814;
    wire N__20811;
    wire N__20804;
    wire N__20803;
    wire N__20800;
    wire N__20797;
    wire N__20796;
    wire N__20793;
    wire N__20790;
    wire N__20787;
    wire N__20782;
    wire N__20779;
    wire N__20776;
    wire N__20773;
    wire N__20768;
    wire N__20767;
    wire N__20764;
    wire N__20763;
    wire N__20760;
    wire N__20757;
    wire N__20754;
    wire N__20751;
    wire N__20748;
    wire N__20745;
    wire N__20742;
    wire N__20737;
    wire N__20734;
    wire N__20731;
    wire N__20726;
    wire N__20723;
    wire N__20720;
    wire N__20717;
    wire N__20714;
    wire N__20711;
    wire N__20708;
    wire N__20705;
    wire N__20702;
    wire N__20699;
    wire N__20696;
    wire N__20693;
    wire N__20692;
    wire N__20689;
    wire N__20688;
    wire N__20685;
    wire N__20682;
    wire N__20679;
    wire N__20674;
    wire N__20671;
    wire N__20666;
    wire N__20663;
    wire N__20660;
    wire N__20657;
    wire N__20654;
    wire N__20651;
    wire N__20648;
    wire N__20647;
    wire N__20644;
    wire N__20643;
    wire N__20640;
    wire N__20637;
    wire N__20634;
    wire N__20631;
    wire N__20626;
    wire N__20623;
    wire N__20620;
    wire N__20615;
    wire N__20612;
    wire N__20611;
    wire N__20610;
    wire N__20609;
    wire N__20608;
    wire N__20607;
    wire N__20606;
    wire N__20603;
    wire N__20600;
    wire N__20599;
    wire N__20598;
    wire N__20597;
    wire N__20596;
    wire N__20595;
    wire N__20592;
    wire N__20589;
    wire N__20588;
    wire N__20587;
    wire N__20586;
    wire N__20585;
    wire N__20582;
    wire N__20581;
    wire N__20580;
    wire N__20579;
    wire N__20578;
    wire N__20573;
    wire N__20570;
    wire N__20567;
    wire N__20564;
    wire N__20561;
    wire N__20558;
    wire N__20557;
    wire N__20554;
    wire N__20551;
    wire N__20544;
    wire N__20539;
    wire N__20532;
    wire N__20527;
    wire N__20524;
    wire N__20519;
    wire N__20516;
    wire N__20507;
    wire N__20486;
    wire N__20483;
    wire N__20482;
    wire N__20479;
    wire N__20476;
    wire N__20473;
    wire N__20470;
    wire N__20469;
    wire N__20466;
    wire N__20463;
    wire N__20460;
    wire N__20453;
    wire N__20450;
    wire N__20449;
    wire N__20446;
    wire N__20443;
    wire N__20438;
    wire N__20437;
    wire N__20434;
    wire N__20431;
    wire N__20426;
    wire N__20425;
    wire N__20422;
    wire N__20419;
    wire N__20416;
    wire N__20415;
    wire N__20412;
    wire N__20409;
    wire N__20406;
    wire N__20399;
    wire N__20396;
    wire N__20393;
    wire N__20390;
    wire N__20387;
    wire N__20386;
    wire N__20385;
    wire N__20382;
    wire N__20379;
    wire N__20376;
    wire N__20369;
    wire N__20366;
    wire N__20363;
    wire N__20360;
    wire N__20357;
    wire N__20354;
    wire N__20353;
    wire N__20352;
    wire N__20349;
    wire N__20346;
    wire N__20343;
    wire N__20340;
    wire N__20337;
    wire N__20334;
    wire N__20331;
    wire N__20328;
    wire N__20321;
    wire N__20318;
    wire N__20315;
    wire N__20312;
    wire N__20309;
    wire N__20306;
    wire N__20303;
    wire N__20300;
    wire N__20297;
    wire N__20294;
    wire N__20291;
    wire N__20288;
    wire N__20285;
    wire N__20282;
    wire N__20281;
    wire N__20278;
    wire N__20275;
    wire N__20274;
    wire N__20269;
    wire N__20266;
    wire N__20263;
    wire N__20260;
    wire N__20257;
    wire N__20254;
    wire N__20249;
    wire N__20248;
    wire N__20245;
    wire N__20244;
    wire N__20241;
    wire N__20238;
    wire N__20235;
    wire N__20230;
    wire N__20227;
    wire N__20224;
    wire N__20219;
    wire N__20216;
    wire N__20213;
    wire N__20210;
    wire N__20207;
    wire N__20206;
    wire N__20203;
    wire N__20200;
    wire N__20197;
    wire N__20194;
    wire N__20189;
    wire N__20186;
    wire N__20183;
    wire N__20180;
    wire N__20177;
    wire N__20174;
    wire N__20171;
    wire N__20168;
    wire N__20165;
    wire N__20162;
    wire N__20159;
    wire N__20156;
    wire N__20155;
    wire N__20152;
    wire N__20151;
    wire N__20148;
    wire N__20145;
    wire N__20142;
    wire N__20139;
    wire N__20132;
    wire N__20131;
    wire N__20130;
    wire N__20127;
    wire N__20124;
    wire N__20121;
    wire N__20118;
    wire N__20115;
    wire N__20112;
    wire N__20107;
    wire N__20104;
    wire N__20101;
    wire N__20096;
    wire N__20093;
    wire N__20090;
    wire N__20087;
    wire N__20084;
    wire N__20081;
    wire N__20078;
    wire N__20075;
    wire N__20072;
    wire N__20071;
    wire N__20070;
    wire N__20067;
    wire N__20064;
    wire N__20061;
    wire N__20056;
    wire N__20053;
    wire N__20050;
    wire N__20045;
    wire N__20042;
    wire N__20039;
    wire N__20036;
    wire N__20033;
    wire N__20030;
    wire N__20027;
    wire N__20024;
    wire N__20023;
    wire N__20022;
    wire N__20019;
    wire N__20016;
    wire N__20013;
    wire N__20006;
    wire N__20003;
    wire N__20000;
    wire N__19997;
    wire N__19996;
    wire N__19993;
    wire N__19990;
    wire N__19987;
    wire N__19984;
    wire N__19983;
    wire N__19980;
    wire N__19977;
    wire N__19974;
    wire N__19967;
    wire N__19966;
    wire N__19965;
    wire N__19964;
    wire N__19963;
    wire N__19960;
    wire N__19959;
    wire N__19958;
    wire N__19955;
    wire N__19954;
    wire N__19953;
    wire N__19952;
    wire N__19949;
    wire N__19948;
    wire N__19945;
    wire N__19944;
    wire N__19943;
    wire N__19936;
    wire N__19935;
    wire N__19934;
    wire N__19931;
    wire N__19930;
    wire N__19925;
    wire N__19920;
    wire N__19915;
    wire N__19908;
    wire N__19905;
    wire N__19902;
    wire N__19895;
    wire N__19892;
    wire N__19877;
    wire N__19874;
    wire N__19873;
    wire N__19870;
    wire N__19869;
    wire N__19866;
    wire N__19863;
    wire N__19860;
    wire N__19853;
    wire N__19850;
    wire N__19847;
    wire N__19844;
    wire N__19843;
    wire N__19842;
    wire N__19839;
    wire N__19836;
    wire N__19833;
    wire N__19826;
    wire N__19823;
    wire N__19820;
    wire N__19817;
    wire N__19814;
    wire N__19811;
    wire N__19808;
    wire N__19805;
    wire N__19802;
    wire N__19801;
    wire N__19798;
    wire N__19795;
    wire N__19792;
    wire N__19787;
    wire N__19784;
    wire N__19783;
    wire N__19780;
    wire N__19777;
    wire N__19774;
    wire N__19769;
    wire N__19766;
    wire N__19763;
    wire N__19760;
    wire N__19757;
    wire N__19754;
    wire N__19751;
    wire N__19748;
    wire N__19747;
    wire N__19744;
    wire N__19741;
    wire N__19736;
    wire N__19733;
    wire N__19732;
    wire N__19731;
    wire N__19728;
    wire N__19725;
    wire N__19722;
    wire N__19719;
    wire N__19712;
    wire N__19709;
    wire N__19706;
    wire N__19703;
    wire N__19702;
    wire N__19701;
    wire N__19698;
    wire N__19693;
    wire N__19690;
    wire N__19685;
    wire N__19682;
    wire N__19679;
    wire N__19676;
    wire N__19673;
    wire N__19670;
    wire N__19669;
    wire N__19668;
    wire N__19665;
    wire N__19662;
    wire N__19659;
    wire N__19656;
    wire N__19651;
    wire N__19646;
    wire N__19643;
    wire N__19640;
    wire N__19637;
    wire N__19634;
    wire N__19633;
    wire N__19630;
    wire N__19627;
    wire N__19624;
    wire N__19621;
    wire N__19616;
    wire N__19615;
    wire N__19612;
    wire N__19609;
    wire N__19604;
    wire N__19603;
    wire N__19600;
    wire N__19597;
    wire N__19594;
    wire N__19589;
    wire N__19586;
    wire N__19583;
    wire N__19580;
    wire N__19577;
    wire N__19574;
    wire N__19571;
    wire N__19568;
    wire N__19565;
    wire N__19562;
    wire N__19559;
    wire N__19556;
    wire N__19553;
    wire N__19550;
    wire N__19549;
    wire N__19546;
    wire N__19543;
    wire N__19540;
    wire N__19539;
    wire N__19536;
    wire N__19533;
    wire N__19530;
    wire N__19523;
    wire N__19520;
    wire N__19519;
    wire N__19516;
    wire N__19513;
    wire N__19512;
    wire N__19509;
    wire N__19506;
    wire N__19503;
    wire N__19500;
    wire N__19497;
    wire N__19494;
    wire N__19487;
    wire N__19484;
    wire N__19483;
    wire N__19480;
    wire N__19477;
    wire N__19474;
    wire N__19471;
    wire N__19466;
    wire N__19463;
    wire N__19460;
    wire N__19457;
    wire N__19454;
    wire N__19451;
    wire N__19448;
    wire N__19445;
    wire N__19442;
    wire N__19439;
    wire N__19438;
    wire N__19435;
    wire N__19432;
    wire N__19431;
    wire N__19428;
    wire N__19425;
    wire N__19422;
    wire N__19419;
    wire N__19416;
    wire N__19409;
    wire N__19406;
    wire N__19403;
    wire N__19400;
    wire N__19399;
    wire N__19396;
    wire N__19395;
    wire N__19392;
    wire N__19389;
    wire N__19386;
    wire N__19383;
    wire N__19378;
    wire N__19373;
    wire N__19370;
    wire N__19367;
    wire N__19364;
    wire N__19361;
    wire N__19360;
    wire N__19357;
    wire N__19354;
    wire N__19353;
    wire N__19350;
    wire N__19347;
    wire N__19344;
    wire N__19337;
    wire N__19336;
    wire N__19333;
    wire N__19330;
    wire N__19327;
    wire N__19324;
    wire N__19321;
    wire N__19316;
    wire N__19313;
    wire N__19310;
    wire N__19309;
    wire N__19308;
    wire N__19305;
    wire N__19302;
    wire N__19297;
    wire N__19292;
    wire N__19289;
    wire N__19286;
    wire N__19283;
    wire N__19280;
    wire N__19277;
    wire N__19274;
    wire N__19271;
    wire N__19268;
    wire N__19267;
    wire N__19266;
    wire N__19263;
    wire N__19262;
    wire N__19261;
    wire N__19260;
    wire N__19259;
    wire N__19258;
    wire N__19257;
    wire N__19256;
    wire N__19255;
    wire N__19254;
    wire N__19253;
    wire N__19250;
    wire N__19247;
    wire N__19244;
    wire N__19241;
    wire N__19240;
    wire N__19239;
    wire N__19236;
    wire N__19233;
    wire N__19230;
    wire N__19227;
    wire N__19226;
    wire N__19225;
    wire N__19224;
    wire N__19221;
    wire N__19218;
    wire N__19215;
    wire N__19212;
    wire N__19211;
    wire N__19208;
    wire N__19201;
    wire N__19194;
    wire N__19193;
    wire N__19188;
    wire N__19179;
    wire N__19168;
    wire N__19165;
    wire N__19162;
    wire N__19157;
    wire N__19154;
    wire N__19139;
    wire N__19136;
    wire N__19135;
    wire N__19132;
    wire N__19131;
    wire N__19128;
    wire N__19125;
    wire N__19122;
    wire N__19115;
    wire N__19112;
    wire N__19111;
    wire N__19110;
    wire N__19107;
    wire N__19102;
    wire N__19099;
    wire N__19094;
    wire N__19091;
    wire N__19090;
    wire N__19089;
    wire N__19086;
    wire N__19083;
    wire N__19080;
    wire N__19073;
    wire N__19070;
    wire N__19067;
    wire N__19064;
    wire N__19063;
    wire N__19062;
    wire N__19059;
    wire N__19056;
    wire N__19053;
    wire N__19050;
    wire N__19043;
    wire N__19040;
    wire N__19037;
    wire N__19034;
    wire N__19031;
    wire N__19028;
    wire N__19025;
    wire N__19022;
    wire N__19021;
    wire N__19018;
    wire N__19017;
    wire N__19014;
    wire N__19011;
    wire N__19008;
    wire N__19005;
    wire N__18998;
    wire N__18995;
    wire N__18992;
    wire N__18989;
    wire N__18986;
    wire N__18983;
    wire N__18980;
    wire N__18979;
    wire N__18976;
    wire N__18975;
    wire N__18972;
    wire N__18969;
    wire N__18964;
    wire N__18959;
    wire N__18956;
    wire N__18953;
    wire N__18950;
    wire N__18947;
    wire N__18946;
    wire N__18945;
    wire N__18942;
    wire N__18937;
    wire N__18934;
    wire N__18929;
    wire N__18926;
    wire N__18923;
    wire N__18920;
    wire N__18917;
    wire N__18914;
    wire N__18911;
    wire N__18910;
    wire N__18907;
    wire N__18906;
    wire N__18903;
    wire N__18900;
    wire N__18897;
    wire N__18894;
    wire N__18887;
    wire N__18884;
    wire N__18881;
    wire N__18878;
    wire N__18875;
    wire N__18872;
    wire N__18869;
    wire N__18866;
    wire N__18863;
    wire N__18862;
    wire N__18859;
    wire N__18856;
    wire N__18855;
    wire N__18852;
    wire N__18849;
    wire N__18846;
    wire N__18839;
    wire N__18836;
    wire N__18833;
    wire N__18830;
    wire N__18827;
    wire N__18824;
    wire N__18821;
    wire N__18818;
    wire N__18815;
    wire N__18812;
    wire N__18809;
    wire N__18806;
    wire N__18805;
    wire N__18804;
    wire N__18801;
    wire N__18796;
    wire N__18791;
    wire N__18788;
    wire N__18785;
    wire N__18782;
    wire N__18781;
    wire N__18778;
    wire N__18777;
    wire N__18774;
    wire N__18771;
    wire N__18768;
    wire N__18761;
    wire N__18758;
    wire N__18757;
    wire N__18756;
    wire N__18753;
    wire N__18750;
    wire N__18747;
    wire N__18744;
    wire N__18739;
    wire N__18736;
    wire N__18731;
    wire N__18728;
    wire N__18725;
    wire N__18722;
    wire N__18719;
    wire N__18718;
    wire N__18717;
    wire N__18714;
    wire N__18709;
    wire N__18706;
    wire N__18701;
    wire N__18698;
    wire N__18695;
    wire N__18694;
    wire N__18693;
    wire N__18690;
    wire N__18687;
    wire N__18684;
    wire N__18677;
    wire N__18674;
    wire N__18671;
    wire N__18668;
    wire N__18665;
    wire N__18662;
    wire N__18659;
    wire N__18656;
    wire N__18655;
    wire N__18654;
    wire N__18649;
    wire N__18646;
    wire N__18643;
    wire N__18640;
    wire N__18635;
    wire N__18632;
    wire N__18629;
    wire N__18626;
    wire N__18623;
    wire N__18622;
    wire N__18621;
    wire N__18616;
    wire N__18613;
    wire N__18610;
    wire N__18607;
    wire N__18604;
    wire N__18601;
    wire N__18596;
    wire N__18593;
    wire N__18590;
    wire N__18587;
    wire N__18586;
    wire N__18583;
    wire N__18580;
    wire N__18577;
    wire N__18572;
    wire N__18569;
    wire N__18566;
    wire N__18563;
    wire N__18560;
    wire N__18557;
    wire N__18554;
    wire N__18551;
    wire N__18550;
    wire N__18547;
    wire N__18546;
    wire N__18543;
    wire N__18540;
    wire N__18537;
    wire N__18534;
    wire N__18527;
    wire N__18524;
    wire N__18521;
    wire N__18518;
    wire N__18515;
    wire N__18512;
    wire N__18511;
    wire N__18508;
    wire N__18505;
    wire N__18504;
    wire N__18501;
    wire N__18498;
    wire N__18495;
    wire N__18490;
    wire N__18485;
    wire N__18482;
    wire N__18479;
    wire N__18476;
    wire N__18473;
    wire N__18472;
    wire N__18469;
    wire N__18466;
    wire N__18463;
    wire N__18460;
    wire N__18459;
    wire N__18454;
    wire N__18451;
    wire N__18446;
    wire N__18443;
    wire N__18440;
    wire N__18437;
    wire N__18434;
    wire N__18433;
    wire N__18430;
    wire N__18427;
    wire N__18424;
    wire N__18421;
    wire N__18416;
    wire N__18413;
    wire N__18410;
    wire N__18409;
    wire N__18406;
    wire N__18403;
    wire N__18402;
    wire N__18397;
    wire N__18394;
    wire N__18389;
    wire N__18386;
    wire N__18383;
    wire N__18382;
    wire N__18379;
    wire N__18376;
    wire N__18373;
    wire N__18370;
    wire N__18369;
    wire N__18366;
    wire N__18363;
    wire N__18360;
    wire N__18353;
    wire N__18350;
    wire N__18347;
    wire N__18344;
    wire N__18341;
    wire N__18340;
    wire N__18339;
    wire N__18338;
    wire N__18337;
    wire N__18336;
    wire N__18333;
    wire N__18332;
    wire N__18331;
    wire N__18328;
    wire N__18327;
    wire N__18326;
    wire N__18323;
    wire N__18320;
    wire N__18319;
    wire N__18316;
    wire N__18315;
    wire N__18314;
    wire N__18313;
    wire N__18304;
    wire N__18299;
    wire N__18296;
    wire N__18285;
    wire N__18282;
    wire N__18279;
    wire N__18278;
    wire N__18273;
    wire N__18268;
    wire N__18261;
    wire N__18258;
    wire N__18251;
    wire N__18248;
    wire N__18247;
    wire N__18244;
    wire N__18241;
    wire N__18236;
    wire N__18233;
    wire N__18230;
    wire N__18227;
    wire N__18224;
    wire N__18221;
    wire N__18218;
    wire N__18215;
    wire N__18212;
    wire N__18209;
    wire N__18206;
    wire N__18203;
    wire N__18202;
    wire N__18199;
    wire N__18196;
    wire N__18193;
    wire N__18190;
    wire N__18185;
    wire N__18182;
    wire N__18179;
    wire N__18176;
    wire N__18173;
    wire N__18170;
    wire N__18167;
    wire N__18164;
    wire N__18161;
    wire N__18158;
    wire N__18155;
    wire N__18152;
    wire N__18149;
    wire N__18146;
    wire N__18143;
    wire N__18140;
    wire N__18139;
    wire N__18136;
    wire N__18133;
    wire N__18132;
    wire N__18129;
    wire N__18126;
    wire N__18123;
    wire N__18116;
    wire N__18113;
    wire N__18110;
    wire N__18107;
    wire N__18104;
    wire N__18101;
    wire N__18098;
    wire N__18095;
    wire N__18094;
    wire N__18091;
    wire N__18088;
    wire N__18085;
    wire N__18082;
    wire N__18077;
    wire N__18074;
    wire N__18071;
    wire N__18068;
    wire N__18065;
    wire N__18062;
    wire N__18059;
    wire N__18056;
    wire N__18053;
    wire N__18050;
    wire N__18047;
    wire N__18044;
    wire N__18041;
    wire N__18038;
    wire N__18035;
    wire N__18034;
    wire N__18033;
    wire N__18030;
    wire N__18025;
    wire N__18020;
    wire N__18017;
    wire N__18014;
    wire N__18011;
    wire N__18008;
    wire N__18005;
    wire N__18002;
    wire N__17999;
    wire N__17996;
    wire N__17993;
    wire N__17990;
    wire N__17987;
    wire N__17984;
    wire N__17981;
    wire N__17978;
    wire N__17975;
    wire N__17972;
    wire N__17969;
    wire N__17966;
    wire N__17963;
    wire N__17960;
    wire N__17957;
    wire N__17954;
    wire N__17951;
    wire N__17950;
    wire N__17947;
    wire N__17944;
    wire N__17941;
    wire N__17938;
    wire N__17933;
    wire N__17930;
    wire N__17927;
    wire N__17924;
    wire N__17921;
    wire N__17918;
    wire N__17915;
    wire N__17914;
    wire N__17911;
    wire N__17908;
    wire N__17905;
    wire N__17900;
    wire N__17897;
    wire N__17894;
    wire N__17891;
    wire N__17888;
    wire N__17885;
    wire N__17882;
    wire N__17879;
    wire N__17876;
    wire N__17873;
    wire N__17870;
    wire N__17867;
    wire N__17864;
    wire N__17861;
    wire N__17858;
    wire N__17855;
    wire N__17852;
    wire N__17849;
    wire N__17846;
    wire N__17843;
    wire N__17840;
    wire N__17837;
    wire N__17834;
    wire N__17831;
    wire N__17828;
    wire N__17825;
    wire N__17822;
    wire N__17819;
    wire N__17816;
    wire N__17813;
    wire N__17810;
    wire N__17807;
    wire N__17804;
    wire N__17801;
    wire N__17798;
    wire N__17795;
    wire N__17792;
    wire N__17789;
    wire N__17786;
    wire N__17783;
    wire N__17780;
    wire N__17777;
    wire N__17774;
    wire N__17771;
    wire N__17768;
    wire N__17765;
    wire N__17762;
    wire N__17759;
    wire N__17756;
    wire N__17753;
    wire N__17750;
    wire N__17747;
    wire N__17744;
    wire N__17741;
    wire N__17738;
    wire N__17735;
    wire N__17732;
    wire N__17729;
    wire N__17726;
    wire N__17723;
    wire N__17720;
    wire N__17717;
    wire N__17714;
    wire N__17713;
    wire N__17710;
    wire N__17707;
    wire N__17706;
    wire N__17703;
    wire N__17700;
    wire N__17697;
    wire N__17690;
    wire N__17687;
    wire N__17684;
    wire N__17681;
    wire N__17680;
    wire N__17677;
    wire N__17674;
    wire N__17671;
    wire N__17668;
    wire N__17665;
    wire N__17662;
    wire N__17657;
    wire N__17654;
    wire N__17651;
    wire N__17648;
    wire N__17645;
    wire N__17642;
    wire N__17639;
    wire N__17636;
    wire N__17633;
    wire N__17630;
    wire N__17627;
    wire N__17624;
    wire N__17621;
    wire N__17618;
    wire N__17615;
    wire N__17612;
    wire N__17609;
    wire N__17606;
    wire N__17603;
    wire N__17600;
    wire N__17597;
    wire N__17594;
    wire N__17591;
    wire N__17588;
    wire N__17585;
    wire N__17582;
    wire N__17579;
    wire N__17576;
    wire N__17573;
    wire N__17570;
    wire N__17567;
    wire N__17564;
    wire N__17561;
    wire N__17558;
    wire N__17555;
    wire N__17552;
    wire N__17549;
    wire N__17546;
    wire N__17543;
    wire N__17540;
    wire N__17537;
    wire N__17534;
    wire N__17531;
    wire N__17528;
    wire N__17525;
    wire N__17522;
    wire N__17519;
    wire N__17518;
    wire N__17515;
    wire N__17512;
    wire N__17509;
    wire N__17506;
    wire N__17501;
    wire N__17498;
    wire N__17495;
    wire N__17492;
    wire N__17491;
    wire N__17488;
    wire N__17487;
    wire N__17484;
    wire N__17481;
    wire N__17478;
    wire N__17473;
    wire N__17470;
    wire N__17465;
    wire N__17462;
    wire N__17459;
    wire N__17458;
    wire N__17457;
    wire N__17454;
    wire N__17451;
    wire N__17448;
    wire N__17441;
    wire N__17438;
    wire N__17437;
    wire N__17434;
    wire N__17431;
    wire N__17430;
    wire N__17427;
    wire N__17424;
    wire N__17421;
    wire N__17416;
    wire N__17411;
    wire N__17408;
    wire N__17405;
    wire N__17402;
    wire N__17399;
    wire N__17396;
    wire N__17393;
    wire N__17390;
    wire N__17389;
    wire N__17386;
    wire N__17383;
    wire N__17380;
    wire N__17377;
    wire N__17376;
    wire N__17371;
    wire N__17368;
    wire N__17363;
    wire N__17362;
    wire N__17359;
    wire N__17356;
    wire N__17353;
    wire N__17350;
    wire N__17345;
    wire N__17342;
    wire N__17339;
    wire N__17336;
    wire N__17333;
    wire N__17330;
    wire N__17327;
    wire N__17324;
    wire N__17323;
    wire N__17320;
    wire N__17319;
    wire N__17316;
    wire N__17313;
    wire N__17310;
    wire N__17303;
    wire N__17300;
    wire N__17297;
    wire N__17294;
    wire N__17291;
    wire N__17288;
    wire N__17285;
    wire N__17282;
    wire N__17279;
    wire N__17276;
    wire N__17273;
    wire N__17270;
    wire N__17267;
    wire N__17264;
    wire N__17261;
    wire N__17258;
    wire N__17255;
    wire N__17254;
    wire N__17251;
    wire N__17248;
    wire N__17247;
    wire N__17244;
    wire N__17241;
    wire N__17238;
    wire N__17231;
    wire N__17228;
    wire N__17225;
    wire N__17222;
    wire N__17221;
    wire N__17220;
    wire N__17219;
    wire N__17218;
    wire N__17217;
    wire N__17214;
    wire N__17213;
    wire N__17212;
    wire N__17211;
    wire N__17210;
    wire N__17207;
    wire N__17204;
    wire N__17203;
    wire N__17202;
    wire N__17199;
    wire N__17198;
    wire N__17195;
    wire N__17194;
    wire N__17191;
    wire N__17188;
    wire N__17185;
    wire N__17180;
    wire N__17171;
    wire N__17160;
    wire N__17147;
    wire N__17144;
    wire N__17141;
    wire N__17138;
    wire N__17135;
    wire N__17132;
    wire N__17129;
    wire N__17126;
    wire N__17123;
    wire N__17122;
    wire N__17121;
    wire N__17118;
    wire N__17115;
    wire N__17112;
    wire N__17109;
    wire N__17104;
    wire N__17101;
    wire N__17098;
    wire N__17093;
    wire N__17090;
    wire N__17087;
    wire N__17084;
    wire N__17081;
    wire N__17080;
    wire N__17077;
    wire N__17074;
    wire N__17071;
    wire N__17066;
    wire N__17063;
    wire N__17060;
    wire N__17057;
    wire N__17054;
    wire N__17051;
    wire N__17050;
    wire N__17047;
    wire N__17046;
    wire N__17043;
    wire N__17040;
    wire N__17037;
    wire N__17030;
    wire N__17027;
    wire N__17024;
    wire N__17021;
    wire N__17018;
    wire N__17015;
    wire N__17012;
    wire N__17009;
    wire N__17006;
    wire N__17003;
    wire N__17002;
    wire N__16999;
    wire N__16996;
    wire N__16993;
    wire N__16990;
    wire N__16985;
    wire N__16982;
    wire N__16981;
    wire N__16980;
    wire N__16977;
    wire N__16972;
    wire N__16967;
    wire N__16964;
    wire N__16961;
    wire N__16958;
    wire N__16957;
    wire N__16954;
    wire N__16953;
    wire N__16950;
    wire N__16947;
    wire N__16942;
    wire N__16937;
    wire N__16934;
    wire N__16931;
    wire N__16928;
    wire N__16925;
    wire N__16922;
    wire N__16919;
    wire N__16916;
    wire N__16915;
    wire N__16912;
    wire N__16909;
    wire N__16908;
    wire N__16905;
    wire N__16902;
    wire N__16899;
    wire N__16892;
    wire N__16891;
    wire N__16888;
    wire N__16885;
    wire N__16884;
    wire N__16881;
    wire N__16878;
    wire N__16875;
    wire N__16868;
    wire N__16865;
    wire N__16862;
    wire N__16859;
    wire N__16856;
    wire N__16855;
    wire N__16852;
    wire N__16849;
    wire N__16846;
    wire N__16843;
    wire N__16842;
    wire N__16839;
    wire N__16836;
    wire N__16833;
    wire N__16826;
    wire N__16823;
    wire N__16820;
    wire N__16817;
    wire N__16814;
    wire N__16811;
    wire N__16810;
    wire N__16809;
    wire N__16806;
    wire N__16803;
    wire N__16800;
    wire N__16797;
    wire N__16790;
    wire N__16787;
    wire N__16784;
    wire N__16781;
    wire N__16778;
    wire N__16775;
    wire N__16772;
    wire N__16769;
    wire N__16766;
    wire N__16763;
    wire N__16762;
    wire N__16761;
    wire N__16758;
    wire N__16755;
    wire N__16752;
    wire N__16747;
    wire N__16744;
    wire N__16741;
    wire N__16736;
    wire N__16733;
    wire N__16730;
    wire N__16727;
    wire N__16724;
    wire N__16721;
    wire N__16718;
    wire N__16715;
    wire N__16712;
    wire N__16709;
    wire N__16708;
    wire N__16707;
    wire N__16704;
    wire N__16701;
    wire N__16698;
    wire N__16695;
    wire N__16692;
    wire N__16685;
    wire N__16682;
    wire N__16679;
    wire N__16676;
    wire N__16675;
    wire N__16674;
    wire N__16671;
    wire N__16666;
    wire N__16663;
    wire N__16660;
    wire N__16655;
    wire N__16652;
    wire N__16649;
    wire N__16646;
    wire N__16643;
    wire N__16640;
    wire N__16637;
    wire N__16636;
    wire N__16633;
    wire N__16630;
    wire N__16629;
    wire N__16626;
    wire N__16621;
    wire N__16616;
    wire N__16613;
    wire N__16610;
    wire N__16607;
    wire N__16604;
    wire N__16603;
    wire N__16602;
    wire N__16601;
    wire N__16600;
    wire N__16599;
    wire N__16598;
    wire N__16597;
    wire N__16594;
    wire N__16593;
    wire N__16592;
    wire N__16591;
    wire N__16588;
    wire N__16583;
    wire N__16580;
    wire N__16575;
    wire N__16572;
    wire N__16569;
    wire N__16562;
    wire N__16547;
    wire N__16546;
    wire N__16543;
    wire N__16540;
    wire N__16537;
    wire N__16534;
    wire N__16531;
    wire N__16526;
    wire N__16523;
    wire N__16522;
    wire N__16519;
    wire N__16516;
    wire N__16513;
    wire N__16510;
    wire N__16507;
    wire N__16504;
    wire N__16499;
    wire N__16498;
    wire N__16495;
    wire N__16492;
    wire N__16489;
    wire N__16486;
    wire N__16485;
    wire N__16482;
    wire N__16479;
    wire N__16476;
    wire N__16469;
    wire N__16466;
    wire N__16463;
    wire N__16460;
    wire N__16457;
    wire N__16456;
    wire N__16453;
    wire N__16450;
    wire N__16447;
    wire N__16444;
    wire N__16439;
    wire N__16436;
    wire N__16433;
    wire N__16430;
    wire N__16427;
    wire N__16426;
    wire N__16423;
    wire N__16420;
    wire N__16417;
    wire N__16414;
    wire N__16413;
    wire N__16410;
    wire N__16407;
    wire N__16404;
    wire N__16397;
    wire N__16396;
    wire N__16393;
    wire N__16390;
    wire N__16387;
    wire N__16386;
    wire N__16383;
    wire N__16380;
    wire N__16377;
    wire N__16370;
    wire N__16369;
    wire N__16368;
    wire N__16367;
    wire N__16366;
    wire N__16365;
    wire N__16364;
    wire N__16361;
    wire N__16358;
    wire N__16355;
    wire N__16354;
    wire N__16353;
    wire N__16350;
    wire N__16347;
    wire N__16346;
    wire N__16343;
    wire N__16340;
    wire N__16339;
    wire N__16336;
    wire N__16333;
    wire N__16328;
    wire N__16319;
    wire N__16312;
    wire N__16309;
    wire N__16298;
    wire N__16295;
    wire N__16292;
    wire N__16289;
    wire N__16288;
    wire N__16285;
    wire N__16282;
    wire N__16277;
    wire N__16274;
    wire N__16271;
    wire N__16268;
    wire N__16265;
    wire N__16262;
    wire N__16259;
    wire N__16258;
    wire N__16255;
    wire N__16252;
    wire N__16247;
    wire N__16244;
    wire N__16241;
    wire N__16238;
    wire N__16237;
    wire N__16234;
    wire N__16231;
    wire N__16230;
    wire N__16227;
    wire N__16224;
    wire N__16221;
    wire N__16214;
    wire N__16211;
    wire N__16208;
    wire N__16205;
    wire N__16204;
    wire N__16203;
    wire N__16200;
    wire N__16197;
    wire N__16194;
    wire N__16191;
    wire N__16188;
    wire N__16181;
    wire N__16178;
    wire N__16175;
    wire N__16172;
    wire N__16169;
    wire N__16166;
    wire N__16165;
    wire N__16162;
    wire N__16159;
    wire N__16154;
    wire N__16151;
    wire N__16148;
    wire N__16145;
    wire N__16142;
    wire N__16139;
    wire N__16136;
    wire N__16135;
    wire N__16132;
    wire N__16129;
    wire N__16124;
    wire N__16121;
    wire N__16118;
    wire N__16115;
    wire N__16114;
    wire N__16111;
    wire N__16108;
    wire N__16107;
    wire N__16104;
    wire N__16101;
    wire N__16098;
    wire N__16091;
    wire N__16090;
    wire N__16087;
    wire N__16084;
    wire N__16083;
    wire N__16080;
    wire N__16077;
    wire N__16074;
    wire N__16067;
    wire N__16064;
    wire N__16061;
    wire N__16058;
    wire N__16055;
    wire N__16052;
    wire N__16051;
    wire N__16050;
    wire N__16047;
    wire N__16044;
    wire N__16041;
    wire N__16038;
    wire N__16035;
    wire N__16032;
    wire N__16025;
    wire N__16022;
    wire N__16021;
    wire N__16018;
    wire N__16015;
    wire N__16014;
    wire N__16011;
    wire N__16008;
    wire N__16005;
    wire N__15998;
    wire N__15995;
    wire N__15992;
    wire N__15989;
    wire N__15986;
    wire N__15983;
    wire N__15982;
    wire N__15979;
    wire N__15978;
    wire N__15977;
    wire N__15974;
    wire N__15973;
    wire N__15972;
    wire N__15967;
    wire N__15964;
    wire N__15963;
    wire N__15962;
    wire N__15961;
    wire N__15960;
    wire N__15959;
    wire N__15956;
    wire N__15951;
    wire N__15948;
    wire N__15941;
    wire N__15936;
    wire N__15935;
    wire N__15932;
    wire N__15931;
    wire N__15928;
    wire N__15925;
    wire N__15920;
    wire N__15917;
    wire N__15910;
    wire N__15899;
    wire N__15898;
    wire N__15897;
    wire N__15894;
    wire N__15891;
    wire N__15888;
    wire N__15885;
    wire N__15878;
    wire N__15875;
    wire N__15872;
    wire N__15869;
    wire N__15868;
    wire N__15865;
    wire N__15862;
    wire N__15859;
    wire N__15858;
    wire N__15855;
    wire N__15852;
    wire N__15849;
    wire N__15846;
    wire N__15839;
    wire N__15836;
    wire N__15833;
    wire N__15830;
    wire N__15829;
    wire N__15826;
    wire N__15823;
    wire N__15820;
    wire N__15819;
    wire N__15816;
    wire N__15813;
    wire N__15810;
    wire N__15807;
    wire N__15804;
    wire N__15801;
    wire N__15794;
    wire N__15793;
    wire N__15790;
    wire N__15787;
    wire N__15784;
    wire N__15781;
    wire N__15780;
    wire N__15777;
    wire N__15774;
    wire N__15771;
    wire N__15768;
    wire N__15761;
    wire N__15758;
    wire N__15755;
    wire N__15752;
    wire N__15751;
    wire N__15750;
    wire N__15747;
    wire N__15744;
    wire N__15741;
    wire N__15738;
    wire N__15731;
    wire N__15728;
    wire N__15727;
    wire N__15724;
    wire N__15721;
    wire N__15718;
    wire N__15717;
    wire N__15712;
    wire N__15709;
    wire N__15706;
    wire N__15701;
    wire N__15698;
    wire N__15695;
    wire N__15692;
    wire N__15689;
    wire N__15686;
    wire N__15685;
    wire N__15684;
    wire N__15681;
    wire N__15678;
    wire N__15675;
    wire N__15668;
    wire N__15665;
    wire N__15662;
    wire N__15659;
    wire N__15656;
    wire N__15653;
    wire N__15652;
    wire N__15649;
    wire N__15646;
    wire N__15643;
    wire N__15640;
    wire N__15635;
    wire N__15632;
    wire N__15629;
    wire N__15626;
    wire N__15623;
    wire N__15620;
    wire N__15617;
    wire N__15616;
    wire N__15613;
    wire N__15610;
    wire N__15609;
    wire N__15606;
    wire N__15603;
    wire N__15600;
    wire N__15597;
    wire N__15594;
    wire N__15587;
    wire N__15584;
    wire N__15583;
    wire N__15580;
    wire N__15579;
    wire N__15576;
    wire N__15573;
    wire N__15570;
    wire N__15565;
    wire N__15560;
    wire N__15557;
    wire N__15554;
    wire N__15551;
    wire N__15548;
    wire N__15547;
    wire N__15544;
    wire N__15541;
    wire N__15538;
    wire N__15537;
    wire N__15534;
    wire N__15531;
    wire N__15528;
    wire N__15521;
    wire N__15520;
    wire N__15519;
    wire N__15518;
    wire N__15517;
    wire N__15514;
    wire N__15513;
    wire N__15512;
    wire N__15509;
    wire N__15506;
    wire N__15505;
    wire N__15504;
    wire N__15501;
    wire N__15500;
    wire N__15499;
    wire N__15498;
    wire N__15495;
    wire N__15494;
    wire N__15489;
    wire N__15484;
    wire N__15479;
    wire N__15472;
    wire N__15469;
    wire N__15462;
    wire N__15457;
    wire N__15446;
    wire N__15443;
    wire N__15440;
    wire N__15437;
    wire N__15434;
    wire N__15431;
    wire N__15430;
    wire N__15427;
    wire N__15424;
    wire N__15419;
    wire N__15418;
    wire N__15415;
    wire N__15412;
    wire N__15409;
    wire N__15406;
    wire N__15401;
    wire N__15398;
    wire N__15395;
    wire N__15392;
    wire N__15389;
    wire N__15386;
    wire N__15383;
    wire N__15380;
    wire N__15377;
    wire N__15374;
    wire N__15371;
    wire N__15370;
    wire N__15369;
    wire N__15366;
    wire N__15363;
    wire N__15360;
    wire N__15357;
    wire N__15354;
    wire N__15347;
    wire N__15344;
    wire N__15341;
    wire N__15338;
    wire N__15335;
    wire N__15334;
    wire N__15331;
    wire N__15328;
    wire N__15327;
    wire N__15324;
    wire N__15321;
    wire N__15318;
    wire N__15315;
    wire N__15312;
    wire N__15309;
    wire N__15306;
    wire N__15301;
    wire N__15296;
    wire N__15293;
    wire N__15290;
    wire N__15287;
    wire N__15284;
    wire N__15283;
    wire N__15280;
    wire N__15277;
    wire N__15276;
    wire N__15273;
    wire N__15270;
    wire N__15267;
    wire N__15262;
    wire N__15259;
    wire N__15256;
    wire N__15253;
    wire N__15250;
    wire N__15247;
    wire N__15242;
    wire N__15239;
    wire N__15236;
    wire N__15233;
    wire N__15230;
    wire N__15227;
    wire N__15224;
    wire N__15223;
    wire N__15220;
    wire N__15217;
    wire N__15214;
    wire N__15211;
    wire N__15206;
    wire N__15203;
    wire N__15200;
    wire N__15197;
    wire N__15194;
    wire N__15191;
    wire N__15188;
    wire N__15187;
    wire N__15184;
    wire N__15181;
    wire N__15180;
    wire N__15175;
    wire N__15172;
    wire N__15169;
    wire N__15164;
    wire N__15161;
    wire N__15158;
    wire N__15155;
    wire N__15152;
    wire N__15149;
    wire N__15148;
    wire N__15145;
    wire N__15144;
    wire N__15141;
    wire N__15138;
    wire N__15135;
    wire N__15132;
    wire N__15125;
    wire N__15122;
    wire N__15119;
    wire N__15116;
    wire N__15113;
    wire N__15112;
    wire N__15109;
    wire N__15106;
    wire N__15103;
    wire N__15100;
    wire N__15097;
    wire N__15096;
    wire N__15093;
    wire N__15090;
    wire N__15087;
    wire N__15080;
    wire N__15077;
    wire N__15074;
    wire N__15071;
    wire N__15068;
    wire N__15067;
    wire N__15064;
    wire N__15061;
    wire N__15058;
    wire N__15055;
    wire N__15052;
    wire N__15051;
    wire N__15048;
    wire N__15045;
    wire N__15042;
    wire N__15035;
    wire N__15032;
    wire N__15029;
    wire N__15026;
    wire N__15023;
    wire N__15020;
    wire N__15019;
    wire N__15016;
    wire N__15013;
    wire N__15010;
    wire N__15007;
    wire N__15006;
    wire N__15003;
    wire N__15000;
    wire N__14997;
    wire N__14994;
    wire N__14991;
    wire N__14988;
    wire N__14981;
    wire N__14978;
    wire N__14975;
    wire N__14972;
    wire N__14969;
    wire N__14968;
    wire N__14965;
    wire N__14962;
    wire N__14959;
    wire N__14958;
    wire N__14955;
    wire N__14952;
    wire N__14949;
    wire N__14942;
    wire N__14939;
    wire N__14936;
    wire N__14933;
    wire N__14930;
    wire N__14927;
    wire N__14924;
    wire N__14921;
    wire N__14918;
    wire N__14915;
    wire N__14914;
    wire N__14911;
    wire N__14910;
    wire N__14907;
    wire N__14904;
    wire N__14901;
    wire N__14894;
    wire N__14891;
    wire N__14888;
    wire N__14885;
    wire N__14882;
    wire N__14879;
    wire N__14878;
    wire N__14875;
    wire N__14874;
    wire N__14871;
    wire N__14868;
    wire N__14865;
    wire N__14858;
    wire N__14855;
    wire N__14852;
    wire N__14849;
    wire N__14846;
    wire N__14843;
    wire N__14840;
    wire N__14837;
    wire N__14834;
    wire N__14831;
    wire N__14828;
    wire N__14825;
    wire N__14822;
    wire N__14819;
    wire N__14816;
    wire N__14813;
    wire N__14810;
    wire N__14807;
    wire N__14804;
    wire N__14801;
    wire N__14800;
    wire N__14799;
    wire N__14794;
    wire N__14791;
    wire N__14786;
    wire N__14783;
    wire N__14782;
    wire N__14781;
    wire N__14776;
    wire N__14773;
    wire N__14768;
    wire N__14765;
    wire N__14764;
    wire N__14761;
    wire N__14760;
    wire N__14755;
    wire N__14752;
    wire N__14747;
    wire N__14744;
    wire N__14743;
    wire N__14742;
    wire N__14737;
    wire N__14734;
    wire N__14729;
    wire N__14726;
    wire N__14723;
    wire N__14722;
    wire N__14719;
    wire N__14716;
    wire N__14711;
    wire N__14708;
    wire N__14705;
    wire N__14702;
    wire N__14699;
    wire N__14696;
    wire N__14693;
    wire N__14690;
    wire N__14687;
    wire N__14684;
    wire N__14681;
    wire N__14678;
    wire N__14675;
    wire N__14672;
    wire N__14669;
    wire N__14666;
    wire N__14663;
    wire N__14660;
    wire N__14657;
    wire N__14654;
    wire N__14651;
    wire N__14648;
    wire N__14645;
    wire N__14642;
    wire N__14639;
    wire N__14636;
    wire N__14633;
    wire N__14630;
    wire N__14627;
    wire N__14624;
    wire N__14621;
    wire N__14618;
    wire N__14615;
    wire N__14612;
    wire N__14609;
    wire N__14606;
    wire N__14603;
    wire N__14600;
    wire N__14597;
    wire N__14594;
    wire N__14591;
    wire N__14588;
    wire N__14585;
    wire N__14582;
    wire N__14579;
    wire N__14576;
    wire N__14573;
    wire N__14570;
    wire N__14567;
    wire N__14564;
    wire N__14561;
    wire N__14558;
    wire N__14557;
    wire N__14556;
    wire N__14553;
    wire N__14550;
    wire N__14547;
    wire N__14544;
    wire N__14541;
    wire N__14538;
    wire N__14531;
    wire N__14528;
    wire N__14525;
    wire N__14522;
    wire N__14519;
    wire N__14516;
    wire N__14515;
    wire N__14512;
    wire N__14509;
    wire N__14506;
    wire N__14503;
    wire N__14500;
    wire N__14497;
    wire N__14492;
    wire N__14489;
    wire N__14486;
    wire N__14483;
    wire N__14480;
    wire N__14479;
    wire N__14478;
    wire N__14475;
    wire N__14470;
    wire N__14467;
    wire N__14462;
    wire N__14459;
    wire N__14456;
    wire N__14453;
    wire N__14450;
    wire N__14447;
    wire N__14444;
    wire N__14441;
    wire N__14440;
    wire N__14437;
    wire N__14436;
    wire N__14433;
    wire N__14430;
    wire N__14427;
    wire N__14424;
    wire N__14419;
    wire N__14414;
    wire N__14411;
    wire N__14408;
    wire N__14405;
    wire N__14402;
    wire N__14399;
    wire N__14398;
    wire N__14395;
    wire N__14392;
    wire N__14387;
    wire N__14384;
    wire N__14381;
    wire N__14378;
    wire N__14375;
    wire N__14372;
    wire N__14369;
    wire N__14366;
    wire N__14363;
    wire N__14360;
    wire N__14357;
    wire N__14354;
    wire N__14351;
    wire N__14348;
    wire N__14345;
    wire N__14344;
    wire N__14343;
    wire N__14340;
    wire N__14335;
    wire N__14332;
    wire N__14327;
    wire N__14324;
    wire N__14321;
    wire N__14318;
    wire N__14315;
    wire N__14314;
    wire N__14311;
    wire N__14308;
    wire N__14305;
    wire N__14302;
    wire N__14299;
    wire N__14296;
    wire N__14295;
    wire N__14290;
    wire N__14287;
    wire N__14282;
    wire N__14279;
    wire N__14276;
    wire N__14273;
    wire N__14272;
    wire N__14269;
    wire N__14266;
    wire N__14263;
    wire N__14262;
    wire N__14257;
    wire N__14254;
    wire N__14249;
    wire N__14246;
    wire N__14245;
    wire N__14242;
    wire N__14239;
    wire N__14234;
    wire N__14231;
    wire N__14228;
    wire N__14225;
    wire N__14224;
    wire N__14221;
    wire N__14218;
    wire N__14215;
    wire N__14210;
    wire N__14207;
    wire N__14204;
    wire N__14201;
    wire N__14198;
    wire N__14195;
    wire N__14192;
    wire N__14189;
    wire N__14186;
    wire N__14185;
    wire N__14182;
    wire N__14179;
    wire N__14178;
    wire N__14175;
    wire N__14172;
    wire N__14169;
    wire N__14164;
    wire N__14159;
    wire N__14156;
    wire N__14155;
    wire N__14152;
    wire N__14149;
    wire N__14146;
    wire N__14145;
    wire N__14142;
    wire N__14139;
    wire N__14136;
    wire N__14129;
    wire N__14128;
    wire N__14127;
    wire N__14124;
    wire N__14121;
    wire N__14118;
    wire N__14115;
    wire N__14112;
    wire N__14109;
    wire N__14104;
    wire N__14099;
    wire N__14096;
    wire N__14093;
    wire N__14090;
    wire N__14087;
    wire N__14084;
    wire N__14081;
    wire N__14078;
    wire N__14075;
    wire N__14072;
    wire N__14069;
    wire N__14068;
    wire N__14065;
    wire N__14064;
    wire N__14061;
    wire N__14058;
    wire N__14055;
    wire N__14052;
    wire N__14045;
    wire N__14042;
    wire N__14039;
    wire N__14036;
    wire N__14035;
    wire N__14034;
    wire N__14031;
    wire N__14028;
    wire N__14025;
    wire N__14022;
    wire N__14019;
    wire N__14012;
    wire N__14011;
    wire N__14008;
    wire N__14005;
    wire N__14004;
    wire N__14001;
    wire N__13998;
    wire N__13995;
    wire N__13988;
    wire N__13985;
    wire N__13982;
    wire N__13979;
    wire N__13978;
    wire N__13975;
    wire N__13974;
    wire N__13971;
    wire N__13968;
    wire N__13965;
    wire N__13958;
    wire N__13955;
    wire N__13952;
    wire N__13951;
    wire N__13950;
    wire N__13949;
    wire N__13946;
    wire N__13943;
    wire N__13940;
    wire N__13939;
    wire N__13938;
    wire N__13937;
    wire N__13936;
    wire N__13935;
    wire N__13932;
    wire N__13931;
    wire N__13928;
    wire N__13917;
    wire N__13908;
    wire N__13901;
    wire N__13898;
    wire N__13897;
    wire N__13894;
    wire N__13891;
    wire N__13886;
    wire N__13885;
    wire N__13884;
    wire N__13881;
    wire N__13878;
    wire N__13875;
    wire N__13872;
    wire N__13869;
    wire N__13862;
    wire N__13859;
    wire N__13856;
    wire N__13853;
    wire N__13850;
    wire N__13847;
    wire N__13844;
    wire N__13843;
    wire N__13840;
    wire N__13837;
    wire N__13834;
    wire N__13831;
    wire N__13826;
    wire N__13823;
    wire N__13820;
    wire N__13817;
    wire N__13814;
    wire N__13813;
    wire N__13810;
    wire N__13807;
    wire N__13804;
    wire N__13801;
    wire N__13796;
    wire N__13793;
    wire N__13792;
    wire N__13791;
    wire N__13788;
    wire N__13785;
    wire N__13782;
    wire N__13777;
    wire N__13772;
    wire N__13769;
    wire N__13766;
    wire N__13763;
    wire N__13760;
    wire N__13757;
    wire N__13756;
    wire N__13753;
    wire N__13750;
    wire N__13747;
    wire N__13744;
    wire N__13743;
    wire N__13738;
    wire N__13735;
    wire N__13730;
    wire N__13727;
    wire N__13724;
    wire N__13721;
    wire N__13720;
    wire N__13719;
    wire N__13716;
    wire N__13713;
    wire N__13710;
    wire N__13705;
    wire N__13702;
    wire N__13699;
    wire N__13694;
    wire N__13691;
    wire N__13688;
    wire N__13685;
    wire N__13682;
    wire N__13679;
    wire N__13678;
    wire N__13675;
    wire N__13674;
    wire N__13671;
    wire N__13668;
    wire N__13665;
    wire N__13658;
    wire N__13655;
    wire N__13652;
    wire N__13649;
    wire N__13646;
    wire N__13643;
    wire N__13640;
    wire N__13637;
    wire N__13636;
    wire N__13633;
    wire N__13632;
    wire N__13629;
    wire N__13626;
    wire N__13623;
    wire N__13616;
    wire N__13613;
    wire N__13610;
    wire N__13607;
    wire N__13604;
    wire N__13601;
    wire N__13598;
    wire N__13595;
    wire N__13592;
    wire N__13589;
    wire N__13586;
    wire N__13585;
    wire N__13584;
    wire N__13581;
    wire N__13578;
    wire N__13575;
    wire N__13570;
    wire N__13565;
    wire N__13562;
    wire N__13559;
    wire N__13556;
    wire N__13553;
    wire N__13550;
    wire N__13547;
    wire N__13544;
    wire N__13541;
    wire N__13538;
    wire N__13535;
    wire N__13532;
    wire N__13531;
    wire N__13528;
    wire N__13525;
    wire N__13520;
    wire N__13517;
    wire N__13514;
    wire N__13511;
    wire N__13508;
    wire N__13505;
    wire N__13502;
    wire N__13499;
    wire N__13496;
    wire N__13493;
    wire N__13490;
    wire N__13487;
    wire N__13484;
    wire N__13481;
    wire N__13478;
    wire N__13475;
    wire N__13474;
    wire N__13471;
    wire N__13470;
    wire N__13467;
    wire N__13464;
    wire N__13461;
    wire N__13454;
    wire N__13451;
    wire N__13448;
    wire N__13445;
    wire N__13442;
    wire N__13439;
    wire N__13436;
    wire N__13433;
    wire N__13430;
    wire N__13429;
    wire N__13426;
    wire N__13423;
    wire N__13418;
    wire N__13415;
    wire N__13414;
    wire N__13413;
    wire N__13408;
    wire N__13405;
    wire N__13400;
    wire N__13397;
    wire N__13394;
    wire N__13391;
    wire N__13388;
    wire N__13385;
    wire N__13382;
    wire N__13381;
    wire N__13376;
    wire N__13375;
    wire N__13372;
    wire N__13369;
    wire N__13364;
    wire N__13361;
    wire N__13360;
    wire N__13359;
    wire N__13356;
    wire N__13351;
    wire N__13348;
    wire N__13343;
    wire N__13340;
    wire N__13337;
    wire N__13334;
    wire N__13331;
    wire N__13328;
    wire N__13325;
    wire N__13324;
    wire N__13321;
    wire N__13320;
    wire N__13317;
    wire N__13314;
    wire N__13311;
    wire N__13304;
    wire N__13301;
    wire N__13298;
    wire N__13295;
    wire N__13292;
    wire N__13289;
    wire N__13288;
    wire N__13285;
    wire N__13284;
    wire N__13281;
    wire N__13278;
    wire N__13273;
    wire N__13268;
    wire N__13265;
    wire N__13262;
    wire N__13259;
    wire N__13256;
    wire N__13255;
    wire N__13254;
    wire N__13251;
    wire N__13248;
    wire N__13245;
    wire N__13242;
    wire N__13239;
    wire N__13232;
    wire N__13229;
    wire N__13226;
    wire N__13223;
    wire N__13220;
    wire N__13217;
    wire N__13216;
    wire N__13213;
    wire N__13210;
    wire N__13209;
    wire N__13206;
    wire N__13201;
    wire N__13196;
    wire N__13193;
    wire N__13190;
    wire N__13187;
    wire N__13184;
    wire N__13181;
    wire N__13178;
    wire N__13175;
    wire N__13172;
    wire N__13171;
    wire N__13168;
    wire N__13165;
    wire N__13160;
    wire N__13157;
    wire N__13154;
    wire N__13151;
    wire N__13148;
    wire N__13145;
    wire N__13142;
    wire N__13139;
    wire N__13136;
    wire N__13133;
    wire N__13130;
    wire N__13127;
    wire N__13124;
    wire N__13121;
    wire N__13118;
    wire N__13117;
    wire N__13116;
    wire N__13115;
    wire N__13114;
    wire N__13113;
    wire N__13110;
    wire N__13107;
    wire N__13104;
    wire N__13103;
    wire N__13102;
    wire N__13101;
    wire N__13100;
    wire N__13097;
    wire N__13094;
    wire N__13091;
    wire N__13090;
    wire N__13087;
    wire N__13076;
    wire N__13073;
    wire N__13064;
    wire N__13055;
    wire N__13052;
    wire N__13051;
    wire N__13050;
    wire N__13047;
    wire N__13044;
    wire N__13041;
    wire N__13036;
    wire N__13031;
    wire N__13028;
    wire N__13025;
    wire N__13022;
    wire N__13019;
    wire N__13016;
    wire N__13013;
    wire N__13010;
    wire N__13009;
    wire N__13006;
    wire N__13003;
    wire N__12998;
    wire N__12995;
    wire N__12992;
    wire N__12989;
    wire N__12986;
    wire N__12983;
    wire N__12980;
    wire N__12977;
    wire N__12976;
    wire N__12975;
    wire N__12972;
    wire N__12969;
    wire N__12966;
    wire N__12959;
    wire N__12956;
    wire N__12953;
    wire N__12950;
    wire N__12947;
    wire N__12946;
    wire N__12943;
    wire N__12940;
    wire N__12937;
    wire N__12934;
    wire N__12929;
    wire N__12928;
    wire N__12927;
    wire N__12926;
    wire N__12923;
    wire N__12920;
    wire N__12917;
    wire N__12916;
    wire N__12915;
    wire N__12912;
    wire N__12911;
    wire N__12908;
    wire N__12899;
    wire N__12894;
    wire N__12887;
    wire N__12884;
    wire N__12881;
    wire N__12878;
    wire N__12875;
    wire N__12872;
    wire N__12869;
    wire N__12866;
    wire N__12863;
    wire N__12860;
    wire N__12857;
    wire N__12854;
    wire N__12851;
    wire N__12848;
    wire N__12845;
    wire N__12842;
    wire N__12839;
    wire N__12836;
    wire N__12833;
    wire N__12832;
    wire N__12829;
    wire N__12828;
    wire N__12825;
    wire N__12822;
    wire N__12819;
    wire N__12812;
    wire N__12809;
    wire N__12806;
    wire N__12803;
    wire N__12800;
    wire N__12797;
    wire N__12794;
    wire N__12793;
    wire N__12792;
    wire N__12789;
    wire N__12784;
    wire N__12781;
    wire N__12776;
    wire N__12773;
    wire N__12770;
    wire N__12767;
    wire N__12766;
    wire N__12765;
    wire N__12762;
    wire N__12759;
    wire N__12756;
    wire N__12753;
    wire N__12746;
    wire N__12743;
    wire N__12742;
    wire N__12739;
    wire N__12736;
    wire N__12733;
    wire N__12728;
    wire N__12727;
    wire N__12726;
    wire N__12723;
    wire N__12720;
    wire N__12715;
    wire N__12712;
    wire N__12709;
    wire N__12704;
    wire N__12701;
    wire N__12698;
    wire N__12695;
    wire N__12692;
    wire N__12689;
    wire N__12686;
    wire N__12685;
    wire N__12682;
    wire N__12681;
    wire N__12678;
    wire N__12675;
    wire N__12672;
    wire N__12665;
    wire N__12662;
    wire N__12661;
    wire N__12660;
    wire N__12657;
    wire N__12654;
    wire N__12651;
    wire N__12648;
    wire N__12645;
    wire N__12638;
    wire N__12635;
    wire N__12632;
    wire N__12629;
    wire N__12626;
    wire N__12623;
    wire N__12620;
    wire N__12617;
    wire N__12616;
    wire N__12611;
    wire N__12608;
    wire N__12607;
    wire N__12606;
    wire N__12605;
    wire N__12602;
    wire N__12601;
    wire N__12600;
    wire N__12599;
    wire N__12598;
    wire N__12595;
    wire N__12590;
    wire N__12587;
    wire N__12578;
    wire N__12575;
    wire N__12566;
    wire N__12563;
    wire N__12560;
    wire N__12557;
    wire N__12554;
    wire N__12551;
    wire N__12548;
    wire N__12545;
    wire N__12542;
    wire N__12539;
    wire N__12536;
    wire N__12533;
    wire N__12530;
    wire N__12527;
    wire N__12524;
    wire N__12521;
    wire N__12518;
    wire N__12515;
    wire N__12512;
    wire N__12511;
    wire N__12508;
    wire N__12507;
    wire N__12504;
    wire N__12501;
    wire N__12498;
    wire N__12491;
    wire N__12488;
    wire N__12487;
    wire N__12484;
    wire N__12481;
    wire N__12478;
    wire N__12473;
    wire N__12472;
    wire N__12471;
    wire N__12470;
    wire N__12467;
    wire N__12466;
    wire N__12463;
    wire N__12460;
    wire N__12459;
    wire N__12456;
    wire N__12453;
    wire N__12450;
    wire N__12443;
    wire N__12434;
    wire N__12431;
    wire N__12428;
    wire N__12425;
    wire N__12422;
    wire N__12419;
    wire N__12416;
    wire N__12413;
    wire N__12410;
    wire N__12407;
    wire N__12404;
    wire N__12401;
    wire N__12398;
    wire N__12397;
    wire N__12394;
    wire N__12393;
    wire N__12390;
    wire N__12387;
    wire N__12384;
    wire N__12377;
    wire N__12374;
    wire N__12371;
    wire N__12368;
    wire N__12365;
    wire N__12362;
    wire N__12359;
    wire N__12356;
    wire N__12353;
    wire N__12350;
    wire N__12347;
    wire N__12344;
    wire N__12341;
    wire N__12338;
    wire N__12335;
    wire N__12334;
    wire N__12331;
    wire N__12330;
    wire N__12327;
    wire N__12324;
    wire N__12321;
    wire N__12314;
    wire N__12311;
    wire N__12308;
    wire N__12307;
    wire N__12306;
    wire N__12303;
    wire N__12300;
    wire N__12297;
    wire N__12292;
    wire N__12287;
    wire N__12284;
    wire N__12281;
    wire N__12278;
    wire N__12275;
    wire N__12272;
    wire N__12271;
    wire N__12268;
    wire N__12267;
    wire N__12264;
    wire N__12261;
    wire N__12258;
    wire N__12251;
    wire N__12248;
    wire N__12245;
    wire N__12242;
    wire N__12239;
    wire N__12236;
    wire N__12233;
    wire N__12230;
    wire N__12229;
    wire N__12228;
    wire N__12225;
    wire N__12222;
    wire N__12219;
    wire N__12216;
    wire N__12209;
    wire N__12206;
    wire N__12205;
    wire N__12202;
    wire N__12199;
    wire N__12194;
    wire N__12191;
    wire N__12188;
    wire N__12187;
    wire N__12184;
    wire N__12181;
    wire N__12178;
    wire N__12175;
    wire N__12172;
    wire N__12167;
    wire N__12166;
    wire N__12165;
    wire N__12162;
    wire N__12159;
    wire N__12156;
    wire N__12149;
    wire N__12146;
    wire N__12143;
    wire N__12140;
    wire N__12137;
    wire N__12134;
    wire N__12131;
    wire N__12130;
    wire N__12127;
    wire N__12124;
    wire N__12119;
    wire N__12116;
    wire N__12113;
    wire N__12110;
    wire N__12107;
    wire N__12104;
    wire N__12101;
    wire N__12098;
    wire N__12095;
    wire N__12094;
    wire N__12091;
    wire N__12090;
    wire N__12087;
    wire N__12084;
    wire N__12081;
    wire N__12074;
    wire N__12071;
    wire N__12068;
    wire N__12065;
    wire N__12062;
    wire N__12059;
    wire N__12056;
    wire N__12053;
    wire N__12050;
    wire N__12047;
    wire N__12044;
    wire N__12043;
    wire N__12040;
    wire N__12037;
    wire N__12034;
    wire N__12031;
    wire N__12028;
    wire N__12025;
    wire N__12020;
    wire N__12017;
    wire N__12014;
    wire N__12011;
    wire N__12008;
    wire N__12005;
    wire N__12004;
    wire N__12001;
    wire N__11998;
    wire N__11995;
    wire N__11990;
    wire N__11987;
    wire N__11984;
    wire N__11983;
    wire N__11982;
    wire N__11979;
    wire N__11976;
    wire N__11973;
    wire N__11970;
    wire N__11967;
    wire N__11960;
    wire N__11957;
    wire N__11954;
    wire N__11951;
    wire N__11948;
    wire N__11945;
    wire N__11942;
    wire N__11939;
    wire N__11936;
    wire N__11935;
    wire N__11930;
    wire N__11927;
    wire N__11924;
    wire N__11921;
    wire N__11920;
    wire N__11919;
    wire N__11916;
    wire N__11913;
    wire N__11910;
    wire N__11903;
    wire N__11902;
    wire N__11899;
    wire N__11896;
    wire N__11893;
    wire N__11888;
    wire N__11885;
    wire N__11882;
    wire N__11879;
    wire N__11876;
    wire N__11873;
    wire N__11870;
    wire N__11867;
    wire N__11864;
    wire N__11863;
    wire N__11862;
    wire N__11859;
    wire N__11856;
    wire N__11851;
    wire N__11846;
    wire N__11843;
    wire N__11840;
    wire N__11837;
    wire N__11834;
    wire N__11831;
    wire N__11828;
    wire N__11825;
    wire N__11822;
    wire N__11819;
    wire N__11816;
    wire N__11813;
    wire N__11812;
    wire N__11809;
    wire N__11808;
    wire N__11805;
    wire N__11802;
    wire N__11799;
    wire N__11792;
    wire N__11789;
    wire N__11786;
    wire N__11783;
    wire N__11780;
    wire N__11777;
    wire N__11774;
    wire N__11771;
    wire N__11768;
    wire N__11765;
    wire N__11762;
    wire N__11759;
    wire N__11756;
    wire N__11753;
    wire N__11750;
    wire N__11747;
    wire N__11744;
    wire N__11741;
    wire N__11738;
    wire N__11735;
    wire N__11732;
    wire N__11731;
    wire N__11728;
    wire N__11727;
    wire N__11724;
    wire N__11721;
    wire N__11718;
    wire N__11711;
    wire N__11708;
    wire N__11705;
    wire N__11702;
    wire N__11699;
    wire N__11696;
    wire N__11693;
    wire N__11690;
    wire N__11687;
    wire N__11684;
    wire N__11681;
    wire N__11678;
    wire N__11675;
    wire N__11672;
    wire N__11669;
    wire N__11666;
    wire N__11663;
    wire N__11660;
    wire N__11657;
    wire N__11654;
    wire N__11651;
    wire N__11648;
    wire N__11645;
    wire N__11642;
    wire N__11639;
    wire N__11636;
    wire N__11633;
    wire N__11630;
    wire N__11627;
    wire N__11624;
    wire N__11621;
    wire N__11618;
    wire N__11615;
    wire N__11612;
    wire N__11609;
    wire N__11606;
    wire N__11603;
    wire N__11600;
    wire N__11597;
    wire N__11594;
    wire N__11591;
    wire N__11588;
    wire N__11585;
    wire N__11582;
    wire N__11579;
    wire N__11576;
    wire N__11573;
    wire N__11570;
    wire N__11567;
    wire N__11564;
    wire N__11561;
    wire N__11558;
    wire N__11555;
    wire N__11552;
    wire N__11549;
    wire N__11546;
    wire N__11543;
    wire N__11540;
    wire N__11537;
    wire N__11536;
    wire N__11535;
    wire N__11532;
    wire N__11529;
    wire N__11526;
    wire N__11521;
    wire N__11516;
    wire N__11513;
    wire N__11510;
    wire N__11507;
    wire N__11504;
    wire N__11501;
    wire N__11498;
    wire N__11495;
    wire N__11492;
    wire N__11489;
    wire N__11486;
    wire N__11483;
    wire N__11480;
    wire N__11477;
    wire N__11474;
    wire N__11471;
    wire N__11468;
    wire N__11465;
    wire N__11462;
    wire N__11459;
    wire N__11456;
    wire N__11453;
    wire N__11450;
    wire N__11447;
    wire N__11444;
    wire N__11441;
    wire N__11438;
    wire N__11435;
    wire N__11432;
    wire N__11429;
    wire N__11426;
    wire N__11423;
    wire N__11420;
    wire N__11417;
    wire N__11414;
    wire N__11411;
    wire N__11408;
    wire N__11405;
    wire N__11402;
    wire N__11399;
    wire N__11396;
    wire N__11393;
    wire N__11390;
    wire N__11387;
    wire N__11384;
    wire N__11381;
    wire N__11378;
    wire N__11375;
    wire N__11372;
    wire N__11369;
    wire N__11366;
    wire N__11363;
    wire N__11360;
    wire N__11357;
    wire N__11354;
    wire N__11351;
    wire N__11348;
    wire N__11345;
    wire N__11342;
    wire N__11339;
    wire N__11336;
    wire N__11333;
    wire N__11330;
    wire N__11327;
    wire N__11324;
    wire N__11321;
    wire N__11318;
    wire N__11315;
    wire N__11312;
    wire N__11309;
    wire N__11306;
    wire N__11303;
    wire N__11300;
    wire N__11297;
    wire N__11294;
    wire N__11291;
    wire N__11288;
    wire N__11285;
    wire N__11282;
    wire N__11279;
    wire N__11276;
    wire N__11273;
    wire N__11270;
    wire N__11267;
    wire N__11264;
    wire N__11261;
    wire N__11258;
    wire N__11255;
    wire N__11252;
    wire N__11249;
    wire N__11246;
    wire N__11243;
    wire N__11240;
    wire N__11237;
    wire N__11234;
    wire N__11231;
    wire N__11230;
    wire N__11227;
    wire N__11226;
    wire N__11223;
    wire N__11220;
    wire N__11217;
    wire N__11212;
    wire N__11207;
    wire N__11204;
    wire N__11201;
    wire N__11198;
    wire N__11197;
    wire N__11192;
    wire N__11191;
    wire N__11188;
    wire N__11185;
    wire N__11182;
    wire N__11177;
    wire N__11174;
    wire N__11171;
    wire N__11168;
    wire N__11165;
    wire N__11162;
    wire N__11159;
    wire N__11156;
    wire N__11153;
    wire N__11150;
    wire N__11147;
    wire N__11144;
    wire N__11141;
    wire N__11138;
    wire N__11137;
    wire N__11136;
    wire N__11133;
    wire N__11128;
    wire N__11123;
    wire N__11120;
    wire N__11117;
    wire N__11114;
    wire N__11111;
    wire N__11108;
    wire N__11105;
    wire N__11102;
    wire N__11099;
    wire N__11096;
    wire CLK_pad_gb_input;
    wire VCCG0;
    wire GNDG0;
    wire bfn_2_17_0_;
    wire \eeprom.n3454 ;
    wire \eeprom.n3455 ;
    wire \eeprom.n3456 ;
    wire \eeprom.n3457 ;
    wire \eeprom.n3458 ;
    wire \eeprom.n3459 ;
    wire \eeprom.n3460 ;
    wire \eeprom.n3461 ;
    wire bfn_2_18_0_;
    wire \eeprom.n3462 ;
    wire \eeprom.n3463 ;
    wire \eeprom.delay_counter_11 ;
    wire \eeprom.n3464 ;
    wire \eeprom.n3465 ;
    wire \eeprom.delay_counter_13 ;
    wire \eeprom.n3466 ;
    wire \eeprom.n3467 ;
    wire \eeprom.n3468 ;
    wire \eeprom.n3469 ;
    wire \eeprom.delay_counter_16 ;
    wire bfn_2_19_0_;
    wire \eeprom.n3470 ;
    wire \eeprom.n3471 ;
    wire \eeprom.n3472 ;
    wire \eeprom.n3473 ;
    wire \eeprom.n3474 ;
    wire \eeprom.n3475 ;
    wire \eeprom.n3476 ;
    wire \eeprom.n3477 ;
    wire bfn_2_20_0_;
    wire \eeprom.n3478 ;
    wire \eeprom.n3479 ;
    wire \eeprom.n3480 ;
    wire \eeprom.n3481 ;
    wire \eeprom.n3482 ;
    wire \eeprom.n3483 ;
    wire \eeprom.n3484 ;
    wire bfn_2_21_0_;
    wire \eeprom.n3786 ;
    wire \eeprom.n31_adj_457 ;
    wire \eeprom.n3787 ;
    wire \eeprom.n3788 ;
    wire \eeprom.n3789 ;
    wire \eeprom.n28_adj_461 ;
    wire \eeprom.n3790 ;
    wire \eeprom.n27_adj_462 ;
    wire \eeprom.n3791 ;
    wire \eeprom.n3792 ;
    wire \eeprom.n3793 ;
    wire bfn_2_22_0_;
    wire \eeprom.n24_adj_463 ;
    wire \eeprom.n3794 ;
    wire \eeprom.n23 ;
    wire \eeprom.n3795 ;
    wire \eeprom.n22_adj_448 ;
    wire \eeprom.n22_adj_447 ;
    wire \eeprom.n3796 ;
    wire \eeprom.n21_adj_440 ;
    wire \eeprom.n3797 ;
    wire \eeprom.n20_adj_431 ;
    wire \eeprom.n20_adj_430 ;
    wire \eeprom.n3798 ;
    wire \eeprom.n3799 ;
    wire \eeprom.n18_adj_427 ;
    wire \eeprom.n3800 ;
    wire \eeprom.n3801 ;
    wire \eeprom.n17_adj_425 ;
    wire \eeprom.n17 ;
    wire bfn_2_23_0_;
    wire \eeprom.n16_adj_424 ;
    wire \eeprom.n3802 ;
    wire \eeprom.n3803 ;
    wire \eeprom.n14_adj_413 ;
    wire \eeprom.n3804 ;
    wire \eeprom.n3805 ;
    wire \eeprom.n3806 ;
    wire \eeprom.n3807 ;
    wire \eeprom.n3808 ;
    wire \eeprom.n3809 ;
    wire bfn_2_24_0_;
    wire \eeprom.n8_adj_407 ;
    wire \eeprom.n3810 ;
    wire \eeprom.n7_adj_405 ;
    wire \eeprom.n3811 ;
    wire \eeprom.n6_adj_403 ;
    wire \eeprom.n3812 ;
    wire \eeprom.n3813 ;
    wire \eeprom.n4_adj_397 ;
    wire \eeprom.n3814 ;
    wire \eeprom.n3_adj_396 ;
    wire \eeprom.n3815 ;
    wire \eeprom.n3816 ;
    wire \eeprom.n14 ;
    wire \eeprom.delay_counter_19 ;
    wire \eeprom.n11_adj_410 ;
    wire bfn_3_17_0_;
    wire \eeprom.n3448 ;
    wire \eeprom.n3449 ;
    wire \eeprom.n3450 ;
    wire \eeprom.n3451 ;
    wire \eeprom.n3452 ;
    wire \eeprom.n3453 ;
    wire \eeprom.n30_adj_458 ;
    wire \eeprom.n26 ;
    wire \eeprom.delay_counter_30 ;
    wire \eeprom.n3 ;
    wire \eeprom.n1341 ;
    wire \eeprom.n1256_cascade_ ;
    wire \eeprom.n5_adj_400 ;
    wire \eeprom.n15_adj_415 ;
    wire \eeprom.n33 ;
    wire \eeprom.delay_counter_25 ;
    wire \eeprom.n8 ;
    wire \eeprom.n1141_cascade_ ;
    wire \eeprom.n2_adj_395 ;
    wire \eeprom.n4399_cascade_ ;
    wire \eeprom.n1343 ;
    wire \eeprom.n1141 ;
    wire \eeprom.n4405_cascade_ ;
    wire \eeprom.delay_counter_28 ;
    wire \eeprom.n5 ;
    wire \eeprom.n1342 ;
    wire \eeprom.n6_adj_402 ;
    wire \eeprom.delay_counter_27 ;
    wire \eeprom.n1139 ;
    wire \eeprom.n25 ;
    wire \eeprom.n9 ;
    wire \eeprom.delay_counter_24 ;
    wire \eeprom.n9_adj_408 ;
    wire \eeprom.n32 ;
    wire \eeprom.delay_counter_26 ;
    wire \eeprom.n7 ;
    wire \eeprom.n1140 ;
    wire \eeprom.delay_counter_29 ;
    wire \eeprom.n4 ;
    wire \eeprom.n1137 ;
    wire \eeprom.n1339 ;
    wire \eeprom.n1137_cascade_ ;
    wire \eeprom.n24_adj_467 ;
    wire \eeprom.delay_counter_9 ;
    wire \eeprom.n33_adj_483 ;
    wire \eeprom.n13_adj_412 ;
    wire \eeprom.n10_adj_409 ;
    wire \eeprom.n19_adj_428 ;
    wire \eeprom.delay_counter_18 ;
    wire \eeprom.n15_adj_414 ;
    wire \eeprom.delay_counter_23 ;
    wire \eeprom.n10 ;
    wire \eeprom.n18_adj_426 ;
    wire \eeprom.delay_counter_15 ;
    wire bfn_3_23_0_;
    wire \eeprom.n3551 ;
    wire \eeprom.n3552 ;
    wire \eeprom.n2383 ;
    wire \eeprom.n3553 ;
    wire \eeprom.n3554 ;
    wire \eeprom.n3555 ;
    wire \eeprom.n3556 ;
    wire \eeprom.n3557 ;
    wire \eeprom.n3558 ;
    wire bfn_3_24_0_;
    wire \eeprom.n3559 ;
    wire \eeprom.n3560 ;
    wire \eeprom.n3561 ;
    wire \eeprom.n2386 ;
    wire \eeprom.n2381 ;
    wire \eeprom.n2384 ;
    wire \eeprom.n2378 ;
    wire \eeprom.n4733 ;
    wire \eeprom.n1340 ;
    wire \eeprom.n1138 ;
    wire \eeprom.n1915_cascade_ ;
    wire \eeprom.n1135 ;
    wire \eeprom.n4405 ;
    wire \eeprom.n1337 ;
    wire \eeprom.n12_adj_411 ;
    wire \eeprom.n25_adj_471 ;
    wire \eeprom.delay_counter_8 ;
    wire \eeprom.delay_counter_17 ;
    wire \eeprom.n16_adj_377 ;
    wire \eeprom.n4734 ;
    wire \eeprom.n1256 ;
    wire bfn_4_19_0_;
    wire \eeprom.n3517 ;
    wire \eeprom.n3518 ;
    wire \eeprom.n3519 ;
    wire \eeprom.n3520 ;
    wire \eeprom.n3521 ;
    wire \eeprom.n3522 ;
    wire \eeprom.n3523 ;
    wire \eeprom.n26_adj_469 ;
    wire \eeprom.delay_counter_7 ;
    wire \eeprom.n1984 ;
    wire \eeprom.n1985 ;
    wire \eeprom.n2017_cascade_ ;
    wire \eeprom.n1917 ;
    wire \eeprom.n4437 ;
    wire \eeprom.n1918 ;
    wire \eeprom.n4441_cascade_ ;
    wire \eeprom.n1912 ;
    wire \eeprom.n1916 ;
    wire \eeprom.n1945_cascade_ ;
    wire \eeprom.n1983 ;
    wire \eeprom.n1981 ;
    wire \eeprom.n1914 ;
    wire \eeprom.n1915 ;
    wire \eeprom.n1982 ;
    wire \eeprom.n2014_cascade_ ;
    wire \eeprom.n4415 ;
    wire \eeprom.n1919 ;
    wire \eeprom.n1986 ;
    wire \eeprom.n1913 ;
    wire \eeprom.n1945 ;
    wire \eeprom.n1980 ;
    wire \eeprom.n4419 ;
    wire \eeprom.n4575_cascade_ ;
    wire \eeprom.n4579 ;
    wire \eeprom.n13 ;
    wire \eeprom.delay_counter_20 ;
    wire \eeprom.n4479_cascade_ ;
    wire \eeprom.n4477 ;
    wire \eeprom.n2385 ;
    wire \eeprom.n2341_cascade_ ;
    wire \eeprom.n2376 ;
    wire \eeprom.n2312 ;
    wire \eeprom.n2312_cascade_ ;
    wire \eeprom.n2379 ;
    wire \eeprom.n2411_cascade_ ;
    wire \eeprom.n4133 ;
    wire \eeprom.n12_adj_472_cascade_ ;
    wire \eeprom.n2382 ;
    wire \eeprom.n2377 ;
    wire \eeprom.n2380 ;
    wire \eeprom.n2341 ;
    wire bfn_4_25_0_;
    wire \eeprom.n2418 ;
    wire \eeprom.n2485 ;
    wire \eeprom.n3562 ;
    wire \eeprom.n2417 ;
    wire \eeprom.n2484 ;
    wire \eeprom.n3563 ;
    wire \eeprom.n2416 ;
    wire \eeprom.n2483 ;
    wire \eeprom.n3564 ;
    wire \eeprom.n2415 ;
    wire \eeprom.n2482 ;
    wire \eeprom.n3565 ;
    wire \eeprom.n2414 ;
    wire \eeprom.n2481 ;
    wire \eeprom.n3566 ;
    wire \eeprom.n3567 ;
    wire \eeprom.n3568 ;
    wire \eeprom.n3569 ;
    wire bfn_4_26_0_;
    wire \eeprom.n3570 ;
    wire \eeprom.n3571 ;
    wire \eeprom.n3572 ;
    wire \eeprom.n2407 ;
    wire \eeprom.n3573 ;
    wire \eeprom.n2410 ;
    wire \eeprom.n2477 ;
    wire \eeprom.n2476 ;
    wire \eeprom.n2409 ;
    wire n4826;
    wire n4825_cascade_;
    wire LED_c;
    wire \eeprom.n23_adj_464 ;
    wire \eeprom.delay_counter_10 ;
    wire \eeprom.n2615_cascade_ ;
    wire \eeprom.n4497_cascade_ ;
    wire \eeprom.n4501_cascade_ ;
    wire \eeprom.n13_adj_474_cascade_ ;
    wire \eeprom.n11_adj_473 ;
    wire \eeprom.n2539_cascade_ ;
    wire \eeprom.delay_counter_14 ;
    wire \eeprom.n19_adj_429 ;
    wire \eeprom.n30 ;
    wire \eeprom.n2114_cascade_ ;
    wire \eeprom.n2411 ;
    wire \eeprom.n2478 ;
    wire \eeprom.n2419 ;
    wire \eeprom.n2486 ;
    wire bfn_5_22_0_;
    wire \eeprom.n2018 ;
    wire \eeprom.n2085 ;
    wire \eeprom.n3524 ;
    wire \eeprom.n3525 ;
    wire \eeprom.n3526 ;
    wire \eeprom.n2015 ;
    wire \eeprom.n2082 ;
    wire \eeprom.n3527 ;
    wire \eeprom.n3528 ;
    wire \eeprom.n2013 ;
    wire \eeprom.n2080 ;
    wire \eeprom.n3529 ;
    wire \eeprom.n3530 ;
    wire \eeprom.n3531 ;
    wire \eeprom.n2011 ;
    wire bfn_5_23_0_;
    wire \eeprom.n2081 ;
    wire \eeprom.n2014 ;
    wire \eeprom.n2012 ;
    wire \eeprom.n2079 ;
    wire \eeprom.n2083 ;
    wire \eeprom.n2016 ;
    wire \eeprom.n7_adj_470 ;
    wire \eeprom.n2019 ;
    wire \eeprom.n2086 ;
    wire \eeprom.n2309 ;
    wire \eeprom.n2319 ;
    wire \eeprom.n4509_cascade_ ;
    wire \eeprom.n8_adj_468 ;
    wire \eeprom.n2310 ;
    wire \eeprom.n6_cascade_ ;
    wire \eeprom.n2242_cascade_ ;
    wire \eeprom.n2044 ;
    wire \eeprom.n2084 ;
    wire \eeprom.n2214_cascade_ ;
    wire \eeprom.n2313 ;
    wire \eeprom.n2313_cascade_ ;
    wire \eeprom.n4505 ;
    wire \eeprom.n11 ;
    wire \eeprom.delay_counter_22 ;
    wire \eeprom.n2315 ;
    wire \eeprom.n2311 ;
    wire \eeprom.n4461 ;
    wire \eeprom.n4463 ;
    wire \eeprom.n4225_cascade_ ;
    wire \eeprom.n2143_cascade_ ;
    wire bfn_5_27_0_;
    wire \eeprom.n2118 ;
    wire \eeprom.n2185 ;
    wire \eeprom.n3532 ;
    wire \eeprom.n2117 ;
    wire \eeprom.n2184 ;
    wire \eeprom.n3533 ;
    wire \eeprom.n2116 ;
    wire \eeprom.n2183 ;
    wire \eeprom.n3534 ;
    wire \eeprom.n2115 ;
    wire \eeprom.n2182 ;
    wire \eeprom.n3535 ;
    wire \eeprom.n2114 ;
    wire \eeprom.n2181 ;
    wire \eeprom.n3536 ;
    wire \eeprom.n3537 ;
    wire \eeprom.n2112 ;
    wire \eeprom.n2179 ;
    wire \eeprom.n3538 ;
    wire \eeprom.n3539 ;
    wire \eeprom.n2111 ;
    wire \eeprom.n2178 ;
    wire bfn_5_28_0_;
    wire \eeprom.n2110 ;
    wire \eeprom.n3540 ;
    wire n26;
    wire bfn_5_29_0_;
    wire n25;
    wire n3485;
    wire n24;
    wire n3486;
    wire n23;
    wire n3487;
    wire n22;
    wire n3488;
    wire n21;
    wire n3489;
    wire n20;
    wire n3490;
    wire n19;
    wire n3491;
    wire n3492;
    wire n18;
    wire bfn_5_30_0_;
    wire n17;
    wire n3493;
    wire n16;
    wire n3494;
    wire n15;
    wire n3495;
    wire n14;
    wire n3496;
    wire n13;
    wire n3497;
    wire n12;
    wire n3498;
    wire n11;
    wire n3499;
    wire n3500;
    wire n10;
    wire bfn_5_31_0_;
    wire n9;
    wire n3501;
    wire n8;
    wire n3502;
    wire n7;
    wire n3503;
    wire n6;
    wire n3504;
    wire blink_counter_21;
    wire n3505;
    wire blink_counter_22;
    wire n3506;
    wire blink_counter_23;
    wire n3507;
    wire n3508;
    wire blink_counter_24;
    wire bfn_5_32_0_;
    wire n3509;
    wire blink_counter_25;
    wire bfn_6_18_0_;
    wire \eeprom.n3587 ;
    wire \eeprom.n3588 ;
    wire \eeprom.n3589 ;
    wire \eeprom.n3590 ;
    wire \eeprom.n3591 ;
    wire \eeprom.n3592 ;
    wire \eeprom.n3593 ;
    wire \eeprom.n3594 ;
    wire bfn_6_19_0_;
    wire \eeprom.n3595 ;
    wire \eeprom.n3596 ;
    wire \eeprom.n3597 ;
    wire \eeprom.n3598 ;
    wire \eeprom.n3599 ;
    wire \eeprom.n3600 ;
    wire \eeprom.n21 ;
    wire \eeprom.delay_counter_12 ;
    wire \eeprom.n29_adj_460 ;
    wire \eeprom.n2609 ;
    wire \eeprom.n2676 ;
    wire \eeprom.n2678 ;
    wire \eeprom.n2611_cascade_ ;
    wire \eeprom.n2519 ;
    wire \eeprom.n2586 ;
    wire bfn_6_21_0_;
    wire \eeprom.n2518 ;
    wire \eeprom.n2585 ;
    wire \eeprom.n3574 ;
    wire \eeprom.n2517 ;
    wire \eeprom.n2584 ;
    wire \eeprom.n3575 ;
    wire \eeprom.n2516 ;
    wire \eeprom.n2583 ;
    wire \eeprom.n3576 ;
    wire \eeprom.n2515 ;
    wire \eeprom.n2582 ;
    wire \eeprom.n3577 ;
    wire \eeprom.n2514 ;
    wire \eeprom.n2581 ;
    wire \eeprom.n3578 ;
    wire \eeprom.n3579 ;
    wire \eeprom.n2579 ;
    wire \eeprom.n3580 ;
    wire \eeprom.n3581 ;
    wire bfn_6_22_0_;
    wire \eeprom.n2510 ;
    wire \eeprom.n2577 ;
    wire \eeprom.n3582 ;
    wire \eeprom.n2509 ;
    wire \eeprom.n2576 ;
    wire \eeprom.n3583 ;
    wire \eeprom.n2508 ;
    wire \eeprom.n2575 ;
    wire \eeprom.n3584 ;
    wire \eeprom.n3585 ;
    wire \eeprom.n2506 ;
    wire \eeprom.n3586 ;
    wire \eeprom.n2412 ;
    wire \eeprom.n2479 ;
    wire \eeprom.n2511 ;
    wire \eeprom.n2578 ;
    wire \eeprom.n2511_cascade_ ;
    wire \eeprom.n12_adj_351 ;
    wire \eeprom.delay_counter_21 ;
    wire \eeprom.n2219_cascade_ ;
    wire \eeprom.n2318 ;
    wire \eeprom.n2580 ;
    wire \eeprom.n2513 ;
    wire \eeprom.n2539 ;
    wire \eeprom.n2574 ;
    wire \eeprom.n2606_cascade_ ;
    wire \eeprom.n2605 ;
    wire \eeprom.n2611 ;
    wire \eeprom.n10_adj_475_cascade_ ;
    wire \eeprom.n2413 ;
    wire \eeprom.n2480 ;
    wire \eeprom.n2512 ;
    wire \eeprom.n2408 ;
    wire \eeprom.n2475 ;
    wire \eeprom.n2440 ;
    wire \eeprom.n2507 ;
    wire \eeprom.n4801 ;
    wire \eeprom.n2017 ;
    wire \eeprom.n4799_cascade_ ;
    wire \eeprom.n4872 ;
    wire \eeprom.n2314 ;
    wire \eeprom.n2316 ;
    wire \eeprom.n2186 ;
    wire \eeprom.n2119 ;
    wire \eeprom.n2218_cascade_ ;
    wire \eeprom.n2317 ;
    wire \eeprom.n4447_cascade_ ;
    wire \eeprom.n4218 ;
    wire \eeprom.n2113 ;
    wire \eeprom.n2143 ;
    wire \eeprom.n2180 ;
    wire \eeprom.n2219 ;
    wire \eeprom.n2286 ;
    wire bfn_6_26_0_;
    wire \eeprom.n2218 ;
    wire \eeprom.n2285 ;
    wire \eeprom.n3541 ;
    wire \eeprom.n2217 ;
    wire \eeprom.n2284 ;
    wire \eeprom.n3542 ;
    wire \eeprom.n2216 ;
    wire \eeprom.n2283 ;
    wire \eeprom.n3543 ;
    wire \eeprom.n2215 ;
    wire \eeprom.n2282 ;
    wire \eeprom.n3544 ;
    wire \eeprom.n2214 ;
    wire \eeprom.n2281 ;
    wire \eeprom.n3545 ;
    wire \eeprom.n2213 ;
    wire \eeprom.n2280 ;
    wire \eeprom.n3546 ;
    wire \eeprom.n2212 ;
    wire \eeprom.n2279 ;
    wire \eeprom.n3547 ;
    wire \eeprom.n3548 ;
    wire \eeprom.n2211 ;
    wire \eeprom.n2278 ;
    wire bfn_6_27_0_;
    wire \eeprom.n2210 ;
    wire \eeprom.n2277 ;
    wire \eeprom.n3549 ;
    wire \eeprom.n2242 ;
    wire \eeprom.n2209 ;
    wire \eeprom.n3550 ;
    wire \eeprom.n2308 ;
    wire \eeprom.n2612 ;
    wire \eeprom.n2679 ;
    wire \eeprom.n2606 ;
    wire \eeprom.n2673 ;
    wire \eeprom.n2680 ;
    wire \eeprom.n2613 ;
    wire \eeprom.n2614 ;
    wire \eeprom.n2681 ;
    wire \eeprom.n2713_cascade_ ;
    wire \eeprom.n4695_cascade_ ;
    wire \eeprom.n16_adj_416_cascade_ ;
    wire \eeprom.n2618 ;
    wire \eeprom.n2685 ;
    wire \eeprom.n2674 ;
    wire \eeprom.n2686 ;
    wire \eeprom.n2619 ;
    wire \eeprom.n2718_cascade_ ;
    wire \eeprom.n4699 ;
    wire \eeprom.n2675 ;
    wire \eeprom.n2682 ;
    wire \eeprom.n2615 ;
    wire \eeprom.n2608 ;
    wire \eeprom.n12 ;
    wire \eeprom.n2607 ;
    wire \eeprom.n16 ;
    wire \eeprom.n2683 ;
    wire \eeprom.n2638_cascade_ ;
    wire \eeprom.n2616 ;
    wire \eeprom.n2617 ;
    wire \eeprom.n2684 ;
    wire \eeprom.n2815_cascade_ ;
    wire \eeprom.n28 ;
    wire \eeprom.n2610 ;
    wire \eeprom.n2677 ;
    wire \eeprom.n2638 ;
    wire \eeprom.n18 ;
    wire \eeprom.n2709_cascade_ ;
    wire \eeprom.n13_adj_417 ;
    wire \eeprom.n2737_cascade_ ;
    wire \eeprom.n2719 ;
    wire \eeprom.n2786 ;
    wire bfn_7_21_0_;
    wire \eeprom.n2718 ;
    wire \eeprom.n2785 ;
    wire \eeprom.n3601 ;
    wire \eeprom.n3602 ;
    wire \eeprom.n2716 ;
    wire \eeprom.n2783 ;
    wire \eeprom.n3603 ;
    wire \eeprom.n3604 ;
    wire \eeprom.n2714 ;
    wire \eeprom.n2781 ;
    wire \eeprom.n3605 ;
    wire \eeprom.n3606 ;
    wire \eeprom.n3607 ;
    wire \eeprom.n3608 ;
    wire bfn_7_22_0_;
    wire \eeprom.n3609 ;
    wire \eeprom.n3610 ;
    wire \eeprom.n3611 ;
    wire \eeprom.n3612 ;
    wire \eeprom.n3613 ;
    wire \eeprom.n3614 ;
    wire \eeprom.n2704 ;
    wire \eeprom.n3615 ;
    wire \eeprom.n2777 ;
    wire \eeprom.n2710 ;
    wire \eeprom.n2778 ;
    wire \eeprom.n2711 ;
    wire \eeprom.n2717 ;
    wire \eeprom.n2784 ;
    wire \eeprom.n2782 ;
    wire \eeprom.n2715 ;
    wire \eeprom.n2713 ;
    wire \eeprom.n2780 ;
    wire bfn_9_17_0_;
    wire \eeprom.n3706 ;
    wire \eeprom.n3707 ;
    wire \eeprom.n3708 ;
    wire \eeprom.n3709 ;
    wire \eeprom.n3710 ;
    wire \eeprom.n3711 ;
    wire \eeprom.n3712 ;
    wire \eeprom.n3713 ;
    wire bfn_9_18_0_;
    wire \eeprom.n3714 ;
    wire \eeprom.n3715 ;
    wire \eeprom.n3716 ;
    wire \eeprom.n3717 ;
    wire \eeprom.n3718 ;
    wire \eeprom.n3719 ;
    wire \eeprom.n3720 ;
    wire \eeprom.n3721 ;
    wire bfn_9_19_0_;
    wire \eeprom.n3722 ;
    wire \eeprom.n3723 ;
    wire \eeprom.n3724 ;
    wire \eeprom.n3725 ;
    wire \eeprom.n3726 ;
    wire bfn_9_20_0_;
    wire \eeprom.n3686 ;
    wire \eeprom.n3687 ;
    wire \eeprom.n3688 ;
    wire \eeprom.n3689 ;
    wire \eeprom.n3281 ;
    wire \eeprom.n3690 ;
    wire \eeprom.n3691 ;
    wire \eeprom.n3692 ;
    wire \eeprom.n3693 ;
    wire bfn_9_21_0_;
    wire \eeprom.n3694 ;
    wire \eeprom.n3695 ;
    wire \eeprom.n3696 ;
    wire \eeprom.n3697 ;
    wire \eeprom.n3698 ;
    wire \eeprom.n3699 ;
    wire \eeprom.n3700 ;
    wire \eeprom.n3701 ;
    wire bfn_9_22_0_;
    wire \eeprom.n3702 ;
    wire \eeprom.n3703 ;
    wire \eeprom.n3704 ;
    wire \eeprom.n3705 ;
    wire \eeprom.n2706 ;
    wire \eeprom.n2773 ;
    wire \eeprom.n2709 ;
    wire \eeprom.n2776 ;
    wire bfn_9_23_0_;
    wire \eeprom.n3616 ;
    wire \eeprom.n3617 ;
    wire \eeprom.n3618 ;
    wire \eeprom.n3619 ;
    wire \eeprom.n3620 ;
    wire \eeprom.n3621 ;
    wire \eeprom.n3622 ;
    wire \eeprom.n3623 ;
    wire bfn_9_24_0_;
    wire \eeprom.n3624 ;
    wire \eeprom.n3625 ;
    wire \eeprom.n3626 ;
    wire \eeprom.n3627 ;
    wire \eeprom.n3628 ;
    wire \eeprom.n3629 ;
    wire \eeprom.n3630 ;
    wire \eeprom.n3631 ;
    wire bfn_9_25_0_;
    wire \eeprom.n2873 ;
    wire \eeprom.n2872 ;
    wire \eeprom.n2904_cascade_ ;
    wire \eeprom.n3286 ;
    wire \eeprom.n3285 ;
    wire \eeprom.n3371 ;
    wire \eeprom.n3282 ;
    wire \eeprom.n3314_cascade_ ;
    wire \eeprom.n3272 ;
    wire \eeprom.n3274 ;
    wire \eeprom.n3273 ;
    wire \eeprom.n3280 ;
    wire \eeprom.n3312 ;
    wire \eeprom.n3379 ;
    wire \eeprom.n3312_cascade_ ;
    wire \eeprom.n3275 ;
    wire \eeprom.n3307 ;
    wire \eeprom.n3374 ;
    wire \eeprom.n3307_cascade_ ;
    wire \eeprom.n28_adj_482_cascade_ ;
    wire \eeprom.n3278 ;
    wire \eeprom.n3232_cascade_ ;
    wire \eeprom.n3367 ;
    wire \eeprom.n3276 ;
    wire \eeprom.n3279 ;
    wire \eeprom.n3271 ;
    wire \eeprom.n3277 ;
    wire \eeprom.n3209 ;
    wire \eeprom.n3369 ;
    wire \eeprom.n27 ;
    wire \eeprom.n3268 ;
    wire \eeprom.n32_adj_480 ;
    wire \eeprom.n3269 ;
    wire \eeprom.n2815 ;
    wire \eeprom.n2882 ;
    wire \eeprom.n2886 ;
    wire \eeprom.n2918_cascade_ ;
    wire \eeprom.n3267 ;
    wire \eeprom.n2705 ;
    wire \eeprom.n2772 ;
    wire \eeprom.n2803 ;
    wire \eeprom.n2804_cascade_ ;
    wire \eeprom.n3270 ;
    wire \eeprom.n2712 ;
    wire \eeprom.n2779 ;
    wire \eeprom.n2707 ;
    wire \eeprom.n2774 ;
    wire \eeprom.n2806 ;
    wire \eeprom.n2806_cascade_ ;
    wire \eeprom.n2805 ;
    wire \eeprom.n18_adj_418 ;
    wire \eeprom.n2708 ;
    wire \eeprom.n2775 ;
    wire \eeprom.n2737 ;
    wire \eeprom.n2807 ;
    wire \eeprom.n2874 ;
    wire \eeprom.n2807_cascade_ ;
    wire \eeprom.n2881 ;
    wire \eeprom.n2913_cascade_ ;
    wire \eeprom.n4529 ;
    wire \eeprom.n2814 ;
    wire \eeprom.n2819 ;
    wire \eeprom.n4533_cascade_ ;
    wire \eeprom.n20 ;
    wire \eeprom.n15_cascade_ ;
    wire \eeprom.n2816 ;
    wire \eeprom.n2836_cascade_ ;
    wire \eeprom.n2883 ;
    wire \eeprom.n2809 ;
    wire \eeprom.n2876 ;
    wire \eeprom.n2804 ;
    wire \eeprom.n2871 ;
    wire \eeprom.n19 ;
    wire \eeprom.n22_cascade_ ;
    wire \eeprom.n2885 ;
    wire \eeprom.n2818 ;
    wire \eeprom.n4703 ;
    wire \eeprom.n2917_cascade_ ;
    wire \eeprom.n4707_cascade_ ;
    wire \eeprom.n15_adj_419 ;
    wire \eeprom.n2875 ;
    wire \eeprom.n2808 ;
    wire \eeprom.n3385 ;
    wire \eeprom.n3283 ;
    wire \eeprom.n3315_cascade_ ;
    wire \eeprom.n3318 ;
    wire \eeprom.n4719_cascade_ ;
    wire \eeprom.n4721 ;
    wire \eeprom.n3304 ;
    wire \eeprom.n4151_cascade_ ;
    wire \eeprom.n3302 ;
    wire \eeprom.n3317 ;
    wire \eeprom.n3384 ;
    wire \eeprom.n3375 ;
    wire \eeprom.n3308 ;
    wire \eeprom.n3407_cascade_ ;
    wire \eeprom.n28_adj_484 ;
    wire \eeprom.n27_adj_486_cascade_ ;
    wire \eeprom.n26_adj_485 ;
    wire \eeprom.n3306 ;
    wire \eeprom.n3331_cascade_ ;
    wire \eeprom.n3373 ;
    wire \eeprom.n3305 ;
    wire \eeprom.n3372 ;
    wire \eeprom.n3376 ;
    wire \eeprom.n3309 ;
    wire \eeprom.n3219 ;
    wire \eeprom.n4615_cascade_ ;
    wire \eeprom.n3218 ;
    wire \eeprom.n21_adj_477 ;
    wire \eeprom.n4611 ;
    wire \eeprom.n3300 ;
    wire \eeprom.n3298 ;
    wire \eeprom.n25_adj_487 ;
    wire \eeprom.n3301 ;
    wire \eeprom.n3368 ;
    wire \eeprom.n3284 ;
    wire \eeprom.n3232 ;
    wire \eeprom.n3210 ;
    wire \eeprom.n3113_cascade_ ;
    wire \eeprom.n3212 ;
    wire \eeprom.n3208 ;
    wire \eeprom.n25_adj_478 ;
    wire \eeprom.n3213 ;
    wire \eeprom.n3116_cascade_ ;
    wire \eeprom.n3215 ;
    wire bfn_11_21_0_;
    wire \eeprom.n2918 ;
    wire \eeprom.n2985 ;
    wire \eeprom.n3632 ;
    wire \eeprom.n3633 ;
    wire \eeprom.n3634 ;
    wire \eeprom.n3635 ;
    wire \eeprom.n3636 ;
    wire \eeprom.n3637 ;
    wire \eeprom.n3638 ;
    wire \eeprom.n3639 ;
    wire bfn_11_22_0_;
    wire \eeprom.n3640 ;
    wire \eeprom.n3641 ;
    wire \eeprom.n3642 ;
    wire \eeprom.n3643 ;
    wire \eeprom.n3644 ;
    wire \eeprom.n3645 ;
    wire \eeprom.n3646 ;
    wire \eeprom.n3647 ;
    wire bfn_11_23_0_;
    wire \eeprom.n2902 ;
    wire \eeprom.n3648 ;
    wire \eeprom.n2906 ;
    wire \eeprom.n2973 ;
    wire \eeprom.n2903 ;
    wire \eeprom.n2970 ;
    wire \eeprom.n2879 ;
    wire \eeprom.n2812 ;
    wire \eeprom.n2880 ;
    wire \eeprom.n2813 ;
    wire \eeprom.n2913 ;
    wire \eeprom.n2980 ;
    wire \eeprom.n2817 ;
    wire \eeprom.n2884 ;
    wire \eeprom.n2877 ;
    wire \eeprom.n2810 ;
    wire \eeprom.n2909_cascade_ ;
    wire \eeprom.n18_adj_420 ;
    wire \eeprom.n2975 ;
    wire \eeprom.n2908 ;
    wire \eeprom.n2878 ;
    wire \eeprom.n2811 ;
    wire \eeprom.n2836 ;
    wire \eeprom.n2915 ;
    wire \eeprom.n2982 ;
    wire \eeprom.n2911 ;
    wire \eeprom.n2978 ;
    wire \eeprom.n2984 ;
    wire \eeprom.n2917 ;
    wire \eeprom.n3315 ;
    wire \eeprom.n3382 ;
    wire \eeprom.n3414_cascade_ ;
    wire \eeprom.n4689_cascade_ ;
    wire \eeprom.n4144_cascade_ ;
    wire \eeprom.n3386 ;
    wire \eeprom.n3319 ;
    wire \eeprom.n3316 ;
    wire \eeprom.n3383 ;
    wire \eeprom.n3314 ;
    wire \eeprom.n3381 ;
    wire \eeprom.n3413_cascade_ ;
    wire \eeprom.n4687 ;
    wire \eeprom.n3378 ;
    wire \eeprom.n3311 ;
    wire \eeprom.n3410_cascade_ ;
    wire \eeprom.n3505_cascade_ ;
    wire \eeprom.n3310 ;
    wire \eeprom.n3377 ;
    wire \eeprom.n3608_adj_451_cascade_ ;
    wire \eeprom.n3313 ;
    wire \eeprom.n3380 ;
    wire \eeprom.n3412_cascade_ ;
    wire \eeprom.n3303 ;
    wire \eeprom.n3370 ;
    wire \eeprom.n3366 ;
    wire \eeprom.n3299 ;
    wire \eeprom.n3331 ;
    wire \eeprom.n3500_cascade_ ;
    wire \eeprom.n3216 ;
    wire \eeprom.n3203 ;
    wire \eeprom.n3217 ;
    wire \eeprom.n18_adj_432_cascade_ ;
    wire \eeprom.n26_adj_466_cascade_ ;
    wire \eeprom.n4711_cascade_ ;
    wire \eeprom.n4715 ;
    wire \eeprom.n3206 ;
    wire \eeprom.n3214 ;
    wire \eeprom.n3119 ;
    wire \eeprom.n3186 ;
    wire bfn_12_22_0_;
    wire \eeprom.n3185 ;
    wire \eeprom.n3667 ;
    wire \eeprom.n3184 ;
    wire \eeprom.n3668 ;
    wire \eeprom.n3116 ;
    wire \eeprom.n3183 ;
    wire \eeprom.n3669 ;
    wire \eeprom.n3182 ;
    wire \eeprom.n3670 ;
    wire \eeprom.n3181 ;
    wire \eeprom.n3671 ;
    wire \eeprom.n3113 ;
    wire \eeprom.n3180 ;
    wire \eeprom.n3672 ;
    wire \eeprom.n3673 ;
    wire \eeprom.n3674 ;
    wire \eeprom.n3178 ;
    wire bfn_12_23_0_;
    wire \eeprom.n3177 ;
    wire \eeprom.n3675 ;
    wire \eeprom.n3176 ;
    wire \eeprom.n3676 ;
    wire \eeprom.n3677 ;
    wire \eeprom.n3174 ;
    wire \eeprom.n3678 ;
    wire \eeprom.n3679 ;
    wire \eeprom.n3680 ;
    wire \eeprom.n3171 ;
    wire \eeprom.n3681 ;
    wire \eeprom.n3682 ;
    wire bfn_12_24_0_;
    wire \eeprom.n3683 ;
    wire \eeprom.n3684 ;
    wire \eeprom.n3685 ;
    wire \eeprom.n2971 ;
    wire \eeprom.n2904 ;
    wire \eeprom.n2977 ;
    wire \eeprom.n2910 ;
    wire \eeprom.n3497_cascade_ ;
    wire \eeprom.n28_adj_493_cascade_ ;
    wire \eeprom.n18_adj_488_cascade_ ;
    wire \eeprom.n29_adj_491 ;
    wire \eeprom.n28_adj_490 ;
    wire \eeprom.n30_adj_489_cascade_ ;
    wire \eeprom.n27_adj_492 ;
    wire \eeprom.n3430_cascade_ ;
    wire \eeprom.n3609_adj_445 ;
    wire \eeprom.n3508_cascade_ ;
    wire \eeprom.n31_adj_496 ;
    wire \eeprom.n29_adj_497 ;
    wire \eeprom.n30_adj_495_cascade_ ;
    wire \eeprom.n32_adj_494 ;
    wire \eeprom.n3606_adj_446_cascade_ ;
    wire \eeprom.n4451_cascade_ ;
    wire \eeprom.n4453 ;
    wire \eeprom.n3599_adj_450_cascade_ ;
    wire \eeprom.n4429 ;
    wire \eeprom.n29 ;
    wire \eeprom.n3600_adj_449 ;
    wire \eeprom.n4581 ;
    wire \eeprom.n3117 ;
    wire \eeprom.n3108 ;
    wire \eeprom.n3175 ;
    wire \eeprom.n3108_cascade_ ;
    wire \eeprom.n3105 ;
    wire \eeprom.n3172 ;
    wire \eeprom.n3105_cascade_ ;
    wire \eeprom.n3204 ;
    wire \eeprom.n3179 ;
    wire \eeprom.n3211 ;
    wire \eeprom.n3115 ;
    wire \eeprom.n3169 ;
    wire \eeprom.n3201 ;
    wire \eeprom.n3207 ;
    wire \eeprom.n3201_cascade_ ;
    wire \eeprom.n24_adj_481 ;
    wire \eeprom.n3114 ;
    wire \eeprom.n2905 ;
    wire \eeprom.n2972 ;
    wire \eeprom.n3118 ;
    wire \eeprom.n3102 ;
    wire \eeprom.n3102_cascade_ ;
    wire \eeprom.n22_adj_465 ;
    wire \eeprom.n3104 ;
    wire \eeprom.n3170 ;
    wire \eeprom.n3202 ;
    wire \eeprom.n3168 ;
    wire \eeprom.n3200 ;
    wire \eeprom.n2983 ;
    wire \eeprom.n2916 ;
    wire \eeprom.n3106 ;
    wire \eeprom.n3173 ;
    wire \eeprom.n3106_cascade_ ;
    wire \eeprom.n3133 ;
    wire \eeprom.n3205 ;
    wire \eeprom.n3205_cascade_ ;
    wire \eeprom.n3199 ;
    wire \eeprom.n16_adj_479 ;
    wire \eeprom.n2907 ;
    wire \eeprom.n2974 ;
    wire \eeprom.n2914 ;
    wire \eeprom.n2981 ;
    wire \eeprom.n3101 ;
    wire bfn_14_17_0_;
    wire \eeprom.n3727 ;
    wire \eeprom.n3728 ;
    wire \eeprom.n3729 ;
    wire \eeprom.n3415 ;
    wire \eeprom.n3482_adj_401 ;
    wire \eeprom.n3730 ;
    wire \eeprom.n3414 ;
    wire \eeprom.n3481_adj_399 ;
    wire \eeprom.n3731 ;
    wire \eeprom.n3413 ;
    wire \eeprom.n3480_adj_398 ;
    wire \eeprom.n3732 ;
    wire \eeprom.n3412 ;
    wire \eeprom.n3479_adj_394 ;
    wire \eeprom.n3733 ;
    wire \eeprom.n3734 ;
    wire \eeprom.n3411 ;
    wire \eeprom.n3478_adj_393 ;
    wire bfn_14_18_0_;
    wire \eeprom.n3410 ;
    wire \eeprom.n3477_adj_392 ;
    wire \eeprom.n3735 ;
    wire \eeprom.n3409 ;
    wire \eeprom.n3476_adj_391 ;
    wire \eeprom.n3736 ;
    wire \eeprom.n3408 ;
    wire \eeprom.n3475_adj_390 ;
    wire \eeprom.n3737 ;
    wire \eeprom.n3407 ;
    wire \eeprom.n3474_adj_389 ;
    wire \eeprom.n3738 ;
    wire \eeprom.n3406 ;
    wire \eeprom.n3473_adj_388 ;
    wire \eeprom.n3739 ;
    wire \eeprom.n3405 ;
    wire \eeprom.n3472_adj_387 ;
    wire \eeprom.n3740 ;
    wire \eeprom.n3741 ;
    wire \eeprom.n3742 ;
    wire \eeprom.n3403 ;
    wire \eeprom.n3470_adj_385 ;
    wire bfn_14_19_0_;
    wire \eeprom.n3402 ;
    wire \eeprom.n3469_adj_384 ;
    wire \eeprom.n3743 ;
    wire \eeprom.n3401 ;
    wire \eeprom.n3468_adj_383 ;
    wire \eeprom.n3744 ;
    wire \eeprom.n3400 ;
    wire \eeprom.n3467_adj_382 ;
    wire \eeprom.n3745 ;
    wire \eeprom.n3399 ;
    wire \eeprom.n3466_adj_381 ;
    wire \eeprom.n3746 ;
    wire \eeprom.n3398 ;
    wire \eeprom.n3465_adj_380 ;
    wire \eeprom.n3747 ;
    wire \eeprom.n3397 ;
    wire \eeprom.n3748 ;
    wire \eeprom.n4583 ;
    wire \eeprom.n31_cascade_ ;
    wire \eeprom.n4433 ;
    wire \eeprom.n3598_adj_452 ;
    wire \eeprom.n31_adj_476 ;
    wire \eeprom.delay_counter_31 ;
    wire \eeprom.n24_adj_459 ;
    wire \eeprom.n4559_cascade_ ;
    wire \eeprom.n4563_cascade_ ;
    wire \eeprom.n21_adj_422 ;
    wire \eeprom.n17_adj_421_cascade_ ;
    wire \eeprom.n24_cascade_ ;
    wire \eeprom.n20_adj_423 ;
    wire \eeprom.n3034_cascade_ ;
    wire \eeprom.n3112 ;
    wire \eeprom.n2912 ;
    wire \eeprom.n2979 ;
    wire \eeprom.n3103 ;
    wire \eeprom.n4137 ;
    wire \eeprom.n3417 ;
    wire \eeprom.n3484_adj_406 ;
    wire \eeprom.n3418 ;
    wire \eeprom.n3485 ;
    wire \eeprom.n3517_adj_374_cascade_ ;
    wire \eeprom.n4729 ;
    wire \eeprom.n3416 ;
    wire \eeprom.n3483_adj_404 ;
    wire \eeprom.n3515_adj_370_cascade_ ;
    wire \eeprom.n4727 ;
    wire \eeprom.n3419 ;
    wire \eeprom.n3486 ;
    wire \eeprom.n3471_adj_386 ;
    wire \eeprom.n3430 ;
    wire \eeprom.n3404 ;
    wire \eeprom.n3615_adj_344_cascade_ ;
    wire \eeprom.n3714_adj_442_cascade_ ;
    wire \eeprom.n3617_adj_346_cascade_ ;
    wire \eeprom.n4619 ;
    wire \eeprom.n4427_cascade_ ;
    wire \eeprom.n3596_adj_454 ;
    wire \eeprom.n28_adj_455_cascade_ ;
    wire \eeprom.n4567 ;
    wire \eeprom.n3628_adj_437_cascade_ ;
    wire \eeprom.n3716_adj_439_cascade_ ;
    wire \eeprom.n3605_adj_453 ;
    wire \eeprom.n3618_adj_350_cascade_ ;
    wire \eeprom.n4623 ;
    wire \eeprom.n4425 ;
    wire \eeprom.delay_counter_0 ;
    wire \eeprom.n1166 ;
    wire bfn_15_20_0_;
    wire \eeprom.delay_counter_1 ;
    wire \eeprom.n3724_adj_335 ;
    wire \eeprom.n3772 ;
    wire \eeprom.delay_counter_2 ;
    wire \eeprom.n3723_adj_334 ;
    wire \eeprom.n3773 ;
    wire \eeprom.delay_counter_3 ;
    wire \eeprom.n3722_adj_433 ;
    wire \eeprom.n3774 ;
    wire \eeprom.delay_counter_4 ;
    wire \eeprom.n3721_adj_434 ;
    wire \eeprom.n3775 ;
    wire \eeprom.delay_counter_5 ;
    wire \eeprom.n3720_adj_435 ;
    wire \eeprom.n3776 ;
    wire \eeprom.delay_counter_6 ;
    wire \eeprom.n3719_adj_436 ;
    wire \eeprom.n3777 ;
    wire \eeprom.n3778 ;
    wire \eeprom.n3779 ;
    wire bfn_15_21_0_;
    wire \eeprom.n4909 ;
    wire \eeprom.n3716_adj_439 ;
    wire \eeprom.n3780 ;
    wire \eeprom.n3781 ;
    wire \eeprom.n4915 ;
    wire \eeprom.n3714_adj_442 ;
    wire \eeprom.n3782 ;
    wire \eeprom.n3783 ;
    wire \eeprom.n4921 ;
    wire \eeprom.n3712_adj_444 ;
    wire \eeprom.n3784 ;
    wire \eeprom.n2 ;
    wire \eeprom.n4924 ;
    wire \eeprom.n3785 ;
    wire \eeprom.n3713_adj_443 ;
    wire \eeprom.n4918 ;
    wire \eeprom.number_of_bytes_7_N_68_5 ;
    wire \eeprom.number_of_bytes_7_N_68_4 ;
    wire \eeprom.number_of_bytes_7_N_68_3 ;
    wire \eeprom.number_of_bytes_7_N_68_6 ;
    wire \eeprom.number_of_bytes_7_N_68_8 ;
    wire \eeprom.n4301_cascade_ ;
    wire \eeprom.number_of_bytes_7_N_68_7 ;
    wire \eeprom.number_of_bytes_7_N_68_9 ;
    wire \eeprom.number_of_bytes_7_N_68_10 ;
    wire \eeprom.n4307_cascade_ ;
    wire \eeprom.number_of_bytes_7_N_68_11 ;
    wire \eeprom.number_of_bytes_7_N_68_12 ;
    wire \eeprom.number_of_bytes_7_N_68_13 ;
    wire \eeprom.n4313_cascade_ ;
    wire \eeprom.number_of_bytes_7_N_68_14 ;
    wire sda_enable;
    wire CLK_N;
    wire \eeprom.number_of_bytes_7_N_68_2 ;
    wire \eeprom.number_of_bytes_7_N_68_0 ;
    wire \eeprom.number_of_bytes_7_N_68_1 ;
    wire \eeprom.n4295 ;
    wire \eeprom.n3111 ;
    wire \eeprom.n3109 ;
    wire \eeprom.n3110 ;
    wire \eeprom.n3107 ;
    wire \eeprom.n2986 ;
    wire \eeprom.n2919 ;
    wire \eeprom.n2909 ;
    wire \eeprom.n2976 ;
    wire \eeprom.n2935 ;
    wire \eeprom.n3519_adj_379 ;
    wire \eeprom.n3586_adj_378 ;
    wire bfn_16_17_0_;
    wire \eeprom.n3518_adj_376 ;
    wire \eeprom.n3585_adj_375 ;
    wire \eeprom.n3749 ;
    wire \eeprom.n3517_adj_374 ;
    wire \eeprom.n3584_adj_373 ;
    wire \eeprom.n3750 ;
    wire \eeprom.n3516_adj_372 ;
    wire \eeprom.n3583_adj_371 ;
    wire \eeprom.n3751 ;
    wire \eeprom.n3515_adj_370 ;
    wire \eeprom.n3582_adj_369 ;
    wire \eeprom.n3752 ;
    wire \eeprom.n3514_adj_368 ;
    wire \eeprom.n3581_adj_367 ;
    wire \eeprom.n3753 ;
    wire \eeprom.n3513_adj_366 ;
    wire \eeprom.n3580_adj_365 ;
    wire \eeprom.n3754 ;
    wire \eeprom.n3512_adj_364 ;
    wire \eeprom.n3579_adj_363 ;
    wire \eeprom.n3755 ;
    wire \eeprom.n3756 ;
    wire \eeprom.n3511_adj_362 ;
    wire \eeprom.n3578_adj_361 ;
    wire bfn_16_18_0_;
    wire \eeprom.n3510_adj_360 ;
    wire \eeprom.n3577_adj_359 ;
    wire \eeprom.n3757 ;
    wire \eeprom.n3509 ;
    wire \eeprom.n3576_adj_358 ;
    wire \eeprom.n3758 ;
    wire \eeprom.n3508 ;
    wire \eeprom.n3575_adj_357 ;
    wire \eeprom.n3759 ;
    wire \eeprom.n3507 ;
    wire \eeprom.n3574_adj_356 ;
    wire \eeprom.n3760 ;
    wire \eeprom.n3506 ;
    wire \eeprom.n3573_adj_355 ;
    wire \eeprom.n3761 ;
    wire \eeprom.n3505 ;
    wire \eeprom.n3572_adj_354 ;
    wire \eeprom.n3762 ;
    wire \eeprom.n3504 ;
    wire \eeprom.n3571_adj_353 ;
    wire \eeprom.n3763 ;
    wire \eeprom.n3764 ;
    wire \eeprom.n3503 ;
    wire \eeprom.n3570_adj_349 ;
    wire bfn_16_19_0_;
    wire \eeprom.n3502 ;
    wire \eeprom.n3569_adj_348 ;
    wire \eeprom.n3765 ;
    wire \eeprom.n3501 ;
    wire \eeprom.n3568_adj_347 ;
    wire \eeprom.n3766 ;
    wire \eeprom.n3500 ;
    wire \eeprom.n3567_adj_341 ;
    wire \eeprom.n3767 ;
    wire \eeprom.n3499 ;
    wire \eeprom.n3566_adj_340 ;
    wire \eeprom.n3768 ;
    wire \eeprom.n3498 ;
    wire \eeprom.n3565_adj_338 ;
    wire \eeprom.n3769 ;
    wire \eeprom.n3497 ;
    wire \eeprom.n3564_adj_337 ;
    wire \eeprom.n3770 ;
    wire \eeprom.n3496 ;
    wire \eeprom.n3529_adj_336 ;
    wire \eeprom.n3771 ;
    wire \eeprom.n4765 ;
    wire bfn_16_20_0_;
    wire \eeprom.n3510 ;
    wire \eeprom.n3617_adj_346 ;
    wire \eeprom.n1351 ;
    wire \eeprom.n3511 ;
    wire \eeprom.n3512 ;
    wire \eeprom.n3615_adj_344 ;
    wire \eeprom.n1349 ;
    wire \eeprom.n3513 ;
    wire \eeprom.n3614_adj_343 ;
    wire \eeprom.n1348 ;
    wire \eeprom.n3514 ;
    wire \eeprom.n3613_adj_342 ;
    wire \eeprom.n1347 ;
    wire \eeprom.n3515 ;
    wire \eeprom.n3612_adj_339 ;
    wire \eeprom.n3516 ;
    wire \eeprom.n1350 ;
    wire \eeprom.n3616_adj_345 ;
    wire \eeprom.n3715_adj_441 ;
    wire \eeprom.n3715_adj_441_cascade_ ;
    wire \eeprom.n4912 ;
    wire \eeprom.n1346 ;
    wire \eeprom.n3711_adj_456 ;
    wire \eeprom.n1352 ;
    wire \eeprom.n3618_adj_350 ;
    wire \eeprom.n3717_adj_438 ;
    wire \eeprom.n3717_adj_438_cascade_ ;
    wire \eeprom.n4906 ;
    wire \eeprom.n1353 ;
    wire \eeprom.n3619_adj_352 ;
    wire \eeprom.n3628_adj_437 ;
    wire \eeprom.n4766 ;
    wire \eeprom.n4766_cascade_ ;
    wire \eeprom.n4903 ;
    wire \eeprom.n3019 ;
    wire \eeprom.n3086 ;
    wire bfn_16_23_0_;
    wire \eeprom.n3018 ;
    wire \eeprom.n3085 ;
    wire \eeprom.n3649 ;
    wire \eeprom.n3017 ;
    wire \eeprom.n3084 ;
    wire \eeprom.n3650 ;
    wire \eeprom.n3016 ;
    wire \eeprom.n3083 ;
    wire \eeprom.n3651 ;
    wire \eeprom.n3015 ;
    wire \eeprom.n3082 ;
    wire \eeprom.n3652 ;
    wire \eeprom.n3014 ;
    wire \eeprom.n3081 ;
    wire \eeprom.n3653 ;
    wire \eeprom.n3013 ;
    wire \eeprom.n3080 ;
    wire \eeprom.n3654 ;
    wire \eeprom.n3012 ;
    wire \eeprom.n3079 ;
    wire \eeprom.n3655 ;
    wire \eeprom.n3656 ;
    wire \eeprom.n3011 ;
    wire \eeprom.n3078 ;
    wire bfn_16_24_0_;
    wire \eeprom.n3010 ;
    wire \eeprom.n3077 ;
    wire \eeprom.n3657 ;
    wire \eeprom.n3009 ;
    wire \eeprom.n3076 ;
    wire \eeprom.n3658 ;
    wire \eeprom.n3008 ;
    wire \eeprom.n3075 ;
    wire \eeprom.n3659 ;
    wire \eeprom.n3007 ;
    wire \eeprom.n3074 ;
    wire \eeprom.n3660 ;
    wire \eeprom.n3006 ;
    wire \eeprom.n3073 ;
    wire \eeprom.n3661 ;
    wire \eeprom.n3005 ;
    wire \eeprom.n3072 ;
    wire \eeprom.n3662 ;
    wire \eeprom.n3004 ;
    wire \eeprom.n3071 ;
    wire \eeprom.n3663 ;
    wire \eeprom.n3664 ;
    wire \eeprom.n3003 ;
    wire \eeprom.n3070 ;
    wire bfn_16_25_0_;
    wire \eeprom.n3002 ;
    wire \eeprom.n3069 ;
    wire \eeprom.n3665 ;
    wire \eeprom.n3001 ;
    wire \eeprom.n3034 ;
    wire \eeprom.n3666 ;
    wire \eeprom.n3100 ;
    wire CONSTANT_ONE_NET;
    wire _gnd_net_;

    defparam CS_CLK_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam CS_CLK_pad_iopad.PULLUP=1'b0;
    IO_PAD CS_CLK_pad_iopad (
            .OE(N__28245),
            .DIN(N__28244),
            .DOUT(N__28243),
            .PACKAGEPIN(CS_CLK));
    defparam CS_CLK_pad_preio.PIN_TYPE=6'b011001;
    defparam CS_CLK_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO CS_CLK_pad_preio (
            .PADOEN(N__28245),
            .PADOUT(N__28244),
            .PADIN(N__28243),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam CS_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam CS_pad_iopad.PULLUP=1'b0;
    IO_PAD CS_pad_iopad (
            .OE(N__28236),
            .DIN(N__28235),
            .DOUT(N__28234),
            .PACKAGEPIN(CS));
    defparam CS_pad_preio.PIN_TYPE=6'b011001;
    defparam CS_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO CS_pad_preio (
            .PADOEN(N__28236),
            .PADOUT(N__28235),
            .PADIN(N__28234),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam DE_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam DE_pad_iopad.PULLUP=1'b0;
    IO_PAD DE_pad_iopad (
            .OE(N__28227),
            .DIN(N__28226),
            .DOUT(N__28225),
            .PACKAGEPIN(DE));
    defparam DE_pad_preio.PIN_TYPE=6'b011001;
    defparam DE_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO DE_pad_preio (
            .PADOEN(N__28227),
            .PADOUT(N__28226),
            .PADIN(N__28225),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam INHA_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam INHA_pad_iopad.PULLUP=1'b0;
    IO_PAD INHA_pad_iopad (
            .OE(N__28218),
            .DIN(N__28217),
            .DOUT(N__28216),
            .PACKAGEPIN(INHA));
    defparam INHA_pad_preio.PIN_TYPE=6'b011001;
    defparam INHA_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO INHA_pad_preio (
            .PADOEN(N__28218),
            .PADOUT(N__28217),
            .PADIN(N__28216),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam INHB_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam INHB_pad_iopad.PULLUP=1'b0;
    IO_PAD INHB_pad_iopad (
            .OE(N__28209),
            .DIN(N__28208),
            .DOUT(N__28207),
            .PACKAGEPIN(INHB));
    defparam INHB_pad_preio.PIN_TYPE=6'b011001;
    defparam INHB_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO INHB_pad_preio (
            .PADOEN(N__28209),
            .PADOUT(N__28208),
            .PADIN(N__28207),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam INHC_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam INHC_pad_iopad.PULLUP=1'b0;
    IO_PAD INHC_pad_iopad (
            .OE(N__28200),
            .DIN(N__28199),
            .DOUT(N__28198),
            .PACKAGEPIN(INHC));
    defparam INHC_pad_preio.PIN_TYPE=6'b011001;
    defparam INHC_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO INHC_pad_preio (
            .PADOEN(N__28200),
            .PADOUT(N__28199),
            .PADIN(N__28198),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam INLA_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam INLA_pad_iopad.PULLUP=1'b0;
    IO_PAD INLA_pad_iopad (
            .OE(N__28191),
            .DIN(N__28190),
            .DOUT(N__28189),
            .PACKAGEPIN(INLA));
    defparam INLA_pad_preio.PIN_TYPE=6'b011001;
    defparam INLA_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO INLA_pad_preio (
            .PADOEN(N__28191),
            .PADOUT(N__28190),
            .PADIN(N__28189),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam INLB_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam INLB_pad_iopad.PULLUP=1'b0;
    IO_PAD INLB_pad_iopad (
            .OE(N__28182),
            .DIN(N__28181),
            .DOUT(N__28180),
            .PACKAGEPIN(INLB));
    defparam INLB_pad_preio.PIN_TYPE=6'b011001;
    defparam INLB_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO INLB_pad_preio (
            .PADOEN(N__28182),
            .PADOUT(N__28181),
            .PADIN(N__28180),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam INLC_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam INLC_pad_iopad.PULLUP=1'b0;
    IO_PAD INLC_pad_iopad (
            .OE(N__28173),
            .DIN(N__28172),
            .DOUT(N__28171),
            .PACKAGEPIN(INLC));
    defparam INLC_pad_preio.PIN_TYPE=6'b011001;
    defparam INLC_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO INLC_pad_preio (
            .PADOEN(N__28173),
            .PADOUT(N__28172),
            .PADIN(N__28171),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam LED_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam LED_pad_iopad.PULLUP=1'b0;
    IO_PAD LED_pad_iopad (
            .OE(N__28164),
            .DIN(N__28163),
            .DOUT(N__28162),
            .PACKAGEPIN(LED));
    defparam LED_pad_preio.PIN_TYPE=6'b011001;
    defparam LED_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO LED_pad_preio (
            .PADOEN(N__28164),
            .PADOUT(N__28163),
            .PADIN(N__28162),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__13496),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam NEOPXL_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam NEOPXL_pad_iopad.PULLUP=1'b0;
    IO_PAD NEOPXL_pad_iopad (
            .OE(N__28155),
            .DIN(N__28154),
            .DOUT(N__28153),
            .PACKAGEPIN(NEOPXL));
    defparam NEOPXL_pad_preio.PIN_TYPE=6'b011001;
    defparam NEOPXL_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO NEOPXL_pad_preio (
            .PADOEN(N__28155),
            .PADOUT(N__28154),
            .PADIN(N__28153),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam TX_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam TX_pad_iopad.PULLUP=1'b0;
    IO_PAD TX_pad_iopad (
            .OE(N__28146),
            .DIN(N__28145),
            .DOUT(N__28144),
            .PACKAGEPIN(TX));
    defparam TX_pad_preio.PIN_TYPE=6'b011001;
    defparam TX_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO TX_pad_preio (
            .PADOEN(N__28146),
            .PADOUT(N__28145),
            .PADIN(N__28144),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam USBPU_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam USBPU_pad_iopad.PULLUP=1'b0;
    IO_PAD USBPU_pad_iopad (
            .OE(N__28137),
            .DIN(N__28136),
            .DOUT(N__28135),
            .PACKAGEPIN(USBPU));
    defparam USBPU_pad_preio.PIN_TYPE=6'b011001;
    defparam USBPU_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO USBPU_pad_preio (
            .PADOEN(N__28137),
            .PADOUT(N__28136),
            .PADIN(N__28135),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam scl_output_iopad.IO_STANDARD="SB_LVCMOS";
    defparam scl_output_iopad.PULLUP=1'b1;
    IO_PAD scl_output_iopad (
            .OE(N__28128),
            .DIN(N__28127),
            .DOUT(N__28126),
            .PACKAGEPIN(SCL));
    defparam scl_output_preio.PIN_TYPE=6'b101001;
    defparam scl_output_preio.NEG_TRIGGER=1'b0;
    PRE_IO scl_output_preio (
            .PADOEN(N__28128),
            .PADOUT(N__28127),
            .PADIN(N__28126),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam sda_output_iopad.IO_STANDARD="SB_LVCMOS";
    defparam sda_output_iopad.PULLUP=1'b1;
    IO_PAD sda_output_iopad (
            .OE(N__28119),
            .DIN(N__28118),
            .DOUT(N__28117),
            .PACKAGEPIN(SDA));
    defparam sda_output_preio.PIN_TYPE=6'b101001;
    defparam sda_output_preio.NEG_TRIGGER=1'b0;
    PRE_IO sda_output_preio (
            .PADOEN(N__28119),
            .PADOUT(N__28118),
            .PADIN(N__28117),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__24374));
    defparam CLK_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam CLK_pad_iopad.PULLUP=1'b0;
    IO_PAD CLK_pad_iopad (
            .OE(N__28110),
            .DIN(N__28109),
            .DOUT(N__28108),
            .PACKAGEPIN(CLK));
    defparam CLK_pad_preio.PIN_TYPE=6'b000001;
    defparam CLK_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO CLK_pad_preio (
            .PADOEN(N__28110),
            .PADOUT(N__28109),
            .PADIN(N__28108),
            .CLOCKENABLE(),
            .DIN0(CLK_pad_gb_input),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    CascadeMux I__6599 (
            .O(N__28091),
            .I(N__28088));
    InMux I__6598 (
            .O(N__28088),
            .I(N__28085));
    LocalMux I__6597 (
            .O(N__28085),
            .I(N__28082));
    Span4Mux_h I__6596 (
            .O(N__28082),
            .I(N__28079));
    Odrv4 I__6595 (
            .O(N__28079),
            .I(\eeprom.n3072 ));
    InMux I__6594 (
            .O(N__28076),
            .I(\eeprom.n3662 ));
    InMux I__6593 (
            .O(N__28073),
            .I(N__28069));
    InMux I__6592 (
            .O(N__28072),
            .I(N__28066));
    LocalMux I__6591 (
            .O(N__28069),
            .I(N__28063));
    LocalMux I__6590 (
            .O(N__28066),
            .I(N__28057));
    Span4Mux_h I__6589 (
            .O(N__28063),
            .I(N__28057));
    InMux I__6588 (
            .O(N__28062),
            .I(N__28054));
    Odrv4 I__6587 (
            .O(N__28057),
            .I(\eeprom.n3004 ));
    LocalMux I__6586 (
            .O(N__28054),
            .I(\eeprom.n3004 ));
    CascadeMux I__6585 (
            .O(N__28049),
            .I(N__28046));
    InMux I__6584 (
            .O(N__28046),
            .I(N__28043));
    LocalMux I__6583 (
            .O(N__28043),
            .I(N__28040));
    Odrv4 I__6582 (
            .O(N__28040),
            .I(\eeprom.n3071 ));
    InMux I__6581 (
            .O(N__28037),
            .I(\eeprom.n3663 ));
    InMux I__6580 (
            .O(N__28034),
            .I(N__28031));
    LocalMux I__6579 (
            .O(N__28031),
            .I(N__28027));
    CascadeMux I__6578 (
            .O(N__28030),
            .I(N__28023));
    Span4Mux_v I__6577 (
            .O(N__28027),
            .I(N__28020));
    InMux I__6576 (
            .O(N__28026),
            .I(N__28015));
    InMux I__6575 (
            .O(N__28023),
            .I(N__28015));
    Odrv4 I__6574 (
            .O(N__28020),
            .I(\eeprom.n3003 ));
    LocalMux I__6573 (
            .O(N__28015),
            .I(\eeprom.n3003 ));
    InMux I__6572 (
            .O(N__28010),
            .I(N__28007));
    LocalMux I__6571 (
            .O(N__28007),
            .I(N__28004));
    Span4Mux_h I__6570 (
            .O(N__28004),
            .I(N__28001));
    Odrv4 I__6569 (
            .O(N__28001),
            .I(\eeprom.n3070 ));
    InMux I__6568 (
            .O(N__27998),
            .I(bfn_16_25_0_));
    InMux I__6567 (
            .O(N__27995),
            .I(N__27991));
    InMux I__6566 (
            .O(N__27994),
            .I(N__27988));
    LocalMux I__6565 (
            .O(N__27991),
            .I(N__27984));
    LocalMux I__6564 (
            .O(N__27988),
            .I(N__27981));
    InMux I__6563 (
            .O(N__27987),
            .I(N__27978));
    Span12Mux_s9_v I__6562 (
            .O(N__27984),
            .I(N__27975));
    Span4Mux_v I__6561 (
            .O(N__27981),
            .I(N__27970));
    LocalMux I__6560 (
            .O(N__27978),
            .I(N__27970));
    Odrv12 I__6559 (
            .O(N__27975),
            .I(\eeprom.n3002 ));
    Odrv4 I__6558 (
            .O(N__27970),
            .I(\eeprom.n3002 ));
    CascadeMux I__6557 (
            .O(N__27965),
            .I(N__27962));
    InMux I__6556 (
            .O(N__27962),
            .I(N__27959));
    LocalMux I__6555 (
            .O(N__27959),
            .I(N__27956));
    Span4Mux_v I__6554 (
            .O(N__27956),
            .I(N__27953));
    Odrv4 I__6553 (
            .O(N__27953),
            .I(\eeprom.n3069 ));
    InMux I__6552 (
            .O(N__27950),
            .I(\eeprom.n3665 ));
    InMux I__6551 (
            .O(N__27947),
            .I(N__27944));
    LocalMux I__6550 (
            .O(N__27944),
            .I(N__27940));
    CascadeMux I__6549 (
            .O(N__27943),
            .I(N__27937));
    Span4Mux_h I__6548 (
            .O(N__27940),
            .I(N__27934));
    InMux I__6547 (
            .O(N__27937),
            .I(N__27931));
    Span4Mux_h I__6546 (
            .O(N__27934),
            .I(N__27928));
    LocalMux I__6545 (
            .O(N__27931),
            .I(N__27925));
    Odrv4 I__6544 (
            .O(N__27928),
            .I(\eeprom.n3001 ));
    Odrv4 I__6543 (
            .O(N__27925),
            .I(\eeprom.n3001 ));
    CascadeMux I__6542 (
            .O(N__27920),
            .I(N__27916));
    CascadeMux I__6541 (
            .O(N__27919),
            .I(N__27912));
    InMux I__6540 (
            .O(N__27916),
            .I(N__27904));
    CascadeMux I__6539 (
            .O(N__27915),
            .I(N__27899));
    InMux I__6538 (
            .O(N__27912),
            .I(N__27894));
    InMux I__6537 (
            .O(N__27911),
            .I(N__27894));
    CascadeMux I__6536 (
            .O(N__27910),
            .I(N__27891));
    CascadeMux I__6535 (
            .O(N__27909),
            .I(N__27883));
    CascadeMux I__6534 (
            .O(N__27908),
            .I(N__27878));
    CascadeMux I__6533 (
            .O(N__27907),
            .I(N__27875));
    LocalMux I__6532 (
            .O(N__27904),
            .I(N__27871));
    InMux I__6531 (
            .O(N__27903),
            .I(N__27864));
    InMux I__6530 (
            .O(N__27902),
            .I(N__27864));
    InMux I__6529 (
            .O(N__27899),
            .I(N__27864));
    LocalMux I__6528 (
            .O(N__27894),
            .I(N__27861));
    InMux I__6527 (
            .O(N__27891),
            .I(N__27856));
    InMux I__6526 (
            .O(N__27890),
            .I(N__27856));
    InMux I__6525 (
            .O(N__27889),
            .I(N__27851));
    InMux I__6524 (
            .O(N__27888),
            .I(N__27851));
    InMux I__6523 (
            .O(N__27887),
            .I(N__27848));
    InMux I__6522 (
            .O(N__27886),
            .I(N__27839));
    InMux I__6521 (
            .O(N__27883),
            .I(N__27839));
    InMux I__6520 (
            .O(N__27882),
            .I(N__27839));
    InMux I__6519 (
            .O(N__27881),
            .I(N__27839));
    InMux I__6518 (
            .O(N__27878),
            .I(N__27832));
    InMux I__6517 (
            .O(N__27875),
            .I(N__27832));
    InMux I__6516 (
            .O(N__27874),
            .I(N__27832));
    Span4Mux_h I__6515 (
            .O(N__27871),
            .I(N__27829));
    LocalMux I__6514 (
            .O(N__27864),
            .I(N__27824));
    Span4Mux_h I__6513 (
            .O(N__27861),
            .I(N__27824));
    LocalMux I__6512 (
            .O(N__27856),
            .I(\eeprom.n3034 ));
    LocalMux I__6511 (
            .O(N__27851),
            .I(\eeprom.n3034 ));
    LocalMux I__6510 (
            .O(N__27848),
            .I(\eeprom.n3034 ));
    LocalMux I__6509 (
            .O(N__27839),
            .I(\eeprom.n3034 ));
    LocalMux I__6508 (
            .O(N__27832),
            .I(\eeprom.n3034 ));
    Odrv4 I__6507 (
            .O(N__27829),
            .I(\eeprom.n3034 ));
    Odrv4 I__6506 (
            .O(N__27824),
            .I(\eeprom.n3034 ));
    InMux I__6505 (
            .O(N__27809),
            .I(\eeprom.n3666 ));
    InMux I__6504 (
            .O(N__27806),
            .I(N__27802));
    InMux I__6503 (
            .O(N__27805),
            .I(N__27799));
    LocalMux I__6502 (
            .O(N__27802),
            .I(N__27794));
    LocalMux I__6501 (
            .O(N__27799),
            .I(N__27794));
    Span4Mux_v I__6500 (
            .O(N__27794),
            .I(N__27791));
    Odrv4 I__6499 (
            .O(N__27791),
            .I(\eeprom.n3100 ));
    CascadeMux I__6498 (
            .O(N__27788),
            .I(N__27770));
    CascadeMux I__6497 (
            .O(N__27787),
            .I(N__27762));
    CascadeMux I__6496 (
            .O(N__27786),
            .I(N__27757));
    CascadeMux I__6495 (
            .O(N__27785),
            .I(N__27739));
    CascadeMux I__6494 (
            .O(N__27784),
            .I(N__27736));
    CascadeMux I__6493 (
            .O(N__27783),
            .I(N__27733));
    InMux I__6492 (
            .O(N__27782),
            .I(N__27716));
    InMux I__6491 (
            .O(N__27781),
            .I(N__27716));
    InMux I__6490 (
            .O(N__27780),
            .I(N__27701));
    InMux I__6489 (
            .O(N__27779),
            .I(N__27701));
    InMux I__6488 (
            .O(N__27778),
            .I(N__27694));
    InMux I__6487 (
            .O(N__27777),
            .I(N__27694));
    InMux I__6486 (
            .O(N__27776),
            .I(N__27694));
    InMux I__6485 (
            .O(N__27775),
            .I(N__27683));
    InMux I__6484 (
            .O(N__27774),
            .I(N__27683));
    InMux I__6483 (
            .O(N__27773),
            .I(N__27683));
    InMux I__6482 (
            .O(N__27770),
            .I(N__27683));
    InMux I__6481 (
            .O(N__27769),
            .I(N__27683));
    CascadeMux I__6480 (
            .O(N__27768),
            .I(N__27680));
    CascadeMux I__6479 (
            .O(N__27767),
            .I(N__27677));
    CascadeMux I__6478 (
            .O(N__27766),
            .I(N__27674));
    CascadeMux I__6477 (
            .O(N__27765),
            .I(N__27671));
    InMux I__6476 (
            .O(N__27762),
            .I(N__27659));
    InMux I__6475 (
            .O(N__27761),
            .I(N__27659));
    InMux I__6474 (
            .O(N__27760),
            .I(N__27659));
    InMux I__6473 (
            .O(N__27757),
            .I(N__27659));
    InMux I__6472 (
            .O(N__27756),
            .I(N__27659));
    InMux I__6471 (
            .O(N__27755),
            .I(N__27654));
    InMux I__6470 (
            .O(N__27754),
            .I(N__27654));
    CascadeMux I__6469 (
            .O(N__27753),
            .I(N__27650));
    CascadeMux I__6468 (
            .O(N__27752),
            .I(N__27644));
    CascadeMux I__6467 (
            .O(N__27751),
            .I(N__27638));
    CascadeMux I__6466 (
            .O(N__27750),
            .I(N__27635));
    InMux I__6465 (
            .O(N__27749),
            .I(N__27630));
    InMux I__6464 (
            .O(N__27748),
            .I(N__27630));
    CascadeMux I__6463 (
            .O(N__27747),
            .I(N__27624));
    CascadeMux I__6462 (
            .O(N__27746),
            .I(N__27621));
    CascadeMux I__6461 (
            .O(N__27745),
            .I(N__27617));
    CascadeMux I__6460 (
            .O(N__27744),
            .I(N__27614));
    CascadeMux I__6459 (
            .O(N__27743),
            .I(N__27608));
    InMux I__6458 (
            .O(N__27742),
            .I(N__27599));
    InMux I__6457 (
            .O(N__27739),
            .I(N__27599));
    InMux I__6456 (
            .O(N__27736),
            .I(N__27596));
    InMux I__6455 (
            .O(N__27733),
            .I(N__27591));
    InMux I__6454 (
            .O(N__27732),
            .I(N__27591));
    InMux I__6453 (
            .O(N__27731),
            .I(N__27583));
    InMux I__6452 (
            .O(N__27730),
            .I(N__27578));
    CascadeMux I__6451 (
            .O(N__27729),
            .I(N__27575));
    InMux I__6450 (
            .O(N__27728),
            .I(N__27570));
    InMux I__6449 (
            .O(N__27727),
            .I(N__27570));
    CascadeMux I__6448 (
            .O(N__27726),
            .I(N__27566));
    CascadeMux I__6447 (
            .O(N__27725),
            .I(N__27561));
    CascadeMux I__6446 (
            .O(N__27724),
            .I(N__27557));
    CascadeMux I__6445 (
            .O(N__27723),
            .I(N__27553));
    CascadeMux I__6444 (
            .O(N__27722),
            .I(N__27550));
    CascadeMux I__6443 (
            .O(N__27721),
            .I(N__27547));
    LocalMux I__6442 (
            .O(N__27716),
            .I(N__27538));
    InMux I__6441 (
            .O(N__27715),
            .I(N__27529));
    InMux I__6440 (
            .O(N__27714),
            .I(N__27529));
    InMux I__6439 (
            .O(N__27713),
            .I(N__27529));
    InMux I__6438 (
            .O(N__27712),
            .I(N__27529));
    InMux I__6437 (
            .O(N__27711),
            .I(N__27520));
    InMux I__6436 (
            .O(N__27710),
            .I(N__27520));
    InMux I__6435 (
            .O(N__27709),
            .I(N__27520));
    InMux I__6434 (
            .O(N__27708),
            .I(N__27520));
    CascadeMux I__6433 (
            .O(N__27707),
            .I(N__27515));
    CascadeMux I__6432 (
            .O(N__27706),
            .I(N__27510));
    LocalMux I__6431 (
            .O(N__27701),
            .I(N__27504));
    LocalMux I__6430 (
            .O(N__27694),
            .I(N__27504));
    LocalMux I__6429 (
            .O(N__27683),
            .I(N__27501));
    InMux I__6428 (
            .O(N__27680),
            .I(N__27490));
    InMux I__6427 (
            .O(N__27677),
            .I(N__27490));
    InMux I__6426 (
            .O(N__27674),
            .I(N__27490));
    InMux I__6425 (
            .O(N__27671),
            .I(N__27490));
    InMux I__6424 (
            .O(N__27670),
            .I(N__27490));
    LocalMux I__6423 (
            .O(N__27659),
            .I(N__27485));
    LocalMux I__6422 (
            .O(N__27654),
            .I(N__27485));
    InMux I__6421 (
            .O(N__27653),
            .I(N__27476));
    InMux I__6420 (
            .O(N__27650),
            .I(N__27476));
    InMux I__6419 (
            .O(N__27649),
            .I(N__27476));
    InMux I__6418 (
            .O(N__27648),
            .I(N__27476));
    InMux I__6417 (
            .O(N__27647),
            .I(N__27467));
    InMux I__6416 (
            .O(N__27644),
            .I(N__27467));
    InMux I__6415 (
            .O(N__27643),
            .I(N__27467));
    InMux I__6414 (
            .O(N__27642),
            .I(N__27467));
    InMux I__6413 (
            .O(N__27641),
            .I(N__27460));
    InMux I__6412 (
            .O(N__27638),
            .I(N__27460));
    InMux I__6411 (
            .O(N__27635),
            .I(N__27460));
    LocalMux I__6410 (
            .O(N__27630),
            .I(N__27456));
    InMux I__6409 (
            .O(N__27629),
            .I(N__27453));
    InMux I__6408 (
            .O(N__27628),
            .I(N__27448));
    InMux I__6407 (
            .O(N__27627),
            .I(N__27448));
    InMux I__6406 (
            .O(N__27624),
            .I(N__27443));
    InMux I__6405 (
            .O(N__27621),
            .I(N__27443));
    InMux I__6404 (
            .O(N__27620),
            .I(N__27436));
    InMux I__6403 (
            .O(N__27617),
            .I(N__27436));
    InMux I__6402 (
            .O(N__27614),
            .I(N__27436));
    InMux I__6401 (
            .O(N__27613),
            .I(N__27431));
    InMux I__6400 (
            .O(N__27612),
            .I(N__27431));
    InMux I__6399 (
            .O(N__27611),
            .I(N__27428));
    InMux I__6398 (
            .O(N__27608),
            .I(N__27423));
    InMux I__6397 (
            .O(N__27607),
            .I(N__27423));
    CascadeMux I__6396 (
            .O(N__27606),
            .I(N__27418));
    CascadeMux I__6395 (
            .O(N__27605),
            .I(N__27415));
    CascadeMux I__6394 (
            .O(N__27604),
            .I(N__27412));
    LocalMux I__6393 (
            .O(N__27599),
            .I(N__27407));
    LocalMux I__6392 (
            .O(N__27596),
            .I(N__27402));
    LocalMux I__6391 (
            .O(N__27591),
            .I(N__27402));
    InMux I__6390 (
            .O(N__27590),
            .I(N__27397));
    InMux I__6389 (
            .O(N__27589),
            .I(N__27397));
    CascadeMux I__6388 (
            .O(N__27588),
            .I(N__27394));
    CascadeMux I__6387 (
            .O(N__27587),
            .I(N__27390));
    CascadeMux I__6386 (
            .O(N__27586),
            .I(N__27387));
    LocalMux I__6385 (
            .O(N__27583),
            .I(N__27378));
    InMux I__6384 (
            .O(N__27582),
            .I(N__27375));
    CascadeMux I__6383 (
            .O(N__27581),
            .I(N__27372));
    LocalMux I__6382 (
            .O(N__27578),
            .I(N__27368));
    InMux I__6381 (
            .O(N__27575),
            .I(N__27365));
    LocalMux I__6380 (
            .O(N__27570),
            .I(N__27362));
    InMux I__6379 (
            .O(N__27569),
            .I(N__27357));
    InMux I__6378 (
            .O(N__27566),
            .I(N__27357));
    InMux I__6377 (
            .O(N__27565),
            .I(N__27348));
    InMux I__6376 (
            .O(N__27564),
            .I(N__27348));
    InMux I__6375 (
            .O(N__27561),
            .I(N__27348));
    InMux I__6374 (
            .O(N__27560),
            .I(N__27348));
    InMux I__6373 (
            .O(N__27557),
            .I(N__27345));
    InMux I__6372 (
            .O(N__27556),
            .I(N__27342));
    InMux I__6371 (
            .O(N__27553),
            .I(N__27335));
    InMux I__6370 (
            .O(N__27550),
            .I(N__27335));
    InMux I__6369 (
            .O(N__27547),
            .I(N__27335));
    CascadeMux I__6368 (
            .O(N__27546),
            .I(N__27327));
    CascadeMux I__6367 (
            .O(N__27545),
            .I(N__27322));
    CascadeMux I__6366 (
            .O(N__27544),
            .I(N__27319));
    CascadeMux I__6365 (
            .O(N__27543),
            .I(N__27315));
    CascadeMux I__6364 (
            .O(N__27542),
            .I(N__27312));
    CascadeMux I__6363 (
            .O(N__27541),
            .I(N__27307));
    Span4Mux_v I__6362 (
            .O(N__27538),
            .I(N__27295));
    LocalMux I__6361 (
            .O(N__27529),
            .I(N__27295));
    LocalMux I__6360 (
            .O(N__27520),
            .I(N__27295));
    InMux I__6359 (
            .O(N__27519),
            .I(N__27290));
    InMux I__6358 (
            .O(N__27518),
            .I(N__27290));
    InMux I__6357 (
            .O(N__27515),
            .I(N__27279));
    InMux I__6356 (
            .O(N__27514),
            .I(N__27279));
    InMux I__6355 (
            .O(N__27513),
            .I(N__27279));
    InMux I__6354 (
            .O(N__27510),
            .I(N__27279));
    InMux I__6353 (
            .O(N__27509),
            .I(N__27279));
    Span4Mux_h I__6352 (
            .O(N__27504),
            .I(N__27272));
    Span4Mux_h I__6351 (
            .O(N__27501),
            .I(N__27272));
    LocalMux I__6350 (
            .O(N__27490),
            .I(N__27272));
    Span4Mux_v I__6349 (
            .O(N__27485),
            .I(N__27263));
    LocalMux I__6348 (
            .O(N__27476),
            .I(N__27263));
    LocalMux I__6347 (
            .O(N__27467),
            .I(N__27263));
    LocalMux I__6346 (
            .O(N__27460),
            .I(N__27263));
    InMux I__6345 (
            .O(N__27459),
            .I(N__27260));
    Span4Mux_v I__6344 (
            .O(N__27456),
            .I(N__27255));
    LocalMux I__6343 (
            .O(N__27453),
            .I(N__27255));
    LocalMux I__6342 (
            .O(N__27448),
            .I(N__27252));
    LocalMux I__6341 (
            .O(N__27443),
            .I(N__27247));
    LocalMux I__6340 (
            .O(N__27436),
            .I(N__27247));
    LocalMux I__6339 (
            .O(N__27431),
            .I(N__27240));
    LocalMux I__6338 (
            .O(N__27428),
            .I(N__27240));
    LocalMux I__6337 (
            .O(N__27423),
            .I(N__27240));
    InMux I__6336 (
            .O(N__27422),
            .I(N__27235));
    InMux I__6335 (
            .O(N__27421),
            .I(N__27235));
    InMux I__6334 (
            .O(N__27418),
            .I(N__27226));
    InMux I__6333 (
            .O(N__27415),
            .I(N__27226));
    InMux I__6332 (
            .O(N__27412),
            .I(N__27226));
    InMux I__6331 (
            .O(N__27411),
            .I(N__27226));
    InMux I__6330 (
            .O(N__27410),
            .I(N__27223));
    Span4Mux_s3_h I__6329 (
            .O(N__27407),
            .I(N__27218));
    Span4Mux_v I__6328 (
            .O(N__27402),
            .I(N__27218));
    LocalMux I__6327 (
            .O(N__27397),
            .I(N__27215));
    InMux I__6326 (
            .O(N__27394),
            .I(N__27206));
    InMux I__6325 (
            .O(N__27393),
            .I(N__27206));
    InMux I__6324 (
            .O(N__27390),
            .I(N__27206));
    InMux I__6323 (
            .O(N__27387),
            .I(N__27206));
    CascadeMux I__6322 (
            .O(N__27386),
            .I(N__27202));
    CascadeMux I__6321 (
            .O(N__27385),
            .I(N__27199));
    CascadeMux I__6320 (
            .O(N__27384),
            .I(N__27196));
    InMux I__6319 (
            .O(N__27383),
            .I(N__27182));
    CascadeMux I__6318 (
            .O(N__27382),
            .I(N__27176));
    CascadeMux I__6317 (
            .O(N__27381),
            .I(N__27171));
    Span4Mux_v I__6316 (
            .O(N__27378),
            .I(N__27166));
    LocalMux I__6315 (
            .O(N__27375),
            .I(N__27166));
    InMux I__6314 (
            .O(N__27372),
            .I(N__27163));
    InMux I__6313 (
            .O(N__27371),
            .I(N__27160));
    Span4Mux_v I__6312 (
            .O(N__27368),
            .I(N__27155));
    LocalMux I__6311 (
            .O(N__27365),
            .I(N__27155));
    Span4Mux_v I__6310 (
            .O(N__27362),
            .I(N__27142));
    LocalMux I__6309 (
            .O(N__27357),
            .I(N__27142));
    LocalMux I__6308 (
            .O(N__27348),
            .I(N__27142));
    LocalMux I__6307 (
            .O(N__27345),
            .I(N__27142));
    LocalMux I__6306 (
            .O(N__27342),
            .I(N__27142));
    LocalMux I__6305 (
            .O(N__27335),
            .I(N__27142));
    CascadeMux I__6304 (
            .O(N__27334),
            .I(N__27139));
    CascadeMux I__6303 (
            .O(N__27333),
            .I(N__27136));
    CascadeMux I__6302 (
            .O(N__27332),
            .I(N__27133));
    CascadeMux I__6301 (
            .O(N__27331),
            .I(N__27130));
    CascadeMux I__6300 (
            .O(N__27330),
            .I(N__27127));
    InMux I__6299 (
            .O(N__27327),
            .I(N__27123));
    InMux I__6298 (
            .O(N__27326),
            .I(N__27118));
    InMux I__6297 (
            .O(N__27325),
            .I(N__27118));
    InMux I__6296 (
            .O(N__27322),
            .I(N__27109));
    InMux I__6295 (
            .O(N__27319),
            .I(N__27109));
    InMux I__6294 (
            .O(N__27318),
            .I(N__27109));
    InMux I__6293 (
            .O(N__27315),
            .I(N__27109));
    InMux I__6292 (
            .O(N__27312),
            .I(N__27106));
    InMux I__6291 (
            .O(N__27311),
            .I(N__27103));
    InMux I__6290 (
            .O(N__27310),
            .I(N__27098));
    InMux I__6289 (
            .O(N__27307),
            .I(N__27098));
    CascadeMux I__6288 (
            .O(N__27306),
            .I(N__27095));
    CascadeMux I__6287 (
            .O(N__27305),
            .I(N__27092));
    CascadeMux I__6286 (
            .O(N__27304),
            .I(N__27088));
    CascadeMux I__6285 (
            .O(N__27303),
            .I(N__27085));
    CascadeMux I__6284 (
            .O(N__27302),
            .I(N__27081));
    Span4Mux_h I__6283 (
            .O(N__27295),
            .I(N__27066));
    LocalMux I__6282 (
            .O(N__27290),
            .I(N__27066));
    LocalMux I__6281 (
            .O(N__27279),
            .I(N__27066));
    Span4Mux_v I__6280 (
            .O(N__27272),
            .I(N__27059));
    Span4Mux_h I__6279 (
            .O(N__27263),
            .I(N__27059));
    LocalMux I__6278 (
            .O(N__27260),
            .I(N__27059));
    Span4Mux_v I__6277 (
            .O(N__27255),
            .I(N__27048));
    Span4Mux_v I__6276 (
            .O(N__27252),
            .I(N__27048));
    Span4Mux_h I__6275 (
            .O(N__27247),
            .I(N__27048));
    Span4Mux_v I__6274 (
            .O(N__27240),
            .I(N__27048));
    LocalMux I__6273 (
            .O(N__27235),
            .I(N__27048));
    LocalMux I__6272 (
            .O(N__27226),
            .I(N__27043));
    LocalMux I__6271 (
            .O(N__27223),
            .I(N__27043));
    Span4Mux_h I__6270 (
            .O(N__27218),
            .I(N__27036));
    Span4Mux_v I__6269 (
            .O(N__27215),
            .I(N__27036));
    LocalMux I__6268 (
            .O(N__27206),
            .I(N__27036));
    InMux I__6267 (
            .O(N__27205),
            .I(N__27031));
    InMux I__6266 (
            .O(N__27202),
            .I(N__27031));
    InMux I__6265 (
            .O(N__27199),
            .I(N__27026));
    InMux I__6264 (
            .O(N__27196),
            .I(N__27026));
    CascadeMux I__6263 (
            .O(N__27195),
            .I(N__27021));
    CascadeMux I__6262 (
            .O(N__27194),
            .I(N__27018));
    CascadeMux I__6261 (
            .O(N__27193),
            .I(N__27013));
    CascadeMux I__6260 (
            .O(N__27192),
            .I(N__27010));
    CascadeMux I__6259 (
            .O(N__27191),
            .I(N__27005));
    CascadeMux I__6258 (
            .O(N__27190),
            .I(N__27002));
    CascadeMux I__6257 (
            .O(N__27189),
            .I(N__26999));
    CascadeMux I__6256 (
            .O(N__27188),
            .I(N__26995));
    CascadeMux I__6255 (
            .O(N__27187),
            .I(N__26992));
    CascadeMux I__6254 (
            .O(N__27186),
            .I(N__26989));
    CascadeMux I__6253 (
            .O(N__27185),
            .I(N__26984));
    LocalMux I__6252 (
            .O(N__27182),
            .I(N__26981));
    InMux I__6251 (
            .O(N__27181),
            .I(N__26978));
    InMux I__6250 (
            .O(N__27180),
            .I(N__26973));
    InMux I__6249 (
            .O(N__27179),
            .I(N__26973));
    InMux I__6248 (
            .O(N__27176),
            .I(N__26964));
    InMux I__6247 (
            .O(N__27175),
            .I(N__26964));
    InMux I__6246 (
            .O(N__27174),
            .I(N__26964));
    InMux I__6245 (
            .O(N__27171),
            .I(N__26964));
    Sp12to4 I__6244 (
            .O(N__27166),
            .I(N__26957));
    LocalMux I__6243 (
            .O(N__27163),
            .I(N__26957));
    LocalMux I__6242 (
            .O(N__27160),
            .I(N__26957));
    Span4Mux_h I__6241 (
            .O(N__27155),
            .I(N__26952));
    Span4Mux_v I__6240 (
            .O(N__27142),
            .I(N__26952));
    InMux I__6239 (
            .O(N__27139),
            .I(N__26947));
    InMux I__6238 (
            .O(N__27136),
            .I(N__26947));
    InMux I__6237 (
            .O(N__27133),
            .I(N__26938));
    InMux I__6236 (
            .O(N__27130),
            .I(N__26938));
    InMux I__6235 (
            .O(N__27127),
            .I(N__26938));
    InMux I__6234 (
            .O(N__27126),
            .I(N__26938));
    LocalMux I__6233 (
            .O(N__27123),
            .I(N__26933));
    LocalMux I__6232 (
            .O(N__27118),
            .I(N__26922));
    LocalMux I__6231 (
            .O(N__27109),
            .I(N__26922));
    LocalMux I__6230 (
            .O(N__27106),
            .I(N__26922));
    LocalMux I__6229 (
            .O(N__27103),
            .I(N__26922));
    LocalMux I__6228 (
            .O(N__27098),
            .I(N__26922));
    InMux I__6227 (
            .O(N__27095),
            .I(N__26919));
    InMux I__6226 (
            .O(N__27092),
            .I(N__26904));
    InMux I__6225 (
            .O(N__27091),
            .I(N__26904));
    InMux I__6224 (
            .O(N__27088),
            .I(N__26904));
    InMux I__6223 (
            .O(N__27085),
            .I(N__26904));
    InMux I__6222 (
            .O(N__27084),
            .I(N__26904));
    InMux I__6221 (
            .O(N__27081),
            .I(N__26904));
    InMux I__6220 (
            .O(N__27080),
            .I(N__26904));
    CascadeMux I__6219 (
            .O(N__27079),
            .I(N__26901));
    CascadeMux I__6218 (
            .O(N__27078),
            .I(N__26898));
    CascadeMux I__6217 (
            .O(N__27077),
            .I(N__26895));
    CascadeMux I__6216 (
            .O(N__27076),
            .I(N__26892));
    CascadeMux I__6215 (
            .O(N__27075),
            .I(N__26889));
    CascadeMux I__6214 (
            .O(N__27074),
            .I(N__26886));
    CascadeMux I__6213 (
            .O(N__27073),
            .I(N__26882));
    Span4Mux_v I__6212 (
            .O(N__27066),
            .I(N__26877));
    Span4Mux_v I__6211 (
            .O(N__27059),
            .I(N__26870));
    Span4Mux_h I__6210 (
            .O(N__27048),
            .I(N__26870));
    Span4Mux_v I__6209 (
            .O(N__27043),
            .I(N__26870));
    Span4Mux_h I__6208 (
            .O(N__27036),
            .I(N__26863));
    LocalMux I__6207 (
            .O(N__27031),
            .I(N__26863));
    LocalMux I__6206 (
            .O(N__27026),
            .I(N__26863));
    InMux I__6205 (
            .O(N__27025),
            .I(N__26858));
    InMux I__6204 (
            .O(N__27024),
            .I(N__26858));
    InMux I__6203 (
            .O(N__27021),
            .I(N__26849));
    InMux I__6202 (
            .O(N__27018),
            .I(N__26849));
    InMux I__6201 (
            .O(N__27017),
            .I(N__26849));
    InMux I__6200 (
            .O(N__27016),
            .I(N__26849));
    InMux I__6199 (
            .O(N__27013),
            .I(N__26840));
    InMux I__6198 (
            .O(N__27010),
            .I(N__26840));
    InMux I__6197 (
            .O(N__27009),
            .I(N__26840));
    InMux I__6196 (
            .O(N__27008),
            .I(N__26840));
    InMux I__6195 (
            .O(N__27005),
            .I(N__26833));
    InMux I__6194 (
            .O(N__27002),
            .I(N__26833));
    InMux I__6193 (
            .O(N__26999),
            .I(N__26833));
    InMux I__6192 (
            .O(N__26998),
            .I(N__26822));
    InMux I__6191 (
            .O(N__26995),
            .I(N__26822));
    InMux I__6190 (
            .O(N__26992),
            .I(N__26822));
    InMux I__6189 (
            .O(N__26989),
            .I(N__26822));
    InMux I__6188 (
            .O(N__26988),
            .I(N__26822));
    InMux I__6187 (
            .O(N__26987),
            .I(N__26817));
    InMux I__6186 (
            .O(N__26984),
            .I(N__26817));
    Span12Mux_v I__6185 (
            .O(N__26981),
            .I(N__26800));
    LocalMux I__6184 (
            .O(N__26978),
            .I(N__26800));
    LocalMux I__6183 (
            .O(N__26973),
            .I(N__26800));
    LocalMux I__6182 (
            .O(N__26964),
            .I(N__26800));
    Span12Mux_s10_v I__6181 (
            .O(N__26957),
            .I(N__26800));
    Sp12to4 I__6180 (
            .O(N__26952),
            .I(N__26800));
    LocalMux I__6179 (
            .O(N__26947),
            .I(N__26800));
    LocalMux I__6178 (
            .O(N__26938),
            .I(N__26800));
    InMux I__6177 (
            .O(N__26937),
            .I(N__26795));
    InMux I__6176 (
            .O(N__26936),
            .I(N__26795));
    Span4Mux_h I__6175 (
            .O(N__26933),
            .I(N__26786));
    Span4Mux_v I__6174 (
            .O(N__26922),
            .I(N__26786));
    LocalMux I__6173 (
            .O(N__26919),
            .I(N__26786));
    LocalMux I__6172 (
            .O(N__26904),
            .I(N__26786));
    InMux I__6171 (
            .O(N__26901),
            .I(N__26779));
    InMux I__6170 (
            .O(N__26898),
            .I(N__26779));
    InMux I__6169 (
            .O(N__26895),
            .I(N__26779));
    InMux I__6168 (
            .O(N__26892),
            .I(N__26768));
    InMux I__6167 (
            .O(N__26889),
            .I(N__26768));
    InMux I__6166 (
            .O(N__26886),
            .I(N__26768));
    InMux I__6165 (
            .O(N__26885),
            .I(N__26768));
    InMux I__6164 (
            .O(N__26882),
            .I(N__26768));
    CascadeMux I__6163 (
            .O(N__26881),
            .I(N__26765));
    CascadeMux I__6162 (
            .O(N__26880),
            .I(N__26761));
    Span4Mux_v I__6161 (
            .O(N__26877),
            .I(N__26756));
    Span4Mux_h I__6160 (
            .O(N__26870),
            .I(N__26756));
    Span4Mux_h I__6159 (
            .O(N__26863),
            .I(N__26753));
    LocalMux I__6158 (
            .O(N__26858),
            .I(N__26740));
    LocalMux I__6157 (
            .O(N__26849),
            .I(N__26740));
    LocalMux I__6156 (
            .O(N__26840),
            .I(N__26740));
    LocalMux I__6155 (
            .O(N__26833),
            .I(N__26740));
    LocalMux I__6154 (
            .O(N__26822),
            .I(N__26740));
    LocalMux I__6153 (
            .O(N__26817),
            .I(N__26740));
    Span12Mux_h I__6152 (
            .O(N__26800),
            .I(N__26735));
    LocalMux I__6151 (
            .O(N__26795),
            .I(N__26735));
    Span4Mux_h I__6150 (
            .O(N__26786),
            .I(N__26728));
    LocalMux I__6149 (
            .O(N__26779),
            .I(N__26728));
    LocalMux I__6148 (
            .O(N__26768),
            .I(N__26728));
    InMux I__6147 (
            .O(N__26765),
            .I(N__26725));
    InMux I__6146 (
            .O(N__26764),
            .I(N__26720));
    InMux I__6145 (
            .O(N__26761),
            .I(N__26720));
    Odrv4 I__6144 (
            .O(N__26756),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__6143 (
            .O(N__26753),
            .I(CONSTANT_ONE_NET));
    Odrv12 I__6142 (
            .O(N__26740),
            .I(CONSTANT_ONE_NET));
    Odrv12 I__6141 (
            .O(N__26735),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__6140 (
            .O(N__26728),
            .I(CONSTANT_ONE_NET));
    LocalMux I__6139 (
            .O(N__26725),
            .I(CONSTANT_ONE_NET));
    LocalMux I__6138 (
            .O(N__26720),
            .I(CONSTANT_ONE_NET));
    CascadeMux I__6137 (
            .O(N__26705),
            .I(N__26700));
    InMux I__6136 (
            .O(N__26704),
            .I(N__26697));
    InMux I__6135 (
            .O(N__26703),
            .I(N__26694));
    InMux I__6134 (
            .O(N__26700),
            .I(N__26691));
    LocalMux I__6133 (
            .O(N__26697),
            .I(N__26684));
    LocalMux I__6132 (
            .O(N__26694),
            .I(N__26684));
    LocalMux I__6131 (
            .O(N__26691),
            .I(N__26684));
    Odrv12 I__6130 (
            .O(N__26684),
            .I(\eeprom.n3012 ));
    InMux I__6129 (
            .O(N__26681),
            .I(N__26678));
    LocalMux I__6128 (
            .O(N__26678),
            .I(\eeprom.n3079 ));
    InMux I__6127 (
            .O(N__26675),
            .I(\eeprom.n3655 ));
    InMux I__6126 (
            .O(N__26672),
            .I(N__26668));
    InMux I__6125 (
            .O(N__26671),
            .I(N__26664));
    LocalMux I__6124 (
            .O(N__26668),
            .I(N__26661));
    InMux I__6123 (
            .O(N__26667),
            .I(N__26658));
    LocalMux I__6122 (
            .O(N__26664),
            .I(\eeprom.n3011 ));
    Odrv4 I__6121 (
            .O(N__26661),
            .I(\eeprom.n3011 ));
    LocalMux I__6120 (
            .O(N__26658),
            .I(\eeprom.n3011 ));
    CascadeMux I__6119 (
            .O(N__26651),
            .I(N__26648));
    InMux I__6118 (
            .O(N__26648),
            .I(N__26645));
    LocalMux I__6117 (
            .O(N__26645),
            .I(\eeprom.n3078 ));
    InMux I__6116 (
            .O(N__26642),
            .I(bfn_16_24_0_));
    InMux I__6115 (
            .O(N__26639),
            .I(N__26636));
    LocalMux I__6114 (
            .O(N__26636),
            .I(N__26631));
    InMux I__6113 (
            .O(N__26635),
            .I(N__26628));
    CascadeMux I__6112 (
            .O(N__26634),
            .I(N__26625));
    Span4Mux_h I__6111 (
            .O(N__26631),
            .I(N__26620));
    LocalMux I__6110 (
            .O(N__26628),
            .I(N__26620));
    InMux I__6109 (
            .O(N__26625),
            .I(N__26617));
    Span4Mux_h I__6108 (
            .O(N__26620),
            .I(N__26614));
    LocalMux I__6107 (
            .O(N__26617),
            .I(N__26611));
    Odrv4 I__6106 (
            .O(N__26614),
            .I(\eeprom.n3010 ));
    Odrv12 I__6105 (
            .O(N__26611),
            .I(\eeprom.n3010 ));
    CascadeMux I__6104 (
            .O(N__26606),
            .I(N__26603));
    InMux I__6103 (
            .O(N__26603),
            .I(N__26600));
    LocalMux I__6102 (
            .O(N__26600),
            .I(\eeprom.n3077 ));
    InMux I__6101 (
            .O(N__26597),
            .I(\eeprom.n3657 ));
    InMux I__6100 (
            .O(N__26594),
            .I(N__26590));
    InMux I__6099 (
            .O(N__26593),
            .I(N__26587));
    LocalMux I__6098 (
            .O(N__26590),
            .I(N__26583));
    LocalMux I__6097 (
            .O(N__26587),
            .I(N__26580));
    InMux I__6096 (
            .O(N__26586),
            .I(N__26577));
    Span4Mux_h I__6095 (
            .O(N__26583),
            .I(N__26574));
    Span4Mux_h I__6094 (
            .O(N__26580),
            .I(N__26571));
    LocalMux I__6093 (
            .O(N__26577),
            .I(N__26568));
    Odrv4 I__6092 (
            .O(N__26574),
            .I(\eeprom.n3009 ));
    Odrv4 I__6091 (
            .O(N__26571),
            .I(\eeprom.n3009 ));
    Odrv12 I__6090 (
            .O(N__26568),
            .I(\eeprom.n3009 ));
    CascadeMux I__6089 (
            .O(N__26561),
            .I(N__26558));
    InMux I__6088 (
            .O(N__26558),
            .I(N__26555));
    LocalMux I__6087 (
            .O(N__26555),
            .I(N__26552));
    Span4Mux_h I__6086 (
            .O(N__26552),
            .I(N__26549));
    Odrv4 I__6085 (
            .O(N__26549),
            .I(\eeprom.n3076 ));
    InMux I__6084 (
            .O(N__26546),
            .I(\eeprom.n3658 ));
    CascadeMux I__6083 (
            .O(N__26543),
            .I(N__26540));
    InMux I__6082 (
            .O(N__26540),
            .I(N__26535));
    InMux I__6081 (
            .O(N__26539),
            .I(N__26532));
    InMux I__6080 (
            .O(N__26538),
            .I(N__26529));
    LocalMux I__6079 (
            .O(N__26535),
            .I(\eeprom.n3008 ));
    LocalMux I__6078 (
            .O(N__26532),
            .I(\eeprom.n3008 ));
    LocalMux I__6077 (
            .O(N__26529),
            .I(\eeprom.n3008 ));
    InMux I__6076 (
            .O(N__26522),
            .I(N__26519));
    LocalMux I__6075 (
            .O(N__26519),
            .I(\eeprom.n3075 ));
    InMux I__6074 (
            .O(N__26516),
            .I(\eeprom.n3659 ));
    InMux I__6073 (
            .O(N__26513),
            .I(N__26508));
    InMux I__6072 (
            .O(N__26512),
            .I(N__26505));
    InMux I__6071 (
            .O(N__26511),
            .I(N__26502));
    LocalMux I__6070 (
            .O(N__26508),
            .I(N__26499));
    LocalMux I__6069 (
            .O(N__26505),
            .I(N__26496));
    LocalMux I__6068 (
            .O(N__26502),
            .I(N__26493));
    Span4Mux_h I__6067 (
            .O(N__26499),
            .I(N__26490));
    Odrv4 I__6066 (
            .O(N__26496),
            .I(\eeprom.n3007 ));
    Odrv12 I__6065 (
            .O(N__26493),
            .I(\eeprom.n3007 ));
    Odrv4 I__6064 (
            .O(N__26490),
            .I(\eeprom.n3007 ));
    CascadeMux I__6063 (
            .O(N__26483),
            .I(N__26480));
    InMux I__6062 (
            .O(N__26480),
            .I(N__26477));
    LocalMux I__6061 (
            .O(N__26477),
            .I(N__26474));
    Odrv4 I__6060 (
            .O(N__26474),
            .I(\eeprom.n3074 ));
    InMux I__6059 (
            .O(N__26471),
            .I(\eeprom.n3660 ));
    InMux I__6058 (
            .O(N__26468),
            .I(N__26464));
    InMux I__6057 (
            .O(N__26467),
            .I(N__26461));
    LocalMux I__6056 (
            .O(N__26464),
            .I(N__26457));
    LocalMux I__6055 (
            .O(N__26461),
            .I(N__26454));
    InMux I__6054 (
            .O(N__26460),
            .I(N__26451));
    Odrv4 I__6053 (
            .O(N__26457),
            .I(\eeprom.n3006 ));
    Odrv4 I__6052 (
            .O(N__26454),
            .I(\eeprom.n3006 ));
    LocalMux I__6051 (
            .O(N__26451),
            .I(\eeprom.n3006 ));
    CascadeMux I__6050 (
            .O(N__26444),
            .I(N__26441));
    InMux I__6049 (
            .O(N__26441),
            .I(N__26438));
    LocalMux I__6048 (
            .O(N__26438),
            .I(N__26435));
    Span4Mux_v I__6047 (
            .O(N__26435),
            .I(N__26432));
    Odrv4 I__6046 (
            .O(N__26432),
            .I(\eeprom.n3073 ));
    InMux I__6045 (
            .O(N__26429),
            .I(\eeprom.n3661 ));
    InMux I__6044 (
            .O(N__26426),
            .I(N__26423));
    LocalMux I__6043 (
            .O(N__26423),
            .I(N__26420));
    Span4Mux_h I__6042 (
            .O(N__26420),
            .I(N__26415));
    InMux I__6041 (
            .O(N__26419),
            .I(N__26410));
    InMux I__6040 (
            .O(N__26418),
            .I(N__26410));
    Span4Mux_h I__6039 (
            .O(N__26415),
            .I(N__26407));
    LocalMux I__6038 (
            .O(N__26410),
            .I(N__26404));
    Odrv4 I__6037 (
            .O(N__26407),
            .I(\eeprom.n3005 ));
    Odrv4 I__6036 (
            .O(N__26404),
            .I(\eeprom.n3005 ));
    CascadeMux I__6035 (
            .O(N__26399),
            .I(\eeprom.n4766_cascade_ ));
    InMux I__6034 (
            .O(N__26396),
            .I(N__26393));
    LocalMux I__6033 (
            .O(N__26393),
            .I(\eeprom.n4903 ));
    InMux I__6032 (
            .O(N__26390),
            .I(N__26387));
    LocalMux I__6031 (
            .O(N__26387),
            .I(N__26382));
    InMux I__6030 (
            .O(N__26386),
            .I(N__26379));
    InMux I__6029 (
            .O(N__26385),
            .I(N__26376));
    Span4Mux_v I__6028 (
            .O(N__26382),
            .I(N__26369));
    LocalMux I__6027 (
            .O(N__26379),
            .I(N__26369));
    LocalMux I__6026 (
            .O(N__26376),
            .I(N__26369));
    Span4Mux_h I__6025 (
            .O(N__26369),
            .I(N__26366));
    Span4Mux_h I__6024 (
            .O(N__26366),
            .I(N__26363));
    Span4Mux_h I__6023 (
            .O(N__26363),
            .I(N__26360));
    Span4Mux_h I__6022 (
            .O(N__26360),
            .I(N__26357));
    Odrv4 I__6021 (
            .O(N__26357),
            .I(\eeprom.n3019 ));
    InMux I__6020 (
            .O(N__26354),
            .I(N__26351));
    LocalMux I__6019 (
            .O(N__26351),
            .I(N__26348));
    Span4Mux_v I__6018 (
            .O(N__26348),
            .I(N__26345));
    Odrv4 I__6017 (
            .O(N__26345),
            .I(\eeprom.n3086 ));
    InMux I__6016 (
            .O(N__26342),
            .I(bfn_16_23_0_));
    InMux I__6015 (
            .O(N__26339),
            .I(N__26336));
    LocalMux I__6014 (
            .O(N__26336),
            .I(N__26332));
    CascadeMux I__6013 (
            .O(N__26335),
            .I(N__26328));
    Span4Mux_h I__6012 (
            .O(N__26332),
            .I(N__26325));
    InMux I__6011 (
            .O(N__26331),
            .I(N__26322));
    InMux I__6010 (
            .O(N__26328),
            .I(N__26319));
    Odrv4 I__6009 (
            .O(N__26325),
            .I(\eeprom.n3018 ));
    LocalMux I__6008 (
            .O(N__26322),
            .I(\eeprom.n3018 ));
    LocalMux I__6007 (
            .O(N__26319),
            .I(\eeprom.n3018 ));
    InMux I__6006 (
            .O(N__26312),
            .I(N__26309));
    LocalMux I__6005 (
            .O(N__26309),
            .I(N__26306));
    Span4Mux_h I__6004 (
            .O(N__26306),
            .I(N__26303));
    Odrv4 I__6003 (
            .O(N__26303),
            .I(\eeprom.n3085 ));
    InMux I__6002 (
            .O(N__26300),
            .I(\eeprom.n3649 ));
    CascadeMux I__6001 (
            .O(N__26297),
            .I(N__26294));
    InMux I__6000 (
            .O(N__26294),
            .I(N__26290));
    InMux I__5999 (
            .O(N__26293),
            .I(N__26287));
    LocalMux I__5998 (
            .O(N__26290),
            .I(N__26284));
    LocalMux I__5997 (
            .O(N__26287),
            .I(N__26278));
    Span4Mux_h I__5996 (
            .O(N__26284),
            .I(N__26278));
    InMux I__5995 (
            .O(N__26283),
            .I(N__26275));
    Span4Mux_h I__5994 (
            .O(N__26278),
            .I(N__26272));
    LocalMux I__5993 (
            .O(N__26275),
            .I(\eeprom.n3017 ));
    Odrv4 I__5992 (
            .O(N__26272),
            .I(\eeprom.n3017 ));
    InMux I__5991 (
            .O(N__26267),
            .I(N__26264));
    LocalMux I__5990 (
            .O(N__26264),
            .I(N__26261));
    Span4Mux_h I__5989 (
            .O(N__26261),
            .I(N__26258));
    Span4Mux_h I__5988 (
            .O(N__26258),
            .I(N__26255));
    Odrv4 I__5987 (
            .O(N__26255),
            .I(\eeprom.n3084 ));
    InMux I__5986 (
            .O(N__26252),
            .I(\eeprom.n3650 ));
    CascadeMux I__5985 (
            .O(N__26249),
            .I(N__26246));
    InMux I__5984 (
            .O(N__26246),
            .I(N__26241));
    InMux I__5983 (
            .O(N__26245),
            .I(N__26238));
    InMux I__5982 (
            .O(N__26244),
            .I(N__26235));
    LocalMux I__5981 (
            .O(N__26241),
            .I(N__26232));
    LocalMux I__5980 (
            .O(N__26238),
            .I(N__26229));
    LocalMux I__5979 (
            .O(N__26235),
            .I(N__26224));
    Span4Mux_h I__5978 (
            .O(N__26232),
            .I(N__26224));
    Span4Mux_h I__5977 (
            .O(N__26229),
            .I(N__26221));
    Span4Mux_h I__5976 (
            .O(N__26224),
            .I(N__26218));
    Odrv4 I__5975 (
            .O(N__26221),
            .I(\eeprom.n3016 ));
    Odrv4 I__5974 (
            .O(N__26218),
            .I(\eeprom.n3016 ));
    CascadeMux I__5973 (
            .O(N__26213),
            .I(N__26210));
    InMux I__5972 (
            .O(N__26210),
            .I(N__26207));
    LocalMux I__5971 (
            .O(N__26207),
            .I(N__26204));
    Span4Mux_h I__5970 (
            .O(N__26204),
            .I(N__26201));
    Odrv4 I__5969 (
            .O(N__26201),
            .I(\eeprom.n3083 ));
    InMux I__5968 (
            .O(N__26198),
            .I(\eeprom.n3651 ));
    CascadeMux I__5967 (
            .O(N__26195),
            .I(N__26192));
    InMux I__5966 (
            .O(N__26192),
            .I(N__26188));
    InMux I__5965 (
            .O(N__26191),
            .I(N__26185));
    LocalMux I__5964 (
            .O(N__26188),
            .I(N__26181));
    LocalMux I__5963 (
            .O(N__26185),
            .I(N__26178));
    InMux I__5962 (
            .O(N__26184),
            .I(N__26175));
    Span4Mux_v I__5961 (
            .O(N__26181),
            .I(N__26172));
    Odrv4 I__5960 (
            .O(N__26178),
            .I(\eeprom.n3015 ));
    LocalMux I__5959 (
            .O(N__26175),
            .I(\eeprom.n3015 ));
    Odrv4 I__5958 (
            .O(N__26172),
            .I(\eeprom.n3015 ));
    InMux I__5957 (
            .O(N__26165),
            .I(N__26162));
    LocalMux I__5956 (
            .O(N__26162),
            .I(N__26159));
    Span4Mux_h I__5955 (
            .O(N__26159),
            .I(N__26156));
    Odrv4 I__5954 (
            .O(N__26156),
            .I(\eeprom.n3082 ));
    InMux I__5953 (
            .O(N__26153),
            .I(\eeprom.n3652 ));
    CascadeMux I__5952 (
            .O(N__26150),
            .I(N__26147));
    InMux I__5951 (
            .O(N__26147),
            .I(N__26142));
    InMux I__5950 (
            .O(N__26146),
            .I(N__26139));
    InMux I__5949 (
            .O(N__26145),
            .I(N__26136));
    LocalMux I__5948 (
            .O(N__26142),
            .I(N__26133));
    LocalMux I__5947 (
            .O(N__26139),
            .I(N__26130));
    LocalMux I__5946 (
            .O(N__26136),
            .I(N__26125));
    Span4Mux_h I__5945 (
            .O(N__26133),
            .I(N__26125));
    Span4Mux_v I__5944 (
            .O(N__26130),
            .I(N__26120));
    Span4Mux_h I__5943 (
            .O(N__26125),
            .I(N__26120));
    Odrv4 I__5942 (
            .O(N__26120),
            .I(\eeprom.n3014 ));
    CascadeMux I__5941 (
            .O(N__26117),
            .I(N__26114));
    InMux I__5940 (
            .O(N__26114),
            .I(N__26111));
    LocalMux I__5939 (
            .O(N__26111),
            .I(N__26108));
    Span4Mux_v I__5938 (
            .O(N__26108),
            .I(N__26105));
    Span4Mux_h I__5937 (
            .O(N__26105),
            .I(N__26102));
    Odrv4 I__5936 (
            .O(N__26102),
            .I(\eeprom.n3081 ));
    InMux I__5935 (
            .O(N__26099),
            .I(\eeprom.n3653 ));
    CascadeMux I__5934 (
            .O(N__26096),
            .I(N__26093));
    InMux I__5933 (
            .O(N__26093),
            .I(N__26089));
    CascadeMux I__5932 (
            .O(N__26092),
            .I(N__26085));
    LocalMux I__5931 (
            .O(N__26089),
            .I(N__26082));
    InMux I__5930 (
            .O(N__26088),
            .I(N__26077));
    InMux I__5929 (
            .O(N__26085),
            .I(N__26077));
    Span4Mux_h I__5928 (
            .O(N__26082),
            .I(N__26074));
    LocalMux I__5927 (
            .O(N__26077),
            .I(\eeprom.n3013 ));
    Odrv4 I__5926 (
            .O(N__26074),
            .I(\eeprom.n3013 ));
    InMux I__5925 (
            .O(N__26069),
            .I(N__26066));
    LocalMux I__5924 (
            .O(N__26066),
            .I(N__26063));
    Odrv4 I__5923 (
            .O(N__26063),
            .I(\eeprom.n3080 ));
    InMux I__5922 (
            .O(N__26060),
            .I(\eeprom.n3654 ));
    InMux I__5921 (
            .O(N__26057),
            .I(N__26052));
    CascadeMux I__5920 (
            .O(N__26056),
            .I(N__26049));
    InMux I__5919 (
            .O(N__26055),
            .I(N__26046));
    LocalMux I__5918 (
            .O(N__26052),
            .I(N__26043));
    InMux I__5917 (
            .O(N__26049),
            .I(N__26040));
    LocalMux I__5916 (
            .O(N__26046),
            .I(\eeprom.n3613_adj_342 ));
    Odrv4 I__5915 (
            .O(N__26043),
            .I(\eeprom.n3613_adj_342 ));
    LocalMux I__5914 (
            .O(N__26040),
            .I(\eeprom.n3613_adj_342 ));
    CascadeMux I__5913 (
            .O(N__26033),
            .I(N__26030));
    InMux I__5912 (
            .O(N__26030),
            .I(N__26027));
    LocalMux I__5911 (
            .O(N__26027),
            .I(N__26024));
    Odrv4 I__5910 (
            .O(N__26024),
            .I(\eeprom.n1347 ));
    InMux I__5909 (
            .O(N__26021),
            .I(\eeprom.n3515 ));
    InMux I__5908 (
            .O(N__26018),
            .I(N__26015));
    LocalMux I__5907 (
            .O(N__26015),
            .I(N__26011));
    InMux I__5906 (
            .O(N__26014),
            .I(N__26008));
    Odrv4 I__5905 (
            .O(N__26011),
            .I(\eeprom.n3612_adj_339 ));
    LocalMux I__5904 (
            .O(N__26008),
            .I(\eeprom.n3612_adj_339 ));
    InMux I__5903 (
            .O(N__26003),
            .I(\eeprom.n3516 ));
    InMux I__5902 (
            .O(N__26000),
            .I(N__25997));
    LocalMux I__5901 (
            .O(N__25997),
            .I(\eeprom.n1350 ));
    InMux I__5900 (
            .O(N__25994),
            .I(N__25990));
    CascadeMux I__5899 (
            .O(N__25993),
            .I(N__25987));
    LocalMux I__5898 (
            .O(N__25990),
            .I(N__25984));
    InMux I__5897 (
            .O(N__25987),
            .I(N__25981));
    Span4Mux_v I__5896 (
            .O(N__25984),
            .I(N__25975));
    LocalMux I__5895 (
            .O(N__25981),
            .I(N__25975));
    InMux I__5894 (
            .O(N__25980),
            .I(N__25972));
    Odrv4 I__5893 (
            .O(N__25975),
            .I(\eeprom.n3616_adj_345 ));
    LocalMux I__5892 (
            .O(N__25972),
            .I(\eeprom.n3616_adj_345 ));
    InMux I__5891 (
            .O(N__25967),
            .I(N__25964));
    LocalMux I__5890 (
            .O(N__25964),
            .I(\eeprom.n3715_adj_441 ));
    CascadeMux I__5889 (
            .O(N__25961),
            .I(\eeprom.n3715_adj_441_cascade_ ));
    InMux I__5888 (
            .O(N__25958),
            .I(N__25955));
    LocalMux I__5887 (
            .O(N__25955),
            .I(\eeprom.n4912 ));
    InMux I__5886 (
            .O(N__25952),
            .I(N__25949));
    LocalMux I__5885 (
            .O(N__25949),
            .I(N__25945));
    InMux I__5884 (
            .O(N__25948),
            .I(N__25942));
    Span4Mux_h I__5883 (
            .O(N__25945),
            .I(N__25939));
    LocalMux I__5882 (
            .O(N__25942),
            .I(\eeprom.n1346 ));
    Odrv4 I__5881 (
            .O(N__25939),
            .I(\eeprom.n1346 ));
    CascadeMux I__5880 (
            .O(N__25934),
            .I(N__25931));
    InMux I__5879 (
            .O(N__25931),
            .I(N__25928));
    LocalMux I__5878 (
            .O(N__25928),
            .I(\eeprom.n3711_adj_456 ));
    InMux I__5877 (
            .O(N__25925),
            .I(N__25922));
    LocalMux I__5876 (
            .O(N__25922),
            .I(\eeprom.n1352 ));
    CascadeMux I__5875 (
            .O(N__25919),
            .I(N__25916));
    InMux I__5874 (
            .O(N__25916),
            .I(N__25913));
    LocalMux I__5873 (
            .O(N__25913),
            .I(N__25909));
    InMux I__5872 (
            .O(N__25912),
            .I(N__25906));
    Odrv4 I__5871 (
            .O(N__25909),
            .I(\eeprom.n3618_adj_350 ));
    LocalMux I__5870 (
            .O(N__25906),
            .I(\eeprom.n3618_adj_350 ));
    CascadeMux I__5869 (
            .O(N__25901),
            .I(N__25898));
    InMux I__5868 (
            .O(N__25898),
            .I(N__25895));
    LocalMux I__5867 (
            .O(N__25895),
            .I(\eeprom.n3717_adj_438 ));
    CascadeMux I__5866 (
            .O(N__25892),
            .I(\eeprom.n3717_adj_438_cascade_ ));
    InMux I__5865 (
            .O(N__25889),
            .I(N__25886));
    LocalMux I__5864 (
            .O(N__25886),
            .I(\eeprom.n4906 ));
    InMux I__5863 (
            .O(N__25883),
            .I(N__25880));
    LocalMux I__5862 (
            .O(N__25880),
            .I(\eeprom.n1353 ));
    InMux I__5861 (
            .O(N__25877),
            .I(N__25872));
    InMux I__5860 (
            .O(N__25876),
            .I(N__25869));
    InMux I__5859 (
            .O(N__25875),
            .I(N__25866));
    LocalMux I__5858 (
            .O(N__25872),
            .I(N__25863));
    LocalMux I__5857 (
            .O(N__25869),
            .I(N__25860));
    LocalMux I__5856 (
            .O(N__25866),
            .I(N__25857));
    Span4Mux_h I__5855 (
            .O(N__25863),
            .I(N__25852));
    Span4Mux_v I__5854 (
            .O(N__25860),
            .I(N__25852));
    Span12Mux_v I__5853 (
            .O(N__25857),
            .I(N__25849));
    Span4Mux_h I__5852 (
            .O(N__25852),
            .I(N__25846));
    Span12Mux_h I__5851 (
            .O(N__25849),
            .I(N__25843));
    Span4Mux_h I__5850 (
            .O(N__25846),
            .I(N__25840));
    Odrv12 I__5849 (
            .O(N__25843),
            .I(\eeprom.n3619_adj_352 ));
    Odrv4 I__5848 (
            .O(N__25840),
            .I(\eeprom.n3619_adj_352 ));
    CascadeMux I__5847 (
            .O(N__25835),
            .I(N__25829));
    CascadeMux I__5846 (
            .O(N__25834),
            .I(N__25826));
    InMux I__5845 (
            .O(N__25833),
            .I(N__25821));
    CascadeMux I__5844 (
            .O(N__25832),
            .I(N__25818));
    InMux I__5843 (
            .O(N__25829),
            .I(N__25807));
    InMux I__5842 (
            .O(N__25826),
            .I(N__25807));
    InMux I__5841 (
            .O(N__25825),
            .I(N__25807));
    InMux I__5840 (
            .O(N__25824),
            .I(N__25807));
    LocalMux I__5839 (
            .O(N__25821),
            .I(N__25804));
    InMux I__5838 (
            .O(N__25818),
            .I(N__25799));
    InMux I__5837 (
            .O(N__25817),
            .I(N__25799));
    InMux I__5836 (
            .O(N__25816),
            .I(N__25796));
    LocalMux I__5835 (
            .O(N__25807),
            .I(N__25793));
    Odrv4 I__5834 (
            .O(N__25804),
            .I(\eeprom.n3628_adj_437 ));
    LocalMux I__5833 (
            .O(N__25799),
            .I(\eeprom.n3628_adj_437 ));
    LocalMux I__5832 (
            .O(N__25796),
            .I(\eeprom.n3628_adj_437 ));
    Odrv4 I__5831 (
            .O(N__25793),
            .I(\eeprom.n3628_adj_437 ));
    CascadeMux I__5830 (
            .O(N__25784),
            .I(N__25781));
    InMux I__5829 (
            .O(N__25781),
            .I(N__25778));
    LocalMux I__5828 (
            .O(N__25778),
            .I(\eeprom.n4766 ));
    InMux I__5827 (
            .O(N__25775),
            .I(N__25772));
    LocalMux I__5826 (
            .O(N__25772),
            .I(\eeprom.n3565_adj_338 ));
    InMux I__5825 (
            .O(N__25769),
            .I(\eeprom.n3769 ));
    CascadeMux I__5824 (
            .O(N__25766),
            .I(N__25763));
    InMux I__5823 (
            .O(N__25763),
            .I(N__25759));
    InMux I__5822 (
            .O(N__25762),
            .I(N__25756));
    LocalMux I__5821 (
            .O(N__25759),
            .I(N__25753));
    LocalMux I__5820 (
            .O(N__25756),
            .I(N__25750));
    Span4Mux_h I__5819 (
            .O(N__25753),
            .I(N__25747));
    Span4Mux_h I__5818 (
            .O(N__25750),
            .I(N__25744));
    Odrv4 I__5817 (
            .O(N__25747),
            .I(\eeprom.n3497 ));
    Odrv4 I__5816 (
            .O(N__25744),
            .I(\eeprom.n3497 ));
    InMux I__5815 (
            .O(N__25739),
            .I(N__25736));
    LocalMux I__5814 (
            .O(N__25736),
            .I(N__25733));
    Span4Mux_h I__5813 (
            .O(N__25733),
            .I(N__25730));
    Odrv4 I__5812 (
            .O(N__25730),
            .I(\eeprom.n3564_adj_337 ));
    InMux I__5811 (
            .O(N__25727),
            .I(\eeprom.n3770 ));
    InMux I__5810 (
            .O(N__25724),
            .I(N__25720));
    InMux I__5809 (
            .O(N__25723),
            .I(N__25717));
    LocalMux I__5808 (
            .O(N__25720),
            .I(N__25714));
    LocalMux I__5807 (
            .O(N__25717),
            .I(N__25711));
    Odrv4 I__5806 (
            .O(N__25714),
            .I(\eeprom.n3496 ));
    Odrv4 I__5805 (
            .O(N__25711),
            .I(\eeprom.n3496 ));
    CascadeMux I__5804 (
            .O(N__25706),
            .I(N__25700));
    CascadeMux I__5803 (
            .O(N__25705),
            .I(N__25697));
    CascadeMux I__5802 (
            .O(N__25704),
            .I(N__25693));
    CascadeMux I__5801 (
            .O(N__25703),
            .I(N__25690));
    InMux I__5800 (
            .O(N__25700),
            .I(N__25686));
    InMux I__5799 (
            .O(N__25697),
            .I(N__25673));
    InMux I__5798 (
            .O(N__25696),
            .I(N__25673));
    InMux I__5797 (
            .O(N__25693),
            .I(N__25665));
    InMux I__5796 (
            .O(N__25690),
            .I(N__25665));
    InMux I__5795 (
            .O(N__25689),
            .I(N__25665));
    LocalMux I__5794 (
            .O(N__25686),
            .I(N__25656));
    InMux I__5793 (
            .O(N__25685),
            .I(N__25649));
    InMux I__5792 (
            .O(N__25684),
            .I(N__25649));
    InMux I__5791 (
            .O(N__25683),
            .I(N__25649));
    InMux I__5790 (
            .O(N__25682),
            .I(N__25642));
    InMux I__5789 (
            .O(N__25681),
            .I(N__25642));
    InMux I__5788 (
            .O(N__25680),
            .I(N__25642));
    InMux I__5787 (
            .O(N__25679),
            .I(N__25637));
    InMux I__5786 (
            .O(N__25678),
            .I(N__25637));
    LocalMux I__5785 (
            .O(N__25673),
            .I(N__25634));
    CascadeMux I__5784 (
            .O(N__25672),
            .I(N__25629));
    LocalMux I__5783 (
            .O(N__25665),
            .I(N__25625));
    InMux I__5782 (
            .O(N__25664),
            .I(N__25616));
    InMux I__5781 (
            .O(N__25663),
            .I(N__25616));
    InMux I__5780 (
            .O(N__25662),
            .I(N__25616));
    InMux I__5779 (
            .O(N__25661),
            .I(N__25616));
    InMux I__5778 (
            .O(N__25660),
            .I(N__25613));
    InMux I__5777 (
            .O(N__25659),
            .I(N__25610));
    Span4Mux_h I__5776 (
            .O(N__25656),
            .I(N__25599));
    LocalMux I__5775 (
            .O(N__25649),
            .I(N__25599));
    LocalMux I__5774 (
            .O(N__25642),
            .I(N__25599));
    LocalMux I__5773 (
            .O(N__25637),
            .I(N__25599));
    Span4Mux_v I__5772 (
            .O(N__25634),
            .I(N__25599));
    InMux I__5771 (
            .O(N__25633),
            .I(N__25590));
    InMux I__5770 (
            .O(N__25632),
            .I(N__25590));
    InMux I__5769 (
            .O(N__25629),
            .I(N__25590));
    InMux I__5768 (
            .O(N__25628),
            .I(N__25590));
    Span4Mux_h I__5767 (
            .O(N__25625),
            .I(N__25587));
    LocalMux I__5766 (
            .O(N__25616),
            .I(\eeprom.n3529_adj_336 ));
    LocalMux I__5765 (
            .O(N__25613),
            .I(\eeprom.n3529_adj_336 ));
    LocalMux I__5764 (
            .O(N__25610),
            .I(\eeprom.n3529_adj_336 ));
    Odrv4 I__5763 (
            .O(N__25599),
            .I(\eeprom.n3529_adj_336 ));
    LocalMux I__5762 (
            .O(N__25590),
            .I(\eeprom.n3529_adj_336 ));
    Odrv4 I__5761 (
            .O(N__25587),
            .I(\eeprom.n3529_adj_336 ));
    InMux I__5760 (
            .O(N__25574),
            .I(\eeprom.n3771 ));
    InMux I__5759 (
            .O(N__25571),
            .I(N__25568));
    LocalMux I__5758 (
            .O(N__25568),
            .I(\eeprom.n4765 ));
    InMux I__5757 (
            .O(N__25565),
            .I(bfn_16_20_0_));
    InMux I__5756 (
            .O(N__25562),
            .I(\eeprom.n3510 ));
    InMux I__5755 (
            .O(N__25559),
            .I(N__25555));
    InMux I__5754 (
            .O(N__25558),
            .I(N__25552));
    LocalMux I__5753 (
            .O(N__25555),
            .I(N__25549));
    LocalMux I__5752 (
            .O(N__25552),
            .I(\eeprom.n3617_adj_346 ));
    Odrv4 I__5751 (
            .O(N__25549),
            .I(\eeprom.n3617_adj_346 ));
    InMux I__5750 (
            .O(N__25544),
            .I(N__25541));
    LocalMux I__5749 (
            .O(N__25541),
            .I(\eeprom.n1351 ));
    InMux I__5748 (
            .O(N__25538),
            .I(\eeprom.n3511 ));
    InMux I__5747 (
            .O(N__25535),
            .I(\eeprom.n3512 ));
    CascadeMux I__5746 (
            .O(N__25532),
            .I(N__25529));
    InMux I__5745 (
            .O(N__25529),
            .I(N__25526));
    LocalMux I__5744 (
            .O(N__25526),
            .I(N__25522));
    InMux I__5743 (
            .O(N__25525),
            .I(N__25519));
    Odrv4 I__5742 (
            .O(N__25522),
            .I(\eeprom.n3615_adj_344 ));
    LocalMux I__5741 (
            .O(N__25519),
            .I(\eeprom.n3615_adj_344 ));
    InMux I__5740 (
            .O(N__25514),
            .I(N__25511));
    LocalMux I__5739 (
            .O(N__25511),
            .I(N__25508));
    Odrv4 I__5738 (
            .O(N__25508),
            .I(\eeprom.n1349 ));
    InMux I__5737 (
            .O(N__25505),
            .I(\eeprom.n3513 ));
    InMux I__5736 (
            .O(N__25502),
            .I(N__25498));
    InMux I__5735 (
            .O(N__25501),
            .I(N__25495));
    LocalMux I__5734 (
            .O(N__25498),
            .I(N__25491));
    LocalMux I__5733 (
            .O(N__25495),
            .I(N__25488));
    InMux I__5732 (
            .O(N__25494),
            .I(N__25485));
    Odrv4 I__5731 (
            .O(N__25491),
            .I(\eeprom.n3614_adj_343 ));
    Odrv4 I__5730 (
            .O(N__25488),
            .I(\eeprom.n3614_adj_343 ));
    LocalMux I__5729 (
            .O(N__25485),
            .I(\eeprom.n3614_adj_343 ));
    InMux I__5728 (
            .O(N__25478),
            .I(N__25475));
    LocalMux I__5727 (
            .O(N__25475),
            .I(N__25472));
    Odrv4 I__5726 (
            .O(N__25472),
            .I(\eeprom.n1348 ));
    InMux I__5725 (
            .O(N__25469),
            .I(\eeprom.n3514 ));
    InMux I__5724 (
            .O(N__25466),
            .I(N__25463));
    LocalMux I__5723 (
            .O(N__25463),
            .I(N__25459));
    InMux I__5722 (
            .O(N__25462),
            .I(N__25456));
    Span4Mux_h I__5721 (
            .O(N__25459),
            .I(N__25453));
    LocalMux I__5720 (
            .O(N__25456),
            .I(N__25450));
    Odrv4 I__5719 (
            .O(N__25453),
            .I(\eeprom.n3505 ));
    Odrv12 I__5718 (
            .O(N__25450),
            .I(\eeprom.n3505 ));
    InMux I__5717 (
            .O(N__25445),
            .I(N__25442));
    LocalMux I__5716 (
            .O(N__25442),
            .I(N__25439));
    Span4Mux_h I__5715 (
            .O(N__25439),
            .I(N__25436));
    Odrv4 I__5714 (
            .O(N__25436),
            .I(\eeprom.n3572_adj_354 ));
    InMux I__5713 (
            .O(N__25433),
            .I(\eeprom.n3762 ));
    InMux I__5712 (
            .O(N__25430),
            .I(N__25426));
    InMux I__5711 (
            .O(N__25429),
            .I(N__25422));
    LocalMux I__5710 (
            .O(N__25426),
            .I(N__25419));
    InMux I__5709 (
            .O(N__25425),
            .I(N__25416));
    LocalMux I__5708 (
            .O(N__25422),
            .I(\eeprom.n3504 ));
    Odrv4 I__5707 (
            .O(N__25419),
            .I(\eeprom.n3504 ));
    LocalMux I__5706 (
            .O(N__25416),
            .I(\eeprom.n3504 ));
    InMux I__5705 (
            .O(N__25409),
            .I(N__25406));
    LocalMux I__5704 (
            .O(N__25406),
            .I(N__25403));
    Span4Mux_h I__5703 (
            .O(N__25403),
            .I(N__25400));
    Odrv4 I__5702 (
            .O(N__25400),
            .I(\eeprom.n3571_adj_353 ));
    InMux I__5701 (
            .O(N__25397),
            .I(\eeprom.n3763 ));
    InMux I__5700 (
            .O(N__25394),
            .I(N__25390));
    InMux I__5699 (
            .O(N__25393),
            .I(N__25386));
    LocalMux I__5698 (
            .O(N__25390),
            .I(N__25383));
    CascadeMux I__5697 (
            .O(N__25389),
            .I(N__25380));
    LocalMux I__5696 (
            .O(N__25386),
            .I(N__25377));
    Span4Mux_h I__5695 (
            .O(N__25383),
            .I(N__25374));
    InMux I__5694 (
            .O(N__25380),
            .I(N__25371));
    Span4Mux_h I__5693 (
            .O(N__25377),
            .I(N__25368));
    Odrv4 I__5692 (
            .O(N__25374),
            .I(\eeprom.n3503 ));
    LocalMux I__5691 (
            .O(N__25371),
            .I(\eeprom.n3503 ));
    Odrv4 I__5690 (
            .O(N__25368),
            .I(\eeprom.n3503 ));
    InMux I__5689 (
            .O(N__25361),
            .I(N__25358));
    LocalMux I__5688 (
            .O(N__25358),
            .I(N__25355));
    Odrv12 I__5687 (
            .O(N__25355),
            .I(\eeprom.n3570_adj_349 ));
    InMux I__5686 (
            .O(N__25352),
            .I(bfn_16_19_0_));
    InMux I__5685 (
            .O(N__25349),
            .I(N__25345));
    InMux I__5684 (
            .O(N__25348),
            .I(N__25342));
    LocalMux I__5683 (
            .O(N__25345),
            .I(N__25336));
    LocalMux I__5682 (
            .O(N__25342),
            .I(N__25336));
    InMux I__5681 (
            .O(N__25341),
            .I(N__25333));
    Odrv4 I__5680 (
            .O(N__25336),
            .I(\eeprom.n3502 ));
    LocalMux I__5679 (
            .O(N__25333),
            .I(\eeprom.n3502 ));
    CascadeMux I__5678 (
            .O(N__25328),
            .I(N__25325));
    InMux I__5677 (
            .O(N__25325),
            .I(N__25322));
    LocalMux I__5676 (
            .O(N__25322),
            .I(\eeprom.n3569_adj_348 ));
    InMux I__5675 (
            .O(N__25319),
            .I(\eeprom.n3765 ));
    InMux I__5674 (
            .O(N__25316),
            .I(N__25313));
    LocalMux I__5673 (
            .O(N__25313),
            .I(N__25309));
    InMux I__5672 (
            .O(N__25312),
            .I(N__25305));
    Span4Mux_h I__5671 (
            .O(N__25309),
            .I(N__25302));
    InMux I__5670 (
            .O(N__25308),
            .I(N__25299));
    LocalMux I__5669 (
            .O(N__25305),
            .I(\eeprom.n3501 ));
    Odrv4 I__5668 (
            .O(N__25302),
            .I(\eeprom.n3501 ));
    LocalMux I__5667 (
            .O(N__25299),
            .I(\eeprom.n3501 ));
    InMux I__5666 (
            .O(N__25292),
            .I(N__25289));
    LocalMux I__5665 (
            .O(N__25289),
            .I(N__25286));
    Span4Mux_h I__5664 (
            .O(N__25286),
            .I(N__25283));
    Odrv4 I__5663 (
            .O(N__25283),
            .I(\eeprom.n3568_adj_347 ));
    InMux I__5662 (
            .O(N__25280),
            .I(\eeprom.n3766 ));
    InMux I__5661 (
            .O(N__25277),
            .I(N__25273));
    CascadeMux I__5660 (
            .O(N__25276),
            .I(N__25270));
    LocalMux I__5659 (
            .O(N__25273),
            .I(N__25267));
    InMux I__5658 (
            .O(N__25270),
            .I(N__25264));
    Span4Mux_v I__5657 (
            .O(N__25267),
            .I(N__25261));
    LocalMux I__5656 (
            .O(N__25264),
            .I(\eeprom.n3500 ));
    Odrv4 I__5655 (
            .O(N__25261),
            .I(\eeprom.n3500 ));
    InMux I__5654 (
            .O(N__25256),
            .I(N__25253));
    LocalMux I__5653 (
            .O(N__25253),
            .I(N__25250));
    Span4Mux_h I__5652 (
            .O(N__25250),
            .I(N__25247));
    Odrv4 I__5651 (
            .O(N__25247),
            .I(\eeprom.n3567_adj_341 ));
    InMux I__5650 (
            .O(N__25244),
            .I(\eeprom.n3767 ));
    InMux I__5649 (
            .O(N__25241),
            .I(N__25236));
    InMux I__5648 (
            .O(N__25240),
            .I(N__25233));
    InMux I__5647 (
            .O(N__25239),
            .I(N__25230));
    LocalMux I__5646 (
            .O(N__25236),
            .I(N__25227));
    LocalMux I__5645 (
            .O(N__25233),
            .I(N__25224));
    LocalMux I__5644 (
            .O(N__25230),
            .I(\eeprom.n3499 ));
    Odrv12 I__5643 (
            .O(N__25227),
            .I(\eeprom.n3499 ));
    Odrv4 I__5642 (
            .O(N__25224),
            .I(\eeprom.n3499 ));
    CascadeMux I__5641 (
            .O(N__25217),
            .I(N__25214));
    InMux I__5640 (
            .O(N__25214),
            .I(N__25211));
    LocalMux I__5639 (
            .O(N__25211),
            .I(N__25208));
    Span4Mux_v I__5638 (
            .O(N__25208),
            .I(N__25205));
    Odrv4 I__5637 (
            .O(N__25205),
            .I(\eeprom.n3566_adj_340 ));
    InMux I__5636 (
            .O(N__25202),
            .I(\eeprom.n3768 ));
    InMux I__5635 (
            .O(N__25199),
            .I(N__25195));
    InMux I__5634 (
            .O(N__25198),
            .I(N__25192));
    LocalMux I__5633 (
            .O(N__25195),
            .I(N__25187));
    LocalMux I__5632 (
            .O(N__25192),
            .I(N__25187));
    Span4Mux_h I__5631 (
            .O(N__25187),
            .I(N__25183));
    InMux I__5630 (
            .O(N__25186),
            .I(N__25180));
    Odrv4 I__5629 (
            .O(N__25183),
            .I(\eeprom.n3498 ));
    LocalMux I__5628 (
            .O(N__25180),
            .I(\eeprom.n3498 ));
    CascadeMux I__5627 (
            .O(N__25175),
            .I(N__25171));
    CascadeMux I__5626 (
            .O(N__25174),
            .I(N__25168));
    InMux I__5625 (
            .O(N__25171),
            .I(N__25165));
    InMux I__5624 (
            .O(N__25168),
            .I(N__25162));
    LocalMux I__5623 (
            .O(N__25165),
            .I(N__25158));
    LocalMux I__5622 (
            .O(N__25162),
            .I(N__25155));
    InMux I__5621 (
            .O(N__25161),
            .I(N__25152));
    Span4Mux_v I__5620 (
            .O(N__25158),
            .I(N__25149));
    Span4Mux_h I__5619 (
            .O(N__25155),
            .I(N__25144));
    LocalMux I__5618 (
            .O(N__25152),
            .I(N__25144));
    Odrv4 I__5617 (
            .O(N__25149),
            .I(\eeprom.n3513_adj_366 ));
    Odrv4 I__5616 (
            .O(N__25144),
            .I(\eeprom.n3513_adj_366 ));
    InMux I__5615 (
            .O(N__25139),
            .I(N__25136));
    LocalMux I__5614 (
            .O(N__25136),
            .I(N__25133));
    Span4Mux_v I__5613 (
            .O(N__25133),
            .I(N__25130));
    Odrv4 I__5612 (
            .O(N__25130),
            .I(\eeprom.n3580_adj_365 ));
    InMux I__5611 (
            .O(N__25127),
            .I(\eeprom.n3754 ));
    CascadeMux I__5610 (
            .O(N__25124),
            .I(N__25120));
    InMux I__5609 (
            .O(N__25123),
            .I(N__25117));
    InMux I__5608 (
            .O(N__25120),
            .I(N__25114));
    LocalMux I__5607 (
            .O(N__25117),
            .I(N__25110));
    LocalMux I__5606 (
            .O(N__25114),
            .I(N__25107));
    InMux I__5605 (
            .O(N__25113),
            .I(N__25104));
    Odrv4 I__5604 (
            .O(N__25110),
            .I(\eeprom.n3512_adj_364 ));
    Odrv4 I__5603 (
            .O(N__25107),
            .I(\eeprom.n3512_adj_364 ));
    LocalMux I__5602 (
            .O(N__25104),
            .I(\eeprom.n3512_adj_364 ));
    CascadeMux I__5601 (
            .O(N__25097),
            .I(N__25094));
    InMux I__5600 (
            .O(N__25094),
            .I(N__25091));
    LocalMux I__5599 (
            .O(N__25091),
            .I(N__25088));
    Span4Mux_h I__5598 (
            .O(N__25088),
            .I(N__25085));
    Odrv4 I__5597 (
            .O(N__25085),
            .I(\eeprom.n3579_adj_363 ));
    InMux I__5596 (
            .O(N__25082),
            .I(\eeprom.n3755 ));
    CascadeMux I__5595 (
            .O(N__25079),
            .I(N__25076));
    InMux I__5594 (
            .O(N__25076),
            .I(N__25073));
    LocalMux I__5593 (
            .O(N__25073),
            .I(N__25068));
    InMux I__5592 (
            .O(N__25072),
            .I(N__25065));
    InMux I__5591 (
            .O(N__25071),
            .I(N__25062));
    Span4Mux_h I__5590 (
            .O(N__25068),
            .I(N__25059));
    LocalMux I__5589 (
            .O(N__25065),
            .I(\eeprom.n3511_adj_362 ));
    LocalMux I__5588 (
            .O(N__25062),
            .I(\eeprom.n3511_adj_362 ));
    Odrv4 I__5587 (
            .O(N__25059),
            .I(\eeprom.n3511_adj_362 ));
    InMux I__5586 (
            .O(N__25052),
            .I(N__25049));
    LocalMux I__5585 (
            .O(N__25049),
            .I(N__25046));
    Span4Mux_h I__5584 (
            .O(N__25046),
            .I(N__25043));
    Odrv4 I__5583 (
            .O(N__25043),
            .I(\eeprom.n3578_adj_361 ));
    InMux I__5582 (
            .O(N__25040),
            .I(bfn_16_18_0_));
    CascadeMux I__5581 (
            .O(N__25037),
            .I(N__25034));
    InMux I__5580 (
            .O(N__25034),
            .I(N__25030));
    CascadeMux I__5579 (
            .O(N__25033),
            .I(N__25027));
    LocalMux I__5578 (
            .O(N__25030),
            .I(N__25023));
    InMux I__5577 (
            .O(N__25027),
            .I(N__25018));
    InMux I__5576 (
            .O(N__25026),
            .I(N__25018));
    Odrv4 I__5575 (
            .O(N__25023),
            .I(\eeprom.n3510_adj_360 ));
    LocalMux I__5574 (
            .O(N__25018),
            .I(\eeprom.n3510_adj_360 ));
    InMux I__5573 (
            .O(N__25013),
            .I(N__25010));
    LocalMux I__5572 (
            .O(N__25010),
            .I(N__25007));
    Span4Mux_h I__5571 (
            .O(N__25007),
            .I(N__25004));
    Odrv4 I__5570 (
            .O(N__25004),
            .I(\eeprom.n3577_adj_359 ));
    InMux I__5569 (
            .O(N__25001),
            .I(\eeprom.n3757 ));
    CascadeMux I__5568 (
            .O(N__24998),
            .I(N__24995));
    InMux I__5567 (
            .O(N__24995),
            .I(N__24991));
    CascadeMux I__5566 (
            .O(N__24994),
            .I(N__24988));
    LocalMux I__5565 (
            .O(N__24991),
            .I(N__24985));
    InMux I__5564 (
            .O(N__24988),
            .I(N__24981));
    Span4Mux_h I__5563 (
            .O(N__24985),
            .I(N__24978));
    InMux I__5562 (
            .O(N__24984),
            .I(N__24975));
    LocalMux I__5561 (
            .O(N__24981),
            .I(\eeprom.n3509 ));
    Odrv4 I__5560 (
            .O(N__24978),
            .I(\eeprom.n3509 ));
    LocalMux I__5559 (
            .O(N__24975),
            .I(\eeprom.n3509 ));
    InMux I__5558 (
            .O(N__24968),
            .I(N__24965));
    LocalMux I__5557 (
            .O(N__24965),
            .I(N__24962));
    Span4Mux_h I__5556 (
            .O(N__24962),
            .I(N__24959));
    Odrv4 I__5555 (
            .O(N__24959),
            .I(\eeprom.n3576_adj_358 ));
    InMux I__5554 (
            .O(N__24956),
            .I(\eeprom.n3758 ));
    CascadeMux I__5553 (
            .O(N__24953),
            .I(N__24950));
    InMux I__5552 (
            .O(N__24950),
            .I(N__24947));
    LocalMux I__5551 (
            .O(N__24947),
            .I(N__24943));
    InMux I__5550 (
            .O(N__24946),
            .I(N__24940));
    Odrv12 I__5549 (
            .O(N__24943),
            .I(\eeprom.n3508 ));
    LocalMux I__5548 (
            .O(N__24940),
            .I(\eeprom.n3508 ));
    InMux I__5547 (
            .O(N__24935),
            .I(N__24932));
    LocalMux I__5546 (
            .O(N__24932),
            .I(N__24929));
    Odrv4 I__5545 (
            .O(N__24929),
            .I(\eeprom.n3575_adj_357 ));
    InMux I__5544 (
            .O(N__24926),
            .I(\eeprom.n3759 ));
    InMux I__5543 (
            .O(N__24923),
            .I(N__24919));
    CascadeMux I__5542 (
            .O(N__24922),
            .I(N__24915));
    LocalMux I__5541 (
            .O(N__24919),
            .I(N__24912));
    InMux I__5540 (
            .O(N__24918),
            .I(N__24907));
    InMux I__5539 (
            .O(N__24915),
            .I(N__24907));
    Odrv4 I__5538 (
            .O(N__24912),
            .I(\eeprom.n3507 ));
    LocalMux I__5537 (
            .O(N__24907),
            .I(\eeprom.n3507 ));
    CascadeMux I__5536 (
            .O(N__24902),
            .I(N__24899));
    InMux I__5535 (
            .O(N__24899),
            .I(N__24896));
    LocalMux I__5534 (
            .O(N__24896),
            .I(N__24893));
    Span4Mux_v I__5533 (
            .O(N__24893),
            .I(N__24890));
    Odrv4 I__5532 (
            .O(N__24890),
            .I(\eeprom.n3574_adj_356 ));
    InMux I__5531 (
            .O(N__24887),
            .I(\eeprom.n3760 ));
    InMux I__5530 (
            .O(N__24884),
            .I(N__24880));
    InMux I__5529 (
            .O(N__24883),
            .I(N__24877));
    LocalMux I__5528 (
            .O(N__24880),
            .I(N__24874));
    LocalMux I__5527 (
            .O(N__24877),
            .I(N__24871));
    Span4Mux_h I__5526 (
            .O(N__24874),
            .I(N__24865));
    Span4Mux_h I__5525 (
            .O(N__24871),
            .I(N__24865));
    InMux I__5524 (
            .O(N__24870),
            .I(N__24862));
    Odrv4 I__5523 (
            .O(N__24865),
            .I(\eeprom.n3506 ));
    LocalMux I__5522 (
            .O(N__24862),
            .I(\eeprom.n3506 ));
    InMux I__5521 (
            .O(N__24857),
            .I(N__24854));
    LocalMux I__5520 (
            .O(N__24854),
            .I(\eeprom.n3573_adj_355 ));
    InMux I__5519 (
            .O(N__24851),
            .I(\eeprom.n3761 ));
    InMux I__5518 (
            .O(N__24848),
            .I(N__24845));
    LocalMux I__5517 (
            .O(N__24845),
            .I(N__24842));
    Span4Mux_v I__5516 (
            .O(N__24842),
            .I(N__24839));
    Odrv4 I__5515 (
            .O(N__24839),
            .I(\eeprom.n2986 ));
    InMux I__5514 (
            .O(N__24836),
            .I(N__24833));
    LocalMux I__5513 (
            .O(N__24833),
            .I(N__24829));
    InMux I__5512 (
            .O(N__24832),
            .I(N__24826));
    Span4Mux_h I__5511 (
            .O(N__24829),
            .I(N__24822));
    LocalMux I__5510 (
            .O(N__24826),
            .I(N__24819));
    InMux I__5509 (
            .O(N__24825),
            .I(N__24816));
    Span4Mux_h I__5508 (
            .O(N__24822),
            .I(N__24811));
    Span4Mux_v I__5507 (
            .O(N__24819),
            .I(N__24811));
    LocalMux I__5506 (
            .O(N__24816),
            .I(N__24808));
    Span4Mux_h I__5505 (
            .O(N__24811),
            .I(N__24803));
    Span4Mux_h I__5504 (
            .O(N__24808),
            .I(N__24803));
    Span4Mux_h I__5503 (
            .O(N__24803),
            .I(N__24800));
    Odrv4 I__5502 (
            .O(N__24800),
            .I(\eeprom.n2919 ));
    CascadeMux I__5501 (
            .O(N__24797),
            .I(N__24793));
    InMux I__5500 (
            .O(N__24796),
            .I(N__24790));
    InMux I__5499 (
            .O(N__24793),
            .I(N__24787));
    LocalMux I__5498 (
            .O(N__24790),
            .I(N__24784));
    LocalMux I__5497 (
            .O(N__24787),
            .I(N__24781));
    Odrv12 I__5496 (
            .O(N__24784),
            .I(\eeprom.n2909 ));
    Odrv4 I__5495 (
            .O(N__24781),
            .I(\eeprom.n2909 ));
    InMux I__5494 (
            .O(N__24776),
            .I(N__24773));
    LocalMux I__5493 (
            .O(N__24773),
            .I(N__24770));
    Span4Mux_v I__5492 (
            .O(N__24770),
            .I(N__24767));
    Odrv4 I__5491 (
            .O(N__24767),
            .I(\eeprom.n2976 ));
    CascadeMux I__5490 (
            .O(N__24764),
            .I(N__24754));
    InMux I__5489 (
            .O(N__24763),
            .I(N__24750));
    InMux I__5488 (
            .O(N__24762),
            .I(N__24747));
    InMux I__5487 (
            .O(N__24761),
            .I(N__24742));
    InMux I__5486 (
            .O(N__24760),
            .I(N__24742));
    CascadeMux I__5485 (
            .O(N__24759),
            .I(N__24738));
    CascadeMux I__5484 (
            .O(N__24758),
            .I(N__24732));
    CascadeMux I__5483 (
            .O(N__24757),
            .I(N__24729));
    InMux I__5482 (
            .O(N__24754),
            .I(N__24722));
    InMux I__5481 (
            .O(N__24753),
            .I(N__24722));
    LocalMux I__5480 (
            .O(N__24750),
            .I(N__24719));
    LocalMux I__5479 (
            .O(N__24747),
            .I(N__24714));
    LocalMux I__5478 (
            .O(N__24742),
            .I(N__24714));
    InMux I__5477 (
            .O(N__24741),
            .I(N__24707));
    InMux I__5476 (
            .O(N__24738),
            .I(N__24707));
    InMux I__5475 (
            .O(N__24737),
            .I(N__24707));
    CascadeMux I__5474 (
            .O(N__24736),
            .I(N__24702));
    InMux I__5473 (
            .O(N__24735),
            .I(N__24698));
    InMux I__5472 (
            .O(N__24732),
            .I(N__24689));
    InMux I__5471 (
            .O(N__24729),
            .I(N__24689));
    InMux I__5470 (
            .O(N__24728),
            .I(N__24689));
    InMux I__5469 (
            .O(N__24727),
            .I(N__24689));
    LocalMux I__5468 (
            .O(N__24722),
            .I(N__24680));
    Span4Mux_v I__5467 (
            .O(N__24719),
            .I(N__24680));
    Span4Mux_h I__5466 (
            .O(N__24714),
            .I(N__24680));
    LocalMux I__5465 (
            .O(N__24707),
            .I(N__24680));
    InMux I__5464 (
            .O(N__24706),
            .I(N__24671));
    InMux I__5463 (
            .O(N__24705),
            .I(N__24671));
    InMux I__5462 (
            .O(N__24702),
            .I(N__24671));
    InMux I__5461 (
            .O(N__24701),
            .I(N__24671));
    LocalMux I__5460 (
            .O(N__24698),
            .I(N__24668));
    LocalMux I__5459 (
            .O(N__24689),
            .I(\eeprom.n2935 ));
    Odrv4 I__5458 (
            .O(N__24680),
            .I(\eeprom.n2935 ));
    LocalMux I__5457 (
            .O(N__24671),
            .I(\eeprom.n2935 ));
    Odrv4 I__5456 (
            .O(N__24668),
            .I(\eeprom.n2935 ));
    InMux I__5455 (
            .O(N__24659),
            .I(N__24655));
    InMux I__5454 (
            .O(N__24658),
            .I(N__24651));
    LocalMux I__5453 (
            .O(N__24655),
            .I(N__24648));
    InMux I__5452 (
            .O(N__24654),
            .I(N__24645));
    LocalMux I__5451 (
            .O(N__24651),
            .I(N__24642));
    Span12Mux_v I__5450 (
            .O(N__24648),
            .I(N__24639));
    LocalMux I__5449 (
            .O(N__24645),
            .I(N__24636));
    Span4Mux_v I__5448 (
            .O(N__24642),
            .I(N__24633));
    Span12Mux_h I__5447 (
            .O(N__24639),
            .I(N__24630));
    Span12Mux_v I__5446 (
            .O(N__24636),
            .I(N__24625));
    Sp12to4 I__5445 (
            .O(N__24633),
            .I(N__24625));
    Odrv12 I__5444 (
            .O(N__24630),
            .I(\eeprom.n3519_adj_379 ));
    Odrv12 I__5443 (
            .O(N__24625),
            .I(\eeprom.n3519_adj_379 ));
    InMux I__5442 (
            .O(N__24620),
            .I(N__24617));
    LocalMux I__5441 (
            .O(N__24617),
            .I(N__24614));
    Span4Mux_h I__5440 (
            .O(N__24614),
            .I(N__24611));
    Odrv4 I__5439 (
            .O(N__24611),
            .I(\eeprom.n3586_adj_378 ));
    InMux I__5438 (
            .O(N__24608),
            .I(bfn_16_17_0_));
    CascadeMux I__5437 (
            .O(N__24605),
            .I(N__24601));
    InMux I__5436 (
            .O(N__24604),
            .I(N__24597));
    InMux I__5435 (
            .O(N__24601),
            .I(N__24594));
    InMux I__5434 (
            .O(N__24600),
            .I(N__24591));
    LocalMux I__5433 (
            .O(N__24597),
            .I(\eeprom.n3518_adj_376 ));
    LocalMux I__5432 (
            .O(N__24594),
            .I(\eeprom.n3518_adj_376 ));
    LocalMux I__5431 (
            .O(N__24591),
            .I(\eeprom.n3518_adj_376 ));
    InMux I__5430 (
            .O(N__24584),
            .I(N__24581));
    LocalMux I__5429 (
            .O(N__24581),
            .I(\eeprom.n3585_adj_375 ));
    InMux I__5428 (
            .O(N__24578),
            .I(\eeprom.n3749 ));
    CascadeMux I__5427 (
            .O(N__24575),
            .I(N__24571));
    InMux I__5426 (
            .O(N__24574),
            .I(N__24568));
    InMux I__5425 (
            .O(N__24571),
            .I(N__24565));
    LocalMux I__5424 (
            .O(N__24568),
            .I(\eeprom.n3517_adj_374 ));
    LocalMux I__5423 (
            .O(N__24565),
            .I(\eeprom.n3517_adj_374 ));
    InMux I__5422 (
            .O(N__24560),
            .I(N__24557));
    LocalMux I__5421 (
            .O(N__24557),
            .I(\eeprom.n3584_adj_373 ));
    InMux I__5420 (
            .O(N__24554),
            .I(\eeprom.n3750 ));
    CascadeMux I__5419 (
            .O(N__24551),
            .I(N__24547));
    CascadeMux I__5418 (
            .O(N__24550),
            .I(N__24544));
    InMux I__5417 (
            .O(N__24547),
            .I(N__24540));
    InMux I__5416 (
            .O(N__24544),
            .I(N__24537));
    InMux I__5415 (
            .O(N__24543),
            .I(N__24534));
    LocalMux I__5414 (
            .O(N__24540),
            .I(\eeprom.n3516_adj_372 ));
    LocalMux I__5413 (
            .O(N__24537),
            .I(\eeprom.n3516_adj_372 ));
    LocalMux I__5412 (
            .O(N__24534),
            .I(\eeprom.n3516_adj_372 ));
    InMux I__5411 (
            .O(N__24527),
            .I(N__24524));
    LocalMux I__5410 (
            .O(N__24524),
            .I(\eeprom.n3583_adj_371 ));
    InMux I__5409 (
            .O(N__24521),
            .I(\eeprom.n3751 ));
    CascadeMux I__5408 (
            .O(N__24518),
            .I(N__24514));
    InMux I__5407 (
            .O(N__24517),
            .I(N__24511));
    InMux I__5406 (
            .O(N__24514),
            .I(N__24508));
    LocalMux I__5405 (
            .O(N__24511),
            .I(\eeprom.n3515_adj_370 ));
    LocalMux I__5404 (
            .O(N__24508),
            .I(\eeprom.n3515_adj_370 ));
    CascadeMux I__5403 (
            .O(N__24503),
            .I(N__24500));
    InMux I__5402 (
            .O(N__24500),
            .I(N__24497));
    LocalMux I__5401 (
            .O(N__24497),
            .I(\eeprom.n3582_adj_369 ));
    InMux I__5400 (
            .O(N__24494),
            .I(\eeprom.n3752 ));
    CascadeMux I__5399 (
            .O(N__24491),
            .I(N__24488));
    InMux I__5398 (
            .O(N__24488),
            .I(N__24484));
    InMux I__5397 (
            .O(N__24487),
            .I(N__24480));
    LocalMux I__5396 (
            .O(N__24484),
            .I(N__24477));
    InMux I__5395 (
            .O(N__24483),
            .I(N__24474));
    LocalMux I__5394 (
            .O(N__24480),
            .I(N__24471));
    Span4Mux_h I__5393 (
            .O(N__24477),
            .I(N__24466));
    LocalMux I__5392 (
            .O(N__24474),
            .I(N__24466));
    Odrv12 I__5391 (
            .O(N__24471),
            .I(\eeprom.n3514_adj_368 ));
    Odrv4 I__5390 (
            .O(N__24466),
            .I(\eeprom.n3514_adj_368 ));
    CascadeMux I__5389 (
            .O(N__24461),
            .I(N__24458));
    InMux I__5388 (
            .O(N__24458),
            .I(N__24455));
    LocalMux I__5387 (
            .O(N__24455),
            .I(N__24452));
    Span4Mux_h I__5386 (
            .O(N__24452),
            .I(N__24449));
    Odrv4 I__5385 (
            .O(N__24449),
            .I(\eeprom.n3581_adj_367 ));
    InMux I__5384 (
            .O(N__24446),
            .I(\eeprom.n3753 ));
    InMux I__5383 (
            .O(N__24443),
            .I(N__24440));
    LocalMux I__5382 (
            .O(N__24440),
            .I(N__24437));
    Odrv12 I__5381 (
            .O(N__24437),
            .I(\eeprom.number_of_bytes_7_N_68_6 ));
    InMux I__5380 (
            .O(N__24434),
            .I(N__24431));
    LocalMux I__5379 (
            .O(N__24431),
            .I(\eeprom.number_of_bytes_7_N_68_8 ));
    CascadeMux I__5378 (
            .O(N__24428),
            .I(\eeprom.n4301_cascade_ ));
    InMux I__5377 (
            .O(N__24425),
            .I(N__24422));
    LocalMux I__5376 (
            .O(N__24422),
            .I(N__24419));
    Odrv4 I__5375 (
            .O(N__24419),
            .I(\eeprom.number_of_bytes_7_N_68_7 ));
    InMux I__5374 (
            .O(N__24416),
            .I(N__24413));
    LocalMux I__5373 (
            .O(N__24413),
            .I(\eeprom.number_of_bytes_7_N_68_9 ));
    InMux I__5372 (
            .O(N__24410),
            .I(N__24407));
    LocalMux I__5371 (
            .O(N__24407),
            .I(\eeprom.number_of_bytes_7_N_68_10 ));
    CascadeMux I__5370 (
            .O(N__24404),
            .I(\eeprom.n4307_cascade_ ));
    InMux I__5369 (
            .O(N__24401),
            .I(N__24398));
    LocalMux I__5368 (
            .O(N__24398),
            .I(\eeprom.number_of_bytes_7_N_68_11 ));
    InMux I__5367 (
            .O(N__24395),
            .I(N__24392));
    LocalMux I__5366 (
            .O(N__24392),
            .I(\eeprom.number_of_bytes_7_N_68_12 ));
    InMux I__5365 (
            .O(N__24389),
            .I(N__24386));
    LocalMux I__5364 (
            .O(N__24386),
            .I(\eeprom.number_of_bytes_7_N_68_13 ));
    CascadeMux I__5363 (
            .O(N__24383),
            .I(\eeprom.n4313_cascade_ ));
    InMux I__5362 (
            .O(N__24380),
            .I(N__24377));
    LocalMux I__5361 (
            .O(N__24377),
            .I(\eeprom.number_of_bytes_7_N_68_14 ));
    IoInMux I__5360 (
            .O(N__24374),
            .I(N__24371));
    LocalMux I__5359 (
            .O(N__24371),
            .I(N__24368));
    IoSpan4Mux I__5358 (
            .O(N__24368),
            .I(N__24365));
    Span4Mux_s3_h I__5357 (
            .O(N__24365),
            .I(N__24362));
    Sp12to4 I__5356 (
            .O(N__24362),
            .I(N__24359));
    Span12Mux_h I__5355 (
            .O(N__24359),
            .I(N__24356));
    Span12Mux_v I__5354 (
            .O(N__24356),
            .I(N__24353));
    Odrv12 I__5353 (
            .O(N__24353),
            .I(sda_enable));
    ClkMux I__5352 (
            .O(N__24350),
            .I(N__24323));
    ClkMux I__5351 (
            .O(N__24349),
            .I(N__24323));
    ClkMux I__5350 (
            .O(N__24348),
            .I(N__24323));
    ClkMux I__5349 (
            .O(N__24347),
            .I(N__24323));
    ClkMux I__5348 (
            .O(N__24346),
            .I(N__24323));
    ClkMux I__5347 (
            .O(N__24345),
            .I(N__24323));
    ClkMux I__5346 (
            .O(N__24344),
            .I(N__24323));
    ClkMux I__5345 (
            .O(N__24343),
            .I(N__24323));
    ClkMux I__5344 (
            .O(N__24342),
            .I(N__24323));
    GlobalMux I__5343 (
            .O(N__24323),
            .I(N__24320));
    gio2CtrlBuf I__5342 (
            .O(N__24320),
            .I(CLK_N));
    InMux I__5341 (
            .O(N__24317),
            .I(N__24314));
    LocalMux I__5340 (
            .O(N__24314),
            .I(N__24311));
    Odrv4 I__5339 (
            .O(N__24311),
            .I(\eeprom.number_of_bytes_7_N_68_2 ));
    InMux I__5338 (
            .O(N__24308),
            .I(N__24305));
    LocalMux I__5337 (
            .O(N__24305),
            .I(N__24302));
    Odrv12 I__5336 (
            .O(N__24302),
            .I(\eeprom.number_of_bytes_7_N_68_0 ));
    InMux I__5335 (
            .O(N__24299),
            .I(N__24296));
    LocalMux I__5334 (
            .O(N__24296),
            .I(N__24293));
    Odrv12 I__5333 (
            .O(N__24293),
            .I(\eeprom.number_of_bytes_7_N_68_1 ));
    InMux I__5332 (
            .O(N__24290),
            .I(N__24287));
    LocalMux I__5331 (
            .O(N__24287),
            .I(\eeprom.n4295 ));
    CascadeMux I__5330 (
            .O(N__24284),
            .I(N__24280));
    InMux I__5329 (
            .O(N__24283),
            .I(N__24277));
    InMux I__5328 (
            .O(N__24280),
            .I(N__24274));
    LocalMux I__5327 (
            .O(N__24277),
            .I(N__24270));
    LocalMux I__5326 (
            .O(N__24274),
            .I(N__24267));
    CascadeMux I__5325 (
            .O(N__24273),
            .I(N__24264));
    Span4Mux_h I__5324 (
            .O(N__24270),
            .I(N__24261));
    Span4Mux_h I__5323 (
            .O(N__24267),
            .I(N__24258));
    InMux I__5322 (
            .O(N__24264),
            .I(N__24255));
    Odrv4 I__5321 (
            .O(N__24261),
            .I(\eeprom.n3111 ));
    Odrv4 I__5320 (
            .O(N__24258),
            .I(\eeprom.n3111 ));
    LocalMux I__5319 (
            .O(N__24255),
            .I(\eeprom.n3111 ));
    InMux I__5318 (
            .O(N__24248),
            .I(N__24245));
    LocalMux I__5317 (
            .O(N__24245),
            .I(N__24241));
    CascadeMux I__5316 (
            .O(N__24244),
            .I(N__24238));
    Span4Mux_v I__5315 (
            .O(N__24241),
            .I(N__24235));
    InMux I__5314 (
            .O(N__24238),
            .I(N__24232));
    Span4Mux_h I__5313 (
            .O(N__24235),
            .I(N__24228));
    LocalMux I__5312 (
            .O(N__24232),
            .I(N__24225));
    InMux I__5311 (
            .O(N__24231),
            .I(N__24222));
    Odrv4 I__5310 (
            .O(N__24228),
            .I(\eeprom.n3109 ));
    Odrv4 I__5309 (
            .O(N__24225),
            .I(\eeprom.n3109 ));
    LocalMux I__5308 (
            .O(N__24222),
            .I(\eeprom.n3109 ));
    InMux I__5307 (
            .O(N__24215),
            .I(N__24212));
    LocalMux I__5306 (
            .O(N__24212),
            .I(N__24209));
    Span4Mux_v I__5305 (
            .O(N__24209),
            .I(N__24205));
    InMux I__5304 (
            .O(N__24208),
            .I(N__24202));
    Span4Mux_h I__5303 (
            .O(N__24205),
            .I(N__24198));
    LocalMux I__5302 (
            .O(N__24202),
            .I(N__24195));
    InMux I__5301 (
            .O(N__24201),
            .I(N__24192));
    Odrv4 I__5300 (
            .O(N__24198),
            .I(\eeprom.n3110 ));
    Odrv4 I__5299 (
            .O(N__24195),
            .I(\eeprom.n3110 ));
    LocalMux I__5298 (
            .O(N__24192),
            .I(\eeprom.n3110 ));
    CascadeMux I__5297 (
            .O(N__24185),
            .I(N__24182));
    InMux I__5296 (
            .O(N__24182),
            .I(N__24179));
    LocalMux I__5295 (
            .O(N__24179),
            .I(N__24175));
    InMux I__5294 (
            .O(N__24178),
            .I(N__24172));
    Span4Mux_h I__5293 (
            .O(N__24175),
            .I(N__24168));
    LocalMux I__5292 (
            .O(N__24172),
            .I(N__24165));
    InMux I__5291 (
            .O(N__24171),
            .I(N__24162));
    Odrv4 I__5290 (
            .O(N__24168),
            .I(\eeprom.n3107 ));
    Odrv4 I__5289 (
            .O(N__24165),
            .I(\eeprom.n3107 ));
    LocalMux I__5288 (
            .O(N__24162),
            .I(\eeprom.n3107 ));
    InMux I__5287 (
            .O(N__24155),
            .I(N__24152));
    LocalMux I__5286 (
            .O(N__24152),
            .I(N__24149));
    Odrv4 I__5285 (
            .O(N__24149),
            .I(\eeprom.n4909 ));
    CascadeMux I__5284 (
            .O(N__24146),
            .I(N__24143));
    InMux I__5283 (
            .O(N__24143),
            .I(N__24140));
    LocalMux I__5282 (
            .O(N__24140),
            .I(N__24137));
    Odrv4 I__5281 (
            .O(N__24137),
            .I(\eeprom.n3716_adj_439 ));
    InMux I__5280 (
            .O(N__24134),
            .I(\eeprom.n3780 ));
    InMux I__5279 (
            .O(N__24131),
            .I(\eeprom.n3781 ));
    InMux I__5278 (
            .O(N__24128),
            .I(N__24125));
    LocalMux I__5277 (
            .O(N__24125),
            .I(N__24122));
    Odrv4 I__5276 (
            .O(N__24122),
            .I(\eeprom.n4915 ));
    CascadeMux I__5275 (
            .O(N__24119),
            .I(N__24116));
    InMux I__5274 (
            .O(N__24116),
            .I(N__24113));
    LocalMux I__5273 (
            .O(N__24113),
            .I(N__24110));
    Odrv4 I__5272 (
            .O(N__24110),
            .I(\eeprom.n3714_adj_442 ));
    InMux I__5271 (
            .O(N__24107),
            .I(\eeprom.n3782 ));
    InMux I__5270 (
            .O(N__24104),
            .I(\eeprom.n3783 ));
    InMux I__5269 (
            .O(N__24101),
            .I(N__24098));
    LocalMux I__5268 (
            .O(N__24098),
            .I(\eeprom.n4921 ));
    CascadeMux I__5267 (
            .O(N__24095),
            .I(N__24092));
    InMux I__5266 (
            .O(N__24092),
            .I(N__24088));
    InMux I__5265 (
            .O(N__24091),
            .I(N__24085));
    LocalMux I__5264 (
            .O(N__24088),
            .I(\eeprom.n3712_adj_444 ));
    LocalMux I__5263 (
            .O(N__24085),
            .I(\eeprom.n3712_adj_444 ));
    InMux I__5262 (
            .O(N__24080),
            .I(\eeprom.n3784 ));
    CascadeMux I__5261 (
            .O(N__24077),
            .I(N__24071));
    CascadeMux I__5260 (
            .O(N__24076),
            .I(N__24067));
    CascadeMux I__5259 (
            .O(N__24075),
            .I(N__24063));
    InMux I__5258 (
            .O(N__24074),
            .I(N__24044));
    InMux I__5257 (
            .O(N__24071),
            .I(N__24044));
    InMux I__5256 (
            .O(N__24070),
            .I(N__24044));
    InMux I__5255 (
            .O(N__24067),
            .I(N__24044));
    InMux I__5254 (
            .O(N__24066),
            .I(N__24044));
    InMux I__5253 (
            .O(N__24063),
            .I(N__24044));
    InMux I__5252 (
            .O(N__24062),
            .I(N__24044));
    CascadeMux I__5251 (
            .O(N__24061),
            .I(N__24038));
    CascadeMux I__5250 (
            .O(N__24060),
            .I(N__24034));
    InMux I__5249 (
            .O(N__24059),
            .I(N__24030));
    LocalMux I__5248 (
            .O(N__24044),
            .I(N__24027));
    InMux I__5247 (
            .O(N__24043),
            .I(N__24024));
    InMux I__5246 (
            .O(N__24042),
            .I(N__24011));
    InMux I__5245 (
            .O(N__24041),
            .I(N__24011));
    InMux I__5244 (
            .O(N__24038),
            .I(N__24011));
    InMux I__5243 (
            .O(N__24037),
            .I(N__24011));
    InMux I__5242 (
            .O(N__24034),
            .I(N__24011));
    InMux I__5241 (
            .O(N__24033),
            .I(N__24011));
    LocalMux I__5240 (
            .O(N__24030),
            .I(N__24008));
    Span4Mux_h I__5239 (
            .O(N__24027),
            .I(N__24005));
    LocalMux I__5238 (
            .O(N__24024),
            .I(N__23999));
    LocalMux I__5237 (
            .O(N__24011),
            .I(N__23999));
    Span12Mux_v I__5236 (
            .O(N__24008),
            .I(N__23996));
    Span4Mux_h I__5235 (
            .O(N__24005),
            .I(N__23993));
    InMux I__5234 (
            .O(N__24004),
            .I(N__23990));
    Span12Mux_h I__5233 (
            .O(N__23999),
            .I(N__23987));
    Span12Mux_h I__5232 (
            .O(N__23996),
            .I(N__23984));
    Span4Mux_h I__5231 (
            .O(N__23993),
            .I(N__23981));
    LocalMux I__5230 (
            .O(N__23990),
            .I(N__23978));
    Odrv12 I__5229 (
            .O(N__23987),
            .I(\eeprom.n2 ));
    Odrv12 I__5228 (
            .O(N__23984),
            .I(\eeprom.n2 ));
    Odrv4 I__5227 (
            .O(N__23981),
            .I(\eeprom.n2 ));
    Odrv4 I__5226 (
            .O(N__23978),
            .I(\eeprom.n2 ));
    InMux I__5225 (
            .O(N__23969),
            .I(N__23966));
    LocalMux I__5224 (
            .O(N__23966),
            .I(\eeprom.n4924 ));
    InMux I__5223 (
            .O(N__23963),
            .I(\eeprom.n3785 ));
    CascadeMux I__5222 (
            .O(N__23960),
            .I(N__23956));
    InMux I__5221 (
            .O(N__23959),
            .I(N__23951));
    InMux I__5220 (
            .O(N__23956),
            .I(N__23951));
    LocalMux I__5219 (
            .O(N__23951),
            .I(\eeprom.n3713_adj_443 ));
    InMux I__5218 (
            .O(N__23948),
            .I(N__23945));
    LocalMux I__5217 (
            .O(N__23945),
            .I(\eeprom.n4918 ));
    InMux I__5216 (
            .O(N__23942),
            .I(N__23939));
    LocalMux I__5215 (
            .O(N__23939),
            .I(N__23936));
    Odrv4 I__5214 (
            .O(N__23936),
            .I(\eeprom.number_of_bytes_7_N_68_5 ));
    InMux I__5213 (
            .O(N__23933),
            .I(N__23930));
    LocalMux I__5212 (
            .O(N__23930),
            .I(N__23927));
    Odrv12 I__5211 (
            .O(N__23927),
            .I(\eeprom.number_of_bytes_7_N_68_4 ));
    CascadeMux I__5210 (
            .O(N__23924),
            .I(N__23921));
    InMux I__5209 (
            .O(N__23921),
            .I(N__23918));
    LocalMux I__5208 (
            .O(N__23918),
            .I(N__23915));
    Odrv12 I__5207 (
            .O(N__23915),
            .I(\eeprom.number_of_bytes_7_N_68_3 ));
    InMux I__5206 (
            .O(N__23912),
            .I(N__23909));
    LocalMux I__5205 (
            .O(N__23909),
            .I(N__23905));
    InMux I__5204 (
            .O(N__23908),
            .I(N__23902));
    Span4Mux_v I__5203 (
            .O(N__23905),
            .I(N__23898));
    LocalMux I__5202 (
            .O(N__23902),
            .I(N__23895));
    InMux I__5201 (
            .O(N__23901),
            .I(N__23892));
    Span4Mux_h I__5200 (
            .O(N__23898),
            .I(N__23886));
    Span4Mux_v I__5199 (
            .O(N__23895),
            .I(N__23886));
    LocalMux I__5198 (
            .O(N__23892),
            .I(N__23883));
    InMux I__5197 (
            .O(N__23891),
            .I(N__23880));
    Sp12to4 I__5196 (
            .O(N__23886),
            .I(N__23877));
    Span4Mux_v I__5195 (
            .O(N__23883),
            .I(N__23874));
    LocalMux I__5194 (
            .O(N__23880),
            .I(\eeprom.delay_counter_1 ));
    Odrv12 I__5193 (
            .O(N__23877),
            .I(\eeprom.delay_counter_1 ));
    Odrv4 I__5192 (
            .O(N__23874),
            .I(\eeprom.delay_counter_1 ));
    InMux I__5191 (
            .O(N__23867),
            .I(N__23864));
    LocalMux I__5190 (
            .O(N__23864),
            .I(N__23861));
    Span12Mux_h I__5189 (
            .O(N__23861),
            .I(N__23858));
    Odrv12 I__5188 (
            .O(N__23858),
            .I(\eeprom.n3724_adj_335 ));
    InMux I__5187 (
            .O(N__23855),
            .I(\eeprom.n3772 ));
    InMux I__5186 (
            .O(N__23852),
            .I(N__23849));
    LocalMux I__5185 (
            .O(N__23849),
            .I(N__23846));
    Span4Mux_v I__5184 (
            .O(N__23846),
            .I(N__23842));
    InMux I__5183 (
            .O(N__23845),
            .I(N__23839));
    Span4Mux_v I__5182 (
            .O(N__23842),
            .I(N__23835));
    LocalMux I__5181 (
            .O(N__23839),
            .I(N__23832));
    CascadeMux I__5180 (
            .O(N__23838),
            .I(N__23829));
    Sp12to4 I__5179 (
            .O(N__23835),
            .I(N__23823));
    Span12Mux_v I__5178 (
            .O(N__23832),
            .I(N__23823));
    InMux I__5177 (
            .O(N__23829),
            .I(N__23820));
    InMux I__5176 (
            .O(N__23828),
            .I(N__23817));
    Span12Mux_h I__5175 (
            .O(N__23823),
            .I(N__23814));
    LocalMux I__5174 (
            .O(N__23820),
            .I(N__23811));
    LocalMux I__5173 (
            .O(N__23817),
            .I(\eeprom.delay_counter_2 ));
    Odrv12 I__5172 (
            .O(N__23814),
            .I(\eeprom.delay_counter_2 ));
    Odrv4 I__5171 (
            .O(N__23811),
            .I(\eeprom.delay_counter_2 ));
    CascadeMux I__5170 (
            .O(N__23804),
            .I(N__23801));
    InMux I__5169 (
            .O(N__23801),
            .I(N__23798));
    LocalMux I__5168 (
            .O(N__23798),
            .I(N__23795));
    Odrv4 I__5167 (
            .O(N__23795),
            .I(\eeprom.n3723_adj_334 ));
    InMux I__5166 (
            .O(N__23792),
            .I(\eeprom.n3773 ));
    InMux I__5165 (
            .O(N__23789),
            .I(N__23785));
    CascadeMux I__5164 (
            .O(N__23788),
            .I(N__23782));
    LocalMux I__5163 (
            .O(N__23785),
            .I(N__23779));
    InMux I__5162 (
            .O(N__23782),
            .I(N__23776));
    Span12Mux_h I__5161 (
            .O(N__23779),
            .I(N__23773));
    LocalMux I__5160 (
            .O(N__23776),
            .I(N__23769));
    Span12Mux_h I__5159 (
            .O(N__23773),
            .I(N__23765));
    InMux I__5158 (
            .O(N__23772),
            .I(N__23762));
    Span4Mux_v I__5157 (
            .O(N__23769),
            .I(N__23759));
    InMux I__5156 (
            .O(N__23768),
            .I(N__23756));
    Odrv12 I__5155 (
            .O(N__23765),
            .I(\eeprom.delay_counter_3 ));
    LocalMux I__5154 (
            .O(N__23762),
            .I(\eeprom.delay_counter_3 ));
    Odrv4 I__5153 (
            .O(N__23759),
            .I(\eeprom.delay_counter_3 ));
    LocalMux I__5152 (
            .O(N__23756),
            .I(\eeprom.delay_counter_3 ));
    InMux I__5151 (
            .O(N__23747),
            .I(N__23744));
    LocalMux I__5150 (
            .O(N__23744),
            .I(N__23741));
    Span4Mux_v I__5149 (
            .O(N__23741),
            .I(N__23738));
    Span4Mux_h I__5148 (
            .O(N__23738),
            .I(N__23735));
    Span4Mux_h I__5147 (
            .O(N__23735),
            .I(N__23732));
    Odrv4 I__5146 (
            .O(N__23732),
            .I(\eeprom.n3722_adj_433 ));
    InMux I__5145 (
            .O(N__23729),
            .I(\eeprom.n3774 ));
    InMux I__5144 (
            .O(N__23726),
            .I(N__23723));
    LocalMux I__5143 (
            .O(N__23723),
            .I(N__23719));
    InMux I__5142 (
            .O(N__23722),
            .I(N__23716));
    Span4Mux_v I__5141 (
            .O(N__23719),
            .I(N__23711));
    LocalMux I__5140 (
            .O(N__23716),
            .I(N__23711));
    Span4Mux_h I__5139 (
            .O(N__23711),
            .I(N__23707));
    InMux I__5138 (
            .O(N__23710),
            .I(N__23704));
    Span4Mux_h I__5137 (
            .O(N__23707),
            .I(N__23698));
    LocalMux I__5136 (
            .O(N__23704),
            .I(N__23698));
    InMux I__5135 (
            .O(N__23703),
            .I(N__23695));
    Span4Mux_h I__5134 (
            .O(N__23698),
            .I(N__23692));
    LocalMux I__5133 (
            .O(N__23695),
            .I(\eeprom.delay_counter_4 ));
    Odrv4 I__5132 (
            .O(N__23692),
            .I(\eeprom.delay_counter_4 ));
    CascadeMux I__5131 (
            .O(N__23687),
            .I(N__23684));
    InMux I__5130 (
            .O(N__23684),
            .I(N__23681));
    LocalMux I__5129 (
            .O(N__23681),
            .I(N__23678));
    Odrv4 I__5128 (
            .O(N__23678),
            .I(\eeprom.n3721_adj_434 ));
    InMux I__5127 (
            .O(N__23675),
            .I(\eeprom.n3775 ));
    InMux I__5126 (
            .O(N__23672),
            .I(N__23669));
    LocalMux I__5125 (
            .O(N__23669),
            .I(N__23666));
    Span4Mux_h I__5124 (
            .O(N__23666),
            .I(N__23662));
    InMux I__5123 (
            .O(N__23665),
            .I(N__23659));
    Span4Mux_h I__5122 (
            .O(N__23662),
            .I(N__23653));
    LocalMux I__5121 (
            .O(N__23659),
            .I(N__23653));
    CascadeMux I__5120 (
            .O(N__23658),
            .I(N__23650));
    Span4Mux_h I__5119 (
            .O(N__23653),
            .I(N__23646));
    InMux I__5118 (
            .O(N__23650),
            .I(N__23643));
    InMux I__5117 (
            .O(N__23649),
            .I(N__23640));
    Span4Mux_h I__5116 (
            .O(N__23646),
            .I(N__23635));
    LocalMux I__5115 (
            .O(N__23643),
            .I(N__23635));
    LocalMux I__5114 (
            .O(N__23640),
            .I(\eeprom.delay_counter_5 ));
    Odrv4 I__5113 (
            .O(N__23635),
            .I(\eeprom.delay_counter_5 ));
    InMux I__5112 (
            .O(N__23630),
            .I(N__23627));
    LocalMux I__5111 (
            .O(N__23627),
            .I(N__23624));
    Odrv12 I__5110 (
            .O(N__23624),
            .I(\eeprom.n3720_adj_435 ));
    InMux I__5109 (
            .O(N__23621),
            .I(\eeprom.n3776 ));
    InMux I__5108 (
            .O(N__23618),
            .I(N__23615));
    LocalMux I__5107 (
            .O(N__23615),
            .I(N__23612));
    Span4Mux_h I__5106 (
            .O(N__23612),
            .I(N__23608));
    InMux I__5105 (
            .O(N__23611),
            .I(N__23605));
    Span4Mux_h I__5104 (
            .O(N__23608),
            .I(N__23600));
    LocalMux I__5103 (
            .O(N__23605),
            .I(N__23600));
    Span4Mux_h I__5102 (
            .O(N__23600),
            .I(N__23596));
    InMux I__5101 (
            .O(N__23599),
            .I(N__23592));
    Span4Mux_h I__5100 (
            .O(N__23596),
            .I(N__23589));
    InMux I__5099 (
            .O(N__23595),
            .I(N__23586));
    LocalMux I__5098 (
            .O(N__23592),
            .I(\eeprom.delay_counter_6 ));
    Odrv4 I__5097 (
            .O(N__23589),
            .I(\eeprom.delay_counter_6 ));
    LocalMux I__5096 (
            .O(N__23586),
            .I(\eeprom.delay_counter_6 ));
    CascadeMux I__5095 (
            .O(N__23579),
            .I(N__23576));
    InMux I__5094 (
            .O(N__23576),
            .I(N__23573));
    LocalMux I__5093 (
            .O(N__23573),
            .I(N__23570));
    Span12Mux_h I__5092 (
            .O(N__23570),
            .I(N__23567));
    Odrv12 I__5091 (
            .O(N__23567),
            .I(\eeprom.n3719_adj_436 ));
    InMux I__5090 (
            .O(N__23564),
            .I(\eeprom.n3777 ));
    InMux I__5089 (
            .O(N__23561),
            .I(\eeprom.n3778 ));
    InMux I__5088 (
            .O(N__23558),
            .I(bfn_15_21_0_));
    CascadeMux I__5087 (
            .O(N__23555),
            .I(\eeprom.n3617_adj_346_cascade_ ));
    InMux I__5086 (
            .O(N__23552),
            .I(N__23549));
    LocalMux I__5085 (
            .O(N__23549),
            .I(\eeprom.n4619 ));
    CascadeMux I__5084 (
            .O(N__23546),
            .I(\eeprom.n4427_cascade_ ));
    InMux I__5083 (
            .O(N__23543),
            .I(N__23540));
    LocalMux I__5082 (
            .O(N__23540),
            .I(\eeprom.n3596_adj_454 ));
    CascadeMux I__5081 (
            .O(N__23537),
            .I(\eeprom.n28_adj_455_cascade_ ));
    InMux I__5080 (
            .O(N__23534),
            .I(N__23531));
    LocalMux I__5079 (
            .O(N__23531),
            .I(\eeprom.n4567 ));
    CascadeMux I__5078 (
            .O(N__23528),
            .I(\eeprom.n3628_adj_437_cascade_ ));
    CascadeMux I__5077 (
            .O(N__23525),
            .I(\eeprom.n3716_adj_439_cascade_ ));
    InMux I__5076 (
            .O(N__23522),
            .I(N__23519));
    LocalMux I__5075 (
            .O(N__23519),
            .I(\eeprom.n3605_adj_453 ));
    CascadeMux I__5074 (
            .O(N__23516),
            .I(\eeprom.n3618_adj_350_cascade_ ));
    InMux I__5073 (
            .O(N__23513),
            .I(N__23510));
    LocalMux I__5072 (
            .O(N__23510),
            .I(\eeprom.n4623 ));
    InMux I__5071 (
            .O(N__23507),
            .I(N__23504));
    LocalMux I__5070 (
            .O(N__23504),
            .I(\eeprom.n4425 ));
    InMux I__5069 (
            .O(N__23501),
            .I(N__23498));
    LocalMux I__5068 (
            .O(N__23498),
            .I(N__23495));
    Span4Mux_v I__5067 (
            .O(N__23495),
            .I(N__23492));
    Span4Mux_h I__5066 (
            .O(N__23492),
            .I(N__23489));
    Span4Mux_h I__5065 (
            .O(N__23489),
            .I(N__23485));
    InMux I__5064 (
            .O(N__23488),
            .I(N__23482));
    Span4Mux_h I__5063 (
            .O(N__23485),
            .I(N__23476));
    LocalMux I__5062 (
            .O(N__23482),
            .I(N__23476));
    InMux I__5061 (
            .O(N__23481),
            .I(N__23472));
    Span4Mux_v I__5060 (
            .O(N__23476),
            .I(N__23469));
    InMux I__5059 (
            .O(N__23475),
            .I(N__23466));
    LocalMux I__5058 (
            .O(N__23472),
            .I(\eeprom.delay_counter_0 ));
    Odrv4 I__5057 (
            .O(N__23469),
            .I(\eeprom.delay_counter_0 ));
    LocalMux I__5056 (
            .O(N__23466),
            .I(\eeprom.delay_counter_0 ));
    CascadeMux I__5055 (
            .O(N__23459),
            .I(N__23456));
    InMux I__5054 (
            .O(N__23456),
            .I(N__23453));
    LocalMux I__5053 (
            .O(N__23453),
            .I(N__23450));
    Span12Mux_v I__5052 (
            .O(N__23450),
            .I(N__23447));
    Span12Mux_h I__5051 (
            .O(N__23447),
            .I(N__23444));
    Odrv12 I__5050 (
            .O(N__23444),
            .I(\eeprom.n1166 ));
    InMux I__5049 (
            .O(N__23441),
            .I(bfn_15_20_0_));
    CascadeMux I__5048 (
            .O(N__23438),
            .I(\eeprom.n3515_adj_370_cascade_ ));
    CascadeMux I__5047 (
            .O(N__23435),
            .I(N__23432));
    InMux I__5046 (
            .O(N__23432),
            .I(N__23429));
    LocalMux I__5045 (
            .O(N__23429),
            .I(\eeprom.n4727 ));
    InMux I__5044 (
            .O(N__23426),
            .I(N__23422));
    InMux I__5043 (
            .O(N__23425),
            .I(N__23418));
    LocalMux I__5042 (
            .O(N__23422),
            .I(N__23415));
    InMux I__5041 (
            .O(N__23421),
            .I(N__23412));
    LocalMux I__5040 (
            .O(N__23418),
            .I(N__23409));
    Span12Mux_v I__5039 (
            .O(N__23415),
            .I(N__23406));
    LocalMux I__5038 (
            .O(N__23412),
            .I(N__23403));
    Span4Mux_v I__5037 (
            .O(N__23409),
            .I(N__23400));
    Span12Mux_h I__5036 (
            .O(N__23406),
            .I(N__23397));
    Span12Mux_v I__5035 (
            .O(N__23403),
            .I(N__23392));
    Sp12to4 I__5034 (
            .O(N__23400),
            .I(N__23392));
    Odrv12 I__5033 (
            .O(N__23397),
            .I(\eeprom.n3419 ));
    Odrv12 I__5032 (
            .O(N__23392),
            .I(\eeprom.n3419 ));
    InMux I__5031 (
            .O(N__23387),
            .I(N__23384));
    LocalMux I__5030 (
            .O(N__23384),
            .I(\eeprom.n3486 ));
    InMux I__5029 (
            .O(N__23381),
            .I(N__23378));
    LocalMux I__5028 (
            .O(N__23378),
            .I(\eeprom.n3471_adj_386 ));
    CascadeMux I__5027 (
            .O(N__23375),
            .I(N__23366));
    InMux I__5026 (
            .O(N__23374),
            .I(N__23354));
    InMux I__5025 (
            .O(N__23373),
            .I(N__23354));
    InMux I__5024 (
            .O(N__23372),
            .I(N__23354));
    CascadeMux I__5023 (
            .O(N__23371),
            .I(N__23349));
    CascadeMux I__5022 (
            .O(N__23370),
            .I(N__23342));
    CascadeMux I__5021 (
            .O(N__23369),
            .I(N__23338));
    InMux I__5020 (
            .O(N__23366),
            .I(N__23333));
    InMux I__5019 (
            .O(N__23365),
            .I(N__23333));
    CascadeMux I__5018 (
            .O(N__23364),
            .I(N__23328));
    CascadeMux I__5017 (
            .O(N__23363),
            .I(N__23325));
    InMux I__5016 (
            .O(N__23362),
            .I(N__23319));
    InMux I__5015 (
            .O(N__23361),
            .I(N__23319));
    LocalMux I__5014 (
            .O(N__23354),
            .I(N__23316));
    InMux I__5013 (
            .O(N__23353),
            .I(N__23313));
    InMux I__5012 (
            .O(N__23352),
            .I(N__23306));
    InMux I__5011 (
            .O(N__23349),
            .I(N__23306));
    InMux I__5010 (
            .O(N__23348),
            .I(N__23306));
    InMux I__5009 (
            .O(N__23347),
            .I(N__23299));
    InMux I__5008 (
            .O(N__23346),
            .I(N__23299));
    InMux I__5007 (
            .O(N__23345),
            .I(N__23299));
    InMux I__5006 (
            .O(N__23342),
            .I(N__23294));
    InMux I__5005 (
            .O(N__23341),
            .I(N__23294));
    InMux I__5004 (
            .O(N__23338),
            .I(N__23291));
    LocalMux I__5003 (
            .O(N__23333),
            .I(N__23288));
    InMux I__5002 (
            .O(N__23332),
            .I(N__23277));
    InMux I__5001 (
            .O(N__23331),
            .I(N__23277));
    InMux I__5000 (
            .O(N__23328),
            .I(N__23277));
    InMux I__4999 (
            .O(N__23325),
            .I(N__23277));
    InMux I__4998 (
            .O(N__23324),
            .I(N__23277));
    LocalMux I__4997 (
            .O(N__23319),
            .I(N__23272));
    Span4Mux_h I__4996 (
            .O(N__23316),
            .I(N__23272));
    LocalMux I__4995 (
            .O(N__23313),
            .I(\eeprom.n3430 ));
    LocalMux I__4994 (
            .O(N__23306),
            .I(\eeprom.n3430 ));
    LocalMux I__4993 (
            .O(N__23299),
            .I(\eeprom.n3430 ));
    LocalMux I__4992 (
            .O(N__23294),
            .I(\eeprom.n3430 ));
    LocalMux I__4991 (
            .O(N__23291),
            .I(\eeprom.n3430 ));
    Odrv4 I__4990 (
            .O(N__23288),
            .I(\eeprom.n3430 ));
    LocalMux I__4989 (
            .O(N__23277),
            .I(\eeprom.n3430 ));
    Odrv4 I__4988 (
            .O(N__23272),
            .I(\eeprom.n3430 ));
    CascadeMux I__4987 (
            .O(N__23255),
            .I(N__23251));
    InMux I__4986 (
            .O(N__23254),
            .I(N__23248));
    InMux I__4985 (
            .O(N__23251),
            .I(N__23245));
    LocalMux I__4984 (
            .O(N__23248),
            .I(N__23239));
    LocalMux I__4983 (
            .O(N__23245),
            .I(N__23239));
    InMux I__4982 (
            .O(N__23244),
            .I(N__23236));
    Odrv12 I__4981 (
            .O(N__23239),
            .I(\eeprom.n3404 ));
    LocalMux I__4980 (
            .O(N__23236),
            .I(\eeprom.n3404 ));
    CascadeMux I__4979 (
            .O(N__23231),
            .I(\eeprom.n3615_adj_344_cascade_ ));
    CascadeMux I__4978 (
            .O(N__23228),
            .I(\eeprom.n3714_adj_442_cascade_ ));
    CascadeMux I__4977 (
            .O(N__23225),
            .I(\eeprom.n3034_cascade_ ));
    InMux I__4976 (
            .O(N__23222),
            .I(N__23217));
    InMux I__4975 (
            .O(N__23221),
            .I(N__23214));
    InMux I__4974 (
            .O(N__23220),
            .I(N__23211));
    LocalMux I__4973 (
            .O(N__23217),
            .I(N__23208));
    LocalMux I__4972 (
            .O(N__23214),
            .I(N__23205));
    LocalMux I__4971 (
            .O(N__23211),
            .I(N__23202));
    Span4Mux_h I__4970 (
            .O(N__23208),
            .I(N__23199));
    Span4Mux_v I__4969 (
            .O(N__23205),
            .I(N__23194));
    Span4Mux_h I__4968 (
            .O(N__23202),
            .I(N__23194));
    Odrv4 I__4967 (
            .O(N__23199),
            .I(\eeprom.n3112 ));
    Odrv4 I__4966 (
            .O(N__23194),
            .I(\eeprom.n3112 ));
    InMux I__4965 (
            .O(N__23189),
            .I(N__23185));
    CascadeMux I__4964 (
            .O(N__23188),
            .I(N__23182));
    LocalMux I__4963 (
            .O(N__23185),
            .I(N__23179));
    InMux I__4962 (
            .O(N__23182),
            .I(N__23175));
    Span4Mux_v I__4961 (
            .O(N__23179),
            .I(N__23172));
    InMux I__4960 (
            .O(N__23178),
            .I(N__23169));
    LocalMux I__4959 (
            .O(N__23175),
            .I(N__23166));
    Odrv4 I__4958 (
            .O(N__23172),
            .I(\eeprom.n2912 ));
    LocalMux I__4957 (
            .O(N__23169),
            .I(\eeprom.n2912 ));
    Odrv4 I__4956 (
            .O(N__23166),
            .I(\eeprom.n2912 ));
    CascadeMux I__4955 (
            .O(N__23159),
            .I(N__23156));
    InMux I__4954 (
            .O(N__23156),
            .I(N__23153));
    LocalMux I__4953 (
            .O(N__23153),
            .I(N__23150));
    Span4Mux_h I__4952 (
            .O(N__23150),
            .I(N__23147));
    Odrv4 I__4951 (
            .O(N__23147),
            .I(\eeprom.n2979 ));
    InMux I__4950 (
            .O(N__23144),
            .I(N__23141));
    LocalMux I__4949 (
            .O(N__23141),
            .I(N__23136));
    InMux I__4948 (
            .O(N__23140),
            .I(N__23131));
    InMux I__4947 (
            .O(N__23139),
            .I(N__23131));
    Odrv4 I__4946 (
            .O(N__23136),
            .I(\eeprom.n3103 ));
    LocalMux I__4945 (
            .O(N__23131),
            .I(\eeprom.n3103 ));
    InMux I__4944 (
            .O(N__23126),
            .I(N__23123));
    LocalMux I__4943 (
            .O(N__23123),
            .I(N__23120));
    Span4Mux_h I__4942 (
            .O(N__23120),
            .I(N__23117));
    Odrv4 I__4941 (
            .O(N__23117),
            .I(\eeprom.n4137 ));
    InMux I__4940 (
            .O(N__23114),
            .I(N__23110));
    CascadeMux I__4939 (
            .O(N__23113),
            .I(N__23107));
    LocalMux I__4938 (
            .O(N__23110),
            .I(N__23103));
    InMux I__4937 (
            .O(N__23107),
            .I(N__23100));
    InMux I__4936 (
            .O(N__23106),
            .I(N__23097));
    Span4Mux_h I__4935 (
            .O(N__23103),
            .I(N__23092));
    LocalMux I__4934 (
            .O(N__23100),
            .I(N__23092));
    LocalMux I__4933 (
            .O(N__23097),
            .I(\eeprom.n3417 ));
    Odrv4 I__4932 (
            .O(N__23092),
            .I(\eeprom.n3417 ));
    CascadeMux I__4931 (
            .O(N__23087),
            .I(N__23084));
    InMux I__4930 (
            .O(N__23084),
            .I(N__23081));
    LocalMux I__4929 (
            .O(N__23081),
            .I(\eeprom.n3484_adj_406 ));
    CascadeMux I__4928 (
            .O(N__23078),
            .I(N__23074));
    InMux I__4927 (
            .O(N__23077),
            .I(N__23070));
    InMux I__4926 (
            .O(N__23074),
            .I(N__23067));
    InMux I__4925 (
            .O(N__23073),
            .I(N__23064));
    LocalMux I__4924 (
            .O(N__23070),
            .I(N__23059));
    LocalMux I__4923 (
            .O(N__23067),
            .I(N__23059));
    LocalMux I__4922 (
            .O(N__23064),
            .I(\eeprom.n3418 ));
    Odrv4 I__4921 (
            .O(N__23059),
            .I(\eeprom.n3418 ));
    CascadeMux I__4920 (
            .O(N__23054),
            .I(N__23051));
    InMux I__4919 (
            .O(N__23051),
            .I(N__23048));
    LocalMux I__4918 (
            .O(N__23048),
            .I(\eeprom.n3485 ));
    CascadeMux I__4917 (
            .O(N__23045),
            .I(\eeprom.n3517_adj_374_cascade_ ));
    InMux I__4916 (
            .O(N__23042),
            .I(N__23039));
    LocalMux I__4915 (
            .O(N__23039),
            .I(\eeprom.n4729 ));
    CascadeMux I__4914 (
            .O(N__23036),
            .I(N__23032));
    InMux I__4913 (
            .O(N__23035),
            .I(N__23028));
    InMux I__4912 (
            .O(N__23032),
            .I(N__23025));
    InMux I__4911 (
            .O(N__23031),
            .I(N__23022));
    LocalMux I__4910 (
            .O(N__23028),
            .I(N__23017));
    LocalMux I__4909 (
            .O(N__23025),
            .I(N__23017));
    LocalMux I__4908 (
            .O(N__23022),
            .I(\eeprom.n3416 ));
    Odrv12 I__4907 (
            .O(N__23017),
            .I(\eeprom.n3416 ));
    CascadeMux I__4906 (
            .O(N__23012),
            .I(N__23009));
    InMux I__4905 (
            .O(N__23009),
            .I(N__23006));
    LocalMux I__4904 (
            .O(N__23006),
            .I(\eeprom.n3483_adj_404 ));
    InMux I__4903 (
            .O(N__23003),
            .I(N__23000));
    LocalMux I__4902 (
            .O(N__23000),
            .I(N__22997));
    Span12Mux_h I__4901 (
            .O(N__22997),
            .I(N__22994));
    Odrv12 I__4900 (
            .O(N__22994),
            .I(\eeprom.n31_adj_476 ));
    InMux I__4899 (
            .O(N__22991),
            .I(N__22987));
    InMux I__4898 (
            .O(N__22990),
            .I(N__22984));
    LocalMux I__4897 (
            .O(N__22987),
            .I(N__22980));
    LocalMux I__4896 (
            .O(N__22984),
            .I(N__22974));
    InMux I__4895 (
            .O(N__22983),
            .I(N__22971));
    Span4Mux_v I__4894 (
            .O(N__22980),
            .I(N__22966));
    InMux I__4893 (
            .O(N__22979),
            .I(N__22963));
    InMux I__4892 (
            .O(N__22978),
            .I(N__22960));
    InMux I__4891 (
            .O(N__22977),
            .I(N__22951));
    Span4Mux_h I__4890 (
            .O(N__22974),
            .I(N__22944));
    LocalMux I__4889 (
            .O(N__22971),
            .I(N__22944));
    InMux I__4888 (
            .O(N__22970),
            .I(N__22939));
    InMux I__4887 (
            .O(N__22969),
            .I(N__22935));
    Span4Mux_h I__4886 (
            .O(N__22966),
            .I(N__22930));
    LocalMux I__4885 (
            .O(N__22963),
            .I(N__22930));
    LocalMux I__4884 (
            .O(N__22960),
            .I(N__22927));
    InMux I__4883 (
            .O(N__22959),
            .I(N__22924));
    InMux I__4882 (
            .O(N__22958),
            .I(N__22917));
    InMux I__4881 (
            .O(N__22957),
            .I(N__22912));
    InMux I__4880 (
            .O(N__22956),
            .I(N__22912));
    InMux I__4879 (
            .O(N__22955),
            .I(N__22907));
    InMux I__4878 (
            .O(N__22954),
            .I(N__22907));
    LocalMux I__4877 (
            .O(N__22951),
            .I(N__22903));
    InMux I__4876 (
            .O(N__22950),
            .I(N__22898));
    InMux I__4875 (
            .O(N__22949),
            .I(N__22898));
    Span4Mux_v I__4874 (
            .O(N__22944),
            .I(N__22895));
    InMux I__4873 (
            .O(N__22943),
            .I(N__22892));
    InMux I__4872 (
            .O(N__22942),
            .I(N__22889));
    LocalMux I__4871 (
            .O(N__22939),
            .I(N__22885));
    InMux I__4870 (
            .O(N__22938),
            .I(N__22882));
    LocalMux I__4869 (
            .O(N__22935),
            .I(N__22879));
    Span4Mux_h I__4868 (
            .O(N__22930),
            .I(N__22874));
    Span4Mux_v I__4867 (
            .O(N__22927),
            .I(N__22874));
    LocalMux I__4866 (
            .O(N__22924),
            .I(N__22871));
    InMux I__4865 (
            .O(N__22923),
            .I(N__22862));
    InMux I__4864 (
            .O(N__22922),
            .I(N__22862));
    InMux I__4863 (
            .O(N__22921),
            .I(N__22862));
    InMux I__4862 (
            .O(N__22920),
            .I(N__22862));
    LocalMux I__4861 (
            .O(N__22917),
            .I(N__22855));
    LocalMux I__4860 (
            .O(N__22912),
            .I(N__22855));
    LocalMux I__4859 (
            .O(N__22907),
            .I(N__22855));
    InMux I__4858 (
            .O(N__22906),
            .I(N__22842));
    Span12Mux_h I__4857 (
            .O(N__22903),
            .I(N__22831));
    LocalMux I__4856 (
            .O(N__22898),
            .I(N__22831));
    Sp12to4 I__4855 (
            .O(N__22895),
            .I(N__22831));
    LocalMux I__4854 (
            .O(N__22892),
            .I(N__22831));
    LocalMux I__4853 (
            .O(N__22889),
            .I(N__22831));
    InMux I__4852 (
            .O(N__22888),
            .I(N__22828));
    Span4Mux_v I__4851 (
            .O(N__22885),
            .I(N__22819));
    LocalMux I__4850 (
            .O(N__22882),
            .I(N__22819));
    Span4Mux_v I__4849 (
            .O(N__22879),
            .I(N__22819));
    Span4Mux_h I__4848 (
            .O(N__22874),
            .I(N__22819));
    Span4Mux_h I__4847 (
            .O(N__22871),
            .I(N__22812));
    LocalMux I__4846 (
            .O(N__22862),
            .I(N__22812));
    Span4Mux_h I__4845 (
            .O(N__22855),
            .I(N__22812));
    InMux I__4844 (
            .O(N__22854),
            .I(N__22803));
    InMux I__4843 (
            .O(N__22853),
            .I(N__22803));
    InMux I__4842 (
            .O(N__22852),
            .I(N__22803));
    InMux I__4841 (
            .O(N__22851),
            .I(N__22803));
    InMux I__4840 (
            .O(N__22850),
            .I(N__22794));
    InMux I__4839 (
            .O(N__22849),
            .I(N__22794));
    InMux I__4838 (
            .O(N__22848),
            .I(N__22794));
    InMux I__4837 (
            .O(N__22847),
            .I(N__22794));
    InMux I__4836 (
            .O(N__22846),
            .I(N__22789));
    InMux I__4835 (
            .O(N__22845),
            .I(N__22789));
    LocalMux I__4834 (
            .O(N__22842),
            .I(\eeprom.delay_counter_31 ));
    Odrv12 I__4833 (
            .O(N__22831),
            .I(\eeprom.delay_counter_31 ));
    LocalMux I__4832 (
            .O(N__22828),
            .I(\eeprom.delay_counter_31 ));
    Odrv4 I__4831 (
            .O(N__22819),
            .I(\eeprom.delay_counter_31 ));
    Odrv4 I__4830 (
            .O(N__22812),
            .I(\eeprom.delay_counter_31 ));
    LocalMux I__4829 (
            .O(N__22803),
            .I(\eeprom.delay_counter_31 ));
    LocalMux I__4828 (
            .O(N__22794),
            .I(\eeprom.delay_counter_31 ));
    LocalMux I__4827 (
            .O(N__22789),
            .I(\eeprom.delay_counter_31 ));
    InMux I__4826 (
            .O(N__22772),
            .I(N__22769));
    LocalMux I__4825 (
            .O(N__22769),
            .I(N__22766));
    Span4Mux_h I__4824 (
            .O(N__22766),
            .I(N__22763));
    Odrv4 I__4823 (
            .O(N__22763),
            .I(\eeprom.n24_adj_459 ));
    CascadeMux I__4822 (
            .O(N__22760),
            .I(\eeprom.n4559_cascade_ ));
    CascadeMux I__4821 (
            .O(N__22757),
            .I(\eeprom.n4563_cascade_ ));
    InMux I__4820 (
            .O(N__22754),
            .I(N__22751));
    LocalMux I__4819 (
            .O(N__22751),
            .I(\eeprom.n21_adj_422 ));
    CascadeMux I__4818 (
            .O(N__22748),
            .I(\eeprom.n17_adj_421_cascade_ ));
    CascadeMux I__4817 (
            .O(N__22745),
            .I(\eeprom.n24_cascade_ ));
    InMux I__4816 (
            .O(N__22742),
            .I(N__22739));
    LocalMux I__4815 (
            .O(N__22739),
            .I(\eeprom.n20_adj_423 ));
    InMux I__4814 (
            .O(N__22736),
            .I(\eeprom.n3747 ));
    InMux I__4813 (
            .O(N__22733),
            .I(N__22729));
    InMux I__4812 (
            .O(N__22732),
            .I(N__22726));
    LocalMux I__4811 (
            .O(N__22729),
            .I(N__22723));
    LocalMux I__4810 (
            .O(N__22726),
            .I(N__22720));
    Span4Mux_h I__4809 (
            .O(N__22723),
            .I(N__22715));
    Span4Mux_v I__4808 (
            .O(N__22720),
            .I(N__22715));
    Odrv4 I__4807 (
            .O(N__22715),
            .I(\eeprom.n3397 ));
    InMux I__4806 (
            .O(N__22712),
            .I(\eeprom.n3748 ));
    CascadeMux I__4805 (
            .O(N__22709),
            .I(N__22706));
    InMux I__4804 (
            .O(N__22706),
            .I(N__22703));
    LocalMux I__4803 (
            .O(N__22703),
            .I(\eeprom.n4583 ));
    CascadeMux I__4802 (
            .O(N__22700),
            .I(\eeprom.n31_cascade_ ));
    InMux I__4801 (
            .O(N__22697),
            .I(N__22694));
    LocalMux I__4800 (
            .O(N__22694),
            .I(\eeprom.n4433 ));
    InMux I__4799 (
            .O(N__22691),
            .I(N__22688));
    LocalMux I__4798 (
            .O(N__22688),
            .I(\eeprom.n3598_adj_452 ));
    CascadeMux I__4797 (
            .O(N__22685),
            .I(N__22681));
    InMux I__4796 (
            .O(N__22684),
            .I(N__22678));
    InMux I__4795 (
            .O(N__22681),
            .I(N__22675));
    LocalMux I__4794 (
            .O(N__22678),
            .I(N__22669));
    LocalMux I__4793 (
            .O(N__22675),
            .I(N__22669));
    InMux I__4792 (
            .O(N__22674),
            .I(N__22666));
    Odrv4 I__4791 (
            .O(N__22669),
            .I(\eeprom.n3405 ));
    LocalMux I__4790 (
            .O(N__22666),
            .I(\eeprom.n3405 ));
    InMux I__4789 (
            .O(N__22661),
            .I(N__22658));
    LocalMux I__4788 (
            .O(N__22658),
            .I(N__22655));
    Odrv4 I__4787 (
            .O(N__22655),
            .I(\eeprom.n3472_adj_387 ));
    InMux I__4786 (
            .O(N__22652),
            .I(\eeprom.n3740 ));
    InMux I__4785 (
            .O(N__22649),
            .I(\eeprom.n3741 ));
    CascadeMux I__4784 (
            .O(N__22646),
            .I(N__22642));
    InMux I__4783 (
            .O(N__22645),
            .I(N__22639));
    InMux I__4782 (
            .O(N__22642),
            .I(N__22636));
    LocalMux I__4781 (
            .O(N__22639),
            .I(N__22630));
    LocalMux I__4780 (
            .O(N__22636),
            .I(N__22630));
    InMux I__4779 (
            .O(N__22635),
            .I(N__22627));
    Span4Mux_v I__4778 (
            .O(N__22630),
            .I(N__22622));
    LocalMux I__4777 (
            .O(N__22627),
            .I(N__22622));
    Odrv4 I__4776 (
            .O(N__22622),
            .I(\eeprom.n3403 ));
    InMux I__4775 (
            .O(N__22619),
            .I(N__22616));
    LocalMux I__4774 (
            .O(N__22616),
            .I(\eeprom.n3470_adj_385 ));
    InMux I__4773 (
            .O(N__22613),
            .I(bfn_14_19_0_));
    InMux I__4772 (
            .O(N__22610),
            .I(N__22607));
    LocalMux I__4771 (
            .O(N__22607),
            .I(N__22602));
    InMux I__4770 (
            .O(N__22606),
            .I(N__22597));
    InMux I__4769 (
            .O(N__22605),
            .I(N__22597));
    Odrv4 I__4768 (
            .O(N__22602),
            .I(\eeprom.n3402 ));
    LocalMux I__4767 (
            .O(N__22597),
            .I(\eeprom.n3402 ));
    CascadeMux I__4766 (
            .O(N__22592),
            .I(N__22589));
    InMux I__4765 (
            .O(N__22589),
            .I(N__22586));
    LocalMux I__4764 (
            .O(N__22586),
            .I(N__22583));
    Span4Mux_h I__4763 (
            .O(N__22583),
            .I(N__22580));
    Odrv4 I__4762 (
            .O(N__22580),
            .I(\eeprom.n3469_adj_384 ));
    InMux I__4761 (
            .O(N__22577),
            .I(\eeprom.n3743 ));
    CascadeMux I__4760 (
            .O(N__22574),
            .I(N__22571));
    InMux I__4759 (
            .O(N__22571),
            .I(N__22567));
    CascadeMux I__4758 (
            .O(N__22570),
            .I(N__22564));
    LocalMux I__4757 (
            .O(N__22567),
            .I(N__22560));
    InMux I__4756 (
            .O(N__22564),
            .I(N__22555));
    InMux I__4755 (
            .O(N__22563),
            .I(N__22555));
    Span4Mux_v I__4754 (
            .O(N__22560),
            .I(N__22552));
    LocalMux I__4753 (
            .O(N__22555),
            .I(N__22549));
    Odrv4 I__4752 (
            .O(N__22552),
            .I(\eeprom.n3401 ));
    Odrv4 I__4751 (
            .O(N__22549),
            .I(\eeprom.n3401 ));
    InMux I__4750 (
            .O(N__22544),
            .I(N__22541));
    LocalMux I__4749 (
            .O(N__22541),
            .I(N__22538));
    Span4Mux_h I__4748 (
            .O(N__22538),
            .I(N__22535));
    Odrv4 I__4747 (
            .O(N__22535),
            .I(\eeprom.n3468_adj_383 ));
    InMux I__4746 (
            .O(N__22532),
            .I(\eeprom.n3744 ));
    CascadeMux I__4745 (
            .O(N__22529),
            .I(N__22525));
    InMux I__4744 (
            .O(N__22528),
            .I(N__22521));
    InMux I__4743 (
            .O(N__22525),
            .I(N__22518));
    CascadeMux I__4742 (
            .O(N__22524),
            .I(N__22515));
    LocalMux I__4741 (
            .O(N__22521),
            .I(N__22510));
    LocalMux I__4740 (
            .O(N__22518),
            .I(N__22510));
    InMux I__4739 (
            .O(N__22515),
            .I(N__22507));
    Odrv12 I__4738 (
            .O(N__22510),
            .I(\eeprom.n3400 ));
    LocalMux I__4737 (
            .O(N__22507),
            .I(\eeprom.n3400 ));
    CascadeMux I__4736 (
            .O(N__22502),
            .I(N__22499));
    InMux I__4735 (
            .O(N__22499),
            .I(N__22496));
    LocalMux I__4734 (
            .O(N__22496),
            .I(\eeprom.n3467_adj_382 ));
    InMux I__4733 (
            .O(N__22493),
            .I(\eeprom.n3745 ));
    CascadeMux I__4732 (
            .O(N__22490),
            .I(N__22486));
    InMux I__4731 (
            .O(N__22489),
            .I(N__22483));
    InMux I__4730 (
            .O(N__22486),
            .I(N__22480));
    LocalMux I__4729 (
            .O(N__22483),
            .I(N__22476));
    LocalMux I__4728 (
            .O(N__22480),
            .I(N__22473));
    InMux I__4727 (
            .O(N__22479),
            .I(N__22470));
    Span4Mux_v I__4726 (
            .O(N__22476),
            .I(N__22463));
    Span4Mux_v I__4725 (
            .O(N__22473),
            .I(N__22463));
    LocalMux I__4724 (
            .O(N__22470),
            .I(N__22463));
    Span4Mux_h I__4723 (
            .O(N__22463),
            .I(N__22460));
    Odrv4 I__4722 (
            .O(N__22460),
            .I(\eeprom.n3399 ));
    InMux I__4721 (
            .O(N__22457),
            .I(N__22454));
    LocalMux I__4720 (
            .O(N__22454),
            .I(N__22451));
    Odrv4 I__4719 (
            .O(N__22451),
            .I(\eeprom.n3466_adj_381 ));
    InMux I__4718 (
            .O(N__22448),
            .I(\eeprom.n3746 ));
    InMux I__4717 (
            .O(N__22445),
            .I(N__22440));
    InMux I__4716 (
            .O(N__22444),
            .I(N__22437));
    CascadeMux I__4715 (
            .O(N__22443),
            .I(N__22434));
    LocalMux I__4714 (
            .O(N__22440),
            .I(N__22431));
    LocalMux I__4713 (
            .O(N__22437),
            .I(N__22428));
    InMux I__4712 (
            .O(N__22434),
            .I(N__22425));
    Odrv4 I__4711 (
            .O(N__22431),
            .I(\eeprom.n3398 ));
    Odrv4 I__4710 (
            .O(N__22428),
            .I(\eeprom.n3398 ));
    LocalMux I__4709 (
            .O(N__22425),
            .I(\eeprom.n3398 ));
    CascadeMux I__4708 (
            .O(N__22418),
            .I(N__22415));
    InMux I__4707 (
            .O(N__22415),
            .I(N__22412));
    LocalMux I__4706 (
            .O(N__22412),
            .I(N__22409));
    Odrv4 I__4705 (
            .O(N__22409),
            .I(\eeprom.n3465_adj_380 ));
    CascadeMux I__4704 (
            .O(N__22406),
            .I(N__22402));
    CascadeMux I__4703 (
            .O(N__22405),
            .I(N__22399));
    InMux I__4702 (
            .O(N__22402),
            .I(N__22396));
    InMux I__4701 (
            .O(N__22399),
            .I(N__22393));
    LocalMux I__4700 (
            .O(N__22396),
            .I(N__22388));
    LocalMux I__4699 (
            .O(N__22393),
            .I(N__22388));
    Odrv4 I__4698 (
            .O(N__22388),
            .I(\eeprom.n3413 ));
    InMux I__4697 (
            .O(N__22385),
            .I(N__22382));
    LocalMux I__4696 (
            .O(N__22382),
            .I(\eeprom.n3480_adj_398 ));
    InMux I__4695 (
            .O(N__22379),
            .I(\eeprom.n3732 ));
    CascadeMux I__4694 (
            .O(N__22376),
            .I(N__22373));
    InMux I__4693 (
            .O(N__22373),
            .I(N__22370));
    LocalMux I__4692 (
            .O(N__22370),
            .I(N__22366));
    InMux I__4691 (
            .O(N__22369),
            .I(N__22363));
    Span4Mux_v I__4690 (
            .O(N__22366),
            .I(N__22360));
    LocalMux I__4689 (
            .O(N__22363),
            .I(\eeprom.n3412 ));
    Odrv4 I__4688 (
            .O(N__22360),
            .I(\eeprom.n3412 ));
    InMux I__4687 (
            .O(N__22355),
            .I(N__22352));
    LocalMux I__4686 (
            .O(N__22352),
            .I(N__22349));
    Span4Mux_h I__4685 (
            .O(N__22349),
            .I(N__22346));
    Odrv4 I__4684 (
            .O(N__22346),
            .I(\eeprom.n3479_adj_394 ));
    InMux I__4683 (
            .O(N__22343),
            .I(\eeprom.n3733 ));
    CascadeMux I__4682 (
            .O(N__22340),
            .I(N__22335));
    InMux I__4681 (
            .O(N__22339),
            .I(N__22332));
    InMux I__4680 (
            .O(N__22338),
            .I(N__22329));
    InMux I__4679 (
            .O(N__22335),
            .I(N__22326));
    LocalMux I__4678 (
            .O(N__22332),
            .I(N__22319));
    LocalMux I__4677 (
            .O(N__22329),
            .I(N__22319));
    LocalMux I__4676 (
            .O(N__22326),
            .I(N__22319));
    Odrv12 I__4675 (
            .O(N__22319),
            .I(\eeprom.n3411 ));
    CascadeMux I__4674 (
            .O(N__22316),
            .I(N__22313));
    InMux I__4673 (
            .O(N__22313),
            .I(N__22310));
    LocalMux I__4672 (
            .O(N__22310),
            .I(\eeprom.n3478_adj_393 ));
    InMux I__4671 (
            .O(N__22307),
            .I(bfn_14_18_0_));
    CascadeMux I__4670 (
            .O(N__22304),
            .I(N__22301));
    InMux I__4669 (
            .O(N__22301),
            .I(N__22298));
    LocalMux I__4668 (
            .O(N__22298),
            .I(N__22294));
    InMux I__4667 (
            .O(N__22297),
            .I(N__22291));
    Odrv4 I__4666 (
            .O(N__22294),
            .I(\eeprom.n3410 ));
    LocalMux I__4665 (
            .O(N__22291),
            .I(\eeprom.n3410 ));
    InMux I__4664 (
            .O(N__22286),
            .I(N__22283));
    LocalMux I__4663 (
            .O(N__22283),
            .I(N__22280));
    Odrv4 I__4662 (
            .O(N__22280),
            .I(\eeprom.n3477_adj_392 ));
    InMux I__4661 (
            .O(N__22277),
            .I(\eeprom.n3735 ));
    CascadeMux I__4660 (
            .O(N__22274),
            .I(N__22271));
    InMux I__4659 (
            .O(N__22271),
            .I(N__22266));
    InMux I__4658 (
            .O(N__22270),
            .I(N__22261));
    InMux I__4657 (
            .O(N__22269),
            .I(N__22261));
    LocalMux I__4656 (
            .O(N__22266),
            .I(N__22258));
    LocalMux I__4655 (
            .O(N__22261),
            .I(\eeprom.n3409 ));
    Odrv4 I__4654 (
            .O(N__22258),
            .I(\eeprom.n3409 ));
    InMux I__4653 (
            .O(N__22253),
            .I(N__22250));
    LocalMux I__4652 (
            .O(N__22250),
            .I(N__22247));
    Odrv4 I__4651 (
            .O(N__22247),
            .I(\eeprom.n3476_adj_391 ));
    InMux I__4650 (
            .O(N__22244),
            .I(\eeprom.n3736 ));
    CascadeMux I__4649 (
            .O(N__22241),
            .I(N__22237));
    InMux I__4648 (
            .O(N__22240),
            .I(N__22234));
    InMux I__4647 (
            .O(N__22237),
            .I(N__22231));
    LocalMux I__4646 (
            .O(N__22234),
            .I(N__22227));
    LocalMux I__4645 (
            .O(N__22231),
            .I(N__22224));
    InMux I__4644 (
            .O(N__22230),
            .I(N__22221));
    Odrv4 I__4643 (
            .O(N__22227),
            .I(\eeprom.n3408 ));
    Odrv12 I__4642 (
            .O(N__22224),
            .I(\eeprom.n3408 ));
    LocalMux I__4641 (
            .O(N__22221),
            .I(\eeprom.n3408 ));
    CascadeMux I__4640 (
            .O(N__22214),
            .I(N__22211));
    InMux I__4639 (
            .O(N__22211),
            .I(N__22208));
    LocalMux I__4638 (
            .O(N__22208),
            .I(N__22205));
    Odrv4 I__4637 (
            .O(N__22205),
            .I(\eeprom.n3475_adj_390 ));
    InMux I__4636 (
            .O(N__22202),
            .I(\eeprom.n3737 ));
    CascadeMux I__4635 (
            .O(N__22199),
            .I(N__22195));
    CascadeMux I__4634 (
            .O(N__22198),
            .I(N__22192));
    InMux I__4633 (
            .O(N__22195),
            .I(N__22189));
    InMux I__4632 (
            .O(N__22192),
            .I(N__22186));
    LocalMux I__4631 (
            .O(N__22189),
            .I(N__22183));
    LocalMux I__4630 (
            .O(N__22186),
            .I(\eeprom.n3407 ));
    Odrv4 I__4629 (
            .O(N__22183),
            .I(\eeprom.n3407 ));
    InMux I__4628 (
            .O(N__22178),
            .I(N__22175));
    LocalMux I__4627 (
            .O(N__22175),
            .I(N__22172));
    Odrv4 I__4626 (
            .O(N__22172),
            .I(\eeprom.n3474_adj_389 ));
    InMux I__4625 (
            .O(N__22169),
            .I(\eeprom.n3738 ));
    CascadeMux I__4624 (
            .O(N__22166),
            .I(N__22162));
    InMux I__4623 (
            .O(N__22165),
            .I(N__22159));
    InMux I__4622 (
            .O(N__22162),
            .I(N__22156));
    LocalMux I__4621 (
            .O(N__22159),
            .I(N__22150));
    LocalMux I__4620 (
            .O(N__22156),
            .I(N__22150));
    InMux I__4619 (
            .O(N__22155),
            .I(N__22147));
    Odrv12 I__4618 (
            .O(N__22150),
            .I(\eeprom.n3406 ));
    LocalMux I__4617 (
            .O(N__22147),
            .I(\eeprom.n3406 ));
    CascadeMux I__4616 (
            .O(N__22142),
            .I(N__22139));
    InMux I__4615 (
            .O(N__22139),
            .I(N__22136));
    LocalMux I__4614 (
            .O(N__22136),
            .I(N__22133));
    Odrv12 I__4613 (
            .O(N__22133),
            .I(\eeprom.n3473_adj_388 ));
    InMux I__4612 (
            .O(N__22130),
            .I(\eeprom.n3739 ));
    InMux I__4611 (
            .O(N__22127),
            .I(N__22122));
    InMux I__4610 (
            .O(N__22126),
            .I(N__22119));
    CascadeMux I__4609 (
            .O(N__22125),
            .I(N__22116));
    LocalMux I__4608 (
            .O(N__22122),
            .I(N__22113));
    LocalMux I__4607 (
            .O(N__22119),
            .I(N__22110));
    InMux I__4606 (
            .O(N__22116),
            .I(N__22107));
    Odrv12 I__4605 (
            .O(N__22113),
            .I(\eeprom.n2907 ));
    Odrv4 I__4604 (
            .O(N__22110),
            .I(\eeprom.n2907 ));
    LocalMux I__4603 (
            .O(N__22107),
            .I(\eeprom.n2907 ));
    CascadeMux I__4602 (
            .O(N__22100),
            .I(N__22097));
    InMux I__4601 (
            .O(N__22097),
            .I(N__22094));
    LocalMux I__4600 (
            .O(N__22094),
            .I(N__22091));
    Span4Mux_v I__4599 (
            .O(N__22091),
            .I(N__22088));
    Odrv4 I__4598 (
            .O(N__22088),
            .I(\eeprom.n2974 ));
    InMux I__4597 (
            .O(N__22085),
            .I(N__22082));
    LocalMux I__4596 (
            .O(N__22082),
            .I(N__22077));
    CascadeMux I__4595 (
            .O(N__22081),
            .I(N__22074));
    InMux I__4594 (
            .O(N__22080),
            .I(N__22071));
    Span4Mux_v I__4593 (
            .O(N__22077),
            .I(N__22068));
    InMux I__4592 (
            .O(N__22074),
            .I(N__22065));
    LocalMux I__4591 (
            .O(N__22071),
            .I(N__22062));
    Odrv4 I__4590 (
            .O(N__22068),
            .I(\eeprom.n2914 ));
    LocalMux I__4589 (
            .O(N__22065),
            .I(\eeprom.n2914 ));
    Odrv12 I__4588 (
            .O(N__22062),
            .I(\eeprom.n2914 ));
    InMux I__4587 (
            .O(N__22055),
            .I(N__22052));
    LocalMux I__4586 (
            .O(N__22052),
            .I(N__22049));
    Span4Mux_h I__4585 (
            .O(N__22049),
            .I(N__22046));
    Odrv4 I__4584 (
            .O(N__22046),
            .I(\eeprom.n2981 ));
    CascadeMux I__4583 (
            .O(N__22043),
            .I(N__22039));
    InMux I__4582 (
            .O(N__22042),
            .I(N__22035));
    InMux I__4581 (
            .O(N__22039),
            .I(N__22030));
    InMux I__4580 (
            .O(N__22038),
            .I(N__22030));
    LocalMux I__4579 (
            .O(N__22035),
            .I(\eeprom.n3101 ));
    LocalMux I__4578 (
            .O(N__22030),
            .I(\eeprom.n3101 ));
    InMux I__4577 (
            .O(N__22025),
            .I(bfn_14_17_0_));
    InMux I__4576 (
            .O(N__22022),
            .I(\eeprom.n3727 ));
    InMux I__4575 (
            .O(N__22019),
            .I(\eeprom.n3728 ));
    InMux I__4574 (
            .O(N__22016),
            .I(\eeprom.n3729 ));
    CascadeMux I__4573 (
            .O(N__22013),
            .I(N__22009));
    CascadeMux I__4572 (
            .O(N__22012),
            .I(N__22006));
    InMux I__4571 (
            .O(N__22009),
            .I(N__22003));
    InMux I__4570 (
            .O(N__22006),
            .I(N__21999));
    LocalMux I__4569 (
            .O(N__22003),
            .I(N__21996));
    InMux I__4568 (
            .O(N__22002),
            .I(N__21993));
    LocalMux I__4567 (
            .O(N__21999),
            .I(\eeprom.n3415 ));
    Odrv4 I__4566 (
            .O(N__21996),
            .I(\eeprom.n3415 ));
    LocalMux I__4565 (
            .O(N__21993),
            .I(\eeprom.n3415 ));
    InMux I__4564 (
            .O(N__21986),
            .I(N__21983));
    LocalMux I__4563 (
            .O(N__21983),
            .I(\eeprom.n3482_adj_401 ));
    InMux I__4562 (
            .O(N__21980),
            .I(\eeprom.n3730 ));
    InMux I__4561 (
            .O(N__21977),
            .I(N__21973));
    InMux I__4560 (
            .O(N__21976),
            .I(N__21970));
    LocalMux I__4559 (
            .O(N__21973),
            .I(N__21967));
    LocalMux I__4558 (
            .O(N__21970),
            .I(\eeprom.n3414 ));
    Odrv4 I__4557 (
            .O(N__21967),
            .I(\eeprom.n3414 ));
    InMux I__4556 (
            .O(N__21962),
            .I(N__21959));
    LocalMux I__4555 (
            .O(N__21959),
            .I(\eeprom.n3481_adj_399 ));
    InMux I__4554 (
            .O(N__21956),
            .I(\eeprom.n3731 ));
    InMux I__4553 (
            .O(N__21953),
            .I(N__21948));
    InMux I__4552 (
            .O(N__21952),
            .I(N__21945));
    InMux I__4551 (
            .O(N__21951),
            .I(N__21942));
    LocalMux I__4550 (
            .O(N__21948),
            .I(N__21937));
    LocalMux I__4549 (
            .O(N__21945),
            .I(N__21937));
    LocalMux I__4548 (
            .O(N__21942),
            .I(\eeprom.n3104 ));
    Odrv4 I__4547 (
            .O(N__21937),
            .I(\eeprom.n3104 ));
    InMux I__4546 (
            .O(N__21932),
            .I(N__21929));
    LocalMux I__4545 (
            .O(N__21929),
            .I(\eeprom.n3170 ));
    InMux I__4544 (
            .O(N__21926),
            .I(N__21922));
    InMux I__4543 (
            .O(N__21925),
            .I(N__21919));
    LocalMux I__4542 (
            .O(N__21922),
            .I(N__21916));
    LocalMux I__4541 (
            .O(N__21919),
            .I(N__21913));
    Span4Mux_h I__4540 (
            .O(N__21916),
            .I(N__21909));
    Span4Mux_h I__4539 (
            .O(N__21913),
            .I(N__21906));
    InMux I__4538 (
            .O(N__21912),
            .I(N__21903));
    Odrv4 I__4537 (
            .O(N__21909),
            .I(\eeprom.n3202 ));
    Odrv4 I__4536 (
            .O(N__21906),
            .I(\eeprom.n3202 ));
    LocalMux I__4535 (
            .O(N__21903),
            .I(\eeprom.n3202 ));
    InMux I__4534 (
            .O(N__21896),
            .I(N__21893));
    LocalMux I__4533 (
            .O(N__21893),
            .I(\eeprom.n3168 ));
    InMux I__4532 (
            .O(N__21890),
            .I(N__21886));
    InMux I__4531 (
            .O(N__21889),
            .I(N__21883));
    LocalMux I__4530 (
            .O(N__21886),
            .I(N__21880));
    LocalMux I__4529 (
            .O(N__21883),
            .I(N__21877));
    Span4Mux_h I__4528 (
            .O(N__21880),
            .I(N__21873));
    Span4Mux_h I__4527 (
            .O(N__21877),
            .I(N__21870));
    InMux I__4526 (
            .O(N__21876),
            .I(N__21867));
    Odrv4 I__4525 (
            .O(N__21873),
            .I(\eeprom.n3200 ));
    Odrv4 I__4524 (
            .O(N__21870),
            .I(\eeprom.n3200 ));
    LocalMux I__4523 (
            .O(N__21867),
            .I(\eeprom.n3200 ));
    InMux I__4522 (
            .O(N__21860),
            .I(N__21857));
    LocalMux I__4521 (
            .O(N__21857),
            .I(N__21854));
    Span4Mux_h I__4520 (
            .O(N__21854),
            .I(N__21851));
    Odrv4 I__4519 (
            .O(N__21851),
            .I(\eeprom.n2983 ));
    CascadeMux I__4518 (
            .O(N__21848),
            .I(N__21845));
    InMux I__4517 (
            .O(N__21845),
            .I(N__21841));
    CascadeMux I__4516 (
            .O(N__21844),
            .I(N__21838));
    LocalMux I__4515 (
            .O(N__21841),
            .I(N__21835));
    InMux I__4514 (
            .O(N__21838),
            .I(N__21832));
    Span4Mux_h I__4513 (
            .O(N__21835),
            .I(N__21826));
    LocalMux I__4512 (
            .O(N__21832),
            .I(N__21826));
    InMux I__4511 (
            .O(N__21831),
            .I(N__21823));
    Odrv4 I__4510 (
            .O(N__21826),
            .I(\eeprom.n2916 ));
    LocalMux I__4509 (
            .O(N__21823),
            .I(\eeprom.n2916 ));
    InMux I__4508 (
            .O(N__21818),
            .I(N__21814));
    InMux I__4507 (
            .O(N__21817),
            .I(N__21811));
    LocalMux I__4506 (
            .O(N__21814),
            .I(N__21808));
    LocalMux I__4505 (
            .O(N__21811),
            .I(\eeprom.n3106 ));
    Odrv4 I__4504 (
            .O(N__21808),
            .I(\eeprom.n3106 ));
    InMux I__4503 (
            .O(N__21803),
            .I(N__21800));
    LocalMux I__4502 (
            .O(N__21800),
            .I(\eeprom.n3173 ));
    CascadeMux I__4501 (
            .O(N__21797),
            .I(\eeprom.n3106_cascade_ ));
    CascadeMux I__4500 (
            .O(N__21794),
            .I(N__21785));
    InMux I__4499 (
            .O(N__21793),
            .I(N__21781));
    CascadeMux I__4498 (
            .O(N__21792),
            .I(N__21778));
    CascadeMux I__4497 (
            .O(N__21791),
            .I(N__21773));
    InMux I__4496 (
            .O(N__21790),
            .I(N__21766));
    InMux I__4495 (
            .O(N__21789),
            .I(N__21766));
    InMux I__4494 (
            .O(N__21788),
            .I(N__21758));
    InMux I__4493 (
            .O(N__21785),
            .I(N__21753));
    InMux I__4492 (
            .O(N__21784),
            .I(N__21753));
    LocalMux I__4491 (
            .O(N__21781),
            .I(N__21750));
    InMux I__4490 (
            .O(N__21778),
            .I(N__21747));
    CascadeMux I__4489 (
            .O(N__21777),
            .I(N__21743));
    InMux I__4488 (
            .O(N__21776),
            .I(N__21738));
    InMux I__4487 (
            .O(N__21773),
            .I(N__21731));
    InMux I__4486 (
            .O(N__21772),
            .I(N__21731));
    InMux I__4485 (
            .O(N__21771),
            .I(N__21731));
    LocalMux I__4484 (
            .O(N__21766),
            .I(N__21728));
    InMux I__4483 (
            .O(N__21765),
            .I(N__21721));
    InMux I__4482 (
            .O(N__21764),
            .I(N__21721));
    InMux I__4481 (
            .O(N__21763),
            .I(N__21721));
    InMux I__4480 (
            .O(N__21762),
            .I(N__21716));
    InMux I__4479 (
            .O(N__21761),
            .I(N__21716));
    LocalMux I__4478 (
            .O(N__21758),
            .I(N__21711));
    LocalMux I__4477 (
            .O(N__21753),
            .I(N__21711));
    Span4Mux_h I__4476 (
            .O(N__21750),
            .I(N__21706));
    LocalMux I__4475 (
            .O(N__21747),
            .I(N__21706));
    InMux I__4474 (
            .O(N__21746),
            .I(N__21697));
    InMux I__4473 (
            .O(N__21743),
            .I(N__21697));
    InMux I__4472 (
            .O(N__21742),
            .I(N__21697));
    InMux I__4471 (
            .O(N__21741),
            .I(N__21697));
    LocalMux I__4470 (
            .O(N__21738),
            .I(\eeprom.n3133 ));
    LocalMux I__4469 (
            .O(N__21731),
            .I(\eeprom.n3133 ));
    Odrv4 I__4468 (
            .O(N__21728),
            .I(\eeprom.n3133 ));
    LocalMux I__4467 (
            .O(N__21721),
            .I(\eeprom.n3133 ));
    LocalMux I__4466 (
            .O(N__21716),
            .I(\eeprom.n3133 ));
    Odrv4 I__4465 (
            .O(N__21711),
            .I(\eeprom.n3133 ));
    Odrv4 I__4464 (
            .O(N__21706),
            .I(\eeprom.n3133 ));
    LocalMux I__4463 (
            .O(N__21697),
            .I(\eeprom.n3133 ));
    InMux I__4462 (
            .O(N__21680),
            .I(N__21677));
    LocalMux I__4461 (
            .O(N__21677),
            .I(N__21673));
    InMux I__4460 (
            .O(N__21676),
            .I(N__21670));
    Span4Mux_v I__4459 (
            .O(N__21673),
            .I(N__21667));
    LocalMux I__4458 (
            .O(N__21670),
            .I(N__21664));
    Span4Mux_h I__4457 (
            .O(N__21667),
            .I(N__21661));
    Span4Mux_h I__4456 (
            .O(N__21664),
            .I(N__21658));
    Odrv4 I__4455 (
            .O(N__21661),
            .I(\eeprom.n3205 ));
    Odrv4 I__4454 (
            .O(N__21658),
            .I(\eeprom.n3205 ));
    CascadeMux I__4453 (
            .O(N__21653),
            .I(\eeprom.n3205_cascade_ ));
    InMux I__4452 (
            .O(N__21650),
            .I(N__21647));
    LocalMux I__4451 (
            .O(N__21647),
            .I(N__21644));
    Span4Mux_v I__4450 (
            .O(N__21644),
            .I(N__21640));
    InMux I__4449 (
            .O(N__21643),
            .I(N__21637));
    Odrv4 I__4448 (
            .O(N__21640),
            .I(\eeprom.n3199 ));
    LocalMux I__4447 (
            .O(N__21637),
            .I(\eeprom.n3199 ));
    InMux I__4446 (
            .O(N__21632),
            .I(N__21629));
    LocalMux I__4445 (
            .O(N__21629),
            .I(N__21626));
    Span4Mux_h I__4444 (
            .O(N__21626),
            .I(N__21623));
    Span4Mux_v I__4443 (
            .O(N__21623),
            .I(N__21620));
    Odrv4 I__4442 (
            .O(N__21620),
            .I(\eeprom.n16_adj_479 ));
    CascadeMux I__4441 (
            .O(N__21617),
            .I(N__21612));
    CascadeMux I__4440 (
            .O(N__21616),
            .I(N__21609));
    CascadeMux I__4439 (
            .O(N__21615),
            .I(N__21606));
    InMux I__4438 (
            .O(N__21612),
            .I(N__21603));
    InMux I__4437 (
            .O(N__21609),
            .I(N__21598));
    InMux I__4436 (
            .O(N__21606),
            .I(N__21598));
    LocalMux I__4435 (
            .O(N__21603),
            .I(\eeprom.n3115 ));
    LocalMux I__4434 (
            .O(N__21598),
            .I(\eeprom.n3115 ));
    InMux I__4433 (
            .O(N__21593),
            .I(N__21590));
    LocalMux I__4432 (
            .O(N__21590),
            .I(N__21587));
    Odrv4 I__4431 (
            .O(N__21587),
            .I(\eeprom.n3169 ));
    InMux I__4430 (
            .O(N__21584),
            .I(N__21581));
    LocalMux I__4429 (
            .O(N__21581),
            .I(N__21577));
    InMux I__4428 (
            .O(N__21580),
            .I(N__21574));
    Span4Mux_h I__4427 (
            .O(N__21577),
            .I(N__21571));
    LocalMux I__4426 (
            .O(N__21574),
            .I(N__21568));
    Odrv4 I__4425 (
            .O(N__21571),
            .I(\eeprom.n3201 ));
    Odrv12 I__4424 (
            .O(N__21568),
            .I(\eeprom.n3201 ));
    InMux I__4423 (
            .O(N__21563),
            .I(N__21560));
    LocalMux I__4422 (
            .O(N__21560),
            .I(N__21556));
    InMux I__4421 (
            .O(N__21559),
            .I(N__21553));
    Span4Mux_h I__4420 (
            .O(N__21556),
            .I(N__21549));
    LocalMux I__4419 (
            .O(N__21553),
            .I(N__21546));
    InMux I__4418 (
            .O(N__21552),
            .I(N__21543));
    Odrv4 I__4417 (
            .O(N__21549),
            .I(\eeprom.n3207 ));
    Odrv12 I__4416 (
            .O(N__21546),
            .I(\eeprom.n3207 ));
    LocalMux I__4415 (
            .O(N__21543),
            .I(\eeprom.n3207 ));
    CascadeMux I__4414 (
            .O(N__21536),
            .I(\eeprom.n3201_cascade_ ));
    InMux I__4413 (
            .O(N__21533),
            .I(N__21530));
    LocalMux I__4412 (
            .O(N__21530),
            .I(N__21527));
    Span4Mux_h I__4411 (
            .O(N__21527),
            .I(N__21524));
    Odrv4 I__4410 (
            .O(N__21524),
            .I(\eeprom.n24_adj_481 ));
    InMux I__4409 (
            .O(N__21521),
            .I(N__21518));
    LocalMux I__4408 (
            .O(N__21518),
            .I(N__21514));
    CascadeMux I__4407 (
            .O(N__21517),
            .I(N__21511));
    Span4Mux_v I__4406 (
            .O(N__21514),
            .I(N__21507));
    InMux I__4405 (
            .O(N__21511),
            .I(N__21504));
    InMux I__4404 (
            .O(N__21510),
            .I(N__21501));
    Odrv4 I__4403 (
            .O(N__21507),
            .I(\eeprom.n3114 ));
    LocalMux I__4402 (
            .O(N__21504),
            .I(\eeprom.n3114 ));
    LocalMux I__4401 (
            .O(N__21501),
            .I(\eeprom.n3114 ));
    InMux I__4400 (
            .O(N__21494),
            .I(N__21490));
    InMux I__4399 (
            .O(N__21493),
            .I(N__21487));
    LocalMux I__4398 (
            .O(N__21490),
            .I(N__21482));
    LocalMux I__4397 (
            .O(N__21487),
            .I(N__21482));
    Span4Mux_h I__4396 (
            .O(N__21482),
            .I(N__21478));
    InMux I__4395 (
            .O(N__21481),
            .I(N__21475));
    Odrv4 I__4394 (
            .O(N__21478),
            .I(\eeprom.n2905 ));
    LocalMux I__4393 (
            .O(N__21475),
            .I(\eeprom.n2905 ));
    CascadeMux I__4392 (
            .O(N__21470),
            .I(N__21467));
    InMux I__4391 (
            .O(N__21467),
            .I(N__21464));
    LocalMux I__4390 (
            .O(N__21464),
            .I(N__21461));
    Odrv4 I__4389 (
            .O(N__21461),
            .I(\eeprom.n2972 ));
    InMux I__4388 (
            .O(N__21458),
            .I(N__21455));
    LocalMux I__4387 (
            .O(N__21455),
            .I(N__21450));
    CascadeMux I__4386 (
            .O(N__21454),
            .I(N__21447));
    CascadeMux I__4385 (
            .O(N__21453),
            .I(N__21444));
    Span4Mux_v I__4384 (
            .O(N__21450),
            .I(N__21441));
    InMux I__4383 (
            .O(N__21447),
            .I(N__21438));
    InMux I__4382 (
            .O(N__21444),
            .I(N__21435));
    Odrv4 I__4381 (
            .O(N__21441),
            .I(\eeprom.n3118 ));
    LocalMux I__4380 (
            .O(N__21438),
            .I(\eeprom.n3118 ));
    LocalMux I__4379 (
            .O(N__21435),
            .I(\eeprom.n3118 ));
    InMux I__4378 (
            .O(N__21428),
            .I(N__21424));
    InMux I__4377 (
            .O(N__21427),
            .I(N__21421));
    LocalMux I__4376 (
            .O(N__21424),
            .I(\eeprom.n3102 ));
    LocalMux I__4375 (
            .O(N__21421),
            .I(\eeprom.n3102 ));
    CascadeMux I__4374 (
            .O(N__21416),
            .I(\eeprom.n3102_cascade_ ));
    InMux I__4373 (
            .O(N__21413),
            .I(N__21410));
    LocalMux I__4372 (
            .O(N__21410),
            .I(N__21407));
    Odrv4 I__4371 (
            .O(N__21407),
            .I(\eeprom.n22_adj_465 ));
    InMux I__4370 (
            .O(N__21404),
            .I(N__21401));
    LocalMux I__4369 (
            .O(N__21401),
            .I(\eeprom.n3600_adj_449 ));
    InMux I__4368 (
            .O(N__21398),
            .I(N__21395));
    LocalMux I__4367 (
            .O(N__21395),
            .I(\eeprom.n4581 ));
    CascadeMux I__4366 (
            .O(N__21392),
            .I(N__21387));
    InMux I__4365 (
            .O(N__21391),
            .I(N__21384));
    InMux I__4364 (
            .O(N__21390),
            .I(N__21381));
    InMux I__4363 (
            .O(N__21387),
            .I(N__21378));
    LocalMux I__4362 (
            .O(N__21384),
            .I(\eeprom.n3117 ));
    LocalMux I__4361 (
            .O(N__21381),
            .I(\eeprom.n3117 ));
    LocalMux I__4360 (
            .O(N__21378),
            .I(\eeprom.n3117 ));
    InMux I__4359 (
            .O(N__21371),
            .I(N__21367));
    InMux I__4358 (
            .O(N__21370),
            .I(N__21364));
    LocalMux I__4357 (
            .O(N__21367),
            .I(N__21361));
    LocalMux I__4356 (
            .O(N__21364),
            .I(\eeprom.n3108 ));
    Odrv4 I__4355 (
            .O(N__21361),
            .I(\eeprom.n3108 ));
    InMux I__4354 (
            .O(N__21356),
            .I(N__21353));
    LocalMux I__4353 (
            .O(N__21353),
            .I(N__21350));
    Odrv4 I__4352 (
            .O(N__21350),
            .I(\eeprom.n3175 ));
    CascadeMux I__4351 (
            .O(N__21347),
            .I(\eeprom.n3108_cascade_ ));
    CascadeMux I__4350 (
            .O(N__21344),
            .I(N__21341));
    InMux I__4349 (
            .O(N__21341),
            .I(N__21337));
    InMux I__4348 (
            .O(N__21340),
            .I(N__21334));
    LocalMux I__4347 (
            .O(N__21337),
            .I(N__21331));
    LocalMux I__4346 (
            .O(N__21334),
            .I(\eeprom.n3105 ));
    Odrv4 I__4345 (
            .O(N__21331),
            .I(\eeprom.n3105 ));
    InMux I__4344 (
            .O(N__21326),
            .I(N__21323));
    LocalMux I__4343 (
            .O(N__21323),
            .I(N__21320));
    Span4Mux_h I__4342 (
            .O(N__21320),
            .I(N__21317));
    Odrv4 I__4341 (
            .O(N__21317),
            .I(\eeprom.n3172 ));
    CascadeMux I__4340 (
            .O(N__21314),
            .I(\eeprom.n3105_cascade_ ));
    InMux I__4339 (
            .O(N__21311),
            .I(N__21307));
    InMux I__4338 (
            .O(N__21310),
            .I(N__21303));
    LocalMux I__4337 (
            .O(N__21307),
            .I(N__21300));
    InMux I__4336 (
            .O(N__21306),
            .I(N__21297));
    LocalMux I__4335 (
            .O(N__21303),
            .I(N__21294));
    Span4Mux_h I__4334 (
            .O(N__21300),
            .I(N__21291));
    LocalMux I__4333 (
            .O(N__21297),
            .I(N__21288));
    Span4Mux_h I__4332 (
            .O(N__21294),
            .I(N__21285));
    Odrv4 I__4331 (
            .O(N__21291),
            .I(\eeprom.n3204 ));
    Odrv12 I__4330 (
            .O(N__21288),
            .I(\eeprom.n3204 ));
    Odrv4 I__4329 (
            .O(N__21285),
            .I(\eeprom.n3204 ));
    CascadeMux I__4328 (
            .O(N__21278),
            .I(N__21275));
    InMux I__4327 (
            .O(N__21275),
            .I(N__21272));
    LocalMux I__4326 (
            .O(N__21272),
            .I(\eeprom.n3179 ));
    InMux I__4325 (
            .O(N__21269),
            .I(N__21266));
    LocalMux I__4324 (
            .O(N__21266),
            .I(N__21261));
    InMux I__4323 (
            .O(N__21265),
            .I(N__21258));
    CascadeMux I__4322 (
            .O(N__21264),
            .I(N__21255));
    Span4Mux_v I__4321 (
            .O(N__21261),
            .I(N__21252));
    LocalMux I__4320 (
            .O(N__21258),
            .I(N__21249));
    InMux I__4319 (
            .O(N__21255),
            .I(N__21246));
    Span4Mux_h I__4318 (
            .O(N__21252),
            .I(N__21241));
    Span4Mux_v I__4317 (
            .O(N__21249),
            .I(N__21241));
    LocalMux I__4316 (
            .O(N__21246),
            .I(N__21238));
    Odrv4 I__4315 (
            .O(N__21241),
            .I(\eeprom.n3211 ));
    Odrv12 I__4314 (
            .O(N__21238),
            .I(\eeprom.n3211 ));
    InMux I__4313 (
            .O(N__21233),
            .I(N__21230));
    LocalMux I__4312 (
            .O(N__21230),
            .I(\eeprom.n31_adj_496 ));
    InMux I__4311 (
            .O(N__21227),
            .I(N__21224));
    LocalMux I__4310 (
            .O(N__21224),
            .I(\eeprom.n29_adj_497 ));
    CascadeMux I__4309 (
            .O(N__21221),
            .I(\eeprom.n30_adj_495_cascade_ ));
    InMux I__4308 (
            .O(N__21218),
            .I(N__21215));
    LocalMux I__4307 (
            .O(N__21215),
            .I(N__21212));
    Odrv4 I__4306 (
            .O(N__21212),
            .I(\eeprom.n32_adj_494 ));
    CascadeMux I__4305 (
            .O(N__21209),
            .I(\eeprom.n3606_adj_446_cascade_ ));
    CascadeMux I__4304 (
            .O(N__21206),
            .I(\eeprom.n4451_cascade_ ));
    InMux I__4303 (
            .O(N__21203),
            .I(N__21200));
    LocalMux I__4302 (
            .O(N__21200),
            .I(\eeprom.n4453 ));
    CascadeMux I__4301 (
            .O(N__21197),
            .I(\eeprom.n3599_adj_450_cascade_ ));
    InMux I__4300 (
            .O(N__21194),
            .I(N__21191));
    LocalMux I__4299 (
            .O(N__21191),
            .I(N__21188));
    Odrv4 I__4298 (
            .O(N__21188),
            .I(\eeprom.n4429 ));
    InMux I__4297 (
            .O(N__21185),
            .I(N__21182));
    LocalMux I__4296 (
            .O(N__21182),
            .I(N__21179));
    Span4Mux_v I__4295 (
            .O(N__21179),
            .I(N__21176));
    Sp12to4 I__4294 (
            .O(N__21176),
            .I(N__21173));
    Odrv12 I__4293 (
            .O(N__21173),
            .I(\eeprom.n29 ));
    CascadeMux I__4292 (
            .O(N__21170),
            .I(\eeprom.n28_adj_493_cascade_ ));
    CascadeMux I__4291 (
            .O(N__21167),
            .I(\eeprom.n18_adj_488_cascade_ ));
    InMux I__4290 (
            .O(N__21164),
            .I(N__21161));
    LocalMux I__4289 (
            .O(N__21161),
            .I(N__21158));
    Odrv4 I__4288 (
            .O(N__21158),
            .I(\eeprom.n29_adj_491 ));
    InMux I__4287 (
            .O(N__21155),
            .I(N__21152));
    LocalMux I__4286 (
            .O(N__21152),
            .I(\eeprom.n28_adj_490 ));
    CascadeMux I__4285 (
            .O(N__21149),
            .I(\eeprom.n30_adj_489_cascade_ ));
    InMux I__4284 (
            .O(N__21146),
            .I(N__21143));
    LocalMux I__4283 (
            .O(N__21143),
            .I(N__21140));
    Odrv4 I__4282 (
            .O(N__21140),
            .I(\eeprom.n27_adj_492 ));
    CascadeMux I__4281 (
            .O(N__21137),
            .I(\eeprom.n3430_cascade_ ));
    InMux I__4280 (
            .O(N__21134),
            .I(N__21131));
    LocalMux I__4279 (
            .O(N__21131),
            .I(\eeprom.n3609_adj_445 ));
    CascadeMux I__4278 (
            .O(N__21128),
            .I(\eeprom.n3508_cascade_ ));
    InMux I__4277 (
            .O(N__21125),
            .I(\eeprom.n3685 ));
    InMux I__4276 (
            .O(N__21122),
            .I(N__21119));
    LocalMux I__4275 (
            .O(N__21119),
            .I(N__21116));
    Odrv4 I__4274 (
            .O(N__21116),
            .I(\eeprom.n2971 ));
    CascadeMux I__4273 (
            .O(N__21113),
            .I(N__21110));
    InMux I__4272 (
            .O(N__21110),
            .I(N__21107));
    LocalMux I__4271 (
            .O(N__21107),
            .I(N__21103));
    InMux I__4270 (
            .O(N__21106),
            .I(N__21100));
    Span4Mux_v I__4269 (
            .O(N__21103),
            .I(N__21095));
    LocalMux I__4268 (
            .O(N__21100),
            .I(N__21095));
    Span4Mux_h I__4267 (
            .O(N__21095),
            .I(N__21092));
    Odrv4 I__4266 (
            .O(N__21092),
            .I(\eeprom.n2904 ));
    InMux I__4265 (
            .O(N__21089),
            .I(N__21086));
    LocalMux I__4264 (
            .O(N__21086),
            .I(N__21083));
    Odrv4 I__4263 (
            .O(N__21083),
            .I(\eeprom.n2977 ));
    CascadeMux I__4262 (
            .O(N__21080),
            .I(N__21077));
    InMux I__4261 (
            .O(N__21077),
            .I(N__21073));
    InMux I__4260 (
            .O(N__21076),
            .I(N__21069));
    LocalMux I__4259 (
            .O(N__21073),
            .I(N__21066));
    InMux I__4258 (
            .O(N__21072),
            .I(N__21063));
    LocalMux I__4257 (
            .O(N__21069),
            .I(\eeprom.n2910 ));
    Odrv4 I__4256 (
            .O(N__21066),
            .I(\eeprom.n2910 ));
    LocalMux I__4255 (
            .O(N__21063),
            .I(\eeprom.n2910 ));
    CascadeMux I__4254 (
            .O(N__21056),
            .I(\eeprom.n3497_cascade_ ));
    CascadeMux I__4253 (
            .O(N__21053),
            .I(N__21050));
    InMux I__4252 (
            .O(N__21050),
            .I(N__21047));
    LocalMux I__4251 (
            .O(N__21047),
            .I(N__21044));
    Span4Mux_v I__4250 (
            .O(N__21044),
            .I(N__21041));
    Odrv4 I__4249 (
            .O(N__21041),
            .I(\eeprom.n3176 ));
    InMux I__4248 (
            .O(N__21038),
            .I(\eeprom.n3676 ));
    InMux I__4247 (
            .O(N__21035),
            .I(\eeprom.n3677 ));
    InMux I__4246 (
            .O(N__21032),
            .I(N__21029));
    LocalMux I__4245 (
            .O(N__21029),
            .I(N__21026));
    Odrv12 I__4244 (
            .O(N__21026),
            .I(\eeprom.n3174 ));
    InMux I__4243 (
            .O(N__21023),
            .I(\eeprom.n3678 ));
    InMux I__4242 (
            .O(N__21020),
            .I(\eeprom.n3679 ));
    InMux I__4241 (
            .O(N__21017),
            .I(\eeprom.n3680 ));
    InMux I__4240 (
            .O(N__21014),
            .I(N__21011));
    LocalMux I__4239 (
            .O(N__21011),
            .I(N__21008));
    Odrv12 I__4238 (
            .O(N__21008),
            .I(\eeprom.n3171 ));
    InMux I__4237 (
            .O(N__21005),
            .I(\eeprom.n3681 ));
    InMux I__4236 (
            .O(N__21002),
            .I(bfn_12_24_0_));
    InMux I__4235 (
            .O(N__20999),
            .I(\eeprom.n3683 ));
    InMux I__4234 (
            .O(N__20996),
            .I(\eeprom.n3684 ));
    CascadeMux I__4233 (
            .O(N__20993),
            .I(N__20990));
    InMux I__4232 (
            .O(N__20990),
            .I(N__20987));
    LocalMux I__4231 (
            .O(N__20987),
            .I(N__20984));
    Odrv4 I__4230 (
            .O(N__20984),
            .I(\eeprom.n3184 ));
    InMux I__4229 (
            .O(N__20981),
            .I(\eeprom.n3668 ));
    CascadeMux I__4228 (
            .O(N__20978),
            .I(N__20975));
    InMux I__4227 (
            .O(N__20975),
            .I(N__20971));
    InMux I__4226 (
            .O(N__20974),
            .I(N__20968));
    LocalMux I__4225 (
            .O(N__20971),
            .I(N__20965));
    LocalMux I__4224 (
            .O(N__20968),
            .I(\eeprom.n3116 ));
    Odrv4 I__4223 (
            .O(N__20965),
            .I(\eeprom.n3116 ));
    InMux I__4222 (
            .O(N__20960),
            .I(N__20957));
    LocalMux I__4221 (
            .O(N__20957),
            .I(N__20954));
    Odrv4 I__4220 (
            .O(N__20954),
            .I(\eeprom.n3183 ));
    InMux I__4219 (
            .O(N__20951),
            .I(\eeprom.n3669 ));
    InMux I__4218 (
            .O(N__20948),
            .I(N__20945));
    LocalMux I__4217 (
            .O(N__20945),
            .I(\eeprom.n3182 ));
    InMux I__4216 (
            .O(N__20942),
            .I(\eeprom.n3670 ));
    CascadeMux I__4215 (
            .O(N__20939),
            .I(N__20936));
    InMux I__4214 (
            .O(N__20936),
            .I(N__20933));
    LocalMux I__4213 (
            .O(N__20933),
            .I(N__20930));
    Odrv4 I__4212 (
            .O(N__20930),
            .I(\eeprom.n3181 ));
    InMux I__4211 (
            .O(N__20927),
            .I(\eeprom.n3671 ));
    CascadeMux I__4210 (
            .O(N__20924),
            .I(N__20921));
    InMux I__4209 (
            .O(N__20921),
            .I(N__20918));
    LocalMux I__4208 (
            .O(N__20918),
            .I(N__20914));
    InMux I__4207 (
            .O(N__20917),
            .I(N__20911));
    Odrv4 I__4206 (
            .O(N__20914),
            .I(\eeprom.n3113 ));
    LocalMux I__4205 (
            .O(N__20911),
            .I(\eeprom.n3113 ));
    InMux I__4204 (
            .O(N__20906),
            .I(N__20903));
    LocalMux I__4203 (
            .O(N__20903),
            .I(N__20900));
    Span4Mux_h I__4202 (
            .O(N__20900),
            .I(N__20897));
    Odrv4 I__4201 (
            .O(N__20897),
            .I(\eeprom.n3180 ));
    InMux I__4200 (
            .O(N__20894),
            .I(\eeprom.n3672 ));
    InMux I__4199 (
            .O(N__20891),
            .I(\eeprom.n3673 ));
    InMux I__4198 (
            .O(N__20888),
            .I(N__20885));
    LocalMux I__4197 (
            .O(N__20885),
            .I(N__20882));
    Span4Mux_h I__4196 (
            .O(N__20882),
            .I(N__20879));
    Odrv4 I__4195 (
            .O(N__20879),
            .I(\eeprom.n3178 ));
    InMux I__4194 (
            .O(N__20876),
            .I(bfn_12_23_0_));
    CascadeMux I__4193 (
            .O(N__20873),
            .I(N__20870));
    InMux I__4192 (
            .O(N__20870),
            .I(N__20867));
    LocalMux I__4191 (
            .O(N__20867),
            .I(N__20864));
    Span4Mux_h I__4190 (
            .O(N__20864),
            .I(N__20861));
    Odrv4 I__4189 (
            .O(N__20861),
            .I(\eeprom.n3177 ));
    InMux I__4188 (
            .O(N__20858),
            .I(\eeprom.n3675 ));
    CascadeMux I__4187 (
            .O(N__20855),
            .I(\eeprom.n18_adj_432_cascade_ ));
    CascadeMux I__4186 (
            .O(N__20852),
            .I(\eeprom.n26_adj_466_cascade_ ));
    CascadeMux I__4185 (
            .O(N__20849),
            .I(\eeprom.n4711_cascade_ ));
    InMux I__4184 (
            .O(N__20846),
            .I(N__20843));
    LocalMux I__4183 (
            .O(N__20843),
            .I(\eeprom.n4715 ));
    CascadeMux I__4182 (
            .O(N__20840),
            .I(N__20837));
    InMux I__4181 (
            .O(N__20837),
            .I(N__20834));
    LocalMux I__4180 (
            .O(N__20834),
            .I(N__20831));
    Span4Mux_v I__4179 (
            .O(N__20831),
            .I(N__20826));
    InMux I__4178 (
            .O(N__20830),
            .I(N__20823));
    CascadeMux I__4177 (
            .O(N__20829),
            .I(N__20820));
    Span4Mux_h I__4176 (
            .O(N__20826),
            .I(N__20817));
    LocalMux I__4175 (
            .O(N__20823),
            .I(N__20814));
    InMux I__4174 (
            .O(N__20820),
            .I(N__20811));
    Odrv4 I__4173 (
            .O(N__20817),
            .I(\eeprom.n3206 ));
    Odrv4 I__4172 (
            .O(N__20814),
            .I(\eeprom.n3206 ));
    LocalMux I__4171 (
            .O(N__20811),
            .I(\eeprom.n3206 ));
    InMux I__4170 (
            .O(N__20804),
            .I(N__20800));
    CascadeMux I__4169 (
            .O(N__20803),
            .I(N__20797));
    LocalMux I__4168 (
            .O(N__20800),
            .I(N__20793));
    InMux I__4167 (
            .O(N__20797),
            .I(N__20790));
    CascadeMux I__4166 (
            .O(N__20796),
            .I(N__20787));
    Span4Mux_v I__4165 (
            .O(N__20793),
            .I(N__20782));
    LocalMux I__4164 (
            .O(N__20790),
            .I(N__20782));
    InMux I__4163 (
            .O(N__20787),
            .I(N__20779));
    Span4Mux_h I__4162 (
            .O(N__20782),
            .I(N__20776));
    LocalMux I__4161 (
            .O(N__20779),
            .I(N__20773));
    Odrv4 I__4160 (
            .O(N__20776),
            .I(\eeprom.n3214 ));
    Odrv4 I__4159 (
            .O(N__20773),
            .I(\eeprom.n3214 ));
    InMux I__4158 (
            .O(N__20768),
            .I(N__20764));
    InMux I__4157 (
            .O(N__20767),
            .I(N__20760));
    LocalMux I__4156 (
            .O(N__20764),
            .I(N__20757));
    InMux I__4155 (
            .O(N__20763),
            .I(N__20754));
    LocalMux I__4154 (
            .O(N__20760),
            .I(N__20751));
    Span4Mux_v I__4153 (
            .O(N__20757),
            .I(N__20748));
    LocalMux I__4152 (
            .O(N__20754),
            .I(N__20745));
    Span4Mux_h I__4151 (
            .O(N__20751),
            .I(N__20742));
    Span4Mux_v I__4150 (
            .O(N__20748),
            .I(N__20737));
    Span4Mux_v I__4149 (
            .O(N__20745),
            .I(N__20737));
    Span4Mux_h I__4148 (
            .O(N__20742),
            .I(N__20734));
    Span4Mux_h I__4147 (
            .O(N__20737),
            .I(N__20731));
    Odrv4 I__4146 (
            .O(N__20734),
            .I(\eeprom.n3119 ));
    Odrv4 I__4145 (
            .O(N__20731),
            .I(\eeprom.n3119 ));
    InMux I__4144 (
            .O(N__20726),
            .I(N__20723));
    LocalMux I__4143 (
            .O(N__20723),
            .I(N__20720));
    Span4Mux_v I__4142 (
            .O(N__20720),
            .I(N__20717));
    Span4Mux_h I__4141 (
            .O(N__20717),
            .I(N__20714));
    Odrv4 I__4140 (
            .O(N__20714),
            .I(\eeprom.n3186 ));
    InMux I__4139 (
            .O(N__20711),
            .I(bfn_12_22_0_));
    CascadeMux I__4138 (
            .O(N__20708),
            .I(N__20705));
    InMux I__4137 (
            .O(N__20705),
            .I(N__20702));
    LocalMux I__4136 (
            .O(N__20702),
            .I(N__20699));
    Odrv4 I__4135 (
            .O(N__20699),
            .I(\eeprom.n3185 ));
    InMux I__4134 (
            .O(N__20696),
            .I(\eeprom.n3667 ));
    CascadeMux I__4133 (
            .O(N__20693),
            .I(N__20689));
    InMux I__4132 (
            .O(N__20692),
            .I(N__20685));
    InMux I__4131 (
            .O(N__20689),
            .I(N__20682));
    InMux I__4130 (
            .O(N__20688),
            .I(N__20679));
    LocalMux I__4129 (
            .O(N__20685),
            .I(N__20674));
    LocalMux I__4128 (
            .O(N__20682),
            .I(N__20674));
    LocalMux I__4127 (
            .O(N__20679),
            .I(N__20671));
    Odrv4 I__4126 (
            .O(N__20674),
            .I(\eeprom.n3303 ));
    Odrv4 I__4125 (
            .O(N__20671),
            .I(\eeprom.n3303 ));
    InMux I__4124 (
            .O(N__20666),
            .I(N__20663));
    LocalMux I__4123 (
            .O(N__20663),
            .I(N__20660));
    Odrv4 I__4122 (
            .O(N__20660),
            .I(\eeprom.n3370 ));
    InMux I__4121 (
            .O(N__20657),
            .I(N__20654));
    LocalMux I__4120 (
            .O(N__20654),
            .I(N__20651));
    Odrv4 I__4119 (
            .O(N__20651),
            .I(\eeprom.n3366 ));
    CascadeMux I__4118 (
            .O(N__20648),
            .I(N__20644));
    CascadeMux I__4117 (
            .O(N__20647),
            .I(N__20640));
    InMux I__4116 (
            .O(N__20644),
            .I(N__20637));
    InMux I__4115 (
            .O(N__20643),
            .I(N__20634));
    InMux I__4114 (
            .O(N__20640),
            .I(N__20631));
    LocalMux I__4113 (
            .O(N__20637),
            .I(N__20626));
    LocalMux I__4112 (
            .O(N__20634),
            .I(N__20626));
    LocalMux I__4111 (
            .O(N__20631),
            .I(N__20623));
    Span4Mux_v I__4110 (
            .O(N__20626),
            .I(N__20620));
    Odrv4 I__4109 (
            .O(N__20623),
            .I(\eeprom.n3299 ));
    Odrv4 I__4108 (
            .O(N__20620),
            .I(\eeprom.n3299 ));
    CascadeMux I__4107 (
            .O(N__20615),
            .I(N__20612));
    InMux I__4106 (
            .O(N__20612),
            .I(N__20603));
    CascadeMux I__4105 (
            .O(N__20611),
            .I(N__20600));
    CascadeMux I__4104 (
            .O(N__20610),
            .I(N__20592));
    CascadeMux I__4103 (
            .O(N__20609),
            .I(N__20589));
    CascadeMux I__4102 (
            .O(N__20608),
            .I(N__20582));
    InMux I__4101 (
            .O(N__20607),
            .I(N__20573));
    InMux I__4100 (
            .O(N__20606),
            .I(N__20573));
    LocalMux I__4099 (
            .O(N__20603),
            .I(N__20570));
    InMux I__4098 (
            .O(N__20600),
            .I(N__20567));
    CascadeMux I__4097 (
            .O(N__20599),
            .I(N__20564));
    CascadeMux I__4096 (
            .O(N__20598),
            .I(N__20561));
    CascadeMux I__4095 (
            .O(N__20597),
            .I(N__20558));
    InMux I__4094 (
            .O(N__20596),
            .I(N__20554));
    InMux I__4093 (
            .O(N__20595),
            .I(N__20551));
    InMux I__4092 (
            .O(N__20592),
            .I(N__20544));
    InMux I__4091 (
            .O(N__20589),
            .I(N__20544));
    InMux I__4090 (
            .O(N__20588),
            .I(N__20544));
    InMux I__4089 (
            .O(N__20587),
            .I(N__20539));
    InMux I__4088 (
            .O(N__20586),
            .I(N__20539));
    InMux I__4087 (
            .O(N__20585),
            .I(N__20532));
    InMux I__4086 (
            .O(N__20582),
            .I(N__20532));
    InMux I__4085 (
            .O(N__20581),
            .I(N__20532));
    InMux I__4084 (
            .O(N__20580),
            .I(N__20527));
    InMux I__4083 (
            .O(N__20579),
            .I(N__20527));
    InMux I__4082 (
            .O(N__20578),
            .I(N__20524));
    LocalMux I__4081 (
            .O(N__20573),
            .I(N__20519));
    Span4Mux_v I__4080 (
            .O(N__20570),
            .I(N__20519));
    LocalMux I__4079 (
            .O(N__20567),
            .I(N__20516));
    InMux I__4078 (
            .O(N__20564),
            .I(N__20507));
    InMux I__4077 (
            .O(N__20561),
            .I(N__20507));
    InMux I__4076 (
            .O(N__20558),
            .I(N__20507));
    InMux I__4075 (
            .O(N__20557),
            .I(N__20507));
    LocalMux I__4074 (
            .O(N__20554),
            .I(\eeprom.n3331 ));
    LocalMux I__4073 (
            .O(N__20551),
            .I(\eeprom.n3331 ));
    LocalMux I__4072 (
            .O(N__20544),
            .I(\eeprom.n3331 ));
    LocalMux I__4071 (
            .O(N__20539),
            .I(\eeprom.n3331 ));
    LocalMux I__4070 (
            .O(N__20532),
            .I(\eeprom.n3331 ));
    LocalMux I__4069 (
            .O(N__20527),
            .I(\eeprom.n3331 ));
    LocalMux I__4068 (
            .O(N__20524),
            .I(\eeprom.n3331 ));
    Odrv4 I__4067 (
            .O(N__20519),
            .I(\eeprom.n3331 ));
    Odrv4 I__4066 (
            .O(N__20516),
            .I(\eeprom.n3331 ));
    LocalMux I__4065 (
            .O(N__20507),
            .I(\eeprom.n3331 ));
    CascadeMux I__4064 (
            .O(N__20486),
            .I(\eeprom.n3500_cascade_ ));
    InMux I__4063 (
            .O(N__20483),
            .I(N__20479));
    CascadeMux I__4062 (
            .O(N__20482),
            .I(N__20476));
    LocalMux I__4061 (
            .O(N__20479),
            .I(N__20473));
    InMux I__4060 (
            .O(N__20476),
            .I(N__20470));
    Span4Mux_h I__4059 (
            .O(N__20473),
            .I(N__20466));
    LocalMux I__4058 (
            .O(N__20470),
            .I(N__20463));
    InMux I__4057 (
            .O(N__20469),
            .I(N__20460));
    Odrv4 I__4056 (
            .O(N__20466),
            .I(\eeprom.n3216 ));
    Odrv4 I__4055 (
            .O(N__20463),
            .I(\eeprom.n3216 ));
    LocalMux I__4054 (
            .O(N__20460),
            .I(\eeprom.n3216 ));
    CascadeMux I__4053 (
            .O(N__20453),
            .I(N__20450));
    InMux I__4052 (
            .O(N__20450),
            .I(N__20446));
    InMux I__4051 (
            .O(N__20449),
            .I(N__20443));
    LocalMux I__4050 (
            .O(N__20446),
            .I(N__20438));
    LocalMux I__4049 (
            .O(N__20443),
            .I(N__20438));
    Span4Mux_h I__4048 (
            .O(N__20438),
            .I(N__20434));
    InMux I__4047 (
            .O(N__20437),
            .I(N__20431));
    Odrv4 I__4046 (
            .O(N__20434),
            .I(\eeprom.n3203 ));
    LocalMux I__4045 (
            .O(N__20431),
            .I(\eeprom.n3203 ));
    CascadeMux I__4044 (
            .O(N__20426),
            .I(N__20422));
    CascadeMux I__4043 (
            .O(N__20425),
            .I(N__20419));
    InMux I__4042 (
            .O(N__20422),
            .I(N__20416));
    InMux I__4041 (
            .O(N__20419),
            .I(N__20412));
    LocalMux I__4040 (
            .O(N__20416),
            .I(N__20409));
    InMux I__4039 (
            .O(N__20415),
            .I(N__20406));
    LocalMux I__4038 (
            .O(N__20412),
            .I(\eeprom.n3217 ));
    Odrv12 I__4037 (
            .O(N__20409),
            .I(\eeprom.n3217 ));
    LocalMux I__4036 (
            .O(N__20406),
            .I(\eeprom.n3217 ));
    CascadeMux I__4035 (
            .O(N__20399),
            .I(\eeprom.n3410_cascade_ ));
    CascadeMux I__4034 (
            .O(N__20396),
            .I(\eeprom.n3505_cascade_ ));
    InMux I__4033 (
            .O(N__20393),
            .I(N__20390));
    LocalMux I__4032 (
            .O(N__20390),
            .I(N__20387));
    Span4Mux_h I__4031 (
            .O(N__20387),
            .I(N__20382));
    InMux I__4030 (
            .O(N__20386),
            .I(N__20379));
    InMux I__4029 (
            .O(N__20385),
            .I(N__20376));
    Odrv4 I__4028 (
            .O(N__20382),
            .I(\eeprom.n3310 ));
    LocalMux I__4027 (
            .O(N__20379),
            .I(\eeprom.n3310 ));
    LocalMux I__4026 (
            .O(N__20376),
            .I(\eeprom.n3310 ));
    CascadeMux I__4025 (
            .O(N__20369),
            .I(N__20366));
    InMux I__4024 (
            .O(N__20366),
            .I(N__20363));
    LocalMux I__4023 (
            .O(N__20363),
            .I(N__20360));
    Odrv4 I__4022 (
            .O(N__20360),
            .I(\eeprom.n3377 ));
    CascadeMux I__4021 (
            .O(N__20357),
            .I(\eeprom.n3608_adj_451_cascade_ ));
    InMux I__4020 (
            .O(N__20354),
            .I(N__20349));
    CascadeMux I__4019 (
            .O(N__20353),
            .I(N__20346));
    InMux I__4018 (
            .O(N__20352),
            .I(N__20343));
    LocalMux I__4017 (
            .O(N__20349),
            .I(N__20340));
    InMux I__4016 (
            .O(N__20346),
            .I(N__20337));
    LocalMux I__4015 (
            .O(N__20343),
            .I(N__20334));
    Span4Mux_h I__4014 (
            .O(N__20340),
            .I(N__20331));
    LocalMux I__4013 (
            .O(N__20337),
            .I(N__20328));
    Odrv12 I__4012 (
            .O(N__20334),
            .I(\eeprom.n3313 ));
    Odrv4 I__4011 (
            .O(N__20331),
            .I(\eeprom.n3313 ));
    Odrv4 I__4010 (
            .O(N__20328),
            .I(\eeprom.n3313 ));
    CascadeMux I__4009 (
            .O(N__20321),
            .I(N__20318));
    InMux I__4008 (
            .O(N__20318),
            .I(N__20315));
    LocalMux I__4007 (
            .O(N__20315),
            .I(N__20312));
    Span4Mux_h I__4006 (
            .O(N__20312),
            .I(N__20309));
    Odrv4 I__4005 (
            .O(N__20309),
            .I(\eeprom.n3380 ));
    CascadeMux I__4004 (
            .O(N__20306),
            .I(\eeprom.n3412_cascade_ ));
    CascadeMux I__4003 (
            .O(N__20303),
            .I(\eeprom.n3414_cascade_ ));
    CascadeMux I__4002 (
            .O(N__20300),
            .I(\eeprom.n4689_cascade_ ));
    CascadeMux I__4001 (
            .O(N__20297),
            .I(\eeprom.n4144_cascade_ ));
    InMux I__4000 (
            .O(N__20294),
            .I(N__20291));
    LocalMux I__3999 (
            .O(N__20291),
            .I(N__20288));
    Span4Mux_h I__3998 (
            .O(N__20288),
            .I(N__20285));
    Odrv4 I__3997 (
            .O(N__20285),
            .I(\eeprom.n3386 ));
    InMux I__3996 (
            .O(N__20282),
            .I(N__20278));
    InMux I__3995 (
            .O(N__20281),
            .I(N__20275));
    LocalMux I__3994 (
            .O(N__20278),
            .I(N__20269));
    LocalMux I__3993 (
            .O(N__20275),
            .I(N__20269));
    InMux I__3992 (
            .O(N__20274),
            .I(N__20266));
    Span4Mux_h I__3991 (
            .O(N__20269),
            .I(N__20263));
    LocalMux I__3990 (
            .O(N__20266),
            .I(N__20260));
    Span4Mux_h I__3989 (
            .O(N__20263),
            .I(N__20257));
    Span4Mux_v I__3988 (
            .O(N__20260),
            .I(N__20254));
    Odrv4 I__3987 (
            .O(N__20257),
            .I(\eeprom.n3319 ));
    Odrv4 I__3986 (
            .O(N__20254),
            .I(\eeprom.n3319 ));
    CascadeMux I__3985 (
            .O(N__20249),
            .I(N__20245));
    InMux I__3984 (
            .O(N__20248),
            .I(N__20241));
    InMux I__3983 (
            .O(N__20245),
            .I(N__20238));
    InMux I__3982 (
            .O(N__20244),
            .I(N__20235));
    LocalMux I__3981 (
            .O(N__20241),
            .I(N__20230));
    LocalMux I__3980 (
            .O(N__20238),
            .I(N__20230));
    LocalMux I__3979 (
            .O(N__20235),
            .I(N__20227));
    Span4Mux_h I__3978 (
            .O(N__20230),
            .I(N__20224));
    Odrv4 I__3977 (
            .O(N__20227),
            .I(\eeprom.n3316 ));
    Odrv4 I__3976 (
            .O(N__20224),
            .I(\eeprom.n3316 ));
    CascadeMux I__3975 (
            .O(N__20219),
            .I(N__20216));
    InMux I__3974 (
            .O(N__20216),
            .I(N__20213));
    LocalMux I__3973 (
            .O(N__20213),
            .I(N__20210));
    Odrv4 I__3972 (
            .O(N__20210),
            .I(\eeprom.n3383 ));
    InMux I__3971 (
            .O(N__20207),
            .I(N__20203));
    CascadeMux I__3970 (
            .O(N__20206),
            .I(N__20200));
    LocalMux I__3969 (
            .O(N__20203),
            .I(N__20197));
    InMux I__3968 (
            .O(N__20200),
            .I(N__20194));
    Odrv12 I__3967 (
            .O(N__20197),
            .I(\eeprom.n3314 ));
    LocalMux I__3966 (
            .O(N__20194),
            .I(\eeprom.n3314 ));
    InMux I__3965 (
            .O(N__20189),
            .I(N__20186));
    LocalMux I__3964 (
            .O(N__20186),
            .I(N__20183));
    Odrv4 I__3963 (
            .O(N__20183),
            .I(\eeprom.n3381 ));
    CascadeMux I__3962 (
            .O(N__20180),
            .I(\eeprom.n3413_cascade_ ));
    InMux I__3961 (
            .O(N__20177),
            .I(N__20174));
    LocalMux I__3960 (
            .O(N__20174),
            .I(\eeprom.n4687 ));
    InMux I__3959 (
            .O(N__20171),
            .I(N__20168));
    LocalMux I__3958 (
            .O(N__20168),
            .I(N__20165));
    Odrv12 I__3957 (
            .O(N__20165),
            .I(\eeprom.n3378 ));
    CascadeMux I__3956 (
            .O(N__20162),
            .I(N__20159));
    InMux I__3955 (
            .O(N__20159),
            .I(N__20156));
    LocalMux I__3954 (
            .O(N__20156),
            .I(N__20152));
    CascadeMux I__3953 (
            .O(N__20155),
            .I(N__20148));
    Span4Mux_h I__3952 (
            .O(N__20152),
            .I(N__20145));
    InMux I__3951 (
            .O(N__20151),
            .I(N__20142));
    InMux I__3950 (
            .O(N__20148),
            .I(N__20139));
    Odrv4 I__3949 (
            .O(N__20145),
            .I(\eeprom.n3311 ));
    LocalMux I__3948 (
            .O(N__20142),
            .I(\eeprom.n3311 ));
    LocalMux I__3947 (
            .O(N__20139),
            .I(\eeprom.n3311 ));
    CascadeMux I__3946 (
            .O(N__20132),
            .I(N__20127));
    CascadeMux I__3945 (
            .O(N__20131),
            .I(N__20124));
    InMux I__3944 (
            .O(N__20130),
            .I(N__20121));
    InMux I__3943 (
            .O(N__20127),
            .I(N__20118));
    InMux I__3942 (
            .O(N__20124),
            .I(N__20115));
    LocalMux I__3941 (
            .O(N__20121),
            .I(N__20112));
    LocalMux I__3940 (
            .O(N__20118),
            .I(N__20107));
    LocalMux I__3939 (
            .O(N__20115),
            .I(N__20107));
    Span4Mux_v I__3938 (
            .O(N__20112),
            .I(N__20104));
    Span4Mux_v I__3937 (
            .O(N__20107),
            .I(N__20101));
    Odrv4 I__3936 (
            .O(N__20104),
            .I(\eeprom.n2817 ));
    Odrv4 I__3935 (
            .O(N__20101),
            .I(\eeprom.n2817 ));
    CascadeMux I__3934 (
            .O(N__20096),
            .I(N__20093));
    InMux I__3933 (
            .O(N__20093),
            .I(N__20090));
    LocalMux I__3932 (
            .O(N__20090),
            .I(N__20087));
    Odrv4 I__3931 (
            .O(N__20087),
            .I(\eeprom.n2884 ));
    CascadeMux I__3930 (
            .O(N__20084),
            .I(N__20081));
    InMux I__3929 (
            .O(N__20081),
            .I(N__20078));
    LocalMux I__3928 (
            .O(N__20078),
            .I(N__20075));
    Odrv4 I__3927 (
            .O(N__20075),
            .I(\eeprom.n2877 ));
    InMux I__3926 (
            .O(N__20072),
            .I(N__20067));
    InMux I__3925 (
            .O(N__20071),
            .I(N__20064));
    InMux I__3924 (
            .O(N__20070),
            .I(N__20061));
    LocalMux I__3923 (
            .O(N__20067),
            .I(N__20056));
    LocalMux I__3922 (
            .O(N__20064),
            .I(N__20056));
    LocalMux I__3921 (
            .O(N__20061),
            .I(N__20053));
    Span4Mux_h I__3920 (
            .O(N__20056),
            .I(N__20050));
    Odrv4 I__3919 (
            .O(N__20053),
            .I(\eeprom.n2810 ));
    Odrv4 I__3918 (
            .O(N__20050),
            .I(\eeprom.n2810 ));
    CascadeMux I__3917 (
            .O(N__20045),
            .I(\eeprom.n2909_cascade_ ));
    InMux I__3916 (
            .O(N__20042),
            .I(N__20039));
    LocalMux I__3915 (
            .O(N__20039),
            .I(\eeprom.n18_adj_420 ));
    CascadeMux I__3914 (
            .O(N__20036),
            .I(N__20033));
    InMux I__3913 (
            .O(N__20033),
            .I(N__20030));
    LocalMux I__3912 (
            .O(N__20030),
            .I(N__20027));
    Odrv4 I__3911 (
            .O(N__20027),
            .I(\eeprom.n2975 ));
    InMux I__3910 (
            .O(N__20024),
            .I(N__20019));
    InMux I__3909 (
            .O(N__20023),
            .I(N__20016));
    InMux I__3908 (
            .O(N__20022),
            .I(N__20013));
    LocalMux I__3907 (
            .O(N__20019),
            .I(\eeprom.n2908 ));
    LocalMux I__3906 (
            .O(N__20016),
            .I(\eeprom.n2908 ));
    LocalMux I__3905 (
            .O(N__20013),
            .I(\eeprom.n2908 ));
    InMux I__3904 (
            .O(N__20006),
            .I(N__20003));
    LocalMux I__3903 (
            .O(N__20003),
            .I(N__20000));
    Odrv4 I__3902 (
            .O(N__20000),
            .I(\eeprom.n2878 ));
    CascadeMux I__3901 (
            .O(N__19997),
            .I(N__19993));
    CascadeMux I__3900 (
            .O(N__19996),
            .I(N__19990));
    InMux I__3899 (
            .O(N__19993),
            .I(N__19987));
    InMux I__3898 (
            .O(N__19990),
            .I(N__19984));
    LocalMux I__3897 (
            .O(N__19987),
            .I(N__19980));
    LocalMux I__3896 (
            .O(N__19984),
            .I(N__19977));
    InMux I__3895 (
            .O(N__19983),
            .I(N__19974));
    Odrv4 I__3894 (
            .O(N__19980),
            .I(\eeprom.n2811 ));
    Odrv4 I__3893 (
            .O(N__19977),
            .I(\eeprom.n2811 ));
    LocalMux I__3892 (
            .O(N__19974),
            .I(\eeprom.n2811 ));
    CascadeMux I__3891 (
            .O(N__19967),
            .I(N__19960));
    CascadeMux I__3890 (
            .O(N__19966),
            .I(N__19955));
    CascadeMux I__3889 (
            .O(N__19965),
            .I(N__19949));
    CascadeMux I__3888 (
            .O(N__19964),
            .I(N__19945));
    InMux I__3887 (
            .O(N__19963),
            .I(N__19936));
    InMux I__3886 (
            .O(N__19960),
            .I(N__19936));
    InMux I__3885 (
            .O(N__19959),
            .I(N__19936));
    CascadeMux I__3884 (
            .O(N__19958),
            .I(N__19931));
    InMux I__3883 (
            .O(N__19955),
            .I(N__19925));
    InMux I__3882 (
            .O(N__19954),
            .I(N__19925));
    InMux I__3881 (
            .O(N__19953),
            .I(N__19920));
    InMux I__3880 (
            .O(N__19952),
            .I(N__19920));
    InMux I__3879 (
            .O(N__19949),
            .I(N__19915));
    InMux I__3878 (
            .O(N__19948),
            .I(N__19915));
    InMux I__3877 (
            .O(N__19945),
            .I(N__19908));
    InMux I__3876 (
            .O(N__19944),
            .I(N__19908));
    InMux I__3875 (
            .O(N__19943),
            .I(N__19908));
    LocalMux I__3874 (
            .O(N__19936),
            .I(N__19905));
    InMux I__3873 (
            .O(N__19935),
            .I(N__19902));
    InMux I__3872 (
            .O(N__19934),
            .I(N__19895));
    InMux I__3871 (
            .O(N__19931),
            .I(N__19895));
    InMux I__3870 (
            .O(N__19930),
            .I(N__19895));
    LocalMux I__3869 (
            .O(N__19925),
            .I(N__19892));
    LocalMux I__3868 (
            .O(N__19920),
            .I(\eeprom.n2836 ));
    LocalMux I__3867 (
            .O(N__19915),
            .I(\eeprom.n2836 ));
    LocalMux I__3866 (
            .O(N__19908),
            .I(\eeprom.n2836 ));
    Odrv4 I__3865 (
            .O(N__19905),
            .I(\eeprom.n2836 ));
    LocalMux I__3864 (
            .O(N__19902),
            .I(\eeprom.n2836 ));
    LocalMux I__3863 (
            .O(N__19895),
            .I(\eeprom.n2836 ));
    Odrv4 I__3862 (
            .O(N__19892),
            .I(\eeprom.n2836 ));
    CascadeMux I__3861 (
            .O(N__19877),
            .I(N__19874));
    InMux I__3860 (
            .O(N__19874),
            .I(N__19870));
    InMux I__3859 (
            .O(N__19873),
            .I(N__19866));
    LocalMux I__3858 (
            .O(N__19870),
            .I(N__19863));
    InMux I__3857 (
            .O(N__19869),
            .I(N__19860));
    LocalMux I__3856 (
            .O(N__19866),
            .I(\eeprom.n2915 ));
    Odrv4 I__3855 (
            .O(N__19863),
            .I(\eeprom.n2915 ));
    LocalMux I__3854 (
            .O(N__19860),
            .I(\eeprom.n2915 ));
    InMux I__3853 (
            .O(N__19853),
            .I(N__19850));
    LocalMux I__3852 (
            .O(N__19850),
            .I(N__19847));
    Odrv12 I__3851 (
            .O(N__19847),
            .I(\eeprom.n2982 ));
    InMux I__3850 (
            .O(N__19844),
            .I(N__19839));
    InMux I__3849 (
            .O(N__19843),
            .I(N__19836));
    InMux I__3848 (
            .O(N__19842),
            .I(N__19833));
    LocalMux I__3847 (
            .O(N__19839),
            .I(\eeprom.n2911 ));
    LocalMux I__3846 (
            .O(N__19836),
            .I(\eeprom.n2911 ));
    LocalMux I__3845 (
            .O(N__19833),
            .I(\eeprom.n2911 ));
    CascadeMux I__3844 (
            .O(N__19826),
            .I(N__19823));
    InMux I__3843 (
            .O(N__19823),
            .I(N__19820));
    LocalMux I__3842 (
            .O(N__19820),
            .I(N__19817));
    Odrv4 I__3841 (
            .O(N__19817),
            .I(\eeprom.n2978 ));
    InMux I__3840 (
            .O(N__19814),
            .I(N__19811));
    LocalMux I__3839 (
            .O(N__19811),
            .I(N__19808));
    Odrv4 I__3838 (
            .O(N__19808),
            .I(\eeprom.n2984 ));
    CascadeMux I__3837 (
            .O(N__19805),
            .I(N__19802));
    InMux I__3836 (
            .O(N__19802),
            .I(N__19798));
    InMux I__3835 (
            .O(N__19801),
            .I(N__19795));
    LocalMux I__3834 (
            .O(N__19798),
            .I(N__19792));
    LocalMux I__3833 (
            .O(N__19795),
            .I(\eeprom.n2917 ));
    Odrv4 I__3832 (
            .O(N__19792),
            .I(\eeprom.n2917 ));
    CascadeMux I__3831 (
            .O(N__19787),
            .I(N__19784));
    InMux I__3830 (
            .O(N__19784),
            .I(N__19780));
    InMux I__3829 (
            .O(N__19783),
            .I(N__19777));
    LocalMux I__3828 (
            .O(N__19780),
            .I(N__19774));
    LocalMux I__3827 (
            .O(N__19777),
            .I(\eeprom.n3315 ));
    Odrv4 I__3826 (
            .O(N__19774),
            .I(\eeprom.n3315 ));
    InMux I__3825 (
            .O(N__19769),
            .I(N__19766));
    LocalMux I__3824 (
            .O(N__19766),
            .I(N__19763));
    Odrv4 I__3823 (
            .O(N__19763),
            .I(\eeprom.n3382 ));
    InMux I__3822 (
            .O(N__19760),
            .I(\eeprom.n3646 ));
    InMux I__3821 (
            .O(N__19757),
            .I(bfn_11_23_0_));
    InMux I__3820 (
            .O(N__19754),
            .I(N__19751));
    LocalMux I__3819 (
            .O(N__19751),
            .I(N__19748));
    Span4Mux_h I__3818 (
            .O(N__19748),
            .I(N__19744));
    InMux I__3817 (
            .O(N__19747),
            .I(N__19741));
    Odrv4 I__3816 (
            .O(N__19744),
            .I(\eeprom.n2902 ));
    LocalMux I__3815 (
            .O(N__19741),
            .I(\eeprom.n2902 ));
    InMux I__3814 (
            .O(N__19736),
            .I(\eeprom.n3648 ));
    InMux I__3813 (
            .O(N__19733),
            .I(N__19728));
    InMux I__3812 (
            .O(N__19732),
            .I(N__19725));
    InMux I__3811 (
            .O(N__19731),
            .I(N__19722));
    LocalMux I__3810 (
            .O(N__19728),
            .I(N__19719));
    LocalMux I__3809 (
            .O(N__19725),
            .I(\eeprom.n2906 ));
    LocalMux I__3808 (
            .O(N__19722),
            .I(\eeprom.n2906 ));
    Odrv4 I__3807 (
            .O(N__19719),
            .I(\eeprom.n2906 ));
    CascadeMux I__3806 (
            .O(N__19712),
            .I(N__19709));
    InMux I__3805 (
            .O(N__19709),
            .I(N__19706));
    LocalMux I__3804 (
            .O(N__19706),
            .I(\eeprom.n2973 ));
    InMux I__3803 (
            .O(N__19703),
            .I(N__19698));
    InMux I__3802 (
            .O(N__19702),
            .I(N__19693));
    InMux I__3801 (
            .O(N__19701),
            .I(N__19693));
    LocalMux I__3800 (
            .O(N__19698),
            .I(N__19690));
    LocalMux I__3799 (
            .O(N__19693),
            .I(\eeprom.n2903 ));
    Odrv4 I__3798 (
            .O(N__19690),
            .I(\eeprom.n2903 ));
    InMux I__3797 (
            .O(N__19685),
            .I(N__19682));
    LocalMux I__3796 (
            .O(N__19682),
            .I(\eeprom.n2970 ));
    InMux I__3795 (
            .O(N__19679),
            .I(N__19676));
    LocalMux I__3794 (
            .O(N__19676),
            .I(N__19673));
    Odrv4 I__3793 (
            .O(N__19673),
            .I(\eeprom.n2879 ));
    InMux I__3792 (
            .O(N__19670),
            .I(N__19665));
    InMux I__3791 (
            .O(N__19669),
            .I(N__19662));
    InMux I__3790 (
            .O(N__19668),
            .I(N__19659));
    LocalMux I__3789 (
            .O(N__19665),
            .I(N__19656));
    LocalMux I__3788 (
            .O(N__19662),
            .I(N__19651));
    LocalMux I__3787 (
            .O(N__19659),
            .I(N__19651));
    Odrv12 I__3786 (
            .O(N__19656),
            .I(\eeprom.n2812 ));
    Odrv4 I__3785 (
            .O(N__19651),
            .I(\eeprom.n2812 ));
    InMux I__3784 (
            .O(N__19646),
            .I(N__19643));
    LocalMux I__3783 (
            .O(N__19643),
            .I(N__19640));
    Odrv4 I__3782 (
            .O(N__19640),
            .I(\eeprom.n2880 ));
    CascadeMux I__3781 (
            .O(N__19637),
            .I(N__19634));
    InMux I__3780 (
            .O(N__19634),
            .I(N__19630));
    CascadeMux I__3779 (
            .O(N__19633),
            .I(N__19627));
    LocalMux I__3778 (
            .O(N__19630),
            .I(N__19624));
    InMux I__3777 (
            .O(N__19627),
            .I(N__19621));
    Span4Mux_h I__3776 (
            .O(N__19624),
            .I(N__19616));
    LocalMux I__3775 (
            .O(N__19621),
            .I(N__19616));
    Span4Mux_h I__3774 (
            .O(N__19616),
            .I(N__19612));
    InMux I__3773 (
            .O(N__19615),
            .I(N__19609));
    Odrv4 I__3772 (
            .O(N__19612),
            .I(\eeprom.n2813 ));
    LocalMux I__3771 (
            .O(N__19609),
            .I(\eeprom.n2813 ));
    InMux I__3770 (
            .O(N__19604),
            .I(N__19600));
    InMux I__3769 (
            .O(N__19603),
            .I(N__19597));
    LocalMux I__3768 (
            .O(N__19600),
            .I(N__19594));
    LocalMux I__3767 (
            .O(N__19597),
            .I(\eeprom.n2913 ));
    Odrv4 I__3766 (
            .O(N__19594),
            .I(\eeprom.n2913 ));
    CascadeMux I__3765 (
            .O(N__19589),
            .I(N__19586));
    InMux I__3764 (
            .O(N__19586),
            .I(N__19583));
    LocalMux I__3763 (
            .O(N__19583),
            .I(N__19580));
    Odrv4 I__3762 (
            .O(N__19580),
            .I(\eeprom.n2980 ));
    InMux I__3761 (
            .O(N__19577),
            .I(\eeprom.n3637 ));
    InMux I__3760 (
            .O(N__19574),
            .I(\eeprom.n3638 ));
    InMux I__3759 (
            .O(N__19571),
            .I(bfn_11_22_0_));
    InMux I__3758 (
            .O(N__19568),
            .I(\eeprom.n3640 ));
    InMux I__3757 (
            .O(N__19565),
            .I(\eeprom.n3641 ));
    InMux I__3756 (
            .O(N__19562),
            .I(\eeprom.n3642 ));
    InMux I__3755 (
            .O(N__19559),
            .I(\eeprom.n3643 ));
    InMux I__3754 (
            .O(N__19556),
            .I(\eeprom.n3644 ));
    InMux I__3753 (
            .O(N__19553),
            .I(\eeprom.n3645 ));
    CascadeMux I__3752 (
            .O(N__19550),
            .I(N__19546));
    InMux I__3751 (
            .O(N__19549),
            .I(N__19543));
    InMux I__3750 (
            .O(N__19546),
            .I(N__19540));
    LocalMux I__3749 (
            .O(N__19543),
            .I(N__19536));
    LocalMux I__3748 (
            .O(N__19540),
            .I(N__19533));
    InMux I__3747 (
            .O(N__19539),
            .I(N__19530));
    Odrv4 I__3746 (
            .O(N__19536),
            .I(\eeprom.n3213 ));
    Odrv4 I__3745 (
            .O(N__19533),
            .I(\eeprom.n3213 ));
    LocalMux I__3744 (
            .O(N__19530),
            .I(\eeprom.n3213 ));
    CascadeMux I__3743 (
            .O(N__19523),
            .I(\eeprom.n3116_cascade_ ));
    InMux I__3742 (
            .O(N__19520),
            .I(N__19516));
    CascadeMux I__3741 (
            .O(N__19519),
            .I(N__19513));
    LocalMux I__3740 (
            .O(N__19516),
            .I(N__19509));
    InMux I__3739 (
            .O(N__19513),
            .I(N__19506));
    CascadeMux I__3738 (
            .O(N__19512),
            .I(N__19503));
    Span4Mux_h I__3737 (
            .O(N__19509),
            .I(N__19500));
    LocalMux I__3736 (
            .O(N__19506),
            .I(N__19497));
    InMux I__3735 (
            .O(N__19503),
            .I(N__19494));
    Odrv4 I__3734 (
            .O(N__19500),
            .I(\eeprom.n3215 ));
    Odrv4 I__3733 (
            .O(N__19497),
            .I(\eeprom.n3215 ));
    LocalMux I__3732 (
            .O(N__19494),
            .I(\eeprom.n3215 ));
    InMux I__3731 (
            .O(N__19487),
            .I(bfn_11_21_0_));
    CascadeMux I__3730 (
            .O(N__19484),
            .I(N__19480));
    InMux I__3729 (
            .O(N__19483),
            .I(N__19477));
    InMux I__3728 (
            .O(N__19480),
            .I(N__19474));
    LocalMux I__3727 (
            .O(N__19477),
            .I(N__19471));
    LocalMux I__3726 (
            .O(N__19474),
            .I(\eeprom.n2918 ));
    Odrv4 I__3725 (
            .O(N__19471),
            .I(\eeprom.n2918 ));
    InMux I__3724 (
            .O(N__19466),
            .I(N__19463));
    LocalMux I__3723 (
            .O(N__19463),
            .I(\eeprom.n2985 ));
    InMux I__3722 (
            .O(N__19460),
            .I(\eeprom.n3632 ));
    InMux I__3721 (
            .O(N__19457),
            .I(\eeprom.n3633 ));
    InMux I__3720 (
            .O(N__19454),
            .I(\eeprom.n3634 ));
    InMux I__3719 (
            .O(N__19451),
            .I(\eeprom.n3635 ));
    InMux I__3718 (
            .O(N__19448),
            .I(\eeprom.n3636 ));
    CascadeMux I__3717 (
            .O(N__19445),
            .I(N__19442));
    InMux I__3716 (
            .O(N__19442),
            .I(N__19439));
    LocalMux I__3715 (
            .O(N__19439),
            .I(N__19435));
    InMux I__3714 (
            .O(N__19438),
            .I(N__19432));
    Span4Mux_v I__3713 (
            .O(N__19435),
            .I(N__19428));
    LocalMux I__3712 (
            .O(N__19432),
            .I(N__19425));
    InMux I__3711 (
            .O(N__19431),
            .I(N__19422));
    Span4Mux_h I__3710 (
            .O(N__19428),
            .I(N__19419));
    Sp12to4 I__3709 (
            .O(N__19425),
            .I(N__19416));
    LocalMux I__3708 (
            .O(N__19422),
            .I(N__19409));
    Sp12to4 I__3707 (
            .O(N__19419),
            .I(N__19409));
    Span12Mux_v I__3706 (
            .O(N__19416),
            .I(N__19409));
    Odrv12 I__3705 (
            .O(N__19409),
            .I(\eeprom.n3219 ));
    CascadeMux I__3704 (
            .O(N__19406),
            .I(\eeprom.n4615_cascade_ ));
    CascadeMux I__3703 (
            .O(N__19403),
            .I(N__19400));
    InMux I__3702 (
            .O(N__19400),
            .I(N__19396));
    CascadeMux I__3701 (
            .O(N__19399),
            .I(N__19392));
    LocalMux I__3700 (
            .O(N__19396),
            .I(N__19389));
    InMux I__3699 (
            .O(N__19395),
            .I(N__19386));
    InMux I__3698 (
            .O(N__19392),
            .I(N__19383));
    Span4Mux_h I__3697 (
            .O(N__19389),
            .I(N__19378));
    LocalMux I__3696 (
            .O(N__19386),
            .I(N__19378));
    LocalMux I__3695 (
            .O(N__19383),
            .I(\eeprom.n3218 ));
    Odrv4 I__3694 (
            .O(N__19378),
            .I(\eeprom.n3218 ));
    InMux I__3693 (
            .O(N__19373),
            .I(N__19370));
    LocalMux I__3692 (
            .O(N__19370),
            .I(\eeprom.n21_adj_477 ));
    InMux I__3691 (
            .O(N__19367),
            .I(N__19364));
    LocalMux I__3690 (
            .O(N__19364),
            .I(\eeprom.n4611 ));
    CascadeMux I__3689 (
            .O(N__19361),
            .I(N__19357));
    CascadeMux I__3688 (
            .O(N__19360),
            .I(N__19354));
    InMux I__3687 (
            .O(N__19357),
            .I(N__19350));
    InMux I__3686 (
            .O(N__19354),
            .I(N__19347));
    InMux I__3685 (
            .O(N__19353),
            .I(N__19344));
    LocalMux I__3684 (
            .O(N__19350),
            .I(\eeprom.n3300 ));
    LocalMux I__3683 (
            .O(N__19347),
            .I(\eeprom.n3300 ));
    LocalMux I__3682 (
            .O(N__19344),
            .I(\eeprom.n3300 ));
    InMux I__3681 (
            .O(N__19337),
            .I(N__19333));
    InMux I__3680 (
            .O(N__19336),
            .I(N__19330));
    LocalMux I__3679 (
            .O(N__19333),
            .I(N__19327));
    LocalMux I__3678 (
            .O(N__19330),
            .I(N__19324));
    Span4Mux_v I__3677 (
            .O(N__19327),
            .I(N__19321));
    Odrv4 I__3676 (
            .O(N__19324),
            .I(\eeprom.n3298 ));
    Odrv4 I__3675 (
            .O(N__19321),
            .I(\eeprom.n3298 ));
    InMux I__3674 (
            .O(N__19316),
            .I(N__19313));
    LocalMux I__3673 (
            .O(N__19313),
            .I(\eeprom.n25_adj_487 ));
    CascadeMux I__3672 (
            .O(N__19310),
            .I(N__19305));
    InMux I__3671 (
            .O(N__19309),
            .I(N__19302));
    InMux I__3670 (
            .O(N__19308),
            .I(N__19297));
    InMux I__3669 (
            .O(N__19305),
            .I(N__19297));
    LocalMux I__3668 (
            .O(N__19302),
            .I(\eeprom.n3301 ));
    LocalMux I__3667 (
            .O(N__19297),
            .I(\eeprom.n3301 ));
    CascadeMux I__3666 (
            .O(N__19292),
            .I(N__19289));
    InMux I__3665 (
            .O(N__19289),
            .I(N__19286));
    LocalMux I__3664 (
            .O(N__19286),
            .I(N__19283));
    Odrv4 I__3663 (
            .O(N__19283),
            .I(\eeprom.n3368 ));
    InMux I__3662 (
            .O(N__19280),
            .I(N__19277));
    LocalMux I__3661 (
            .O(N__19277),
            .I(N__19274));
    Span4Mux_h I__3660 (
            .O(N__19274),
            .I(N__19271));
    Odrv4 I__3659 (
            .O(N__19271),
            .I(\eeprom.n3284 ));
    CascadeMux I__3658 (
            .O(N__19268),
            .I(N__19263));
    InMux I__3657 (
            .O(N__19267),
            .I(N__19250));
    InMux I__3656 (
            .O(N__19266),
            .I(N__19247));
    InMux I__3655 (
            .O(N__19263),
            .I(N__19244));
    CascadeMux I__3654 (
            .O(N__19262),
            .I(N__19241));
    CascadeMux I__3653 (
            .O(N__19261),
            .I(N__19236));
    CascadeMux I__3652 (
            .O(N__19260),
            .I(N__19233));
    CascadeMux I__3651 (
            .O(N__19259),
            .I(N__19230));
    CascadeMux I__3650 (
            .O(N__19258),
            .I(N__19227));
    CascadeMux I__3649 (
            .O(N__19257),
            .I(N__19221));
    CascadeMux I__3648 (
            .O(N__19256),
            .I(N__19218));
    CascadeMux I__3647 (
            .O(N__19255),
            .I(N__19215));
    CascadeMux I__3646 (
            .O(N__19254),
            .I(N__19212));
    InMux I__3645 (
            .O(N__19253),
            .I(N__19208));
    LocalMux I__3644 (
            .O(N__19250),
            .I(N__19201));
    LocalMux I__3643 (
            .O(N__19247),
            .I(N__19201));
    LocalMux I__3642 (
            .O(N__19244),
            .I(N__19201));
    InMux I__3641 (
            .O(N__19241),
            .I(N__19194));
    InMux I__3640 (
            .O(N__19240),
            .I(N__19194));
    InMux I__3639 (
            .O(N__19239),
            .I(N__19194));
    InMux I__3638 (
            .O(N__19236),
            .I(N__19188));
    InMux I__3637 (
            .O(N__19233),
            .I(N__19188));
    InMux I__3636 (
            .O(N__19230),
            .I(N__19179));
    InMux I__3635 (
            .O(N__19227),
            .I(N__19179));
    InMux I__3634 (
            .O(N__19226),
            .I(N__19179));
    InMux I__3633 (
            .O(N__19225),
            .I(N__19179));
    InMux I__3632 (
            .O(N__19224),
            .I(N__19168));
    InMux I__3631 (
            .O(N__19221),
            .I(N__19168));
    InMux I__3630 (
            .O(N__19218),
            .I(N__19168));
    InMux I__3629 (
            .O(N__19215),
            .I(N__19168));
    InMux I__3628 (
            .O(N__19212),
            .I(N__19168));
    InMux I__3627 (
            .O(N__19211),
            .I(N__19165));
    LocalMux I__3626 (
            .O(N__19208),
            .I(N__19162));
    Span4Mux_v I__3625 (
            .O(N__19201),
            .I(N__19157));
    LocalMux I__3624 (
            .O(N__19194),
            .I(N__19157));
    InMux I__3623 (
            .O(N__19193),
            .I(N__19154));
    LocalMux I__3622 (
            .O(N__19188),
            .I(\eeprom.n3232 ));
    LocalMux I__3621 (
            .O(N__19179),
            .I(\eeprom.n3232 ));
    LocalMux I__3620 (
            .O(N__19168),
            .I(\eeprom.n3232 ));
    LocalMux I__3619 (
            .O(N__19165),
            .I(\eeprom.n3232 ));
    Odrv4 I__3618 (
            .O(N__19162),
            .I(\eeprom.n3232 ));
    Odrv4 I__3617 (
            .O(N__19157),
            .I(\eeprom.n3232 ));
    LocalMux I__3616 (
            .O(N__19154),
            .I(\eeprom.n3232 ));
    InMux I__3615 (
            .O(N__19139),
            .I(N__19136));
    LocalMux I__3614 (
            .O(N__19136),
            .I(N__19132));
    InMux I__3613 (
            .O(N__19135),
            .I(N__19128));
    Span4Mux_h I__3612 (
            .O(N__19132),
            .I(N__19125));
    InMux I__3611 (
            .O(N__19131),
            .I(N__19122));
    LocalMux I__3610 (
            .O(N__19128),
            .I(\eeprom.n3210 ));
    Odrv4 I__3609 (
            .O(N__19125),
            .I(\eeprom.n3210 ));
    LocalMux I__3608 (
            .O(N__19122),
            .I(\eeprom.n3210 ));
    CascadeMux I__3607 (
            .O(N__19115),
            .I(\eeprom.n3113_cascade_ ));
    InMux I__3606 (
            .O(N__19112),
            .I(N__19107));
    InMux I__3605 (
            .O(N__19111),
            .I(N__19102));
    InMux I__3604 (
            .O(N__19110),
            .I(N__19102));
    LocalMux I__3603 (
            .O(N__19107),
            .I(N__19099));
    LocalMux I__3602 (
            .O(N__19102),
            .I(\eeprom.n3212 ));
    Odrv4 I__3601 (
            .O(N__19099),
            .I(\eeprom.n3212 ));
    InMux I__3600 (
            .O(N__19094),
            .I(N__19091));
    LocalMux I__3599 (
            .O(N__19091),
            .I(N__19086));
    InMux I__3598 (
            .O(N__19090),
            .I(N__19083));
    InMux I__3597 (
            .O(N__19089),
            .I(N__19080));
    Odrv4 I__3596 (
            .O(N__19086),
            .I(\eeprom.n3208 ));
    LocalMux I__3595 (
            .O(N__19083),
            .I(\eeprom.n3208 ));
    LocalMux I__3594 (
            .O(N__19080),
            .I(\eeprom.n3208 ));
    CascadeMux I__3593 (
            .O(N__19073),
            .I(N__19070));
    InMux I__3592 (
            .O(N__19070),
            .I(N__19067));
    LocalMux I__3591 (
            .O(N__19067),
            .I(\eeprom.n25_adj_478 ));
    CascadeMux I__3590 (
            .O(N__19064),
            .I(N__19059));
    InMux I__3589 (
            .O(N__19063),
            .I(N__19056));
    InMux I__3588 (
            .O(N__19062),
            .I(N__19053));
    InMux I__3587 (
            .O(N__19059),
            .I(N__19050));
    LocalMux I__3586 (
            .O(N__19056),
            .I(\eeprom.n3317 ));
    LocalMux I__3585 (
            .O(N__19053),
            .I(\eeprom.n3317 ));
    LocalMux I__3584 (
            .O(N__19050),
            .I(\eeprom.n3317 ));
    CascadeMux I__3583 (
            .O(N__19043),
            .I(N__19040));
    InMux I__3582 (
            .O(N__19040),
            .I(N__19037));
    LocalMux I__3581 (
            .O(N__19037),
            .I(N__19034));
    Odrv4 I__3580 (
            .O(N__19034),
            .I(\eeprom.n3384 ));
    InMux I__3579 (
            .O(N__19031),
            .I(N__19028));
    LocalMux I__3578 (
            .O(N__19028),
            .I(N__19025));
    Odrv4 I__3577 (
            .O(N__19025),
            .I(\eeprom.n3375 ));
    InMux I__3576 (
            .O(N__19022),
            .I(N__19018));
    CascadeMux I__3575 (
            .O(N__19021),
            .I(N__19014));
    LocalMux I__3574 (
            .O(N__19018),
            .I(N__19011));
    InMux I__3573 (
            .O(N__19017),
            .I(N__19008));
    InMux I__3572 (
            .O(N__19014),
            .I(N__19005));
    Odrv4 I__3571 (
            .O(N__19011),
            .I(\eeprom.n3308 ));
    LocalMux I__3570 (
            .O(N__19008),
            .I(\eeprom.n3308 ));
    LocalMux I__3569 (
            .O(N__19005),
            .I(\eeprom.n3308 ));
    CascadeMux I__3568 (
            .O(N__18998),
            .I(\eeprom.n3407_cascade_ ));
    InMux I__3567 (
            .O(N__18995),
            .I(N__18992));
    LocalMux I__3566 (
            .O(N__18992),
            .I(\eeprom.n28_adj_484 ));
    CascadeMux I__3565 (
            .O(N__18989),
            .I(\eeprom.n27_adj_486_cascade_ ));
    InMux I__3564 (
            .O(N__18986),
            .I(N__18983));
    LocalMux I__3563 (
            .O(N__18983),
            .I(\eeprom.n26_adj_485 ));
    CascadeMux I__3562 (
            .O(N__18980),
            .I(N__18976));
    CascadeMux I__3561 (
            .O(N__18979),
            .I(N__18972));
    InMux I__3560 (
            .O(N__18976),
            .I(N__18969));
    InMux I__3559 (
            .O(N__18975),
            .I(N__18964));
    InMux I__3558 (
            .O(N__18972),
            .I(N__18964));
    LocalMux I__3557 (
            .O(N__18969),
            .I(\eeprom.n3306 ));
    LocalMux I__3556 (
            .O(N__18964),
            .I(\eeprom.n3306 ));
    CascadeMux I__3555 (
            .O(N__18959),
            .I(\eeprom.n3331_cascade_ ));
    InMux I__3554 (
            .O(N__18956),
            .I(N__18953));
    LocalMux I__3553 (
            .O(N__18953),
            .I(N__18950));
    Odrv4 I__3552 (
            .O(N__18950),
            .I(\eeprom.n3373 ));
    CascadeMux I__3551 (
            .O(N__18947),
            .I(N__18942));
    InMux I__3550 (
            .O(N__18946),
            .I(N__18937));
    InMux I__3549 (
            .O(N__18945),
            .I(N__18937));
    InMux I__3548 (
            .O(N__18942),
            .I(N__18934));
    LocalMux I__3547 (
            .O(N__18937),
            .I(\eeprom.n3305 ));
    LocalMux I__3546 (
            .O(N__18934),
            .I(\eeprom.n3305 ));
    InMux I__3545 (
            .O(N__18929),
            .I(N__18926));
    LocalMux I__3544 (
            .O(N__18926),
            .I(N__18923));
    Odrv4 I__3543 (
            .O(N__18923),
            .I(\eeprom.n3372 ));
    InMux I__3542 (
            .O(N__18920),
            .I(N__18917));
    LocalMux I__3541 (
            .O(N__18917),
            .I(N__18914));
    Odrv4 I__3540 (
            .O(N__18914),
            .I(\eeprom.n3376 ));
    CascadeMux I__3539 (
            .O(N__18911),
            .I(N__18907));
    CascadeMux I__3538 (
            .O(N__18910),
            .I(N__18903));
    InMux I__3537 (
            .O(N__18907),
            .I(N__18900));
    InMux I__3536 (
            .O(N__18906),
            .I(N__18897));
    InMux I__3535 (
            .O(N__18903),
            .I(N__18894));
    LocalMux I__3534 (
            .O(N__18900),
            .I(\eeprom.n3309 ));
    LocalMux I__3533 (
            .O(N__18897),
            .I(\eeprom.n3309 ));
    LocalMux I__3532 (
            .O(N__18894),
            .I(\eeprom.n3309 ));
    InMux I__3531 (
            .O(N__18887),
            .I(N__18884));
    LocalMux I__3530 (
            .O(N__18884),
            .I(\eeprom.n4703 ));
    CascadeMux I__3529 (
            .O(N__18881),
            .I(\eeprom.n2917_cascade_ ));
    CascadeMux I__3528 (
            .O(N__18878),
            .I(\eeprom.n4707_cascade_ ));
    InMux I__3527 (
            .O(N__18875),
            .I(N__18872));
    LocalMux I__3526 (
            .O(N__18872),
            .I(\eeprom.n15_adj_419 ));
    InMux I__3525 (
            .O(N__18869),
            .I(N__18866));
    LocalMux I__3524 (
            .O(N__18866),
            .I(\eeprom.n2875 ));
    InMux I__3523 (
            .O(N__18863),
            .I(N__18859));
    InMux I__3522 (
            .O(N__18862),
            .I(N__18856));
    LocalMux I__3521 (
            .O(N__18859),
            .I(N__18852));
    LocalMux I__3520 (
            .O(N__18856),
            .I(N__18849));
    InMux I__3519 (
            .O(N__18855),
            .I(N__18846));
    Odrv4 I__3518 (
            .O(N__18852),
            .I(\eeprom.n2808 ));
    Odrv4 I__3517 (
            .O(N__18849),
            .I(\eeprom.n2808 ));
    LocalMux I__3516 (
            .O(N__18846),
            .I(\eeprom.n2808 ));
    CascadeMux I__3515 (
            .O(N__18839),
            .I(N__18836));
    InMux I__3514 (
            .O(N__18836),
            .I(N__18833));
    LocalMux I__3513 (
            .O(N__18833),
            .I(N__18830));
    Odrv4 I__3512 (
            .O(N__18830),
            .I(\eeprom.n3385 ));
    CascadeMux I__3511 (
            .O(N__18827),
            .I(N__18824));
    InMux I__3510 (
            .O(N__18824),
            .I(N__18821));
    LocalMux I__3509 (
            .O(N__18821),
            .I(N__18818));
    Span4Mux_h I__3508 (
            .O(N__18818),
            .I(N__18815));
    Odrv4 I__3507 (
            .O(N__18815),
            .I(\eeprom.n3283 ));
    CascadeMux I__3506 (
            .O(N__18812),
            .I(\eeprom.n3315_cascade_ ));
    CascadeMux I__3505 (
            .O(N__18809),
            .I(N__18806));
    InMux I__3504 (
            .O(N__18806),
            .I(N__18801));
    InMux I__3503 (
            .O(N__18805),
            .I(N__18796));
    InMux I__3502 (
            .O(N__18804),
            .I(N__18796));
    LocalMux I__3501 (
            .O(N__18801),
            .I(\eeprom.n3318 ));
    LocalMux I__3500 (
            .O(N__18796),
            .I(\eeprom.n3318 ));
    CascadeMux I__3499 (
            .O(N__18791),
            .I(\eeprom.n4719_cascade_ ));
    InMux I__3498 (
            .O(N__18788),
            .I(N__18785));
    LocalMux I__3497 (
            .O(N__18785),
            .I(\eeprom.n4721 ));
    CascadeMux I__3496 (
            .O(N__18782),
            .I(N__18778));
    InMux I__3495 (
            .O(N__18781),
            .I(N__18774));
    InMux I__3494 (
            .O(N__18778),
            .I(N__18771));
    InMux I__3493 (
            .O(N__18777),
            .I(N__18768));
    LocalMux I__3492 (
            .O(N__18774),
            .I(\eeprom.n3304 ));
    LocalMux I__3491 (
            .O(N__18771),
            .I(\eeprom.n3304 ));
    LocalMux I__3490 (
            .O(N__18768),
            .I(\eeprom.n3304 ));
    CascadeMux I__3489 (
            .O(N__18761),
            .I(\eeprom.n4151_cascade_ ));
    InMux I__3488 (
            .O(N__18758),
            .I(N__18753));
    InMux I__3487 (
            .O(N__18757),
            .I(N__18750));
    InMux I__3486 (
            .O(N__18756),
            .I(N__18747));
    LocalMux I__3485 (
            .O(N__18753),
            .I(N__18744));
    LocalMux I__3484 (
            .O(N__18750),
            .I(N__18739));
    LocalMux I__3483 (
            .O(N__18747),
            .I(N__18739));
    Span4Mux_v I__3482 (
            .O(N__18744),
            .I(N__18736));
    Odrv4 I__3481 (
            .O(N__18739),
            .I(\eeprom.n3302 ));
    Odrv4 I__3480 (
            .O(N__18736),
            .I(\eeprom.n3302 ));
    InMux I__3479 (
            .O(N__18731),
            .I(N__18728));
    LocalMux I__3478 (
            .O(N__18728),
            .I(N__18725));
    Span4Mux_h I__3477 (
            .O(N__18725),
            .I(N__18722));
    Odrv4 I__3476 (
            .O(N__18722),
            .I(\eeprom.n4529 ));
    CascadeMux I__3475 (
            .O(N__18719),
            .I(N__18714));
    InMux I__3474 (
            .O(N__18718),
            .I(N__18709));
    InMux I__3473 (
            .O(N__18717),
            .I(N__18709));
    InMux I__3472 (
            .O(N__18714),
            .I(N__18706));
    LocalMux I__3471 (
            .O(N__18709),
            .I(N__18701));
    LocalMux I__3470 (
            .O(N__18706),
            .I(N__18701));
    Odrv4 I__3469 (
            .O(N__18701),
            .I(\eeprom.n2814 ));
    InMux I__3468 (
            .O(N__18698),
            .I(N__18695));
    LocalMux I__3467 (
            .O(N__18695),
            .I(N__18690));
    InMux I__3466 (
            .O(N__18694),
            .I(N__18687));
    InMux I__3465 (
            .O(N__18693),
            .I(N__18684));
    Span4Mux_v I__3464 (
            .O(N__18690),
            .I(N__18677));
    LocalMux I__3463 (
            .O(N__18687),
            .I(N__18677));
    LocalMux I__3462 (
            .O(N__18684),
            .I(N__18677));
    Span4Mux_h I__3461 (
            .O(N__18677),
            .I(N__18674));
    Span4Mux_h I__3460 (
            .O(N__18674),
            .I(N__18671));
    Odrv4 I__3459 (
            .O(N__18671),
            .I(\eeprom.n2819 ));
    CascadeMux I__3458 (
            .O(N__18668),
            .I(\eeprom.n4533_cascade_ ));
    InMux I__3457 (
            .O(N__18665),
            .I(N__18662));
    LocalMux I__3456 (
            .O(N__18662),
            .I(\eeprom.n20 ));
    CascadeMux I__3455 (
            .O(N__18659),
            .I(\eeprom.n15_cascade_ ));
    InMux I__3454 (
            .O(N__18656),
            .I(N__18649));
    InMux I__3453 (
            .O(N__18655),
            .I(N__18649));
    CascadeMux I__3452 (
            .O(N__18654),
            .I(N__18646));
    LocalMux I__3451 (
            .O(N__18649),
            .I(N__18643));
    InMux I__3450 (
            .O(N__18646),
            .I(N__18640));
    Span4Mux_h I__3449 (
            .O(N__18643),
            .I(N__18635));
    LocalMux I__3448 (
            .O(N__18640),
            .I(N__18635));
    Odrv4 I__3447 (
            .O(N__18635),
            .I(\eeprom.n2816 ));
    CascadeMux I__3446 (
            .O(N__18632),
            .I(\eeprom.n2836_cascade_ ));
    InMux I__3445 (
            .O(N__18629),
            .I(N__18626));
    LocalMux I__3444 (
            .O(N__18626),
            .I(\eeprom.n2883 ));
    InMux I__3443 (
            .O(N__18623),
            .I(N__18616));
    InMux I__3442 (
            .O(N__18622),
            .I(N__18616));
    InMux I__3441 (
            .O(N__18621),
            .I(N__18613));
    LocalMux I__3440 (
            .O(N__18616),
            .I(N__18610));
    LocalMux I__3439 (
            .O(N__18613),
            .I(N__18607));
    Span4Mux_h I__3438 (
            .O(N__18610),
            .I(N__18604));
    Span4Mux_h I__3437 (
            .O(N__18607),
            .I(N__18601));
    Odrv4 I__3436 (
            .O(N__18604),
            .I(\eeprom.n2809 ));
    Odrv4 I__3435 (
            .O(N__18601),
            .I(\eeprom.n2809 ));
    CascadeMux I__3434 (
            .O(N__18596),
            .I(N__18593));
    InMux I__3433 (
            .O(N__18593),
            .I(N__18590));
    LocalMux I__3432 (
            .O(N__18590),
            .I(\eeprom.n2876 ));
    InMux I__3431 (
            .O(N__18587),
            .I(N__18583));
    InMux I__3430 (
            .O(N__18586),
            .I(N__18580));
    LocalMux I__3429 (
            .O(N__18583),
            .I(N__18577));
    LocalMux I__3428 (
            .O(N__18580),
            .I(\eeprom.n2804 ));
    Odrv4 I__3427 (
            .O(N__18577),
            .I(\eeprom.n2804 ));
    InMux I__3426 (
            .O(N__18572),
            .I(N__18569));
    LocalMux I__3425 (
            .O(N__18569),
            .I(\eeprom.n2871 ));
    InMux I__3424 (
            .O(N__18566),
            .I(N__18563));
    LocalMux I__3423 (
            .O(N__18563),
            .I(\eeprom.n19 ));
    CascadeMux I__3422 (
            .O(N__18560),
            .I(\eeprom.n22_cascade_ ));
    InMux I__3421 (
            .O(N__18557),
            .I(N__18554));
    LocalMux I__3420 (
            .O(N__18554),
            .I(\eeprom.n2885 ));
    CascadeMux I__3419 (
            .O(N__18551),
            .I(N__18547));
    CascadeMux I__3418 (
            .O(N__18550),
            .I(N__18543));
    InMux I__3417 (
            .O(N__18547),
            .I(N__18540));
    InMux I__3416 (
            .O(N__18546),
            .I(N__18537));
    InMux I__3415 (
            .O(N__18543),
            .I(N__18534));
    LocalMux I__3414 (
            .O(N__18540),
            .I(N__18527));
    LocalMux I__3413 (
            .O(N__18537),
            .I(N__18527));
    LocalMux I__3412 (
            .O(N__18534),
            .I(N__18527));
    Span4Mux_v I__3411 (
            .O(N__18527),
            .I(N__18524));
    Odrv4 I__3410 (
            .O(N__18524),
            .I(\eeprom.n2818 ));
    InMux I__3409 (
            .O(N__18521),
            .I(N__18518));
    LocalMux I__3408 (
            .O(N__18518),
            .I(\eeprom.n3270 ));
    InMux I__3407 (
            .O(N__18515),
            .I(N__18512));
    LocalMux I__3406 (
            .O(N__18512),
            .I(N__18508));
    CascadeMux I__3405 (
            .O(N__18511),
            .I(N__18505));
    Span4Mux_h I__3404 (
            .O(N__18508),
            .I(N__18501));
    InMux I__3403 (
            .O(N__18505),
            .I(N__18498));
    InMux I__3402 (
            .O(N__18504),
            .I(N__18495));
    Sp12to4 I__3401 (
            .O(N__18501),
            .I(N__18490));
    LocalMux I__3400 (
            .O(N__18498),
            .I(N__18490));
    LocalMux I__3399 (
            .O(N__18495),
            .I(\eeprom.n2712 ));
    Odrv12 I__3398 (
            .O(N__18490),
            .I(\eeprom.n2712 ));
    InMux I__3397 (
            .O(N__18485),
            .I(N__18482));
    LocalMux I__3396 (
            .O(N__18482),
            .I(N__18479));
    Span4Mux_h I__3395 (
            .O(N__18479),
            .I(N__18476));
    Odrv4 I__3394 (
            .O(N__18476),
            .I(\eeprom.n2779 ));
    InMux I__3393 (
            .O(N__18473),
            .I(N__18469));
    CascadeMux I__3392 (
            .O(N__18472),
            .I(N__18466));
    LocalMux I__3391 (
            .O(N__18469),
            .I(N__18463));
    InMux I__3390 (
            .O(N__18466),
            .I(N__18460));
    Span4Mux_h I__3389 (
            .O(N__18463),
            .I(N__18454));
    LocalMux I__3388 (
            .O(N__18460),
            .I(N__18454));
    InMux I__3387 (
            .O(N__18459),
            .I(N__18451));
    Odrv4 I__3386 (
            .O(N__18454),
            .I(\eeprom.n2707 ));
    LocalMux I__3385 (
            .O(N__18451),
            .I(\eeprom.n2707 ));
    CascadeMux I__3384 (
            .O(N__18446),
            .I(N__18443));
    InMux I__3383 (
            .O(N__18443),
            .I(N__18440));
    LocalMux I__3382 (
            .O(N__18440),
            .I(N__18437));
    Odrv4 I__3381 (
            .O(N__18437),
            .I(\eeprom.n2774 ));
    InMux I__3380 (
            .O(N__18434),
            .I(N__18430));
    CascadeMux I__3379 (
            .O(N__18433),
            .I(N__18427));
    LocalMux I__3378 (
            .O(N__18430),
            .I(N__18424));
    InMux I__3377 (
            .O(N__18427),
            .I(N__18421));
    Span4Mux_h I__3376 (
            .O(N__18424),
            .I(N__18416));
    LocalMux I__3375 (
            .O(N__18421),
            .I(N__18416));
    Odrv4 I__3374 (
            .O(N__18416),
            .I(\eeprom.n2806 ));
    CascadeMux I__3373 (
            .O(N__18413),
            .I(\eeprom.n2806_cascade_ ));
    InMux I__3372 (
            .O(N__18410),
            .I(N__18406));
    InMux I__3371 (
            .O(N__18409),
            .I(N__18403));
    LocalMux I__3370 (
            .O(N__18406),
            .I(N__18397));
    LocalMux I__3369 (
            .O(N__18403),
            .I(N__18397));
    InMux I__3368 (
            .O(N__18402),
            .I(N__18394));
    Odrv4 I__3367 (
            .O(N__18397),
            .I(\eeprom.n2805 ));
    LocalMux I__3366 (
            .O(N__18394),
            .I(\eeprom.n2805 ));
    InMux I__3365 (
            .O(N__18389),
            .I(N__18386));
    LocalMux I__3364 (
            .O(N__18386),
            .I(\eeprom.n18_adj_418 ));
    InMux I__3363 (
            .O(N__18383),
            .I(N__18379));
    CascadeMux I__3362 (
            .O(N__18382),
            .I(N__18376));
    LocalMux I__3361 (
            .O(N__18379),
            .I(N__18373));
    InMux I__3360 (
            .O(N__18376),
            .I(N__18370));
    Span4Mux_v I__3359 (
            .O(N__18373),
            .I(N__18366));
    LocalMux I__3358 (
            .O(N__18370),
            .I(N__18363));
    InMux I__3357 (
            .O(N__18369),
            .I(N__18360));
    Odrv4 I__3356 (
            .O(N__18366),
            .I(\eeprom.n2708 ));
    Odrv4 I__3355 (
            .O(N__18363),
            .I(\eeprom.n2708 ));
    LocalMux I__3354 (
            .O(N__18360),
            .I(\eeprom.n2708 ));
    CascadeMux I__3353 (
            .O(N__18353),
            .I(N__18350));
    InMux I__3352 (
            .O(N__18350),
            .I(N__18347));
    LocalMux I__3351 (
            .O(N__18347),
            .I(N__18344));
    Odrv4 I__3350 (
            .O(N__18344),
            .I(\eeprom.n2775 ));
    CascadeMux I__3349 (
            .O(N__18341),
            .I(N__18333));
    CascadeMux I__3348 (
            .O(N__18340),
            .I(N__18328));
    CascadeMux I__3347 (
            .O(N__18339),
            .I(N__18323));
    CascadeMux I__3346 (
            .O(N__18338),
            .I(N__18320));
    CascadeMux I__3345 (
            .O(N__18337),
            .I(N__18316));
    InMux I__3344 (
            .O(N__18336),
            .I(N__18304));
    InMux I__3343 (
            .O(N__18333),
            .I(N__18304));
    InMux I__3342 (
            .O(N__18332),
            .I(N__18304));
    InMux I__3341 (
            .O(N__18331),
            .I(N__18304));
    InMux I__3340 (
            .O(N__18328),
            .I(N__18299));
    InMux I__3339 (
            .O(N__18327),
            .I(N__18299));
    InMux I__3338 (
            .O(N__18326),
            .I(N__18296));
    InMux I__3337 (
            .O(N__18323),
            .I(N__18285));
    InMux I__3336 (
            .O(N__18320),
            .I(N__18285));
    InMux I__3335 (
            .O(N__18319),
            .I(N__18285));
    InMux I__3334 (
            .O(N__18316),
            .I(N__18285));
    InMux I__3333 (
            .O(N__18315),
            .I(N__18285));
    CascadeMux I__3332 (
            .O(N__18314),
            .I(N__18282));
    CascadeMux I__3331 (
            .O(N__18313),
            .I(N__18279));
    LocalMux I__3330 (
            .O(N__18304),
            .I(N__18273));
    LocalMux I__3329 (
            .O(N__18299),
            .I(N__18273));
    LocalMux I__3328 (
            .O(N__18296),
            .I(N__18268));
    LocalMux I__3327 (
            .O(N__18285),
            .I(N__18268));
    InMux I__3326 (
            .O(N__18282),
            .I(N__18261));
    InMux I__3325 (
            .O(N__18279),
            .I(N__18261));
    InMux I__3324 (
            .O(N__18278),
            .I(N__18261));
    Span4Mux_h I__3323 (
            .O(N__18273),
            .I(N__18258));
    Odrv4 I__3322 (
            .O(N__18268),
            .I(\eeprom.n2737 ));
    LocalMux I__3321 (
            .O(N__18261),
            .I(\eeprom.n2737 ));
    Odrv4 I__3320 (
            .O(N__18258),
            .I(\eeprom.n2737 ));
    InMux I__3319 (
            .O(N__18251),
            .I(N__18248));
    LocalMux I__3318 (
            .O(N__18248),
            .I(N__18244));
    InMux I__3317 (
            .O(N__18247),
            .I(N__18241));
    Odrv4 I__3316 (
            .O(N__18244),
            .I(\eeprom.n2807 ));
    LocalMux I__3315 (
            .O(N__18241),
            .I(\eeprom.n2807 ));
    InMux I__3314 (
            .O(N__18236),
            .I(N__18233));
    LocalMux I__3313 (
            .O(N__18233),
            .I(N__18230));
    Odrv4 I__3312 (
            .O(N__18230),
            .I(\eeprom.n2874 ));
    CascadeMux I__3311 (
            .O(N__18227),
            .I(\eeprom.n2807_cascade_ ));
    CascadeMux I__3310 (
            .O(N__18224),
            .I(N__18221));
    InMux I__3309 (
            .O(N__18221),
            .I(N__18218));
    LocalMux I__3308 (
            .O(N__18218),
            .I(\eeprom.n2881 ));
    CascadeMux I__3307 (
            .O(N__18215),
            .I(\eeprom.n2913_cascade_ ));
    InMux I__3306 (
            .O(N__18212),
            .I(N__18209));
    LocalMux I__3305 (
            .O(N__18209),
            .I(N__18206));
    Odrv4 I__3304 (
            .O(N__18206),
            .I(\eeprom.n3269 ));
    InMux I__3303 (
            .O(N__18203),
            .I(N__18199));
    CascadeMux I__3302 (
            .O(N__18202),
            .I(N__18196));
    LocalMux I__3301 (
            .O(N__18199),
            .I(N__18193));
    InMux I__3300 (
            .O(N__18196),
            .I(N__18190));
    Span4Mux_v I__3299 (
            .O(N__18193),
            .I(N__18185));
    LocalMux I__3298 (
            .O(N__18190),
            .I(N__18185));
    Span4Mux_h I__3297 (
            .O(N__18185),
            .I(N__18182));
    Odrv4 I__3296 (
            .O(N__18182),
            .I(\eeprom.n2815 ));
    CascadeMux I__3295 (
            .O(N__18179),
            .I(N__18176));
    InMux I__3294 (
            .O(N__18176),
            .I(N__18173));
    LocalMux I__3293 (
            .O(N__18173),
            .I(N__18170));
    Odrv4 I__3292 (
            .O(N__18170),
            .I(\eeprom.n2882 ));
    InMux I__3291 (
            .O(N__18167),
            .I(N__18164));
    LocalMux I__3290 (
            .O(N__18164),
            .I(N__18161));
    Span4Mux_h I__3289 (
            .O(N__18161),
            .I(N__18158));
    Odrv4 I__3288 (
            .O(N__18158),
            .I(\eeprom.n2886 ));
    CascadeMux I__3287 (
            .O(N__18155),
            .I(\eeprom.n2918_cascade_ ));
    CascadeMux I__3286 (
            .O(N__18152),
            .I(N__18149));
    InMux I__3285 (
            .O(N__18149),
            .I(N__18146));
    LocalMux I__3284 (
            .O(N__18146),
            .I(\eeprom.n3267 ));
    InMux I__3283 (
            .O(N__18143),
            .I(N__18140));
    LocalMux I__3282 (
            .O(N__18140),
            .I(N__18136));
    InMux I__3281 (
            .O(N__18139),
            .I(N__18133));
    Span4Mux_v I__3280 (
            .O(N__18136),
            .I(N__18129));
    LocalMux I__3279 (
            .O(N__18133),
            .I(N__18126));
    InMux I__3278 (
            .O(N__18132),
            .I(N__18123));
    Odrv4 I__3277 (
            .O(N__18129),
            .I(\eeprom.n2705 ));
    Odrv12 I__3276 (
            .O(N__18126),
            .I(\eeprom.n2705 ));
    LocalMux I__3275 (
            .O(N__18123),
            .I(\eeprom.n2705 ));
    CascadeMux I__3274 (
            .O(N__18116),
            .I(N__18113));
    InMux I__3273 (
            .O(N__18113),
            .I(N__18110));
    LocalMux I__3272 (
            .O(N__18110),
            .I(N__18107));
    Span4Mux_h I__3271 (
            .O(N__18107),
            .I(N__18104));
    Odrv4 I__3270 (
            .O(N__18104),
            .I(\eeprom.n2772 ));
    CascadeMux I__3269 (
            .O(N__18101),
            .I(N__18098));
    InMux I__3268 (
            .O(N__18098),
            .I(N__18095));
    LocalMux I__3267 (
            .O(N__18095),
            .I(N__18091));
    InMux I__3266 (
            .O(N__18094),
            .I(N__18088));
    Span4Mux_h I__3265 (
            .O(N__18091),
            .I(N__18085));
    LocalMux I__3264 (
            .O(N__18088),
            .I(N__18082));
    Odrv4 I__3263 (
            .O(N__18085),
            .I(\eeprom.n2803 ));
    Odrv12 I__3262 (
            .O(N__18082),
            .I(\eeprom.n2803 ));
    CascadeMux I__3261 (
            .O(N__18077),
            .I(\eeprom.n2804_cascade_ ));
    InMux I__3260 (
            .O(N__18074),
            .I(N__18071));
    LocalMux I__3259 (
            .O(N__18071),
            .I(N__18068));
    Odrv4 I__3258 (
            .O(N__18068),
            .I(\eeprom.n3276 ));
    CascadeMux I__3257 (
            .O(N__18065),
            .I(N__18062));
    InMux I__3256 (
            .O(N__18062),
            .I(N__18059));
    LocalMux I__3255 (
            .O(N__18059),
            .I(\eeprom.n3279 ));
    InMux I__3254 (
            .O(N__18056),
            .I(N__18053));
    LocalMux I__3253 (
            .O(N__18053),
            .I(N__18050));
    Odrv4 I__3252 (
            .O(N__18050),
            .I(\eeprom.n3271 ));
    CascadeMux I__3251 (
            .O(N__18047),
            .I(N__18044));
    InMux I__3250 (
            .O(N__18044),
            .I(N__18041));
    LocalMux I__3249 (
            .O(N__18041),
            .I(N__18038));
    Odrv4 I__3248 (
            .O(N__18038),
            .I(\eeprom.n3277 ));
    InMux I__3247 (
            .O(N__18035),
            .I(N__18030));
    InMux I__3246 (
            .O(N__18034),
            .I(N__18025));
    InMux I__3245 (
            .O(N__18033),
            .I(N__18025));
    LocalMux I__3244 (
            .O(N__18030),
            .I(\eeprom.n3209 ));
    LocalMux I__3243 (
            .O(N__18025),
            .I(\eeprom.n3209 ));
    InMux I__3242 (
            .O(N__18020),
            .I(N__18017));
    LocalMux I__3241 (
            .O(N__18017),
            .I(\eeprom.n3369 ));
    InMux I__3240 (
            .O(N__18014),
            .I(N__18011));
    LocalMux I__3239 (
            .O(N__18011),
            .I(N__18008));
    Span4Mux_h I__3238 (
            .O(N__18008),
            .I(N__18005));
    Span4Mux_h I__3237 (
            .O(N__18005),
            .I(N__18002));
    Span4Mux_h I__3236 (
            .O(N__18002),
            .I(N__17999));
    Odrv4 I__3235 (
            .O(N__17999),
            .I(\eeprom.n27 ));
    InMux I__3234 (
            .O(N__17996),
            .I(N__17993));
    LocalMux I__3233 (
            .O(N__17993),
            .I(N__17990));
    Odrv4 I__3232 (
            .O(N__17990),
            .I(\eeprom.n3268 ));
    InMux I__3231 (
            .O(N__17987),
            .I(N__17984));
    LocalMux I__3230 (
            .O(N__17984),
            .I(N__17981));
    Span4Mux_v I__3229 (
            .O(N__17981),
            .I(N__17978));
    Span4Mux_h I__3228 (
            .O(N__17978),
            .I(N__17975));
    Span4Mux_h I__3227 (
            .O(N__17975),
            .I(N__17972));
    Odrv4 I__3226 (
            .O(N__17972),
            .I(\eeprom.n32_adj_480 ));
    InMux I__3225 (
            .O(N__17969),
            .I(N__17966));
    LocalMux I__3224 (
            .O(N__17966),
            .I(N__17963));
    Odrv4 I__3223 (
            .O(N__17963),
            .I(\eeprom.n3273 ));
    InMux I__3222 (
            .O(N__17960),
            .I(N__17957));
    LocalMux I__3221 (
            .O(N__17957),
            .I(N__17954));
    Odrv4 I__3220 (
            .O(N__17954),
            .I(\eeprom.n3280 ));
    CascadeMux I__3219 (
            .O(N__17951),
            .I(N__17947));
    CascadeMux I__3218 (
            .O(N__17950),
            .I(N__17944));
    InMux I__3217 (
            .O(N__17947),
            .I(N__17941));
    InMux I__3216 (
            .O(N__17944),
            .I(N__17938));
    LocalMux I__3215 (
            .O(N__17941),
            .I(\eeprom.n3312 ));
    LocalMux I__3214 (
            .O(N__17938),
            .I(\eeprom.n3312 ));
    InMux I__3213 (
            .O(N__17933),
            .I(N__17930));
    LocalMux I__3212 (
            .O(N__17930),
            .I(\eeprom.n3379 ));
    CascadeMux I__3211 (
            .O(N__17927),
            .I(\eeprom.n3312_cascade_ ));
    InMux I__3210 (
            .O(N__17924),
            .I(N__17921));
    LocalMux I__3209 (
            .O(N__17921),
            .I(N__17918));
    Odrv4 I__3208 (
            .O(N__17918),
            .I(\eeprom.n3275 ));
    CascadeMux I__3207 (
            .O(N__17915),
            .I(N__17911));
    InMux I__3206 (
            .O(N__17914),
            .I(N__17908));
    InMux I__3205 (
            .O(N__17911),
            .I(N__17905));
    LocalMux I__3204 (
            .O(N__17908),
            .I(\eeprom.n3307 ));
    LocalMux I__3203 (
            .O(N__17905),
            .I(\eeprom.n3307 ));
    InMux I__3202 (
            .O(N__17900),
            .I(N__17897));
    LocalMux I__3201 (
            .O(N__17897),
            .I(\eeprom.n3374 ));
    CascadeMux I__3200 (
            .O(N__17894),
            .I(\eeprom.n3307_cascade_ ));
    CascadeMux I__3199 (
            .O(N__17891),
            .I(\eeprom.n28_adj_482_cascade_ ));
    InMux I__3198 (
            .O(N__17888),
            .I(N__17885));
    LocalMux I__3197 (
            .O(N__17885),
            .I(N__17882));
    Odrv4 I__3196 (
            .O(N__17882),
            .I(\eeprom.n3278 ));
    CascadeMux I__3195 (
            .O(N__17879),
            .I(\eeprom.n3232_cascade_ ));
    InMux I__3194 (
            .O(N__17876),
            .I(N__17873));
    LocalMux I__3193 (
            .O(N__17873),
            .I(\eeprom.n3367 ));
    CascadeMux I__3192 (
            .O(N__17870),
            .I(\eeprom.n2904_cascade_ ));
    CascadeMux I__3191 (
            .O(N__17867),
            .I(N__17864));
    InMux I__3190 (
            .O(N__17864),
            .I(N__17861));
    LocalMux I__3189 (
            .O(N__17861),
            .I(N__17858));
    Span4Mux_h I__3188 (
            .O(N__17858),
            .I(N__17855));
    Odrv4 I__3187 (
            .O(N__17855),
            .I(\eeprom.n3286 ));
    InMux I__3186 (
            .O(N__17852),
            .I(N__17849));
    LocalMux I__3185 (
            .O(N__17849),
            .I(N__17846));
    Odrv4 I__3184 (
            .O(N__17846),
            .I(\eeprom.n3285 ));
    CascadeMux I__3183 (
            .O(N__17843),
            .I(N__17840));
    InMux I__3182 (
            .O(N__17840),
            .I(N__17837));
    LocalMux I__3181 (
            .O(N__17837),
            .I(\eeprom.n3371 ));
    InMux I__3180 (
            .O(N__17834),
            .I(N__17831));
    LocalMux I__3179 (
            .O(N__17831),
            .I(N__17828));
    Odrv4 I__3178 (
            .O(N__17828),
            .I(\eeprom.n3282 ));
    CascadeMux I__3177 (
            .O(N__17825),
            .I(\eeprom.n3314_cascade_ ));
    InMux I__3176 (
            .O(N__17822),
            .I(N__17819));
    LocalMux I__3175 (
            .O(N__17819),
            .I(N__17816));
    Span4Mux_h I__3174 (
            .O(N__17816),
            .I(N__17813));
    Odrv4 I__3173 (
            .O(N__17813),
            .I(\eeprom.n3272 ));
    InMux I__3172 (
            .O(N__17810),
            .I(N__17807));
    LocalMux I__3171 (
            .O(N__17807),
            .I(N__17804));
    Odrv4 I__3170 (
            .O(N__17804),
            .I(\eeprom.n3274 ));
    InMux I__3169 (
            .O(N__17801),
            .I(\eeprom.n3625 ));
    InMux I__3168 (
            .O(N__17798),
            .I(\eeprom.n3626 ));
    InMux I__3167 (
            .O(N__17795),
            .I(\eeprom.n3627 ));
    InMux I__3166 (
            .O(N__17792),
            .I(\eeprom.n3628 ));
    InMux I__3165 (
            .O(N__17789),
            .I(\eeprom.n3629 ));
    InMux I__3164 (
            .O(N__17786),
            .I(\eeprom.n3630 ));
    InMux I__3163 (
            .O(N__17783),
            .I(bfn_9_25_0_));
    InMux I__3162 (
            .O(N__17780),
            .I(N__17777));
    LocalMux I__3161 (
            .O(N__17777),
            .I(\eeprom.n2873 ));
    CascadeMux I__3160 (
            .O(N__17774),
            .I(N__17771));
    InMux I__3159 (
            .O(N__17771),
            .I(N__17768));
    LocalMux I__3158 (
            .O(N__17768),
            .I(\eeprom.n2872 ));
    InMux I__3157 (
            .O(N__17765),
            .I(bfn_9_23_0_));
    InMux I__3156 (
            .O(N__17762),
            .I(\eeprom.n3616 ));
    InMux I__3155 (
            .O(N__17759),
            .I(\eeprom.n3617 ));
    InMux I__3154 (
            .O(N__17756),
            .I(\eeprom.n3618 ));
    InMux I__3153 (
            .O(N__17753),
            .I(\eeprom.n3619 ));
    InMux I__3152 (
            .O(N__17750),
            .I(\eeprom.n3620 ));
    InMux I__3151 (
            .O(N__17747),
            .I(\eeprom.n3621 ));
    InMux I__3150 (
            .O(N__17744),
            .I(\eeprom.n3622 ));
    InMux I__3149 (
            .O(N__17741),
            .I(bfn_9_24_0_));
    InMux I__3148 (
            .O(N__17738),
            .I(\eeprom.n3624 ));
    InMux I__3147 (
            .O(N__17735),
            .I(\eeprom.n3700 ));
    InMux I__3146 (
            .O(N__17732),
            .I(bfn_9_22_0_));
    InMux I__3145 (
            .O(N__17729),
            .I(\eeprom.n3702 ));
    InMux I__3144 (
            .O(N__17726),
            .I(\eeprom.n3703 ));
    InMux I__3143 (
            .O(N__17723),
            .I(\eeprom.n3704 ));
    InMux I__3142 (
            .O(N__17720),
            .I(\eeprom.n3705 ));
    InMux I__3141 (
            .O(N__17717),
            .I(N__17714));
    LocalMux I__3140 (
            .O(N__17714),
            .I(N__17710));
    InMux I__3139 (
            .O(N__17713),
            .I(N__17707));
    Span4Mux_v I__3138 (
            .O(N__17710),
            .I(N__17703));
    LocalMux I__3137 (
            .O(N__17707),
            .I(N__17700));
    InMux I__3136 (
            .O(N__17706),
            .I(N__17697));
    Odrv4 I__3135 (
            .O(N__17703),
            .I(\eeprom.n2706 ));
    Odrv12 I__3134 (
            .O(N__17700),
            .I(\eeprom.n2706 ));
    LocalMux I__3133 (
            .O(N__17697),
            .I(\eeprom.n2706 ));
    InMux I__3132 (
            .O(N__17690),
            .I(N__17687));
    LocalMux I__3131 (
            .O(N__17687),
            .I(N__17684));
    Odrv4 I__3130 (
            .O(N__17684),
            .I(\eeprom.n2773 ));
    InMux I__3129 (
            .O(N__17681),
            .I(N__17677));
    CascadeMux I__3128 (
            .O(N__17680),
            .I(N__17674));
    LocalMux I__3127 (
            .O(N__17677),
            .I(N__17671));
    InMux I__3126 (
            .O(N__17674),
            .I(N__17668));
    Span4Mux_h I__3125 (
            .O(N__17671),
            .I(N__17665));
    LocalMux I__3124 (
            .O(N__17668),
            .I(N__17662));
    Odrv4 I__3123 (
            .O(N__17665),
            .I(\eeprom.n2709 ));
    Odrv4 I__3122 (
            .O(N__17662),
            .I(\eeprom.n2709 ));
    CascadeMux I__3121 (
            .O(N__17657),
            .I(N__17654));
    InMux I__3120 (
            .O(N__17654),
            .I(N__17651));
    LocalMux I__3119 (
            .O(N__17651),
            .I(N__17648));
    Odrv4 I__3118 (
            .O(N__17648),
            .I(\eeprom.n2776 ));
    InMux I__3117 (
            .O(N__17645),
            .I(\eeprom.n3690 ));
    InMux I__3116 (
            .O(N__17642),
            .I(\eeprom.n3691 ));
    InMux I__3115 (
            .O(N__17639),
            .I(\eeprom.n3692 ));
    InMux I__3114 (
            .O(N__17636),
            .I(bfn_9_21_0_));
    InMux I__3113 (
            .O(N__17633),
            .I(\eeprom.n3694 ));
    InMux I__3112 (
            .O(N__17630),
            .I(\eeprom.n3695 ));
    InMux I__3111 (
            .O(N__17627),
            .I(\eeprom.n3696 ));
    InMux I__3110 (
            .O(N__17624),
            .I(\eeprom.n3697 ));
    InMux I__3109 (
            .O(N__17621),
            .I(\eeprom.n3698 ));
    InMux I__3108 (
            .O(N__17618),
            .I(\eeprom.n3699 ));
    InMux I__3107 (
            .O(N__17615),
            .I(\eeprom.n3724 ));
    InMux I__3106 (
            .O(N__17612),
            .I(\eeprom.n3725 ));
    InMux I__3105 (
            .O(N__17609),
            .I(\eeprom.n3726 ));
    InMux I__3104 (
            .O(N__17606),
            .I(bfn_9_20_0_));
    InMux I__3103 (
            .O(N__17603),
            .I(\eeprom.n3686 ));
    InMux I__3102 (
            .O(N__17600),
            .I(\eeprom.n3687 ));
    InMux I__3101 (
            .O(N__17597),
            .I(\eeprom.n3688 ));
    InMux I__3100 (
            .O(N__17594),
            .I(\eeprom.n3689 ));
    CascadeMux I__3099 (
            .O(N__17591),
            .I(N__17588));
    InMux I__3098 (
            .O(N__17588),
            .I(N__17585));
    LocalMux I__3097 (
            .O(N__17585),
            .I(\eeprom.n3281 ));
    InMux I__3096 (
            .O(N__17582),
            .I(\eeprom.n3715 ));
    InMux I__3095 (
            .O(N__17579),
            .I(\eeprom.n3716 ));
    InMux I__3094 (
            .O(N__17576),
            .I(\eeprom.n3717 ));
    InMux I__3093 (
            .O(N__17573),
            .I(\eeprom.n3718 ));
    InMux I__3092 (
            .O(N__17570),
            .I(\eeprom.n3719 ));
    InMux I__3091 (
            .O(N__17567),
            .I(\eeprom.n3720 ));
    InMux I__3090 (
            .O(N__17564),
            .I(bfn_9_19_0_));
    InMux I__3089 (
            .O(N__17561),
            .I(\eeprom.n3722 ));
    InMux I__3088 (
            .O(N__17558),
            .I(\eeprom.n3723 ));
    InMux I__3087 (
            .O(N__17555),
            .I(\eeprom.n3706 ));
    InMux I__3086 (
            .O(N__17552),
            .I(\eeprom.n3707 ));
    InMux I__3085 (
            .O(N__17549),
            .I(\eeprom.n3708 ));
    InMux I__3084 (
            .O(N__17546),
            .I(\eeprom.n3709 ));
    InMux I__3083 (
            .O(N__17543),
            .I(\eeprom.n3710 ));
    InMux I__3082 (
            .O(N__17540),
            .I(\eeprom.n3711 ));
    InMux I__3081 (
            .O(N__17537),
            .I(\eeprom.n3712 ));
    InMux I__3080 (
            .O(N__17534),
            .I(bfn_9_18_0_));
    InMux I__3079 (
            .O(N__17531),
            .I(\eeprom.n3714 ));
    InMux I__3078 (
            .O(N__17528),
            .I(\eeprom.n3613 ));
    InMux I__3077 (
            .O(N__17525),
            .I(\eeprom.n3614 ));
    CascadeMux I__3076 (
            .O(N__17522),
            .I(N__17519));
    InMux I__3075 (
            .O(N__17519),
            .I(N__17515));
    CascadeMux I__3074 (
            .O(N__17518),
            .I(N__17512));
    LocalMux I__3073 (
            .O(N__17515),
            .I(N__17509));
    InMux I__3072 (
            .O(N__17512),
            .I(N__17506));
    Odrv4 I__3071 (
            .O(N__17509),
            .I(\eeprom.n2704 ));
    LocalMux I__3070 (
            .O(N__17506),
            .I(\eeprom.n2704 ));
    InMux I__3069 (
            .O(N__17501),
            .I(\eeprom.n3615 ));
    InMux I__3068 (
            .O(N__17498),
            .I(N__17495));
    LocalMux I__3067 (
            .O(N__17495),
            .I(\eeprom.n2777 ));
    CascadeMux I__3066 (
            .O(N__17492),
            .I(N__17488));
    InMux I__3065 (
            .O(N__17491),
            .I(N__17484));
    InMux I__3064 (
            .O(N__17488),
            .I(N__17481));
    InMux I__3063 (
            .O(N__17487),
            .I(N__17478));
    LocalMux I__3062 (
            .O(N__17484),
            .I(N__17473));
    LocalMux I__3061 (
            .O(N__17481),
            .I(N__17473));
    LocalMux I__3060 (
            .O(N__17478),
            .I(N__17470));
    Odrv4 I__3059 (
            .O(N__17473),
            .I(\eeprom.n2710 ));
    Odrv4 I__3058 (
            .O(N__17470),
            .I(\eeprom.n2710 ));
    InMux I__3057 (
            .O(N__17465),
            .I(N__17462));
    LocalMux I__3056 (
            .O(N__17462),
            .I(\eeprom.n2778 ));
    InMux I__3055 (
            .O(N__17459),
            .I(N__17454));
    InMux I__3054 (
            .O(N__17458),
            .I(N__17451));
    InMux I__3053 (
            .O(N__17457),
            .I(N__17448));
    LocalMux I__3052 (
            .O(N__17454),
            .I(N__17441));
    LocalMux I__3051 (
            .O(N__17451),
            .I(N__17441));
    LocalMux I__3050 (
            .O(N__17448),
            .I(N__17441));
    Odrv12 I__3049 (
            .O(N__17441),
            .I(\eeprom.n2711 ));
    InMux I__3048 (
            .O(N__17438),
            .I(N__17434));
    CascadeMux I__3047 (
            .O(N__17437),
            .I(N__17431));
    LocalMux I__3046 (
            .O(N__17434),
            .I(N__17427));
    InMux I__3045 (
            .O(N__17431),
            .I(N__17424));
    InMux I__3044 (
            .O(N__17430),
            .I(N__17421));
    Span4Mux_v I__3043 (
            .O(N__17427),
            .I(N__17416));
    LocalMux I__3042 (
            .O(N__17424),
            .I(N__17416));
    LocalMux I__3041 (
            .O(N__17421),
            .I(\eeprom.n2717 ));
    Odrv4 I__3040 (
            .O(N__17416),
            .I(\eeprom.n2717 ));
    CascadeMux I__3039 (
            .O(N__17411),
            .I(N__17408));
    InMux I__3038 (
            .O(N__17408),
            .I(N__17405));
    LocalMux I__3037 (
            .O(N__17405),
            .I(N__17402));
    Odrv4 I__3036 (
            .O(N__17402),
            .I(\eeprom.n2784 ));
    InMux I__3035 (
            .O(N__17399),
            .I(N__17396));
    LocalMux I__3034 (
            .O(N__17396),
            .I(N__17393));
    Odrv4 I__3033 (
            .O(N__17393),
            .I(\eeprom.n2782 ));
    InMux I__3032 (
            .O(N__17390),
            .I(N__17386));
    CascadeMux I__3031 (
            .O(N__17389),
            .I(N__17383));
    LocalMux I__3030 (
            .O(N__17386),
            .I(N__17380));
    InMux I__3029 (
            .O(N__17383),
            .I(N__17377));
    Span4Mux_v I__3028 (
            .O(N__17380),
            .I(N__17371));
    LocalMux I__3027 (
            .O(N__17377),
            .I(N__17371));
    InMux I__3026 (
            .O(N__17376),
            .I(N__17368));
    Odrv4 I__3025 (
            .O(N__17371),
            .I(\eeprom.n2715 ));
    LocalMux I__3024 (
            .O(N__17368),
            .I(\eeprom.n2715 ));
    InMux I__3023 (
            .O(N__17363),
            .I(N__17359));
    CascadeMux I__3022 (
            .O(N__17362),
            .I(N__17356));
    LocalMux I__3021 (
            .O(N__17359),
            .I(N__17353));
    InMux I__3020 (
            .O(N__17356),
            .I(N__17350));
    Span4Mux_v I__3019 (
            .O(N__17353),
            .I(N__17345));
    LocalMux I__3018 (
            .O(N__17350),
            .I(N__17345));
    Odrv4 I__3017 (
            .O(N__17345),
            .I(\eeprom.n2713 ));
    CascadeMux I__3016 (
            .O(N__17342),
            .I(N__17339));
    InMux I__3015 (
            .O(N__17339),
            .I(N__17336));
    LocalMux I__3014 (
            .O(N__17336),
            .I(N__17333));
    Odrv4 I__3013 (
            .O(N__17333),
            .I(\eeprom.n2780 ));
    InMux I__3012 (
            .O(N__17330),
            .I(bfn_9_17_0_));
    CascadeMux I__3011 (
            .O(N__17327),
            .I(N__17324));
    InMux I__3010 (
            .O(N__17324),
            .I(N__17320));
    InMux I__3009 (
            .O(N__17323),
            .I(N__17316));
    LocalMux I__3008 (
            .O(N__17320),
            .I(N__17313));
    InMux I__3007 (
            .O(N__17319),
            .I(N__17310));
    LocalMux I__3006 (
            .O(N__17316),
            .I(\eeprom.n2714 ));
    Odrv4 I__3005 (
            .O(N__17313),
            .I(\eeprom.n2714 ));
    LocalMux I__3004 (
            .O(N__17310),
            .I(\eeprom.n2714 ));
    InMux I__3003 (
            .O(N__17303),
            .I(N__17300));
    LocalMux I__3002 (
            .O(N__17300),
            .I(\eeprom.n2781 ));
    InMux I__3001 (
            .O(N__17297),
            .I(\eeprom.n3605 ));
    InMux I__3000 (
            .O(N__17294),
            .I(\eeprom.n3606 ));
    InMux I__2999 (
            .O(N__17291),
            .I(\eeprom.n3607 ));
    InMux I__2998 (
            .O(N__17288),
            .I(bfn_7_22_0_));
    InMux I__2997 (
            .O(N__17285),
            .I(\eeprom.n3609 ));
    InMux I__2996 (
            .O(N__17282),
            .I(\eeprom.n3610 ));
    InMux I__2995 (
            .O(N__17279),
            .I(\eeprom.n3611 ));
    InMux I__2994 (
            .O(N__17276),
            .I(\eeprom.n3612 ));
    InMux I__2993 (
            .O(N__17273),
            .I(N__17270));
    LocalMux I__2992 (
            .O(N__17270),
            .I(N__17267));
    Span4Mux_v I__2991 (
            .O(N__17267),
            .I(N__17264));
    Span4Mux_h I__2990 (
            .O(N__17264),
            .I(N__17261));
    Odrv4 I__2989 (
            .O(N__17261),
            .I(\eeprom.n28 ));
    InMux I__2988 (
            .O(N__17258),
            .I(N__17255));
    LocalMux I__2987 (
            .O(N__17255),
            .I(N__17251));
    InMux I__2986 (
            .O(N__17254),
            .I(N__17248));
    Span4Mux_h I__2985 (
            .O(N__17251),
            .I(N__17244));
    LocalMux I__2984 (
            .O(N__17248),
            .I(N__17241));
    InMux I__2983 (
            .O(N__17247),
            .I(N__17238));
    Odrv4 I__2982 (
            .O(N__17244),
            .I(\eeprom.n2610 ));
    Odrv12 I__2981 (
            .O(N__17241),
            .I(\eeprom.n2610 ));
    LocalMux I__2980 (
            .O(N__17238),
            .I(\eeprom.n2610 ));
    CascadeMux I__2979 (
            .O(N__17231),
            .I(N__17228));
    InMux I__2978 (
            .O(N__17228),
            .I(N__17225));
    LocalMux I__2977 (
            .O(N__17225),
            .I(\eeprom.n2677 ));
    InMux I__2976 (
            .O(N__17222),
            .I(N__17214));
    CascadeMux I__2975 (
            .O(N__17221),
            .I(N__17207));
    CascadeMux I__2974 (
            .O(N__17220),
            .I(N__17204));
    CascadeMux I__2973 (
            .O(N__17219),
            .I(N__17199));
    CascadeMux I__2972 (
            .O(N__17218),
            .I(N__17195));
    InMux I__2971 (
            .O(N__17217),
            .I(N__17191));
    LocalMux I__2970 (
            .O(N__17214),
            .I(N__17188));
    InMux I__2969 (
            .O(N__17213),
            .I(N__17185));
    InMux I__2968 (
            .O(N__17212),
            .I(N__17180));
    InMux I__2967 (
            .O(N__17211),
            .I(N__17180));
    InMux I__2966 (
            .O(N__17210),
            .I(N__17171));
    InMux I__2965 (
            .O(N__17207),
            .I(N__17171));
    InMux I__2964 (
            .O(N__17204),
            .I(N__17171));
    InMux I__2963 (
            .O(N__17203),
            .I(N__17171));
    InMux I__2962 (
            .O(N__17202),
            .I(N__17160));
    InMux I__2961 (
            .O(N__17199),
            .I(N__17160));
    InMux I__2960 (
            .O(N__17198),
            .I(N__17160));
    InMux I__2959 (
            .O(N__17195),
            .I(N__17160));
    InMux I__2958 (
            .O(N__17194),
            .I(N__17160));
    LocalMux I__2957 (
            .O(N__17191),
            .I(\eeprom.n2638 ));
    Odrv4 I__2956 (
            .O(N__17188),
            .I(\eeprom.n2638 ));
    LocalMux I__2955 (
            .O(N__17185),
            .I(\eeprom.n2638 ));
    LocalMux I__2954 (
            .O(N__17180),
            .I(\eeprom.n2638 ));
    LocalMux I__2953 (
            .O(N__17171),
            .I(\eeprom.n2638 ));
    LocalMux I__2952 (
            .O(N__17160),
            .I(\eeprom.n2638 ));
    InMux I__2951 (
            .O(N__17147),
            .I(N__17144));
    LocalMux I__2950 (
            .O(N__17144),
            .I(N__17141));
    Odrv4 I__2949 (
            .O(N__17141),
            .I(\eeprom.n18 ));
    CascadeMux I__2948 (
            .O(N__17138),
            .I(\eeprom.n2709_cascade_ ));
    InMux I__2947 (
            .O(N__17135),
            .I(N__17132));
    LocalMux I__2946 (
            .O(N__17132),
            .I(\eeprom.n13_adj_417 ));
    CascadeMux I__2945 (
            .O(N__17129),
            .I(\eeprom.n2737_cascade_ ));
    InMux I__2944 (
            .O(N__17126),
            .I(N__17123));
    LocalMux I__2943 (
            .O(N__17123),
            .I(N__17118));
    InMux I__2942 (
            .O(N__17122),
            .I(N__17115));
    InMux I__2941 (
            .O(N__17121),
            .I(N__17112));
    Span4Mux_h I__2940 (
            .O(N__17118),
            .I(N__17109));
    LocalMux I__2939 (
            .O(N__17115),
            .I(N__17104));
    LocalMux I__2938 (
            .O(N__17112),
            .I(N__17104));
    Span4Mux_h I__2937 (
            .O(N__17109),
            .I(N__17101));
    Span12Mux_v I__2936 (
            .O(N__17104),
            .I(N__17098));
    Odrv4 I__2935 (
            .O(N__17101),
            .I(\eeprom.n2719 ));
    Odrv12 I__2934 (
            .O(N__17098),
            .I(\eeprom.n2719 ));
    InMux I__2933 (
            .O(N__17093),
            .I(N__17090));
    LocalMux I__2932 (
            .O(N__17090),
            .I(\eeprom.n2786 ));
    InMux I__2931 (
            .O(N__17087),
            .I(bfn_7_21_0_));
    CascadeMux I__2930 (
            .O(N__17084),
            .I(N__17081));
    InMux I__2929 (
            .O(N__17081),
            .I(N__17077));
    InMux I__2928 (
            .O(N__17080),
            .I(N__17074));
    LocalMux I__2927 (
            .O(N__17077),
            .I(N__17071));
    LocalMux I__2926 (
            .O(N__17074),
            .I(\eeprom.n2718 ));
    Odrv4 I__2925 (
            .O(N__17071),
            .I(\eeprom.n2718 ));
    InMux I__2924 (
            .O(N__17066),
            .I(N__17063));
    LocalMux I__2923 (
            .O(N__17063),
            .I(\eeprom.n2785 ));
    InMux I__2922 (
            .O(N__17060),
            .I(\eeprom.n3601 ));
    InMux I__2921 (
            .O(N__17057),
            .I(\eeprom.n3602 ));
    CascadeMux I__2920 (
            .O(N__17054),
            .I(N__17051));
    InMux I__2919 (
            .O(N__17051),
            .I(N__17047));
    InMux I__2918 (
            .O(N__17050),
            .I(N__17043));
    LocalMux I__2917 (
            .O(N__17047),
            .I(N__17040));
    InMux I__2916 (
            .O(N__17046),
            .I(N__17037));
    LocalMux I__2915 (
            .O(N__17043),
            .I(\eeprom.n2716 ));
    Odrv4 I__2914 (
            .O(N__17040),
            .I(\eeprom.n2716 ));
    LocalMux I__2913 (
            .O(N__17037),
            .I(\eeprom.n2716 ));
    InMux I__2912 (
            .O(N__17030),
            .I(N__17027));
    LocalMux I__2911 (
            .O(N__17027),
            .I(\eeprom.n2783 ));
    InMux I__2910 (
            .O(N__17024),
            .I(\eeprom.n3603 ));
    InMux I__2909 (
            .O(N__17021),
            .I(\eeprom.n3604 ));
    CascadeMux I__2908 (
            .O(N__17018),
            .I(N__17015));
    InMux I__2907 (
            .O(N__17015),
            .I(N__17012));
    LocalMux I__2906 (
            .O(N__17012),
            .I(\eeprom.n2675 ));
    InMux I__2905 (
            .O(N__17009),
            .I(N__17006));
    LocalMux I__2904 (
            .O(N__17006),
            .I(\eeprom.n2682 ));
    InMux I__2903 (
            .O(N__17003),
            .I(N__16999));
    CascadeMux I__2902 (
            .O(N__17002),
            .I(N__16996));
    LocalMux I__2901 (
            .O(N__16999),
            .I(N__16993));
    InMux I__2900 (
            .O(N__16996),
            .I(N__16990));
    Odrv12 I__2899 (
            .O(N__16993),
            .I(\eeprom.n2615 ));
    LocalMux I__2898 (
            .O(N__16990),
            .I(\eeprom.n2615 ));
    CascadeMux I__2897 (
            .O(N__16985),
            .I(N__16982));
    InMux I__2896 (
            .O(N__16982),
            .I(N__16977));
    InMux I__2895 (
            .O(N__16981),
            .I(N__16972));
    InMux I__2894 (
            .O(N__16980),
            .I(N__16972));
    LocalMux I__2893 (
            .O(N__16977),
            .I(\eeprom.n2608 ));
    LocalMux I__2892 (
            .O(N__16972),
            .I(\eeprom.n2608 ));
    InMux I__2891 (
            .O(N__16967),
            .I(N__16964));
    LocalMux I__2890 (
            .O(N__16964),
            .I(N__16961));
    Odrv4 I__2889 (
            .O(N__16961),
            .I(\eeprom.n12 ));
    CascadeMux I__2888 (
            .O(N__16958),
            .I(N__16954));
    CascadeMux I__2887 (
            .O(N__16957),
            .I(N__16950));
    InMux I__2886 (
            .O(N__16954),
            .I(N__16947));
    InMux I__2885 (
            .O(N__16953),
            .I(N__16942));
    InMux I__2884 (
            .O(N__16950),
            .I(N__16942));
    LocalMux I__2883 (
            .O(N__16947),
            .I(\eeprom.n2607 ));
    LocalMux I__2882 (
            .O(N__16942),
            .I(\eeprom.n2607 ));
    InMux I__2881 (
            .O(N__16937),
            .I(N__16934));
    LocalMux I__2880 (
            .O(N__16934),
            .I(N__16931));
    Span4Mux_v I__2879 (
            .O(N__16931),
            .I(N__16928));
    Odrv4 I__2878 (
            .O(N__16928),
            .I(\eeprom.n16 ));
    InMux I__2877 (
            .O(N__16925),
            .I(N__16922));
    LocalMux I__2876 (
            .O(N__16922),
            .I(\eeprom.n2683 ));
    CascadeMux I__2875 (
            .O(N__16919),
            .I(\eeprom.n2638_cascade_ ));
    InMux I__2874 (
            .O(N__16916),
            .I(N__16912));
    CascadeMux I__2873 (
            .O(N__16915),
            .I(N__16909));
    LocalMux I__2872 (
            .O(N__16912),
            .I(N__16905));
    InMux I__2871 (
            .O(N__16909),
            .I(N__16902));
    InMux I__2870 (
            .O(N__16908),
            .I(N__16899));
    Odrv4 I__2869 (
            .O(N__16905),
            .I(\eeprom.n2616 ));
    LocalMux I__2868 (
            .O(N__16902),
            .I(\eeprom.n2616 ));
    LocalMux I__2867 (
            .O(N__16899),
            .I(\eeprom.n2616 ));
    InMux I__2866 (
            .O(N__16892),
            .I(N__16888));
    CascadeMux I__2865 (
            .O(N__16891),
            .I(N__16885));
    LocalMux I__2864 (
            .O(N__16888),
            .I(N__16881));
    InMux I__2863 (
            .O(N__16885),
            .I(N__16878));
    InMux I__2862 (
            .O(N__16884),
            .I(N__16875));
    Odrv4 I__2861 (
            .O(N__16881),
            .I(\eeprom.n2617 ));
    LocalMux I__2860 (
            .O(N__16878),
            .I(\eeprom.n2617 ));
    LocalMux I__2859 (
            .O(N__16875),
            .I(\eeprom.n2617 ));
    CascadeMux I__2858 (
            .O(N__16868),
            .I(N__16865));
    InMux I__2857 (
            .O(N__16865),
            .I(N__16862));
    LocalMux I__2856 (
            .O(N__16862),
            .I(\eeprom.n2684 ));
    CascadeMux I__2855 (
            .O(N__16859),
            .I(\eeprom.n2815_cascade_ ));
    InMux I__2854 (
            .O(N__16856),
            .I(N__16852));
    CascadeMux I__2853 (
            .O(N__16855),
            .I(N__16849));
    LocalMux I__2852 (
            .O(N__16852),
            .I(N__16846));
    InMux I__2851 (
            .O(N__16849),
            .I(N__16843));
    Span4Mux_h I__2850 (
            .O(N__16846),
            .I(N__16839));
    LocalMux I__2849 (
            .O(N__16843),
            .I(N__16836));
    InMux I__2848 (
            .O(N__16842),
            .I(N__16833));
    Odrv4 I__2847 (
            .O(N__16839),
            .I(\eeprom.n2614 ));
    Odrv4 I__2846 (
            .O(N__16836),
            .I(\eeprom.n2614 ));
    LocalMux I__2845 (
            .O(N__16833),
            .I(\eeprom.n2614 ));
    InMux I__2844 (
            .O(N__16826),
            .I(N__16823));
    LocalMux I__2843 (
            .O(N__16823),
            .I(\eeprom.n2681 ));
    CascadeMux I__2842 (
            .O(N__16820),
            .I(\eeprom.n2713_cascade_ ));
    CascadeMux I__2841 (
            .O(N__16817),
            .I(\eeprom.n4695_cascade_ ));
    CascadeMux I__2840 (
            .O(N__16814),
            .I(\eeprom.n16_adj_416_cascade_ ));
    CascadeMux I__2839 (
            .O(N__16811),
            .I(N__16806));
    InMux I__2838 (
            .O(N__16810),
            .I(N__16803));
    InMux I__2837 (
            .O(N__16809),
            .I(N__16800));
    InMux I__2836 (
            .O(N__16806),
            .I(N__16797));
    LocalMux I__2835 (
            .O(N__16803),
            .I(\eeprom.n2618 ));
    LocalMux I__2834 (
            .O(N__16800),
            .I(\eeprom.n2618 ));
    LocalMux I__2833 (
            .O(N__16797),
            .I(\eeprom.n2618 ));
    CascadeMux I__2832 (
            .O(N__16790),
            .I(N__16787));
    InMux I__2831 (
            .O(N__16787),
            .I(N__16784));
    LocalMux I__2830 (
            .O(N__16784),
            .I(\eeprom.n2685 ));
    InMux I__2829 (
            .O(N__16781),
            .I(N__16778));
    LocalMux I__2828 (
            .O(N__16778),
            .I(\eeprom.n2674 ));
    InMux I__2827 (
            .O(N__16775),
            .I(N__16772));
    LocalMux I__2826 (
            .O(N__16772),
            .I(N__16769));
    Span4Mux_h I__2825 (
            .O(N__16769),
            .I(N__16766));
    Odrv4 I__2824 (
            .O(N__16766),
            .I(\eeprom.n2686 ));
    InMux I__2823 (
            .O(N__16763),
            .I(N__16758));
    InMux I__2822 (
            .O(N__16762),
            .I(N__16755));
    InMux I__2821 (
            .O(N__16761),
            .I(N__16752));
    LocalMux I__2820 (
            .O(N__16758),
            .I(N__16747));
    LocalMux I__2819 (
            .O(N__16755),
            .I(N__16747));
    LocalMux I__2818 (
            .O(N__16752),
            .I(N__16744));
    Span4Mux_h I__2817 (
            .O(N__16747),
            .I(N__16741));
    Odrv4 I__2816 (
            .O(N__16744),
            .I(\eeprom.n2619 ));
    Odrv4 I__2815 (
            .O(N__16741),
            .I(\eeprom.n2619 ));
    CascadeMux I__2814 (
            .O(N__16736),
            .I(\eeprom.n2718_cascade_ ));
    InMux I__2813 (
            .O(N__16733),
            .I(N__16730));
    LocalMux I__2812 (
            .O(N__16730),
            .I(\eeprom.n4699 ));
    CascadeMux I__2811 (
            .O(N__16727),
            .I(N__16724));
    InMux I__2810 (
            .O(N__16724),
            .I(N__16721));
    LocalMux I__2809 (
            .O(N__16721),
            .I(N__16718));
    Span4Mux_h I__2808 (
            .O(N__16718),
            .I(N__16715));
    Odrv4 I__2807 (
            .O(N__16715),
            .I(\eeprom.n2280 ));
    InMux I__2806 (
            .O(N__16712),
            .I(\eeprom.n3546 ));
    CascadeMux I__2805 (
            .O(N__16709),
            .I(N__16704));
    InMux I__2804 (
            .O(N__16708),
            .I(N__16701));
    InMux I__2803 (
            .O(N__16707),
            .I(N__16698));
    InMux I__2802 (
            .O(N__16704),
            .I(N__16695));
    LocalMux I__2801 (
            .O(N__16701),
            .I(N__16692));
    LocalMux I__2800 (
            .O(N__16698),
            .I(\eeprom.n2212 ));
    LocalMux I__2799 (
            .O(N__16695),
            .I(\eeprom.n2212 ));
    Odrv4 I__2798 (
            .O(N__16692),
            .I(\eeprom.n2212 ));
    InMux I__2797 (
            .O(N__16685),
            .I(N__16682));
    LocalMux I__2796 (
            .O(N__16682),
            .I(\eeprom.n2279 ));
    InMux I__2795 (
            .O(N__16679),
            .I(\eeprom.n3547 ));
    CascadeMux I__2794 (
            .O(N__16676),
            .I(N__16671));
    InMux I__2793 (
            .O(N__16675),
            .I(N__16666));
    InMux I__2792 (
            .O(N__16674),
            .I(N__16666));
    InMux I__2791 (
            .O(N__16671),
            .I(N__16663));
    LocalMux I__2790 (
            .O(N__16666),
            .I(N__16660));
    LocalMux I__2789 (
            .O(N__16663),
            .I(\eeprom.n2211 ));
    Odrv4 I__2788 (
            .O(N__16660),
            .I(\eeprom.n2211 ));
    CascadeMux I__2787 (
            .O(N__16655),
            .I(N__16652));
    InMux I__2786 (
            .O(N__16652),
            .I(N__16649));
    LocalMux I__2785 (
            .O(N__16649),
            .I(N__16646));
    Span4Mux_h I__2784 (
            .O(N__16646),
            .I(N__16643));
    Odrv4 I__2783 (
            .O(N__16643),
            .I(\eeprom.n2278 ));
    InMux I__2782 (
            .O(N__16640),
            .I(bfn_6_27_0_));
    InMux I__2781 (
            .O(N__16637),
            .I(N__16633));
    CascadeMux I__2780 (
            .O(N__16636),
            .I(N__16630));
    LocalMux I__2779 (
            .O(N__16633),
            .I(N__16626));
    InMux I__2778 (
            .O(N__16630),
            .I(N__16621));
    InMux I__2777 (
            .O(N__16629),
            .I(N__16621));
    Odrv4 I__2776 (
            .O(N__16626),
            .I(\eeprom.n2210 ));
    LocalMux I__2775 (
            .O(N__16621),
            .I(\eeprom.n2210 ));
    InMux I__2774 (
            .O(N__16616),
            .I(N__16613));
    LocalMux I__2773 (
            .O(N__16613),
            .I(N__16610));
    Odrv4 I__2772 (
            .O(N__16610),
            .I(\eeprom.n2277 ));
    InMux I__2771 (
            .O(N__16607),
            .I(\eeprom.n3549 ));
    InMux I__2770 (
            .O(N__16604),
            .I(N__16594));
    InMux I__2769 (
            .O(N__16603),
            .I(N__16588));
    InMux I__2768 (
            .O(N__16602),
            .I(N__16583));
    InMux I__2767 (
            .O(N__16601),
            .I(N__16583));
    InMux I__2766 (
            .O(N__16600),
            .I(N__16580));
    InMux I__2765 (
            .O(N__16599),
            .I(N__16575));
    InMux I__2764 (
            .O(N__16598),
            .I(N__16575));
    InMux I__2763 (
            .O(N__16597),
            .I(N__16572));
    LocalMux I__2762 (
            .O(N__16594),
            .I(N__16569));
    InMux I__2761 (
            .O(N__16593),
            .I(N__16562));
    InMux I__2760 (
            .O(N__16592),
            .I(N__16562));
    InMux I__2759 (
            .O(N__16591),
            .I(N__16562));
    LocalMux I__2758 (
            .O(N__16588),
            .I(\eeprom.n2242 ));
    LocalMux I__2757 (
            .O(N__16583),
            .I(\eeprom.n2242 ));
    LocalMux I__2756 (
            .O(N__16580),
            .I(\eeprom.n2242 ));
    LocalMux I__2755 (
            .O(N__16575),
            .I(\eeprom.n2242 ));
    LocalMux I__2754 (
            .O(N__16572),
            .I(\eeprom.n2242 ));
    Odrv4 I__2753 (
            .O(N__16569),
            .I(\eeprom.n2242 ));
    LocalMux I__2752 (
            .O(N__16562),
            .I(\eeprom.n2242 ));
    InMux I__2751 (
            .O(N__16547),
            .I(N__16543));
    CascadeMux I__2750 (
            .O(N__16546),
            .I(N__16540));
    LocalMux I__2749 (
            .O(N__16543),
            .I(N__16537));
    InMux I__2748 (
            .O(N__16540),
            .I(N__16534));
    Span4Mux_h I__2747 (
            .O(N__16537),
            .I(N__16531));
    LocalMux I__2746 (
            .O(N__16534),
            .I(\eeprom.n2209 ));
    Odrv4 I__2745 (
            .O(N__16531),
            .I(\eeprom.n2209 ));
    InMux I__2744 (
            .O(N__16526),
            .I(\eeprom.n3550 ));
    InMux I__2743 (
            .O(N__16523),
            .I(N__16519));
    InMux I__2742 (
            .O(N__16522),
            .I(N__16516));
    LocalMux I__2741 (
            .O(N__16519),
            .I(N__16513));
    LocalMux I__2740 (
            .O(N__16516),
            .I(N__16510));
    Span4Mux_h I__2739 (
            .O(N__16513),
            .I(N__16507));
    Span4Mux_h I__2738 (
            .O(N__16510),
            .I(N__16504));
    Odrv4 I__2737 (
            .O(N__16507),
            .I(\eeprom.n2308 ));
    Odrv4 I__2736 (
            .O(N__16504),
            .I(\eeprom.n2308 ));
    InMux I__2735 (
            .O(N__16499),
            .I(N__16495));
    CascadeMux I__2734 (
            .O(N__16498),
            .I(N__16492));
    LocalMux I__2733 (
            .O(N__16495),
            .I(N__16489));
    InMux I__2732 (
            .O(N__16492),
            .I(N__16486));
    Span4Mux_v I__2731 (
            .O(N__16489),
            .I(N__16482));
    LocalMux I__2730 (
            .O(N__16486),
            .I(N__16479));
    InMux I__2729 (
            .O(N__16485),
            .I(N__16476));
    Odrv4 I__2728 (
            .O(N__16482),
            .I(\eeprom.n2612 ));
    Odrv12 I__2727 (
            .O(N__16479),
            .I(\eeprom.n2612 ));
    LocalMux I__2726 (
            .O(N__16476),
            .I(\eeprom.n2612 ));
    CascadeMux I__2725 (
            .O(N__16469),
            .I(N__16466));
    InMux I__2724 (
            .O(N__16466),
            .I(N__16463));
    LocalMux I__2723 (
            .O(N__16463),
            .I(\eeprom.n2679 ));
    InMux I__2722 (
            .O(N__16460),
            .I(N__16457));
    LocalMux I__2721 (
            .O(N__16457),
            .I(N__16453));
    InMux I__2720 (
            .O(N__16456),
            .I(N__16450));
    Span4Mux_v I__2719 (
            .O(N__16453),
            .I(N__16447));
    LocalMux I__2718 (
            .O(N__16450),
            .I(N__16444));
    Odrv4 I__2717 (
            .O(N__16447),
            .I(\eeprom.n2606 ));
    Odrv12 I__2716 (
            .O(N__16444),
            .I(\eeprom.n2606 ));
    InMux I__2715 (
            .O(N__16439),
            .I(N__16436));
    LocalMux I__2714 (
            .O(N__16436),
            .I(\eeprom.n2673 ));
    InMux I__2713 (
            .O(N__16433),
            .I(N__16430));
    LocalMux I__2712 (
            .O(N__16430),
            .I(\eeprom.n2680 ));
    InMux I__2711 (
            .O(N__16427),
            .I(N__16423));
    CascadeMux I__2710 (
            .O(N__16426),
            .I(N__16420));
    LocalMux I__2709 (
            .O(N__16423),
            .I(N__16417));
    InMux I__2708 (
            .O(N__16420),
            .I(N__16414));
    Span4Mux_v I__2707 (
            .O(N__16417),
            .I(N__16410));
    LocalMux I__2706 (
            .O(N__16414),
            .I(N__16407));
    InMux I__2705 (
            .O(N__16413),
            .I(N__16404));
    Odrv4 I__2704 (
            .O(N__16410),
            .I(\eeprom.n2613 ));
    Odrv4 I__2703 (
            .O(N__16407),
            .I(\eeprom.n2613 ));
    LocalMux I__2702 (
            .O(N__16404),
            .I(\eeprom.n2613 ));
    CascadeMux I__2701 (
            .O(N__16397),
            .I(N__16393));
    InMux I__2700 (
            .O(N__16396),
            .I(N__16390));
    InMux I__2699 (
            .O(N__16393),
            .I(N__16387));
    LocalMux I__2698 (
            .O(N__16390),
            .I(N__16383));
    LocalMux I__2697 (
            .O(N__16387),
            .I(N__16380));
    InMux I__2696 (
            .O(N__16386),
            .I(N__16377));
    Odrv4 I__2695 (
            .O(N__16383),
            .I(\eeprom.n2113 ));
    Odrv12 I__2694 (
            .O(N__16380),
            .I(\eeprom.n2113 ));
    LocalMux I__2693 (
            .O(N__16377),
            .I(\eeprom.n2113 ));
    CascadeMux I__2692 (
            .O(N__16370),
            .I(N__16361));
    InMux I__2691 (
            .O(N__16369),
            .I(N__16358));
    CascadeMux I__2690 (
            .O(N__16368),
            .I(N__16355));
    CascadeMux I__2689 (
            .O(N__16367),
            .I(N__16350));
    CascadeMux I__2688 (
            .O(N__16366),
            .I(N__16347));
    CascadeMux I__2687 (
            .O(N__16365),
            .I(N__16343));
    CascadeMux I__2686 (
            .O(N__16364),
            .I(N__16340));
    InMux I__2685 (
            .O(N__16361),
            .I(N__16336));
    LocalMux I__2684 (
            .O(N__16358),
            .I(N__16333));
    InMux I__2683 (
            .O(N__16355),
            .I(N__16328));
    InMux I__2682 (
            .O(N__16354),
            .I(N__16328));
    InMux I__2681 (
            .O(N__16353),
            .I(N__16319));
    InMux I__2680 (
            .O(N__16350),
            .I(N__16319));
    InMux I__2679 (
            .O(N__16347),
            .I(N__16319));
    InMux I__2678 (
            .O(N__16346),
            .I(N__16319));
    InMux I__2677 (
            .O(N__16343),
            .I(N__16312));
    InMux I__2676 (
            .O(N__16340),
            .I(N__16312));
    InMux I__2675 (
            .O(N__16339),
            .I(N__16312));
    LocalMux I__2674 (
            .O(N__16336),
            .I(N__16309));
    Odrv4 I__2673 (
            .O(N__16333),
            .I(\eeprom.n2143 ));
    LocalMux I__2672 (
            .O(N__16328),
            .I(\eeprom.n2143 ));
    LocalMux I__2671 (
            .O(N__16319),
            .I(\eeprom.n2143 ));
    LocalMux I__2670 (
            .O(N__16312),
            .I(\eeprom.n2143 ));
    Odrv4 I__2669 (
            .O(N__16309),
            .I(\eeprom.n2143 ));
    InMux I__2668 (
            .O(N__16298),
            .I(N__16295));
    LocalMux I__2667 (
            .O(N__16295),
            .I(N__16292));
    Odrv4 I__2666 (
            .O(N__16292),
            .I(\eeprom.n2180 ));
    InMux I__2665 (
            .O(N__16289),
            .I(N__16285));
    InMux I__2664 (
            .O(N__16288),
            .I(N__16282));
    LocalMux I__2663 (
            .O(N__16285),
            .I(N__16277));
    LocalMux I__2662 (
            .O(N__16282),
            .I(N__16277));
    Odrv4 I__2661 (
            .O(N__16277),
            .I(\eeprom.n2219 ));
    InMux I__2660 (
            .O(N__16274),
            .I(N__16271));
    LocalMux I__2659 (
            .O(N__16271),
            .I(N__16268));
    Odrv12 I__2658 (
            .O(N__16268),
            .I(\eeprom.n2286 ));
    InMux I__2657 (
            .O(N__16265),
            .I(bfn_6_26_0_));
    CascadeMux I__2656 (
            .O(N__16262),
            .I(N__16259));
    InMux I__2655 (
            .O(N__16259),
            .I(N__16255));
    InMux I__2654 (
            .O(N__16258),
            .I(N__16252));
    LocalMux I__2653 (
            .O(N__16255),
            .I(\eeprom.n2218 ));
    LocalMux I__2652 (
            .O(N__16252),
            .I(\eeprom.n2218 ));
    InMux I__2651 (
            .O(N__16247),
            .I(N__16244));
    LocalMux I__2650 (
            .O(N__16244),
            .I(\eeprom.n2285 ));
    InMux I__2649 (
            .O(N__16241),
            .I(\eeprom.n3541 ));
    CascadeMux I__2648 (
            .O(N__16238),
            .I(N__16234));
    CascadeMux I__2647 (
            .O(N__16237),
            .I(N__16231));
    InMux I__2646 (
            .O(N__16234),
            .I(N__16227));
    InMux I__2645 (
            .O(N__16231),
            .I(N__16224));
    InMux I__2644 (
            .O(N__16230),
            .I(N__16221));
    LocalMux I__2643 (
            .O(N__16227),
            .I(\eeprom.n2217 ));
    LocalMux I__2642 (
            .O(N__16224),
            .I(\eeprom.n2217 ));
    LocalMux I__2641 (
            .O(N__16221),
            .I(\eeprom.n2217 ));
    InMux I__2640 (
            .O(N__16214),
            .I(N__16211));
    LocalMux I__2639 (
            .O(N__16211),
            .I(\eeprom.n2284 ));
    InMux I__2638 (
            .O(N__16208),
            .I(\eeprom.n3542 ));
    CascadeMux I__2637 (
            .O(N__16205),
            .I(N__16200));
    CascadeMux I__2636 (
            .O(N__16204),
            .I(N__16197));
    InMux I__2635 (
            .O(N__16203),
            .I(N__16194));
    InMux I__2634 (
            .O(N__16200),
            .I(N__16191));
    InMux I__2633 (
            .O(N__16197),
            .I(N__16188));
    LocalMux I__2632 (
            .O(N__16194),
            .I(\eeprom.n2216 ));
    LocalMux I__2631 (
            .O(N__16191),
            .I(\eeprom.n2216 ));
    LocalMux I__2630 (
            .O(N__16188),
            .I(\eeprom.n2216 ));
    CascadeMux I__2629 (
            .O(N__16181),
            .I(N__16178));
    InMux I__2628 (
            .O(N__16178),
            .I(N__16175));
    LocalMux I__2627 (
            .O(N__16175),
            .I(\eeprom.n2283 ));
    InMux I__2626 (
            .O(N__16172),
            .I(\eeprom.n3543 ));
    CascadeMux I__2625 (
            .O(N__16169),
            .I(N__16166));
    InMux I__2624 (
            .O(N__16166),
            .I(N__16162));
    InMux I__2623 (
            .O(N__16165),
            .I(N__16159));
    LocalMux I__2622 (
            .O(N__16162),
            .I(\eeprom.n2215 ));
    LocalMux I__2621 (
            .O(N__16159),
            .I(\eeprom.n2215 ));
    CascadeMux I__2620 (
            .O(N__16154),
            .I(N__16151));
    InMux I__2619 (
            .O(N__16151),
            .I(N__16148));
    LocalMux I__2618 (
            .O(N__16148),
            .I(N__16145));
    Odrv4 I__2617 (
            .O(N__16145),
            .I(\eeprom.n2282 ));
    InMux I__2616 (
            .O(N__16142),
            .I(\eeprom.n3544 ));
    CascadeMux I__2615 (
            .O(N__16139),
            .I(N__16136));
    InMux I__2614 (
            .O(N__16136),
            .I(N__16132));
    InMux I__2613 (
            .O(N__16135),
            .I(N__16129));
    LocalMux I__2612 (
            .O(N__16132),
            .I(\eeprom.n2214 ));
    LocalMux I__2611 (
            .O(N__16129),
            .I(\eeprom.n2214 ));
    InMux I__2610 (
            .O(N__16124),
            .I(N__16121));
    LocalMux I__2609 (
            .O(N__16121),
            .I(\eeprom.n2281 ));
    InMux I__2608 (
            .O(N__16118),
            .I(\eeprom.n3545 ));
    InMux I__2607 (
            .O(N__16115),
            .I(N__16111));
    CascadeMux I__2606 (
            .O(N__16114),
            .I(N__16108));
    LocalMux I__2605 (
            .O(N__16111),
            .I(N__16104));
    InMux I__2604 (
            .O(N__16108),
            .I(N__16101));
    InMux I__2603 (
            .O(N__16107),
            .I(N__16098));
    Odrv4 I__2602 (
            .O(N__16104),
            .I(\eeprom.n2213 ));
    LocalMux I__2601 (
            .O(N__16101),
            .I(\eeprom.n2213 ));
    LocalMux I__2600 (
            .O(N__16098),
            .I(\eeprom.n2213 ));
    InMux I__2599 (
            .O(N__16091),
            .I(N__16087));
    CascadeMux I__2598 (
            .O(N__16090),
            .I(N__16084));
    LocalMux I__2597 (
            .O(N__16087),
            .I(N__16080));
    InMux I__2596 (
            .O(N__16084),
            .I(N__16077));
    InMux I__2595 (
            .O(N__16083),
            .I(N__16074));
    Odrv12 I__2594 (
            .O(N__16080),
            .I(\eeprom.n2413 ));
    LocalMux I__2593 (
            .O(N__16077),
            .I(\eeprom.n2413 ));
    LocalMux I__2592 (
            .O(N__16074),
            .I(\eeprom.n2413 ));
    CascadeMux I__2591 (
            .O(N__16067),
            .I(N__16064));
    InMux I__2590 (
            .O(N__16064),
            .I(N__16061));
    LocalMux I__2589 (
            .O(N__16061),
            .I(N__16058));
    Span4Mux_h I__2588 (
            .O(N__16058),
            .I(N__16055));
    Odrv4 I__2587 (
            .O(N__16055),
            .I(\eeprom.n2480 ));
    InMux I__2586 (
            .O(N__16052),
            .I(N__16047));
    CascadeMux I__2585 (
            .O(N__16051),
            .I(N__16044));
    InMux I__2584 (
            .O(N__16050),
            .I(N__16041));
    LocalMux I__2583 (
            .O(N__16047),
            .I(N__16038));
    InMux I__2582 (
            .O(N__16044),
            .I(N__16035));
    LocalMux I__2581 (
            .O(N__16041),
            .I(N__16032));
    Span4Mux_h I__2580 (
            .O(N__16038),
            .I(N__16025));
    LocalMux I__2579 (
            .O(N__16035),
            .I(N__16025));
    Span4Mux_h I__2578 (
            .O(N__16032),
            .I(N__16025));
    Odrv4 I__2577 (
            .O(N__16025),
            .I(\eeprom.n2512 ));
    InMux I__2576 (
            .O(N__16022),
            .I(N__16018));
    InMux I__2575 (
            .O(N__16021),
            .I(N__16015));
    LocalMux I__2574 (
            .O(N__16018),
            .I(N__16011));
    LocalMux I__2573 (
            .O(N__16015),
            .I(N__16008));
    InMux I__2572 (
            .O(N__16014),
            .I(N__16005));
    Odrv12 I__2571 (
            .O(N__16011),
            .I(\eeprom.n2408 ));
    Odrv4 I__2570 (
            .O(N__16008),
            .I(\eeprom.n2408 ));
    LocalMux I__2569 (
            .O(N__16005),
            .I(\eeprom.n2408 ));
    CascadeMux I__2568 (
            .O(N__15998),
            .I(N__15995));
    InMux I__2567 (
            .O(N__15995),
            .I(N__15992));
    LocalMux I__2566 (
            .O(N__15992),
            .I(N__15989));
    Span4Mux_v I__2565 (
            .O(N__15989),
            .I(N__15986));
    Odrv4 I__2564 (
            .O(N__15986),
            .I(\eeprom.n2475 ));
    CascadeMux I__2563 (
            .O(N__15983),
            .I(N__15979));
    InMux I__2562 (
            .O(N__15982),
            .I(N__15974));
    InMux I__2561 (
            .O(N__15979),
            .I(N__15967));
    InMux I__2560 (
            .O(N__15978),
            .I(N__15967));
    CascadeMux I__2559 (
            .O(N__15977),
            .I(N__15964));
    LocalMux I__2558 (
            .O(N__15974),
            .I(N__15956));
    InMux I__2557 (
            .O(N__15973),
            .I(N__15951));
    InMux I__2556 (
            .O(N__15972),
            .I(N__15951));
    LocalMux I__2555 (
            .O(N__15967),
            .I(N__15948));
    InMux I__2554 (
            .O(N__15964),
            .I(N__15941));
    InMux I__2553 (
            .O(N__15963),
            .I(N__15941));
    InMux I__2552 (
            .O(N__15962),
            .I(N__15941));
    InMux I__2551 (
            .O(N__15961),
            .I(N__15936));
    InMux I__2550 (
            .O(N__15960),
            .I(N__15936));
    CascadeMux I__2549 (
            .O(N__15959),
            .I(N__15932));
    Span4Mux_h I__2548 (
            .O(N__15956),
            .I(N__15928));
    LocalMux I__2547 (
            .O(N__15951),
            .I(N__15925));
    Span4Mux_v I__2546 (
            .O(N__15948),
            .I(N__15920));
    LocalMux I__2545 (
            .O(N__15941),
            .I(N__15920));
    LocalMux I__2544 (
            .O(N__15936),
            .I(N__15917));
    InMux I__2543 (
            .O(N__15935),
            .I(N__15910));
    InMux I__2542 (
            .O(N__15932),
            .I(N__15910));
    InMux I__2541 (
            .O(N__15931),
            .I(N__15910));
    Odrv4 I__2540 (
            .O(N__15928),
            .I(\eeprom.n2440 ));
    Odrv4 I__2539 (
            .O(N__15925),
            .I(\eeprom.n2440 ));
    Odrv4 I__2538 (
            .O(N__15920),
            .I(\eeprom.n2440 ));
    Odrv4 I__2537 (
            .O(N__15917),
            .I(\eeprom.n2440 ));
    LocalMux I__2536 (
            .O(N__15910),
            .I(\eeprom.n2440 ));
    InMux I__2535 (
            .O(N__15899),
            .I(N__15894));
    InMux I__2534 (
            .O(N__15898),
            .I(N__15891));
    InMux I__2533 (
            .O(N__15897),
            .I(N__15888));
    LocalMux I__2532 (
            .O(N__15894),
            .I(N__15885));
    LocalMux I__2531 (
            .O(N__15891),
            .I(N__15878));
    LocalMux I__2530 (
            .O(N__15888),
            .I(N__15878));
    Span4Mux_h I__2529 (
            .O(N__15885),
            .I(N__15878));
    Odrv4 I__2528 (
            .O(N__15878),
            .I(\eeprom.n2507 ));
    InMux I__2527 (
            .O(N__15875),
            .I(N__15872));
    LocalMux I__2526 (
            .O(N__15872),
            .I(\eeprom.n4801 ));
    InMux I__2525 (
            .O(N__15869),
            .I(N__15865));
    CascadeMux I__2524 (
            .O(N__15868),
            .I(N__15862));
    LocalMux I__2523 (
            .O(N__15865),
            .I(N__15859));
    InMux I__2522 (
            .O(N__15862),
            .I(N__15855));
    Span4Mux_v I__2521 (
            .O(N__15859),
            .I(N__15852));
    InMux I__2520 (
            .O(N__15858),
            .I(N__15849));
    LocalMux I__2519 (
            .O(N__15855),
            .I(N__15846));
    Odrv4 I__2518 (
            .O(N__15852),
            .I(\eeprom.n2017 ));
    LocalMux I__2517 (
            .O(N__15849),
            .I(\eeprom.n2017 ));
    Odrv4 I__2516 (
            .O(N__15846),
            .I(\eeprom.n2017 ));
    CascadeMux I__2515 (
            .O(N__15839),
            .I(\eeprom.n4799_cascade_ ));
    InMux I__2514 (
            .O(N__15836),
            .I(N__15833));
    LocalMux I__2513 (
            .O(N__15833),
            .I(\eeprom.n4872 ));
    CascadeMux I__2512 (
            .O(N__15830),
            .I(N__15826));
    CascadeMux I__2511 (
            .O(N__15829),
            .I(N__15823));
    InMux I__2510 (
            .O(N__15826),
            .I(N__15820));
    InMux I__2509 (
            .O(N__15823),
            .I(N__15816));
    LocalMux I__2508 (
            .O(N__15820),
            .I(N__15813));
    CascadeMux I__2507 (
            .O(N__15819),
            .I(N__15810));
    LocalMux I__2506 (
            .O(N__15816),
            .I(N__15807));
    Span4Mux_h I__2505 (
            .O(N__15813),
            .I(N__15804));
    InMux I__2504 (
            .O(N__15810),
            .I(N__15801));
    Odrv4 I__2503 (
            .O(N__15807),
            .I(\eeprom.n2314 ));
    Odrv4 I__2502 (
            .O(N__15804),
            .I(\eeprom.n2314 ));
    LocalMux I__2501 (
            .O(N__15801),
            .I(\eeprom.n2314 ));
    CascadeMux I__2500 (
            .O(N__15794),
            .I(N__15790));
    InMux I__2499 (
            .O(N__15793),
            .I(N__15787));
    InMux I__2498 (
            .O(N__15790),
            .I(N__15784));
    LocalMux I__2497 (
            .O(N__15787),
            .I(N__15781));
    LocalMux I__2496 (
            .O(N__15784),
            .I(N__15777));
    Span4Mux_h I__2495 (
            .O(N__15781),
            .I(N__15774));
    InMux I__2494 (
            .O(N__15780),
            .I(N__15771));
    Span4Mux_h I__2493 (
            .O(N__15777),
            .I(N__15768));
    Odrv4 I__2492 (
            .O(N__15774),
            .I(\eeprom.n2316 ));
    LocalMux I__2491 (
            .O(N__15771),
            .I(\eeprom.n2316 ));
    Odrv4 I__2490 (
            .O(N__15768),
            .I(\eeprom.n2316 ));
    InMux I__2489 (
            .O(N__15761),
            .I(N__15758));
    LocalMux I__2488 (
            .O(N__15758),
            .I(N__15755));
    Odrv4 I__2487 (
            .O(N__15755),
            .I(\eeprom.n2186 ));
    InMux I__2486 (
            .O(N__15752),
            .I(N__15747));
    InMux I__2485 (
            .O(N__15751),
            .I(N__15744));
    InMux I__2484 (
            .O(N__15750),
            .I(N__15741));
    LocalMux I__2483 (
            .O(N__15747),
            .I(N__15738));
    LocalMux I__2482 (
            .O(N__15744),
            .I(\eeprom.n2119 ));
    LocalMux I__2481 (
            .O(N__15741),
            .I(\eeprom.n2119 ));
    Odrv4 I__2480 (
            .O(N__15738),
            .I(\eeprom.n2119 ));
    CascadeMux I__2479 (
            .O(N__15731),
            .I(\eeprom.n2218_cascade_ ));
    CascadeMux I__2478 (
            .O(N__15728),
            .I(N__15724));
    InMux I__2477 (
            .O(N__15727),
            .I(N__15721));
    InMux I__2476 (
            .O(N__15724),
            .I(N__15718));
    LocalMux I__2475 (
            .O(N__15721),
            .I(N__15712));
    LocalMux I__2474 (
            .O(N__15718),
            .I(N__15712));
    InMux I__2473 (
            .O(N__15717),
            .I(N__15709));
    Span4Mux_v I__2472 (
            .O(N__15712),
            .I(N__15706));
    LocalMux I__2471 (
            .O(N__15709),
            .I(\eeprom.n2317 ));
    Odrv4 I__2470 (
            .O(N__15706),
            .I(\eeprom.n2317 ));
    CascadeMux I__2469 (
            .O(N__15701),
            .I(\eeprom.n4447_cascade_ ));
    InMux I__2468 (
            .O(N__15698),
            .I(N__15695));
    LocalMux I__2467 (
            .O(N__15695),
            .I(\eeprom.n4218 ));
    InMux I__2466 (
            .O(N__15692),
            .I(N__15689));
    LocalMux I__2465 (
            .O(N__15689),
            .I(N__15686));
    Span4Mux_h I__2464 (
            .O(N__15686),
            .I(N__15681));
    InMux I__2463 (
            .O(N__15685),
            .I(N__15678));
    InMux I__2462 (
            .O(N__15684),
            .I(N__15675));
    Odrv4 I__2461 (
            .O(N__15681),
            .I(\eeprom.n2412 ));
    LocalMux I__2460 (
            .O(N__15678),
            .I(\eeprom.n2412 ));
    LocalMux I__2459 (
            .O(N__15675),
            .I(\eeprom.n2412 ));
    CascadeMux I__2458 (
            .O(N__15668),
            .I(N__15665));
    InMux I__2457 (
            .O(N__15665),
            .I(N__15662));
    LocalMux I__2456 (
            .O(N__15662),
            .I(N__15659));
    Span4Mux_h I__2455 (
            .O(N__15659),
            .I(N__15656));
    Odrv4 I__2454 (
            .O(N__15656),
            .I(\eeprom.n2479 ));
    InMux I__2453 (
            .O(N__15653),
            .I(N__15649));
    CascadeMux I__2452 (
            .O(N__15652),
            .I(N__15646));
    LocalMux I__2451 (
            .O(N__15649),
            .I(N__15643));
    InMux I__2450 (
            .O(N__15646),
            .I(N__15640));
    Odrv4 I__2449 (
            .O(N__15643),
            .I(\eeprom.n2511 ));
    LocalMux I__2448 (
            .O(N__15640),
            .I(\eeprom.n2511 ));
    InMux I__2447 (
            .O(N__15635),
            .I(N__15632));
    LocalMux I__2446 (
            .O(N__15632),
            .I(\eeprom.n2578 ));
    CascadeMux I__2445 (
            .O(N__15629),
            .I(\eeprom.n2511_cascade_ ));
    InMux I__2444 (
            .O(N__15626),
            .I(N__15623));
    LocalMux I__2443 (
            .O(N__15623),
            .I(N__15620));
    Odrv12 I__2442 (
            .O(N__15620),
            .I(\eeprom.n12_adj_351 ));
    InMux I__2441 (
            .O(N__15617),
            .I(N__15613));
    InMux I__2440 (
            .O(N__15616),
            .I(N__15610));
    LocalMux I__2439 (
            .O(N__15613),
            .I(N__15606));
    LocalMux I__2438 (
            .O(N__15610),
            .I(N__15603));
    InMux I__2437 (
            .O(N__15609),
            .I(N__15600));
    Span4Mux_v I__2436 (
            .O(N__15606),
            .I(N__15597));
    Span4Mux_h I__2435 (
            .O(N__15603),
            .I(N__15594));
    LocalMux I__2434 (
            .O(N__15600),
            .I(\eeprom.delay_counter_21 ));
    Odrv4 I__2433 (
            .O(N__15597),
            .I(\eeprom.delay_counter_21 ));
    Odrv4 I__2432 (
            .O(N__15594),
            .I(\eeprom.delay_counter_21 ));
    CascadeMux I__2431 (
            .O(N__15587),
            .I(\eeprom.n2219_cascade_ ));
    CascadeMux I__2430 (
            .O(N__15584),
            .I(N__15580));
    InMux I__2429 (
            .O(N__15583),
            .I(N__15576));
    InMux I__2428 (
            .O(N__15580),
            .I(N__15573));
    InMux I__2427 (
            .O(N__15579),
            .I(N__15570));
    LocalMux I__2426 (
            .O(N__15576),
            .I(N__15565));
    LocalMux I__2425 (
            .O(N__15573),
            .I(N__15565));
    LocalMux I__2424 (
            .O(N__15570),
            .I(\eeprom.n2318 ));
    Odrv4 I__2423 (
            .O(N__15565),
            .I(\eeprom.n2318 ));
    InMux I__2422 (
            .O(N__15560),
            .I(N__15557));
    LocalMux I__2421 (
            .O(N__15557),
            .I(N__15554));
    Odrv4 I__2420 (
            .O(N__15554),
            .I(\eeprom.n2580 ));
    CascadeMux I__2419 (
            .O(N__15551),
            .I(N__15548));
    InMux I__2418 (
            .O(N__15548),
            .I(N__15544));
    InMux I__2417 (
            .O(N__15547),
            .I(N__15541));
    LocalMux I__2416 (
            .O(N__15544),
            .I(N__15538));
    LocalMux I__2415 (
            .O(N__15541),
            .I(N__15534));
    Span4Mux_h I__2414 (
            .O(N__15538),
            .I(N__15531));
    InMux I__2413 (
            .O(N__15537),
            .I(N__15528));
    Odrv4 I__2412 (
            .O(N__15534),
            .I(\eeprom.n2513 ));
    Odrv4 I__2411 (
            .O(N__15531),
            .I(\eeprom.n2513 ));
    LocalMux I__2410 (
            .O(N__15528),
            .I(\eeprom.n2513 ));
    CascadeMux I__2409 (
            .O(N__15521),
            .I(N__15514));
    CascadeMux I__2408 (
            .O(N__15520),
            .I(N__15509));
    CascadeMux I__2407 (
            .O(N__15519),
            .I(N__15506));
    CascadeMux I__2406 (
            .O(N__15518),
            .I(N__15501));
    CascadeMux I__2405 (
            .O(N__15517),
            .I(N__15495));
    InMux I__2404 (
            .O(N__15514),
            .I(N__15489));
    InMux I__2403 (
            .O(N__15513),
            .I(N__15489));
    InMux I__2402 (
            .O(N__15512),
            .I(N__15484));
    InMux I__2401 (
            .O(N__15509),
            .I(N__15484));
    InMux I__2400 (
            .O(N__15506),
            .I(N__15479));
    InMux I__2399 (
            .O(N__15505),
            .I(N__15479));
    InMux I__2398 (
            .O(N__15504),
            .I(N__15472));
    InMux I__2397 (
            .O(N__15501),
            .I(N__15472));
    InMux I__2396 (
            .O(N__15500),
            .I(N__15472));
    InMux I__2395 (
            .O(N__15499),
            .I(N__15469));
    InMux I__2394 (
            .O(N__15498),
            .I(N__15462));
    InMux I__2393 (
            .O(N__15495),
            .I(N__15462));
    InMux I__2392 (
            .O(N__15494),
            .I(N__15462));
    LocalMux I__2391 (
            .O(N__15489),
            .I(N__15457));
    LocalMux I__2390 (
            .O(N__15484),
            .I(N__15457));
    LocalMux I__2389 (
            .O(N__15479),
            .I(\eeprom.n2539 ));
    LocalMux I__2388 (
            .O(N__15472),
            .I(\eeprom.n2539 ));
    LocalMux I__2387 (
            .O(N__15469),
            .I(\eeprom.n2539 ));
    LocalMux I__2386 (
            .O(N__15462),
            .I(\eeprom.n2539 ));
    Odrv4 I__2385 (
            .O(N__15457),
            .I(\eeprom.n2539 ));
    InMux I__2384 (
            .O(N__15446),
            .I(N__15443));
    LocalMux I__2383 (
            .O(N__15443),
            .I(\eeprom.n2574 ));
    CascadeMux I__2382 (
            .O(N__15440),
            .I(\eeprom.n2606_cascade_ ));
    CascadeMux I__2381 (
            .O(N__15437),
            .I(N__15434));
    InMux I__2380 (
            .O(N__15434),
            .I(N__15431));
    LocalMux I__2379 (
            .O(N__15431),
            .I(N__15427));
    InMux I__2378 (
            .O(N__15430),
            .I(N__15424));
    Odrv4 I__2377 (
            .O(N__15427),
            .I(\eeprom.n2605 ));
    LocalMux I__2376 (
            .O(N__15424),
            .I(\eeprom.n2605 ));
    CascadeMux I__2375 (
            .O(N__15419),
            .I(N__15415));
    InMux I__2374 (
            .O(N__15418),
            .I(N__15412));
    InMux I__2373 (
            .O(N__15415),
            .I(N__15409));
    LocalMux I__2372 (
            .O(N__15412),
            .I(N__15406));
    LocalMux I__2371 (
            .O(N__15409),
            .I(\eeprom.n2611 ));
    Odrv4 I__2370 (
            .O(N__15406),
            .I(\eeprom.n2611 ));
    CascadeMux I__2369 (
            .O(N__15401),
            .I(\eeprom.n10_adj_475_cascade_ ));
    InMux I__2368 (
            .O(N__15398),
            .I(N__15395));
    LocalMux I__2367 (
            .O(N__15395),
            .I(\eeprom.n2581 ));
    InMux I__2366 (
            .O(N__15392),
            .I(\eeprom.n3578 ));
    InMux I__2365 (
            .O(N__15389),
            .I(\eeprom.n3579 ));
    CascadeMux I__2364 (
            .O(N__15386),
            .I(N__15383));
    InMux I__2363 (
            .O(N__15383),
            .I(N__15380));
    LocalMux I__2362 (
            .O(N__15380),
            .I(\eeprom.n2579 ));
    InMux I__2361 (
            .O(N__15377),
            .I(\eeprom.n3580 ));
    InMux I__2360 (
            .O(N__15374),
            .I(bfn_6_22_0_));
    CascadeMux I__2359 (
            .O(N__15371),
            .I(N__15366));
    CascadeMux I__2358 (
            .O(N__15370),
            .I(N__15363));
    InMux I__2357 (
            .O(N__15369),
            .I(N__15360));
    InMux I__2356 (
            .O(N__15366),
            .I(N__15357));
    InMux I__2355 (
            .O(N__15363),
            .I(N__15354));
    LocalMux I__2354 (
            .O(N__15360),
            .I(\eeprom.n2510 ));
    LocalMux I__2353 (
            .O(N__15357),
            .I(\eeprom.n2510 ));
    LocalMux I__2352 (
            .O(N__15354),
            .I(\eeprom.n2510 ));
    InMux I__2351 (
            .O(N__15347),
            .I(N__15344));
    LocalMux I__2350 (
            .O(N__15344),
            .I(N__15341));
    Odrv4 I__2349 (
            .O(N__15341),
            .I(\eeprom.n2577 ));
    InMux I__2348 (
            .O(N__15338),
            .I(\eeprom.n3582 ));
    InMux I__2347 (
            .O(N__15335),
            .I(N__15331));
    CascadeMux I__2346 (
            .O(N__15334),
            .I(N__15328));
    LocalMux I__2345 (
            .O(N__15331),
            .I(N__15324));
    InMux I__2344 (
            .O(N__15328),
            .I(N__15321));
    InMux I__2343 (
            .O(N__15327),
            .I(N__15318));
    Span4Mux_h I__2342 (
            .O(N__15324),
            .I(N__15315));
    LocalMux I__2341 (
            .O(N__15321),
            .I(N__15312));
    LocalMux I__2340 (
            .O(N__15318),
            .I(N__15309));
    Span4Mux_v I__2339 (
            .O(N__15315),
            .I(N__15306));
    Span4Mux_h I__2338 (
            .O(N__15312),
            .I(N__15301));
    Span4Mux_v I__2337 (
            .O(N__15309),
            .I(N__15301));
    Odrv4 I__2336 (
            .O(N__15306),
            .I(\eeprom.n2509 ));
    Odrv4 I__2335 (
            .O(N__15301),
            .I(\eeprom.n2509 ));
    InMux I__2334 (
            .O(N__15296),
            .I(N__15293));
    LocalMux I__2333 (
            .O(N__15293),
            .I(N__15290));
    Odrv4 I__2332 (
            .O(N__15290),
            .I(\eeprom.n2576 ));
    InMux I__2331 (
            .O(N__15287),
            .I(\eeprom.n3583 ));
    InMux I__2330 (
            .O(N__15284),
            .I(N__15280));
    CascadeMux I__2329 (
            .O(N__15283),
            .I(N__15277));
    LocalMux I__2328 (
            .O(N__15280),
            .I(N__15273));
    InMux I__2327 (
            .O(N__15277),
            .I(N__15270));
    CascadeMux I__2326 (
            .O(N__15276),
            .I(N__15267));
    Span4Mux_v I__2325 (
            .O(N__15273),
            .I(N__15262));
    LocalMux I__2324 (
            .O(N__15270),
            .I(N__15262));
    InMux I__2323 (
            .O(N__15267),
            .I(N__15259));
    Span4Mux_h I__2322 (
            .O(N__15262),
            .I(N__15256));
    LocalMux I__2321 (
            .O(N__15259),
            .I(N__15253));
    Span4Mux_v I__2320 (
            .O(N__15256),
            .I(N__15250));
    Span4Mux_v I__2319 (
            .O(N__15253),
            .I(N__15247));
    Odrv4 I__2318 (
            .O(N__15250),
            .I(\eeprom.n2508 ));
    Odrv4 I__2317 (
            .O(N__15247),
            .I(\eeprom.n2508 ));
    CascadeMux I__2316 (
            .O(N__15242),
            .I(N__15239));
    InMux I__2315 (
            .O(N__15239),
            .I(N__15236));
    LocalMux I__2314 (
            .O(N__15236),
            .I(N__15233));
    Odrv4 I__2313 (
            .O(N__15233),
            .I(\eeprom.n2575 ));
    InMux I__2312 (
            .O(N__15230),
            .I(\eeprom.n3584 ));
    InMux I__2311 (
            .O(N__15227),
            .I(\eeprom.n3585 ));
    InMux I__2310 (
            .O(N__15224),
            .I(N__15220));
    InMux I__2309 (
            .O(N__15223),
            .I(N__15217));
    LocalMux I__2308 (
            .O(N__15220),
            .I(N__15214));
    LocalMux I__2307 (
            .O(N__15217),
            .I(N__15211));
    Span4Mux_h I__2306 (
            .O(N__15214),
            .I(N__15206));
    Span4Mux_v I__2305 (
            .O(N__15211),
            .I(N__15206));
    Odrv4 I__2304 (
            .O(N__15206),
            .I(\eeprom.n2506 ));
    InMux I__2303 (
            .O(N__15203),
            .I(\eeprom.n3586 ));
    InMux I__2302 (
            .O(N__15200),
            .I(N__15197));
    LocalMux I__2301 (
            .O(N__15197),
            .I(\eeprom.n2678 ));
    CascadeMux I__2300 (
            .O(N__15194),
            .I(\eeprom.n2611_cascade_ ));
    InMux I__2299 (
            .O(N__15191),
            .I(N__15188));
    LocalMux I__2298 (
            .O(N__15188),
            .I(N__15184));
    InMux I__2297 (
            .O(N__15187),
            .I(N__15181));
    Span4Mux_v I__2296 (
            .O(N__15184),
            .I(N__15175));
    LocalMux I__2295 (
            .O(N__15181),
            .I(N__15175));
    InMux I__2294 (
            .O(N__15180),
            .I(N__15172));
    Span4Mux_h I__2293 (
            .O(N__15175),
            .I(N__15169));
    LocalMux I__2292 (
            .O(N__15172),
            .I(\eeprom.n2519 ));
    Odrv4 I__2291 (
            .O(N__15169),
            .I(\eeprom.n2519 ));
    InMux I__2290 (
            .O(N__15164),
            .I(N__15161));
    LocalMux I__2289 (
            .O(N__15161),
            .I(N__15158));
    Odrv4 I__2288 (
            .O(N__15158),
            .I(\eeprom.n2586 ));
    InMux I__2287 (
            .O(N__15155),
            .I(bfn_6_21_0_));
    CascadeMux I__2286 (
            .O(N__15152),
            .I(N__15149));
    InMux I__2285 (
            .O(N__15149),
            .I(N__15145));
    CascadeMux I__2284 (
            .O(N__15148),
            .I(N__15141));
    LocalMux I__2283 (
            .O(N__15145),
            .I(N__15138));
    InMux I__2282 (
            .O(N__15144),
            .I(N__15135));
    InMux I__2281 (
            .O(N__15141),
            .I(N__15132));
    Odrv4 I__2280 (
            .O(N__15138),
            .I(\eeprom.n2518 ));
    LocalMux I__2279 (
            .O(N__15135),
            .I(\eeprom.n2518 ));
    LocalMux I__2278 (
            .O(N__15132),
            .I(\eeprom.n2518 ));
    InMux I__2277 (
            .O(N__15125),
            .I(N__15122));
    LocalMux I__2276 (
            .O(N__15122),
            .I(N__15119));
    Odrv4 I__2275 (
            .O(N__15119),
            .I(\eeprom.n2585 ));
    InMux I__2274 (
            .O(N__15116),
            .I(\eeprom.n3574 ));
    CascadeMux I__2273 (
            .O(N__15113),
            .I(N__15109));
    InMux I__2272 (
            .O(N__15112),
            .I(N__15106));
    InMux I__2271 (
            .O(N__15109),
            .I(N__15103));
    LocalMux I__2270 (
            .O(N__15106),
            .I(N__15100));
    LocalMux I__2269 (
            .O(N__15103),
            .I(N__15097));
    Span4Mux_v I__2268 (
            .O(N__15100),
            .I(N__15093));
    Span4Mux_h I__2267 (
            .O(N__15097),
            .I(N__15090));
    InMux I__2266 (
            .O(N__15096),
            .I(N__15087));
    Odrv4 I__2265 (
            .O(N__15093),
            .I(\eeprom.n2517 ));
    Odrv4 I__2264 (
            .O(N__15090),
            .I(\eeprom.n2517 ));
    LocalMux I__2263 (
            .O(N__15087),
            .I(\eeprom.n2517 ));
    InMux I__2262 (
            .O(N__15080),
            .I(N__15077));
    LocalMux I__2261 (
            .O(N__15077),
            .I(N__15074));
    Odrv4 I__2260 (
            .O(N__15074),
            .I(\eeprom.n2584 ));
    InMux I__2259 (
            .O(N__15071),
            .I(\eeprom.n3575 ));
    CascadeMux I__2258 (
            .O(N__15068),
            .I(N__15064));
    InMux I__2257 (
            .O(N__15067),
            .I(N__15061));
    InMux I__2256 (
            .O(N__15064),
            .I(N__15058));
    LocalMux I__2255 (
            .O(N__15061),
            .I(N__15055));
    LocalMux I__2254 (
            .O(N__15058),
            .I(N__15052));
    Span4Mux_v I__2253 (
            .O(N__15055),
            .I(N__15048));
    Span4Mux_h I__2252 (
            .O(N__15052),
            .I(N__15045));
    InMux I__2251 (
            .O(N__15051),
            .I(N__15042));
    Odrv4 I__2250 (
            .O(N__15048),
            .I(\eeprom.n2516 ));
    Odrv4 I__2249 (
            .O(N__15045),
            .I(\eeprom.n2516 ));
    LocalMux I__2248 (
            .O(N__15042),
            .I(\eeprom.n2516 ));
    CascadeMux I__2247 (
            .O(N__15035),
            .I(N__15032));
    InMux I__2246 (
            .O(N__15032),
            .I(N__15029));
    LocalMux I__2245 (
            .O(N__15029),
            .I(N__15026));
    Odrv4 I__2244 (
            .O(N__15026),
            .I(\eeprom.n2583 ));
    InMux I__2243 (
            .O(N__15023),
            .I(\eeprom.n3576 ));
    CascadeMux I__2242 (
            .O(N__15020),
            .I(N__15016));
    CascadeMux I__2241 (
            .O(N__15019),
            .I(N__15013));
    InMux I__2240 (
            .O(N__15016),
            .I(N__15010));
    InMux I__2239 (
            .O(N__15013),
            .I(N__15007));
    LocalMux I__2238 (
            .O(N__15010),
            .I(N__15003));
    LocalMux I__2237 (
            .O(N__15007),
            .I(N__15000));
    CascadeMux I__2236 (
            .O(N__15006),
            .I(N__14997));
    Span4Mux_h I__2235 (
            .O(N__15003),
            .I(N__14994));
    Span4Mux_h I__2234 (
            .O(N__15000),
            .I(N__14991));
    InMux I__2233 (
            .O(N__14997),
            .I(N__14988));
    Odrv4 I__2232 (
            .O(N__14994),
            .I(\eeprom.n2515 ));
    Odrv4 I__2231 (
            .O(N__14991),
            .I(\eeprom.n2515 ));
    LocalMux I__2230 (
            .O(N__14988),
            .I(\eeprom.n2515 ));
    InMux I__2229 (
            .O(N__14981),
            .I(N__14978));
    LocalMux I__2228 (
            .O(N__14978),
            .I(\eeprom.n2582 ));
    InMux I__2227 (
            .O(N__14975),
            .I(\eeprom.n3577 ));
    CascadeMux I__2226 (
            .O(N__14972),
            .I(N__14969));
    InMux I__2225 (
            .O(N__14969),
            .I(N__14965));
    InMux I__2224 (
            .O(N__14968),
            .I(N__14962));
    LocalMux I__2223 (
            .O(N__14965),
            .I(N__14959));
    LocalMux I__2222 (
            .O(N__14962),
            .I(N__14955));
    Span4Mux_h I__2221 (
            .O(N__14959),
            .I(N__14952));
    InMux I__2220 (
            .O(N__14958),
            .I(N__14949));
    Odrv4 I__2219 (
            .O(N__14955),
            .I(\eeprom.n2514 ));
    Odrv4 I__2218 (
            .O(N__14952),
            .I(\eeprom.n2514 ));
    LocalMux I__2217 (
            .O(N__14949),
            .I(\eeprom.n2514 ));
    InMux I__2216 (
            .O(N__14942),
            .I(\eeprom.n3597 ));
    InMux I__2215 (
            .O(N__14939),
            .I(\eeprom.n3598 ));
    InMux I__2214 (
            .O(N__14936),
            .I(\eeprom.n3599 ));
    InMux I__2213 (
            .O(N__14933),
            .I(\eeprom.n3600 ));
    InMux I__2212 (
            .O(N__14930),
            .I(N__14927));
    LocalMux I__2211 (
            .O(N__14927),
            .I(N__14924));
    Span4Mux_v I__2210 (
            .O(N__14924),
            .I(N__14921));
    Odrv4 I__2209 (
            .O(N__14921),
            .I(\eeprom.n21 ));
    InMux I__2208 (
            .O(N__14918),
            .I(N__14915));
    LocalMux I__2207 (
            .O(N__14915),
            .I(N__14911));
    InMux I__2206 (
            .O(N__14914),
            .I(N__14907));
    Span4Mux_h I__2205 (
            .O(N__14911),
            .I(N__14904));
    InMux I__2204 (
            .O(N__14910),
            .I(N__14901));
    LocalMux I__2203 (
            .O(N__14907),
            .I(\eeprom.delay_counter_12 ));
    Odrv4 I__2202 (
            .O(N__14904),
            .I(\eeprom.delay_counter_12 ));
    LocalMux I__2201 (
            .O(N__14901),
            .I(\eeprom.delay_counter_12 ));
    CascadeMux I__2200 (
            .O(N__14894),
            .I(N__14891));
    InMux I__2199 (
            .O(N__14891),
            .I(N__14888));
    LocalMux I__2198 (
            .O(N__14888),
            .I(N__14885));
    Span4Mux_h I__2197 (
            .O(N__14885),
            .I(N__14882));
    Odrv4 I__2196 (
            .O(N__14882),
            .I(\eeprom.n29_adj_460 ));
    CascadeMux I__2195 (
            .O(N__14879),
            .I(N__14875));
    InMux I__2194 (
            .O(N__14878),
            .I(N__14871));
    InMux I__2193 (
            .O(N__14875),
            .I(N__14868));
    InMux I__2192 (
            .O(N__14874),
            .I(N__14865));
    LocalMux I__2191 (
            .O(N__14871),
            .I(\eeprom.n2609 ));
    LocalMux I__2190 (
            .O(N__14868),
            .I(\eeprom.n2609 ));
    LocalMux I__2189 (
            .O(N__14865),
            .I(\eeprom.n2609 ));
    CascadeMux I__2188 (
            .O(N__14858),
            .I(N__14855));
    InMux I__2187 (
            .O(N__14855),
            .I(N__14852));
    LocalMux I__2186 (
            .O(N__14852),
            .I(\eeprom.n2676 ));
    InMux I__2185 (
            .O(N__14849),
            .I(\eeprom.n3588 ));
    InMux I__2184 (
            .O(N__14846),
            .I(\eeprom.n3589 ));
    InMux I__2183 (
            .O(N__14843),
            .I(\eeprom.n3590 ));
    InMux I__2182 (
            .O(N__14840),
            .I(\eeprom.n3591 ));
    InMux I__2181 (
            .O(N__14837),
            .I(\eeprom.n3592 ));
    InMux I__2180 (
            .O(N__14834),
            .I(\eeprom.n3593 ));
    InMux I__2179 (
            .O(N__14831),
            .I(bfn_6_19_0_));
    InMux I__2178 (
            .O(N__14828),
            .I(\eeprom.n3595 ));
    InMux I__2177 (
            .O(N__14825),
            .I(\eeprom.n3596 ));
    InMux I__2176 (
            .O(N__14822),
            .I(N__14819));
    LocalMux I__2175 (
            .O(N__14819),
            .I(n7));
    InMux I__2174 (
            .O(N__14816),
            .I(n3503));
    InMux I__2173 (
            .O(N__14813),
            .I(N__14810));
    LocalMux I__2172 (
            .O(N__14810),
            .I(n6));
    InMux I__2171 (
            .O(N__14807),
            .I(n3504));
    CascadeMux I__2170 (
            .O(N__14804),
            .I(N__14801));
    InMux I__2169 (
            .O(N__14801),
            .I(N__14794));
    InMux I__2168 (
            .O(N__14800),
            .I(N__14794));
    InMux I__2167 (
            .O(N__14799),
            .I(N__14791));
    LocalMux I__2166 (
            .O(N__14794),
            .I(blink_counter_21));
    LocalMux I__2165 (
            .O(N__14791),
            .I(blink_counter_21));
    InMux I__2164 (
            .O(N__14786),
            .I(n3505));
    InMux I__2163 (
            .O(N__14783),
            .I(N__14776));
    InMux I__2162 (
            .O(N__14782),
            .I(N__14776));
    InMux I__2161 (
            .O(N__14781),
            .I(N__14773));
    LocalMux I__2160 (
            .O(N__14776),
            .I(blink_counter_22));
    LocalMux I__2159 (
            .O(N__14773),
            .I(blink_counter_22));
    InMux I__2158 (
            .O(N__14768),
            .I(n3506));
    CascadeMux I__2157 (
            .O(N__14765),
            .I(N__14761));
    InMux I__2156 (
            .O(N__14764),
            .I(N__14755));
    InMux I__2155 (
            .O(N__14761),
            .I(N__14755));
    InMux I__2154 (
            .O(N__14760),
            .I(N__14752));
    LocalMux I__2153 (
            .O(N__14755),
            .I(blink_counter_23));
    LocalMux I__2152 (
            .O(N__14752),
            .I(blink_counter_23));
    InMux I__2151 (
            .O(N__14747),
            .I(n3507));
    InMux I__2150 (
            .O(N__14744),
            .I(N__14737));
    InMux I__2149 (
            .O(N__14743),
            .I(N__14737));
    InMux I__2148 (
            .O(N__14742),
            .I(N__14734));
    LocalMux I__2147 (
            .O(N__14737),
            .I(blink_counter_24));
    LocalMux I__2146 (
            .O(N__14734),
            .I(blink_counter_24));
    InMux I__2145 (
            .O(N__14729),
            .I(bfn_5_32_0_));
    InMux I__2144 (
            .O(N__14726),
            .I(n3509));
    InMux I__2143 (
            .O(N__14723),
            .I(N__14719));
    InMux I__2142 (
            .O(N__14722),
            .I(N__14716));
    LocalMux I__2141 (
            .O(N__14719),
            .I(blink_counter_25));
    LocalMux I__2140 (
            .O(N__14716),
            .I(blink_counter_25));
    InMux I__2139 (
            .O(N__14711),
            .I(bfn_6_18_0_));
    InMux I__2138 (
            .O(N__14708),
            .I(\eeprom.n3587 ));
    InMux I__2137 (
            .O(N__14705),
            .I(N__14702));
    LocalMux I__2136 (
            .O(N__14702),
            .I(n15));
    InMux I__2135 (
            .O(N__14699),
            .I(n3495));
    InMux I__2134 (
            .O(N__14696),
            .I(N__14693));
    LocalMux I__2133 (
            .O(N__14693),
            .I(n14));
    InMux I__2132 (
            .O(N__14690),
            .I(n3496));
    InMux I__2131 (
            .O(N__14687),
            .I(N__14684));
    LocalMux I__2130 (
            .O(N__14684),
            .I(n13));
    InMux I__2129 (
            .O(N__14681),
            .I(n3497));
    InMux I__2128 (
            .O(N__14678),
            .I(N__14675));
    LocalMux I__2127 (
            .O(N__14675),
            .I(n12));
    InMux I__2126 (
            .O(N__14672),
            .I(n3498));
    InMux I__2125 (
            .O(N__14669),
            .I(N__14666));
    LocalMux I__2124 (
            .O(N__14666),
            .I(n11));
    InMux I__2123 (
            .O(N__14663),
            .I(n3499));
    InMux I__2122 (
            .O(N__14660),
            .I(N__14657));
    LocalMux I__2121 (
            .O(N__14657),
            .I(n10));
    InMux I__2120 (
            .O(N__14654),
            .I(bfn_5_31_0_));
    InMux I__2119 (
            .O(N__14651),
            .I(N__14648));
    LocalMux I__2118 (
            .O(N__14648),
            .I(n9));
    InMux I__2117 (
            .O(N__14645),
            .I(n3501));
    InMux I__2116 (
            .O(N__14642),
            .I(N__14639));
    LocalMux I__2115 (
            .O(N__14639),
            .I(n8));
    InMux I__2114 (
            .O(N__14636),
            .I(n3502));
    InMux I__2113 (
            .O(N__14633),
            .I(N__14630));
    LocalMux I__2112 (
            .O(N__14630),
            .I(n23));
    InMux I__2111 (
            .O(N__14627),
            .I(n3487));
    InMux I__2110 (
            .O(N__14624),
            .I(N__14621));
    LocalMux I__2109 (
            .O(N__14621),
            .I(n22));
    InMux I__2108 (
            .O(N__14618),
            .I(n3488));
    InMux I__2107 (
            .O(N__14615),
            .I(N__14612));
    LocalMux I__2106 (
            .O(N__14612),
            .I(n21));
    InMux I__2105 (
            .O(N__14609),
            .I(n3489));
    InMux I__2104 (
            .O(N__14606),
            .I(N__14603));
    LocalMux I__2103 (
            .O(N__14603),
            .I(n20));
    InMux I__2102 (
            .O(N__14600),
            .I(n3490));
    InMux I__2101 (
            .O(N__14597),
            .I(N__14594));
    LocalMux I__2100 (
            .O(N__14594),
            .I(n19));
    InMux I__2099 (
            .O(N__14591),
            .I(n3491));
    InMux I__2098 (
            .O(N__14588),
            .I(N__14585));
    LocalMux I__2097 (
            .O(N__14585),
            .I(n18));
    InMux I__2096 (
            .O(N__14582),
            .I(bfn_5_30_0_));
    InMux I__2095 (
            .O(N__14579),
            .I(N__14576));
    LocalMux I__2094 (
            .O(N__14576),
            .I(n17));
    InMux I__2093 (
            .O(N__14573),
            .I(n3493));
    InMux I__2092 (
            .O(N__14570),
            .I(N__14567));
    LocalMux I__2091 (
            .O(N__14567),
            .I(n16));
    InMux I__2090 (
            .O(N__14564),
            .I(n3494));
    CascadeMux I__2089 (
            .O(N__14561),
            .I(N__14558));
    InMux I__2088 (
            .O(N__14558),
            .I(N__14553));
    InMux I__2087 (
            .O(N__14557),
            .I(N__14550));
    CascadeMux I__2086 (
            .O(N__14556),
            .I(N__14547));
    LocalMux I__2085 (
            .O(N__14553),
            .I(N__14544));
    LocalMux I__2084 (
            .O(N__14550),
            .I(N__14541));
    InMux I__2083 (
            .O(N__14547),
            .I(N__14538));
    Odrv4 I__2082 (
            .O(N__14544),
            .I(\eeprom.n2115 ));
    Odrv12 I__2081 (
            .O(N__14541),
            .I(\eeprom.n2115 ));
    LocalMux I__2080 (
            .O(N__14538),
            .I(\eeprom.n2115 ));
    InMux I__2079 (
            .O(N__14531),
            .I(N__14528));
    LocalMux I__2078 (
            .O(N__14528),
            .I(N__14525));
    Odrv4 I__2077 (
            .O(N__14525),
            .I(\eeprom.n2182 ));
    InMux I__2076 (
            .O(N__14522),
            .I(\eeprom.n3535 ));
    InMux I__2075 (
            .O(N__14519),
            .I(N__14516));
    LocalMux I__2074 (
            .O(N__14516),
            .I(N__14512));
    InMux I__2073 (
            .O(N__14515),
            .I(N__14509));
    Span4Mux_v I__2072 (
            .O(N__14512),
            .I(N__14506));
    LocalMux I__2071 (
            .O(N__14509),
            .I(N__14503));
    Span4Mux_v I__2070 (
            .O(N__14506),
            .I(N__14500));
    Span4Mux_v I__2069 (
            .O(N__14503),
            .I(N__14497));
    Odrv4 I__2068 (
            .O(N__14500),
            .I(\eeprom.n2114 ));
    Odrv4 I__2067 (
            .O(N__14497),
            .I(\eeprom.n2114 ));
    InMux I__2066 (
            .O(N__14492),
            .I(N__14489));
    LocalMux I__2065 (
            .O(N__14489),
            .I(\eeprom.n2181 ));
    InMux I__2064 (
            .O(N__14486),
            .I(\eeprom.n3536 ));
    InMux I__2063 (
            .O(N__14483),
            .I(\eeprom.n3537 ));
    CascadeMux I__2062 (
            .O(N__14480),
            .I(N__14475));
    InMux I__2061 (
            .O(N__14479),
            .I(N__14470));
    InMux I__2060 (
            .O(N__14478),
            .I(N__14470));
    InMux I__2059 (
            .O(N__14475),
            .I(N__14467));
    LocalMux I__2058 (
            .O(N__14470),
            .I(N__14462));
    LocalMux I__2057 (
            .O(N__14467),
            .I(N__14462));
    Span4Mux_v I__2056 (
            .O(N__14462),
            .I(N__14459));
    Odrv4 I__2055 (
            .O(N__14459),
            .I(\eeprom.n2112 ));
    CascadeMux I__2054 (
            .O(N__14456),
            .I(N__14453));
    InMux I__2053 (
            .O(N__14453),
            .I(N__14450));
    LocalMux I__2052 (
            .O(N__14450),
            .I(\eeprom.n2179 ));
    InMux I__2051 (
            .O(N__14447),
            .I(\eeprom.n3538 ));
    CascadeMux I__2050 (
            .O(N__14444),
            .I(N__14441));
    InMux I__2049 (
            .O(N__14441),
            .I(N__14437));
    InMux I__2048 (
            .O(N__14440),
            .I(N__14433));
    LocalMux I__2047 (
            .O(N__14437),
            .I(N__14430));
    InMux I__2046 (
            .O(N__14436),
            .I(N__14427));
    LocalMux I__2045 (
            .O(N__14433),
            .I(N__14424));
    Span4Mux_v I__2044 (
            .O(N__14430),
            .I(N__14419));
    LocalMux I__2043 (
            .O(N__14427),
            .I(N__14419));
    Odrv4 I__2042 (
            .O(N__14424),
            .I(\eeprom.n2111 ));
    Odrv4 I__2041 (
            .O(N__14419),
            .I(\eeprom.n2111 ));
    InMux I__2040 (
            .O(N__14414),
            .I(N__14411));
    LocalMux I__2039 (
            .O(N__14411),
            .I(N__14408));
    Odrv4 I__2038 (
            .O(N__14408),
            .I(\eeprom.n2178 ));
    InMux I__2037 (
            .O(N__14405),
            .I(bfn_5_28_0_));
    InMux I__2036 (
            .O(N__14402),
            .I(N__14399));
    LocalMux I__2035 (
            .O(N__14399),
            .I(N__14395));
    InMux I__2034 (
            .O(N__14398),
            .I(N__14392));
    Span4Mux_v I__2033 (
            .O(N__14395),
            .I(N__14387));
    LocalMux I__2032 (
            .O(N__14392),
            .I(N__14387));
    Span4Mux_v I__2031 (
            .O(N__14387),
            .I(N__14384));
    Odrv4 I__2030 (
            .O(N__14384),
            .I(\eeprom.n2110 ));
    InMux I__2029 (
            .O(N__14381),
            .I(\eeprom.n3540 ));
    InMux I__2028 (
            .O(N__14378),
            .I(N__14375));
    LocalMux I__2027 (
            .O(N__14375),
            .I(n26));
    InMux I__2026 (
            .O(N__14372),
            .I(bfn_5_29_0_));
    InMux I__2025 (
            .O(N__14369),
            .I(N__14366));
    LocalMux I__2024 (
            .O(N__14366),
            .I(n25));
    InMux I__2023 (
            .O(N__14363),
            .I(n3485));
    InMux I__2022 (
            .O(N__14360),
            .I(N__14357));
    LocalMux I__2021 (
            .O(N__14357),
            .I(n24));
    InMux I__2020 (
            .O(N__14354),
            .I(n3486));
    CascadeMux I__2019 (
            .O(N__14351),
            .I(\eeprom.n2143_cascade_ ));
    InMux I__2018 (
            .O(N__14348),
            .I(bfn_5_27_0_));
    CascadeMux I__2017 (
            .O(N__14345),
            .I(N__14340));
    InMux I__2016 (
            .O(N__14344),
            .I(N__14335));
    InMux I__2015 (
            .O(N__14343),
            .I(N__14335));
    InMux I__2014 (
            .O(N__14340),
            .I(N__14332));
    LocalMux I__2013 (
            .O(N__14335),
            .I(N__14327));
    LocalMux I__2012 (
            .O(N__14332),
            .I(N__14327));
    Odrv12 I__2011 (
            .O(N__14327),
            .I(\eeprom.n2118 ));
    InMux I__2010 (
            .O(N__14324),
            .I(N__14321));
    LocalMux I__2009 (
            .O(N__14321),
            .I(\eeprom.n2185 ));
    InMux I__2008 (
            .O(N__14318),
            .I(\eeprom.n3532 ));
    CascadeMux I__2007 (
            .O(N__14315),
            .I(N__14311));
    CascadeMux I__2006 (
            .O(N__14314),
            .I(N__14308));
    InMux I__2005 (
            .O(N__14311),
            .I(N__14305));
    InMux I__2004 (
            .O(N__14308),
            .I(N__14302));
    LocalMux I__2003 (
            .O(N__14305),
            .I(N__14299));
    LocalMux I__2002 (
            .O(N__14302),
            .I(N__14296));
    Span4Mux_v I__2001 (
            .O(N__14299),
            .I(N__14290));
    Span4Mux_v I__2000 (
            .O(N__14296),
            .I(N__14290));
    InMux I__1999 (
            .O(N__14295),
            .I(N__14287));
    Odrv4 I__1998 (
            .O(N__14290),
            .I(\eeprom.n2117 ));
    LocalMux I__1997 (
            .O(N__14287),
            .I(\eeprom.n2117 ));
    InMux I__1996 (
            .O(N__14282),
            .I(N__14279));
    LocalMux I__1995 (
            .O(N__14279),
            .I(\eeprom.n2184 ));
    InMux I__1994 (
            .O(N__14276),
            .I(\eeprom.n3533 ));
    CascadeMux I__1993 (
            .O(N__14273),
            .I(N__14269));
    InMux I__1992 (
            .O(N__14272),
            .I(N__14266));
    InMux I__1991 (
            .O(N__14269),
            .I(N__14263));
    LocalMux I__1990 (
            .O(N__14266),
            .I(N__14257));
    LocalMux I__1989 (
            .O(N__14263),
            .I(N__14257));
    InMux I__1988 (
            .O(N__14262),
            .I(N__14254));
    Odrv12 I__1987 (
            .O(N__14257),
            .I(\eeprom.n2116 ));
    LocalMux I__1986 (
            .O(N__14254),
            .I(\eeprom.n2116 ));
    InMux I__1985 (
            .O(N__14249),
            .I(N__14246));
    LocalMux I__1984 (
            .O(N__14246),
            .I(N__14242));
    InMux I__1983 (
            .O(N__14245),
            .I(N__14239));
    Odrv4 I__1982 (
            .O(N__14242),
            .I(\eeprom.n2183 ));
    LocalMux I__1981 (
            .O(N__14239),
            .I(\eeprom.n2183 ));
    InMux I__1980 (
            .O(N__14234),
            .I(\eeprom.n3534 ));
    CascadeMux I__1979 (
            .O(N__14231),
            .I(\eeprom.n2214_cascade_ ));
    InMux I__1978 (
            .O(N__14228),
            .I(N__14225));
    LocalMux I__1977 (
            .O(N__14225),
            .I(N__14221));
    InMux I__1976 (
            .O(N__14224),
            .I(N__14218));
    Span4Mux_v I__1975 (
            .O(N__14221),
            .I(N__14215));
    LocalMux I__1974 (
            .O(N__14218),
            .I(\eeprom.n2313 ));
    Odrv4 I__1973 (
            .O(N__14215),
            .I(\eeprom.n2313 ));
    CascadeMux I__1972 (
            .O(N__14210),
            .I(\eeprom.n2313_cascade_ ));
    InMux I__1971 (
            .O(N__14207),
            .I(N__14204));
    LocalMux I__1970 (
            .O(N__14204),
            .I(\eeprom.n4505 ));
    InMux I__1969 (
            .O(N__14201),
            .I(N__14198));
    LocalMux I__1968 (
            .O(N__14198),
            .I(N__14195));
    Span4Mux_h I__1967 (
            .O(N__14195),
            .I(N__14192));
    Odrv4 I__1966 (
            .O(N__14192),
            .I(\eeprom.n11 ));
    InMux I__1965 (
            .O(N__14189),
            .I(N__14186));
    LocalMux I__1964 (
            .O(N__14186),
            .I(N__14182));
    InMux I__1963 (
            .O(N__14185),
            .I(N__14179));
    Span4Mux_v I__1962 (
            .O(N__14182),
            .I(N__14175));
    LocalMux I__1961 (
            .O(N__14179),
            .I(N__14172));
    InMux I__1960 (
            .O(N__14178),
            .I(N__14169));
    Span4Mux_h I__1959 (
            .O(N__14175),
            .I(N__14164));
    Span4Mux_v I__1958 (
            .O(N__14172),
            .I(N__14164));
    LocalMux I__1957 (
            .O(N__14169),
            .I(\eeprom.delay_counter_22 ));
    Odrv4 I__1956 (
            .O(N__14164),
            .I(\eeprom.delay_counter_22 ));
    CascadeMux I__1955 (
            .O(N__14159),
            .I(N__14156));
    InMux I__1954 (
            .O(N__14156),
            .I(N__14152));
    CascadeMux I__1953 (
            .O(N__14155),
            .I(N__14149));
    LocalMux I__1952 (
            .O(N__14152),
            .I(N__14146));
    InMux I__1951 (
            .O(N__14149),
            .I(N__14142));
    Span4Mux_h I__1950 (
            .O(N__14146),
            .I(N__14139));
    InMux I__1949 (
            .O(N__14145),
            .I(N__14136));
    LocalMux I__1948 (
            .O(N__14142),
            .I(\eeprom.n2315 ));
    Odrv4 I__1947 (
            .O(N__14139),
            .I(\eeprom.n2315 ));
    LocalMux I__1946 (
            .O(N__14136),
            .I(\eeprom.n2315 ));
    CascadeMux I__1945 (
            .O(N__14129),
            .I(N__14124));
    CascadeMux I__1944 (
            .O(N__14128),
            .I(N__14121));
    InMux I__1943 (
            .O(N__14127),
            .I(N__14118));
    InMux I__1942 (
            .O(N__14124),
            .I(N__14115));
    InMux I__1941 (
            .O(N__14121),
            .I(N__14112));
    LocalMux I__1940 (
            .O(N__14118),
            .I(N__14109));
    LocalMux I__1939 (
            .O(N__14115),
            .I(N__14104));
    LocalMux I__1938 (
            .O(N__14112),
            .I(N__14104));
    Span4Mux_s3_h I__1937 (
            .O(N__14109),
            .I(N__14099));
    Span4Mux_v I__1936 (
            .O(N__14104),
            .I(N__14099));
    Odrv4 I__1935 (
            .O(N__14099),
            .I(\eeprom.n2311 ));
    CascadeMux I__1934 (
            .O(N__14096),
            .I(N__14093));
    InMux I__1933 (
            .O(N__14093),
            .I(N__14090));
    LocalMux I__1932 (
            .O(N__14090),
            .I(N__14087));
    Odrv4 I__1931 (
            .O(N__14087),
            .I(\eeprom.n4461 ));
    InMux I__1930 (
            .O(N__14084),
            .I(N__14081));
    LocalMux I__1929 (
            .O(N__14081),
            .I(N__14078));
    Odrv12 I__1928 (
            .O(N__14078),
            .I(\eeprom.n4463 ));
    CascadeMux I__1927 (
            .O(N__14075),
            .I(\eeprom.n4225_cascade_ ));
    InMux I__1926 (
            .O(N__14072),
            .I(N__14069));
    LocalMux I__1925 (
            .O(N__14069),
            .I(N__14065));
    InMux I__1924 (
            .O(N__14068),
            .I(N__14061));
    Span12Mux_s10_v I__1923 (
            .O(N__14065),
            .I(N__14058));
    InMux I__1922 (
            .O(N__14064),
            .I(N__14055));
    LocalMux I__1921 (
            .O(N__14061),
            .I(N__14052));
    Odrv12 I__1920 (
            .O(N__14058),
            .I(\eeprom.n2019 ));
    LocalMux I__1919 (
            .O(N__14055),
            .I(\eeprom.n2019 ));
    Odrv12 I__1918 (
            .O(N__14052),
            .I(\eeprom.n2019 ));
    CascadeMux I__1917 (
            .O(N__14045),
            .I(N__14042));
    InMux I__1916 (
            .O(N__14042),
            .I(N__14039));
    LocalMux I__1915 (
            .O(N__14039),
            .I(\eeprom.n2086 ));
    InMux I__1914 (
            .O(N__14036),
            .I(N__14031));
    CascadeMux I__1913 (
            .O(N__14035),
            .I(N__14028));
    InMux I__1912 (
            .O(N__14034),
            .I(N__14025));
    LocalMux I__1911 (
            .O(N__14031),
            .I(N__14022));
    InMux I__1910 (
            .O(N__14028),
            .I(N__14019));
    LocalMux I__1909 (
            .O(N__14025),
            .I(\eeprom.n2309 ));
    Odrv4 I__1908 (
            .O(N__14022),
            .I(\eeprom.n2309 ));
    LocalMux I__1907 (
            .O(N__14019),
            .I(\eeprom.n2309 ));
    InMux I__1906 (
            .O(N__14012),
            .I(N__14008));
    InMux I__1905 (
            .O(N__14011),
            .I(N__14005));
    LocalMux I__1904 (
            .O(N__14008),
            .I(N__14001));
    LocalMux I__1903 (
            .O(N__14005),
            .I(N__13998));
    InMux I__1902 (
            .O(N__14004),
            .I(N__13995));
    Odrv4 I__1901 (
            .O(N__14001),
            .I(\eeprom.n2319 ));
    Odrv4 I__1900 (
            .O(N__13998),
            .I(\eeprom.n2319 ));
    LocalMux I__1899 (
            .O(N__13995),
            .I(\eeprom.n2319 ));
    CascadeMux I__1898 (
            .O(N__13988),
            .I(\eeprom.n4509_cascade_ ));
    InMux I__1897 (
            .O(N__13985),
            .I(N__13982));
    LocalMux I__1896 (
            .O(N__13982),
            .I(\eeprom.n8_adj_468 ));
    InMux I__1895 (
            .O(N__13979),
            .I(N__13975));
    InMux I__1894 (
            .O(N__13978),
            .I(N__13971));
    LocalMux I__1893 (
            .O(N__13975),
            .I(N__13968));
    InMux I__1892 (
            .O(N__13974),
            .I(N__13965));
    LocalMux I__1891 (
            .O(N__13971),
            .I(\eeprom.n2310 ));
    Odrv4 I__1890 (
            .O(N__13968),
            .I(\eeprom.n2310 ));
    LocalMux I__1889 (
            .O(N__13965),
            .I(\eeprom.n2310 ));
    CascadeMux I__1888 (
            .O(N__13958),
            .I(\eeprom.n6_cascade_ ));
    CascadeMux I__1887 (
            .O(N__13955),
            .I(\eeprom.n2242_cascade_ ));
    InMux I__1886 (
            .O(N__13952),
            .I(N__13946));
    CascadeMux I__1885 (
            .O(N__13951),
            .I(N__13943));
    CascadeMux I__1884 (
            .O(N__13950),
            .I(N__13940));
    CascadeMux I__1883 (
            .O(N__13949),
            .I(N__13932));
    LocalMux I__1882 (
            .O(N__13946),
            .I(N__13928));
    InMux I__1881 (
            .O(N__13943),
            .I(N__13917));
    InMux I__1880 (
            .O(N__13940),
            .I(N__13917));
    InMux I__1879 (
            .O(N__13939),
            .I(N__13917));
    InMux I__1878 (
            .O(N__13938),
            .I(N__13917));
    InMux I__1877 (
            .O(N__13937),
            .I(N__13917));
    InMux I__1876 (
            .O(N__13936),
            .I(N__13908));
    InMux I__1875 (
            .O(N__13935),
            .I(N__13908));
    InMux I__1874 (
            .O(N__13932),
            .I(N__13908));
    InMux I__1873 (
            .O(N__13931),
            .I(N__13908));
    Odrv4 I__1872 (
            .O(N__13928),
            .I(\eeprom.n2044 ));
    LocalMux I__1871 (
            .O(N__13917),
            .I(\eeprom.n2044 ));
    LocalMux I__1870 (
            .O(N__13908),
            .I(\eeprom.n2044 ));
    InMux I__1869 (
            .O(N__13901),
            .I(N__13898));
    LocalMux I__1868 (
            .O(N__13898),
            .I(N__13894));
    InMux I__1867 (
            .O(N__13897),
            .I(N__13891));
    Odrv4 I__1866 (
            .O(N__13894),
            .I(\eeprom.n2084 ));
    LocalMux I__1865 (
            .O(N__13891),
            .I(\eeprom.n2084 ));
    CascadeMux I__1864 (
            .O(N__13886),
            .I(N__13881));
    CascadeMux I__1863 (
            .O(N__13885),
            .I(N__13878));
    InMux I__1862 (
            .O(N__13884),
            .I(N__13875));
    InMux I__1861 (
            .O(N__13881),
            .I(N__13872));
    InMux I__1860 (
            .O(N__13878),
            .I(N__13869));
    LocalMux I__1859 (
            .O(N__13875),
            .I(\eeprom.n2013 ));
    LocalMux I__1858 (
            .O(N__13872),
            .I(\eeprom.n2013 ));
    LocalMux I__1857 (
            .O(N__13869),
            .I(\eeprom.n2013 ));
    CascadeMux I__1856 (
            .O(N__13862),
            .I(N__13859));
    InMux I__1855 (
            .O(N__13859),
            .I(N__13856));
    LocalMux I__1854 (
            .O(N__13856),
            .I(\eeprom.n2080 ));
    InMux I__1853 (
            .O(N__13853),
            .I(\eeprom.n3529 ));
    InMux I__1852 (
            .O(N__13850),
            .I(\eeprom.n3530 ));
    InMux I__1851 (
            .O(N__13847),
            .I(N__13844));
    LocalMux I__1850 (
            .O(N__13844),
            .I(N__13840));
    InMux I__1849 (
            .O(N__13843),
            .I(N__13837));
    Span4Mux_v I__1848 (
            .O(N__13840),
            .I(N__13834));
    LocalMux I__1847 (
            .O(N__13837),
            .I(N__13831));
    Odrv4 I__1846 (
            .O(N__13834),
            .I(\eeprom.n2011 ));
    Odrv4 I__1845 (
            .O(N__13831),
            .I(\eeprom.n2011 ));
    InMux I__1844 (
            .O(N__13826),
            .I(bfn_5_23_0_));
    InMux I__1843 (
            .O(N__13823),
            .I(N__13820));
    LocalMux I__1842 (
            .O(N__13820),
            .I(\eeprom.n2081 ));
    CascadeMux I__1841 (
            .O(N__13817),
            .I(N__13814));
    InMux I__1840 (
            .O(N__13814),
            .I(N__13810));
    CascadeMux I__1839 (
            .O(N__13813),
            .I(N__13807));
    LocalMux I__1838 (
            .O(N__13810),
            .I(N__13804));
    InMux I__1837 (
            .O(N__13807),
            .I(N__13801));
    Odrv4 I__1836 (
            .O(N__13804),
            .I(\eeprom.n2014 ));
    LocalMux I__1835 (
            .O(N__13801),
            .I(\eeprom.n2014 ));
    InMux I__1834 (
            .O(N__13796),
            .I(N__13793));
    LocalMux I__1833 (
            .O(N__13793),
            .I(N__13788));
    InMux I__1832 (
            .O(N__13792),
            .I(N__13785));
    InMux I__1831 (
            .O(N__13791),
            .I(N__13782));
    Span4Mux_h I__1830 (
            .O(N__13788),
            .I(N__13777));
    LocalMux I__1829 (
            .O(N__13785),
            .I(N__13777));
    LocalMux I__1828 (
            .O(N__13782),
            .I(\eeprom.n2012 ));
    Odrv4 I__1827 (
            .O(N__13777),
            .I(\eeprom.n2012 ));
    InMux I__1826 (
            .O(N__13772),
            .I(N__13769));
    LocalMux I__1825 (
            .O(N__13769),
            .I(\eeprom.n2079 ));
    InMux I__1824 (
            .O(N__13766),
            .I(N__13763));
    LocalMux I__1823 (
            .O(N__13763),
            .I(\eeprom.n2083 ));
    CascadeMux I__1822 (
            .O(N__13760),
            .I(N__13757));
    InMux I__1821 (
            .O(N__13757),
            .I(N__13753));
    CascadeMux I__1820 (
            .O(N__13756),
            .I(N__13750));
    LocalMux I__1819 (
            .O(N__13753),
            .I(N__13747));
    InMux I__1818 (
            .O(N__13750),
            .I(N__13744));
    Span4Mux_v I__1817 (
            .O(N__13747),
            .I(N__13738));
    LocalMux I__1816 (
            .O(N__13744),
            .I(N__13738));
    InMux I__1815 (
            .O(N__13743),
            .I(N__13735));
    Odrv4 I__1814 (
            .O(N__13738),
            .I(\eeprom.n2016 ));
    LocalMux I__1813 (
            .O(N__13735),
            .I(\eeprom.n2016 ));
    InMux I__1812 (
            .O(N__13730),
            .I(N__13727));
    LocalMux I__1811 (
            .O(N__13727),
            .I(\eeprom.n7_adj_470 ));
    InMux I__1810 (
            .O(N__13724),
            .I(N__13721));
    LocalMux I__1809 (
            .O(N__13721),
            .I(N__13716));
    InMux I__1808 (
            .O(N__13720),
            .I(N__13713));
    InMux I__1807 (
            .O(N__13719),
            .I(N__13710));
    Span4Mux_v I__1806 (
            .O(N__13716),
            .I(N__13705));
    LocalMux I__1805 (
            .O(N__13713),
            .I(N__13705));
    LocalMux I__1804 (
            .O(N__13710),
            .I(N__13702));
    Span4Mux_h I__1803 (
            .O(N__13705),
            .I(N__13699));
    Odrv4 I__1802 (
            .O(N__13702),
            .I(\eeprom.n2419 ));
    Odrv4 I__1801 (
            .O(N__13699),
            .I(\eeprom.n2419 ));
    InMux I__1800 (
            .O(N__13694),
            .I(N__13691));
    LocalMux I__1799 (
            .O(N__13691),
            .I(N__13688));
    Span4Mux_v I__1798 (
            .O(N__13688),
            .I(N__13685));
    Odrv4 I__1797 (
            .O(N__13685),
            .I(\eeprom.n2486 ));
    InMux I__1796 (
            .O(N__13682),
            .I(bfn_5_22_0_));
    CascadeMux I__1795 (
            .O(N__13679),
            .I(N__13675));
    InMux I__1794 (
            .O(N__13678),
            .I(N__13671));
    InMux I__1793 (
            .O(N__13675),
            .I(N__13668));
    InMux I__1792 (
            .O(N__13674),
            .I(N__13665));
    LocalMux I__1791 (
            .O(N__13671),
            .I(\eeprom.n2018 ));
    LocalMux I__1790 (
            .O(N__13668),
            .I(\eeprom.n2018 ));
    LocalMux I__1789 (
            .O(N__13665),
            .I(\eeprom.n2018 ));
    CascadeMux I__1788 (
            .O(N__13658),
            .I(N__13655));
    InMux I__1787 (
            .O(N__13655),
            .I(N__13652));
    LocalMux I__1786 (
            .O(N__13652),
            .I(\eeprom.n2085 ));
    InMux I__1785 (
            .O(N__13649),
            .I(\eeprom.n3524 ));
    InMux I__1784 (
            .O(N__13646),
            .I(\eeprom.n3525 ));
    InMux I__1783 (
            .O(N__13643),
            .I(\eeprom.n3526 ));
    CascadeMux I__1782 (
            .O(N__13640),
            .I(N__13637));
    InMux I__1781 (
            .O(N__13637),
            .I(N__13633));
    InMux I__1780 (
            .O(N__13636),
            .I(N__13629));
    LocalMux I__1779 (
            .O(N__13633),
            .I(N__13626));
    InMux I__1778 (
            .O(N__13632),
            .I(N__13623));
    LocalMux I__1777 (
            .O(N__13629),
            .I(\eeprom.n2015 ));
    Odrv4 I__1776 (
            .O(N__13626),
            .I(\eeprom.n2015 ));
    LocalMux I__1775 (
            .O(N__13623),
            .I(\eeprom.n2015 ));
    CascadeMux I__1774 (
            .O(N__13616),
            .I(N__13613));
    InMux I__1773 (
            .O(N__13613),
            .I(N__13610));
    LocalMux I__1772 (
            .O(N__13610),
            .I(\eeprom.n2082 ));
    InMux I__1771 (
            .O(N__13607),
            .I(\eeprom.n3527 ));
    InMux I__1770 (
            .O(N__13604),
            .I(\eeprom.n3528 ));
    CascadeMux I__1769 (
            .O(N__13601),
            .I(\eeprom.n13_adj_474_cascade_ ));
    InMux I__1768 (
            .O(N__13598),
            .I(N__13595));
    LocalMux I__1767 (
            .O(N__13595),
            .I(\eeprom.n11_adj_473 ));
    CascadeMux I__1766 (
            .O(N__13592),
            .I(\eeprom.n2539_cascade_ ));
    InMux I__1765 (
            .O(N__13589),
            .I(N__13586));
    LocalMux I__1764 (
            .O(N__13586),
            .I(N__13581));
    InMux I__1763 (
            .O(N__13585),
            .I(N__13578));
    InMux I__1762 (
            .O(N__13584),
            .I(N__13575));
    Span4Mux_h I__1761 (
            .O(N__13581),
            .I(N__13570));
    LocalMux I__1760 (
            .O(N__13578),
            .I(N__13570));
    LocalMux I__1759 (
            .O(N__13575),
            .I(N__13565));
    Span4Mux_v I__1758 (
            .O(N__13570),
            .I(N__13565));
    Odrv4 I__1757 (
            .O(N__13565),
            .I(\eeprom.delay_counter_14 ));
    CascadeMux I__1756 (
            .O(N__13562),
            .I(N__13559));
    InMux I__1755 (
            .O(N__13559),
            .I(N__13556));
    LocalMux I__1754 (
            .O(N__13556),
            .I(N__13553));
    Span4Mux_h I__1753 (
            .O(N__13553),
            .I(N__13550));
    Odrv4 I__1752 (
            .O(N__13550),
            .I(\eeprom.n19_adj_429 ));
    InMux I__1751 (
            .O(N__13547),
            .I(N__13544));
    LocalMux I__1750 (
            .O(N__13544),
            .I(N__13541));
    Odrv12 I__1749 (
            .O(N__13541),
            .I(\eeprom.n30 ));
    CascadeMux I__1748 (
            .O(N__13538),
            .I(\eeprom.n2114_cascade_ ));
    InMux I__1747 (
            .O(N__13535),
            .I(N__13532));
    LocalMux I__1746 (
            .O(N__13532),
            .I(N__13528));
    InMux I__1745 (
            .O(N__13531),
            .I(N__13525));
    Span4Mux_v I__1744 (
            .O(N__13528),
            .I(N__13520));
    LocalMux I__1743 (
            .O(N__13525),
            .I(N__13520));
    Odrv4 I__1742 (
            .O(N__13520),
            .I(\eeprom.n2411 ));
    InMux I__1741 (
            .O(N__13517),
            .I(N__13514));
    LocalMux I__1740 (
            .O(N__13514),
            .I(N__13511));
    Span4Mux_v I__1739 (
            .O(N__13511),
            .I(N__13508));
    Odrv4 I__1738 (
            .O(N__13508),
            .I(\eeprom.n2478 ));
    InMux I__1737 (
            .O(N__13505),
            .I(N__13502));
    LocalMux I__1736 (
            .O(N__13502),
            .I(n4826));
    CascadeMux I__1735 (
            .O(N__13499),
            .I(n4825_cascade_));
    IoInMux I__1734 (
            .O(N__13496),
            .I(N__13493));
    LocalMux I__1733 (
            .O(N__13493),
            .I(N__13490));
    Odrv4 I__1732 (
            .O(N__13490),
            .I(LED_c));
    InMux I__1731 (
            .O(N__13487),
            .I(N__13484));
    LocalMux I__1730 (
            .O(N__13484),
            .I(N__13481));
    Span4Mux_h I__1729 (
            .O(N__13481),
            .I(N__13478));
    Odrv4 I__1728 (
            .O(N__13478),
            .I(\eeprom.n23_adj_464 ));
    InMux I__1727 (
            .O(N__13475),
            .I(N__13471));
    InMux I__1726 (
            .O(N__13474),
            .I(N__13467));
    LocalMux I__1725 (
            .O(N__13471),
            .I(N__13464));
    InMux I__1724 (
            .O(N__13470),
            .I(N__13461));
    LocalMux I__1723 (
            .O(N__13467),
            .I(\eeprom.delay_counter_10 ));
    Odrv4 I__1722 (
            .O(N__13464),
            .I(\eeprom.delay_counter_10 ));
    LocalMux I__1721 (
            .O(N__13461),
            .I(\eeprom.delay_counter_10 ));
    CascadeMux I__1720 (
            .O(N__13454),
            .I(\eeprom.n2615_cascade_ ));
    CascadeMux I__1719 (
            .O(N__13451),
            .I(\eeprom.n4497_cascade_ ));
    CascadeMux I__1718 (
            .O(N__13448),
            .I(\eeprom.n4501_cascade_ ));
    InMux I__1717 (
            .O(N__13445),
            .I(bfn_4_26_0_));
    InMux I__1716 (
            .O(N__13442),
            .I(\eeprom.n3570 ));
    InMux I__1715 (
            .O(N__13439),
            .I(\eeprom.n3571 ));
    InMux I__1714 (
            .O(N__13436),
            .I(\eeprom.n3572 ));
    InMux I__1713 (
            .O(N__13433),
            .I(N__13430));
    LocalMux I__1712 (
            .O(N__13430),
            .I(N__13426));
    InMux I__1711 (
            .O(N__13429),
            .I(N__13423));
    Odrv4 I__1710 (
            .O(N__13426),
            .I(\eeprom.n2407 ));
    LocalMux I__1709 (
            .O(N__13423),
            .I(\eeprom.n2407 ));
    InMux I__1708 (
            .O(N__13418),
            .I(\eeprom.n3573 ));
    InMux I__1707 (
            .O(N__13415),
            .I(N__13408));
    InMux I__1706 (
            .O(N__13414),
            .I(N__13408));
    InMux I__1705 (
            .O(N__13413),
            .I(N__13405));
    LocalMux I__1704 (
            .O(N__13408),
            .I(\eeprom.n2410 ));
    LocalMux I__1703 (
            .O(N__13405),
            .I(\eeprom.n2410 ));
    CascadeMux I__1702 (
            .O(N__13400),
            .I(N__13397));
    InMux I__1701 (
            .O(N__13397),
            .I(N__13394));
    LocalMux I__1700 (
            .O(N__13394),
            .I(\eeprom.n2477 ));
    InMux I__1699 (
            .O(N__13391),
            .I(N__13388));
    LocalMux I__1698 (
            .O(N__13388),
            .I(\eeprom.n2476 ));
    CascadeMux I__1697 (
            .O(N__13385),
            .I(N__13382));
    InMux I__1696 (
            .O(N__13382),
            .I(N__13376));
    InMux I__1695 (
            .O(N__13381),
            .I(N__13376));
    LocalMux I__1694 (
            .O(N__13376),
            .I(N__13372));
    InMux I__1693 (
            .O(N__13375),
            .I(N__13369));
    Odrv4 I__1692 (
            .O(N__13372),
            .I(\eeprom.n2409 ));
    LocalMux I__1691 (
            .O(N__13369),
            .I(\eeprom.n2409 ));
    InMux I__1690 (
            .O(N__13364),
            .I(bfn_4_25_0_));
    CascadeMux I__1689 (
            .O(N__13361),
            .I(N__13356));
    InMux I__1688 (
            .O(N__13360),
            .I(N__13351));
    InMux I__1687 (
            .O(N__13359),
            .I(N__13351));
    InMux I__1686 (
            .O(N__13356),
            .I(N__13348));
    LocalMux I__1685 (
            .O(N__13351),
            .I(\eeprom.n2418 ));
    LocalMux I__1684 (
            .O(N__13348),
            .I(\eeprom.n2418 ));
    CascadeMux I__1683 (
            .O(N__13343),
            .I(N__13340));
    InMux I__1682 (
            .O(N__13340),
            .I(N__13337));
    LocalMux I__1681 (
            .O(N__13337),
            .I(N__13334));
    Odrv4 I__1680 (
            .O(N__13334),
            .I(\eeprom.n2485 ));
    InMux I__1679 (
            .O(N__13331),
            .I(\eeprom.n3562 ));
    CascadeMux I__1678 (
            .O(N__13328),
            .I(N__13325));
    InMux I__1677 (
            .O(N__13325),
            .I(N__13321));
    InMux I__1676 (
            .O(N__13324),
            .I(N__13317));
    LocalMux I__1675 (
            .O(N__13321),
            .I(N__13314));
    InMux I__1674 (
            .O(N__13320),
            .I(N__13311));
    LocalMux I__1673 (
            .O(N__13317),
            .I(\eeprom.n2417 ));
    Odrv4 I__1672 (
            .O(N__13314),
            .I(\eeprom.n2417 ));
    LocalMux I__1671 (
            .O(N__13311),
            .I(\eeprom.n2417 ));
    CascadeMux I__1670 (
            .O(N__13304),
            .I(N__13301));
    InMux I__1669 (
            .O(N__13301),
            .I(N__13298));
    LocalMux I__1668 (
            .O(N__13298),
            .I(N__13295));
    Odrv4 I__1667 (
            .O(N__13295),
            .I(\eeprom.n2484 ));
    InMux I__1666 (
            .O(N__13292),
            .I(\eeprom.n3563 ));
    CascadeMux I__1665 (
            .O(N__13289),
            .I(N__13285));
    CascadeMux I__1664 (
            .O(N__13288),
            .I(N__13281));
    InMux I__1663 (
            .O(N__13285),
            .I(N__13278));
    InMux I__1662 (
            .O(N__13284),
            .I(N__13273));
    InMux I__1661 (
            .O(N__13281),
            .I(N__13273));
    LocalMux I__1660 (
            .O(N__13278),
            .I(\eeprom.n2416 ));
    LocalMux I__1659 (
            .O(N__13273),
            .I(\eeprom.n2416 ));
    InMux I__1658 (
            .O(N__13268),
            .I(N__13265));
    LocalMux I__1657 (
            .O(N__13265),
            .I(N__13262));
    Odrv4 I__1656 (
            .O(N__13262),
            .I(\eeprom.n2483 ));
    InMux I__1655 (
            .O(N__13259),
            .I(\eeprom.n3564 ));
    InMux I__1654 (
            .O(N__13256),
            .I(N__13251));
    CascadeMux I__1653 (
            .O(N__13255),
            .I(N__13248));
    InMux I__1652 (
            .O(N__13254),
            .I(N__13245));
    LocalMux I__1651 (
            .O(N__13251),
            .I(N__13242));
    InMux I__1650 (
            .O(N__13248),
            .I(N__13239));
    LocalMux I__1649 (
            .O(N__13245),
            .I(\eeprom.n2415 ));
    Odrv4 I__1648 (
            .O(N__13242),
            .I(\eeprom.n2415 ));
    LocalMux I__1647 (
            .O(N__13239),
            .I(\eeprom.n2415 ));
    CascadeMux I__1646 (
            .O(N__13232),
            .I(N__13229));
    InMux I__1645 (
            .O(N__13229),
            .I(N__13226));
    LocalMux I__1644 (
            .O(N__13226),
            .I(N__13223));
    Odrv4 I__1643 (
            .O(N__13223),
            .I(\eeprom.n2482 ));
    InMux I__1642 (
            .O(N__13220),
            .I(\eeprom.n3565 ));
    CascadeMux I__1641 (
            .O(N__13217),
            .I(N__13213));
    CascadeMux I__1640 (
            .O(N__13216),
            .I(N__13210));
    InMux I__1639 (
            .O(N__13213),
            .I(N__13206));
    InMux I__1638 (
            .O(N__13210),
            .I(N__13201));
    InMux I__1637 (
            .O(N__13209),
            .I(N__13201));
    LocalMux I__1636 (
            .O(N__13206),
            .I(\eeprom.n2414 ));
    LocalMux I__1635 (
            .O(N__13201),
            .I(\eeprom.n2414 ));
    InMux I__1634 (
            .O(N__13196),
            .I(N__13193));
    LocalMux I__1633 (
            .O(N__13193),
            .I(N__13190));
    Odrv4 I__1632 (
            .O(N__13190),
            .I(\eeprom.n2481 ));
    InMux I__1631 (
            .O(N__13187),
            .I(\eeprom.n3566 ));
    InMux I__1630 (
            .O(N__13184),
            .I(\eeprom.n3567 ));
    InMux I__1629 (
            .O(N__13181),
            .I(\eeprom.n3568 ));
    InMux I__1628 (
            .O(N__13178),
            .I(N__13175));
    LocalMux I__1627 (
            .O(N__13175),
            .I(\eeprom.n2376 ));
    InMux I__1626 (
            .O(N__13172),
            .I(N__13168));
    InMux I__1625 (
            .O(N__13171),
            .I(N__13165));
    LocalMux I__1624 (
            .O(N__13168),
            .I(\eeprom.n2312 ));
    LocalMux I__1623 (
            .O(N__13165),
            .I(\eeprom.n2312 ));
    CascadeMux I__1622 (
            .O(N__13160),
            .I(\eeprom.n2312_cascade_ ));
    InMux I__1621 (
            .O(N__13157),
            .I(N__13154));
    LocalMux I__1620 (
            .O(N__13154),
            .I(\eeprom.n2379 ));
    CascadeMux I__1619 (
            .O(N__13151),
            .I(\eeprom.n2411_cascade_ ));
    InMux I__1618 (
            .O(N__13148),
            .I(N__13145));
    LocalMux I__1617 (
            .O(N__13145),
            .I(\eeprom.n4133 ));
    CascadeMux I__1616 (
            .O(N__13142),
            .I(\eeprom.n12_adj_472_cascade_ ));
    InMux I__1615 (
            .O(N__13139),
            .I(N__13136));
    LocalMux I__1614 (
            .O(N__13136),
            .I(\eeprom.n2382 ));
    InMux I__1613 (
            .O(N__13133),
            .I(N__13130));
    LocalMux I__1612 (
            .O(N__13130),
            .I(\eeprom.n2377 ));
    CascadeMux I__1611 (
            .O(N__13127),
            .I(N__13124));
    InMux I__1610 (
            .O(N__13124),
            .I(N__13121));
    LocalMux I__1609 (
            .O(N__13121),
            .I(\eeprom.n2380 ));
    InMux I__1608 (
            .O(N__13118),
            .I(N__13110));
    CascadeMux I__1607 (
            .O(N__13117),
            .I(N__13107));
    CascadeMux I__1606 (
            .O(N__13116),
            .I(N__13104));
    CascadeMux I__1605 (
            .O(N__13115),
            .I(N__13097));
    CascadeMux I__1604 (
            .O(N__13114),
            .I(N__13094));
    CascadeMux I__1603 (
            .O(N__13113),
            .I(N__13091));
    LocalMux I__1602 (
            .O(N__13110),
            .I(N__13087));
    InMux I__1601 (
            .O(N__13107),
            .I(N__13076));
    InMux I__1600 (
            .O(N__13104),
            .I(N__13076));
    InMux I__1599 (
            .O(N__13103),
            .I(N__13076));
    InMux I__1598 (
            .O(N__13102),
            .I(N__13076));
    InMux I__1597 (
            .O(N__13101),
            .I(N__13076));
    InMux I__1596 (
            .O(N__13100),
            .I(N__13073));
    InMux I__1595 (
            .O(N__13097),
            .I(N__13064));
    InMux I__1594 (
            .O(N__13094),
            .I(N__13064));
    InMux I__1593 (
            .O(N__13091),
            .I(N__13064));
    InMux I__1592 (
            .O(N__13090),
            .I(N__13064));
    Odrv4 I__1591 (
            .O(N__13087),
            .I(\eeprom.n2341 ));
    LocalMux I__1590 (
            .O(N__13076),
            .I(\eeprom.n2341 ));
    LocalMux I__1589 (
            .O(N__13073),
            .I(\eeprom.n2341 ));
    LocalMux I__1588 (
            .O(N__13064),
            .I(\eeprom.n2341 ));
    InMux I__1587 (
            .O(N__13055),
            .I(N__13052));
    LocalMux I__1586 (
            .O(N__13052),
            .I(N__13047));
    InMux I__1585 (
            .O(N__13051),
            .I(N__13044));
    InMux I__1584 (
            .O(N__13050),
            .I(N__13041));
    Span4Mux_h I__1583 (
            .O(N__13047),
            .I(N__13036));
    LocalMux I__1582 (
            .O(N__13044),
            .I(N__13036));
    LocalMux I__1581 (
            .O(N__13041),
            .I(\eeprom.delay_counter_20 ));
    Odrv4 I__1580 (
            .O(N__13036),
            .I(\eeprom.delay_counter_20 ));
    CascadeMux I__1579 (
            .O(N__13031),
            .I(\eeprom.n4479_cascade_ ));
    InMux I__1578 (
            .O(N__13028),
            .I(N__13025));
    LocalMux I__1577 (
            .O(N__13025),
            .I(\eeprom.n4477 ));
    InMux I__1576 (
            .O(N__13022),
            .I(N__13019));
    LocalMux I__1575 (
            .O(N__13019),
            .I(\eeprom.n2385 ));
    CascadeMux I__1574 (
            .O(N__13016),
            .I(\eeprom.n2341_cascade_ ));
    InMux I__1573 (
            .O(N__13013),
            .I(N__13010));
    LocalMux I__1572 (
            .O(N__13010),
            .I(N__13006));
    InMux I__1571 (
            .O(N__13009),
            .I(N__13003));
    Odrv12 I__1570 (
            .O(N__13006),
            .I(\eeprom.n1915 ));
    LocalMux I__1569 (
            .O(N__13003),
            .I(\eeprom.n1915 ));
    CascadeMux I__1568 (
            .O(N__12998),
            .I(N__12995));
    InMux I__1567 (
            .O(N__12995),
            .I(N__12992));
    LocalMux I__1566 (
            .O(N__12992),
            .I(N__12989));
    Odrv4 I__1565 (
            .O(N__12989),
            .I(\eeprom.n1982 ));
    CascadeMux I__1564 (
            .O(N__12986),
            .I(\eeprom.n2014_cascade_ ));
    InMux I__1563 (
            .O(N__12983),
            .I(N__12980));
    LocalMux I__1562 (
            .O(N__12980),
            .I(\eeprom.n4415 ));
    InMux I__1561 (
            .O(N__12977),
            .I(N__12972));
    InMux I__1560 (
            .O(N__12976),
            .I(N__12969));
    InMux I__1559 (
            .O(N__12975),
            .I(N__12966));
    LocalMux I__1558 (
            .O(N__12972),
            .I(\eeprom.n1919 ));
    LocalMux I__1557 (
            .O(N__12969),
            .I(\eeprom.n1919 ));
    LocalMux I__1556 (
            .O(N__12966),
            .I(\eeprom.n1919 ));
    CascadeMux I__1555 (
            .O(N__12959),
            .I(N__12956));
    InMux I__1554 (
            .O(N__12956),
            .I(N__12953));
    LocalMux I__1553 (
            .O(N__12953),
            .I(N__12950));
    Odrv4 I__1552 (
            .O(N__12950),
            .I(\eeprom.n1986 ));
    InMux I__1551 (
            .O(N__12947),
            .I(N__12943));
    CascadeMux I__1550 (
            .O(N__12946),
            .I(N__12940));
    LocalMux I__1549 (
            .O(N__12943),
            .I(N__12937));
    InMux I__1548 (
            .O(N__12940),
            .I(N__12934));
    Odrv4 I__1547 (
            .O(N__12937),
            .I(\eeprom.n1913 ));
    LocalMux I__1546 (
            .O(N__12934),
            .I(\eeprom.n1913 ));
    CascadeMux I__1545 (
            .O(N__12929),
            .I(N__12923));
    CascadeMux I__1544 (
            .O(N__12928),
            .I(N__12920));
    CascadeMux I__1543 (
            .O(N__12927),
            .I(N__12917));
    CascadeMux I__1542 (
            .O(N__12926),
            .I(N__12912));
    InMux I__1541 (
            .O(N__12923),
            .I(N__12908));
    InMux I__1540 (
            .O(N__12920),
            .I(N__12899));
    InMux I__1539 (
            .O(N__12917),
            .I(N__12899));
    InMux I__1538 (
            .O(N__12916),
            .I(N__12899));
    InMux I__1537 (
            .O(N__12915),
            .I(N__12899));
    InMux I__1536 (
            .O(N__12912),
            .I(N__12894));
    InMux I__1535 (
            .O(N__12911),
            .I(N__12894));
    LocalMux I__1534 (
            .O(N__12908),
            .I(\eeprom.n1945 ));
    LocalMux I__1533 (
            .O(N__12899),
            .I(\eeprom.n1945 ));
    LocalMux I__1532 (
            .O(N__12894),
            .I(\eeprom.n1945 ));
    InMux I__1531 (
            .O(N__12887),
            .I(N__12884));
    LocalMux I__1530 (
            .O(N__12884),
            .I(N__12881));
    Odrv4 I__1529 (
            .O(N__12881),
            .I(\eeprom.n1980 ));
    InMux I__1528 (
            .O(N__12878),
            .I(N__12875));
    LocalMux I__1527 (
            .O(N__12875),
            .I(\eeprom.n4419 ));
    CascadeMux I__1526 (
            .O(N__12872),
            .I(\eeprom.n4575_cascade_ ));
    InMux I__1525 (
            .O(N__12869),
            .I(N__12866));
    LocalMux I__1524 (
            .O(N__12866),
            .I(\eeprom.n4579 ));
    InMux I__1523 (
            .O(N__12863),
            .I(N__12860));
    LocalMux I__1522 (
            .O(N__12860),
            .I(N__12857));
    Span4Mux_h I__1521 (
            .O(N__12857),
            .I(N__12854));
    Odrv4 I__1520 (
            .O(N__12854),
            .I(\eeprom.n13 ));
    InMux I__1519 (
            .O(N__12851),
            .I(\eeprom.n3523 ));
    InMux I__1518 (
            .O(N__12848),
            .I(N__12845));
    LocalMux I__1517 (
            .O(N__12845),
            .I(N__12842));
    Span4Mux_v I__1516 (
            .O(N__12842),
            .I(N__12839));
    Odrv4 I__1515 (
            .O(N__12839),
            .I(\eeprom.n26_adj_469 ));
    InMux I__1514 (
            .O(N__12836),
            .I(N__12833));
    LocalMux I__1513 (
            .O(N__12833),
            .I(N__12829));
    InMux I__1512 (
            .O(N__12832),
            .I(N__12825));
    Span4Mux_v I__1511 (
            .O(N__12829),
            .I(N__12822));
    InMux I__1510 (
            .O(N__12828),
            .I(N__12819));
    LocalMux I__1509 (
            .O(N__12825),
            .I(\eeprom.delay_counter_7 ));
    Odrv4 I__1508 (
            .O(N__12822),
            .I(\eeprom.delay_counter_7 ));
    LocalMux I__1507 (
            .O(N__12819),
            .I(\eeprom.delay_counter_7 ));
    CascadeMux I__1506 (
            .O(N__12812),
            .I(N__12809));
    InMux I__1505 (
            .O(N__12809),
            .I(N__12806));
    LocalMux I__1504 (
            .O(N__12806),
            .I(\eeprom.n1984 ));
    InMux I__1503 (
            .O(N__12803),
            .I(N__12800));
    LocalMux I__1502 (
            .O(N__12800),
            .I(\eeprom.n1985 ));
    CascadeMux I__1501 (
            .O(N__12797),
            .I(\eeprom.n2017_cascade_ ));
    CascadeMux I__1500 (
            .O(N__12794),
            .I(N__12789));
    InMux I__1499 (
            .O(N__12793),
            .I(N__12784));
    InMux I__1498 (
            .O(N__12792),
            .I(N__12784));
    InMux I__1497 (
            .O(N__12789),
            .I(N__12781));
    LocalMux I__1496 (
            .O(N__12784),
            .I(\eeprom.n1917 ));
    LocalMux I__1495 (
            .O(N__12781),
            .I(\eeprom.n1917 ));
    InMux I__1494 (
            .O(N__12776),
            .I(N__12773));
    LocalMux I__1493 (
            .O(N__12773),
            .I(N__12770));
    Odrv4 I__1492 (
            .O(N__12770),
            .I(\eeprom.n4437 ));
    CascadeMux I__1491 (
            .O(N__12767),
            .I(N__12762));
    InMux I__1490 (
            .O(N__12766),
            .I(N__12759));
    InMux I__1489 (
            .O(N__12765),
            .I(N__12756));
    InMux I__1488 (
            .O(N__12762),
            .I(N__12753));
    LocalMux I__1487 (
            .O(N__12759),
            .I(\eeprom.n1918 ));
    LocalMux I__1486 (
            .O(N__12756),
            .I(\eeprom.n1918 ));
    LocalMux I__1485 (
            .O(N__12753),
            .I(\eeprom.n1918 ));
    CascadeMux I__1484 (
            .O(N__12746),
            .I(\eeprom.n4441_cascade_ ));
    InMux I__1483 (
            .O(N__12743),
            .I(N__12739));
    InMux I__1482 (
            .O(N__12742),
            .I(N__12736));
    LocalMux I__1481 (
            .O(N__12739),
            .I(N__12733));
    LocalMux I__1480 (
            .O(N__12736),
            .I(\eeprom.n1912 ));
    Odrv4 I__1479 (
            .O(N__12733),
            .I(\eeprom.n1912 ));
    CascadeMux I__1478 (
            .O(N__12728),
            .I(N__12723));
    CascadeMux I__1477 (
            .O(N__12727),
            .I(N__12720));
    InMux I__1476 (
            .O(N__12726),
            .I(N__12715));
    InMux I__1475 (
            .O(N__12723),
            .I(N__12715));
    InMux I__1474 (
            .O(N__12720),
            .I(N__12712));
    LocalMux I__1473 (
            .O(N__12715),
            .I(N__12709));
    LocalMux I__1472 (
            .O(N__12712),
            .I(\eeprom.n1916 ));
    Odrv4 I__1471 (
            .O(N__12709),
            .I(\eeprom.n1916 ));
    CascadeMux I__1470 (
            .O(N__12704),
            .I(\eeprom.n1945_cascade_ ));
    InMux I__1469 (
            .O(N__12701),
            .I(N__12698));
    LocalMux I__1468 (
            .O(N__12698),
            .I(\eeprom.n1983 ));
    InMux I__1467 (
            .O(N__12695),
            .I(N__12692));
    LocalMux I__1466 (
            .O(N__12692),
            .I(N__12689));
    Odrv4 I__1465 (
            .O(N__12689),
            .I(\eeprom.n1981 ));
    CascadeMux I__1464 (
            .O(N__12686),
            .I(N__12682));
    InMux I__1463 (
            .O(N__12685),
            .I(N__12678));
    InMux I__1462 (
            .O(N__12682),
            .I(N__12675));
    InMux I__1461 (
            .O(N__12681),
            .I(N__12672));
    LocalMux I__1460 (
            .O(N__12678),
            .I(\eeprom.n1914 ));
    LocalMux I__1459 (
            .O(N__12675),
            .I(\eeprom.n1914 ));
    LocalMux I__1458 (
            .O(N__12672),
            .I(\eeprom.n1914 ));
    InMux I__1457 (
            .O(N__12665),
            .I(N__12662));
    LocalMux I__1456 (
            .O(N__12662),
            .I(N__12657));
    InMux I__1455 (
            .O(N__12661),
            .I(N__12654));
    InMux I__1454 (
            .O(N__12660),
            .I(N__12651));
    Span4Mux_v I__1453 (
            .O(N__12657),
            .I(N__12648));
    LocalMux I__1452 (
            .O(N__12654),
            .I(N__12645));
    LocalMux I__1451 (
            .O(N__12651),
            .I(N__12638));
    Span4Mux_h I__1450 (
            .O(N__12648),
            .I(N__12638));
    Span4Mux_v I__1449 (
            .O(N__12645),
            .I(N__12638));
    Odrv4 I__1448 (
            .O(N__12638),
            .I(\eeprom.delay_counter_17 ));
    InMux I__1447 (
            .O(N__12635),
            .I(N__12632));
    LocalMux I__1446 (
            .O(N__12632),
            .I(N__12629));
    Span4Mux_v I__1445 (
            .O(N__12629),
            .I(N__12626));
    Span4Mux_v I__1444 (
            .O(N__12626),
            .I(N__12623));
    Odrv4 I__1443 (
            .O(N__12623),
            .I(\eeprom.n16_adj_377 ));
    CascadeMux I__1442 (
            .O(N__12620),
            .I(N__12617));
    InMux I__1441 (
            .O(N__12617),
            .I(N__12611));
    InMux I__1440 (
            .O(N__12616),
            .I(N__12611));
    LocalMux I__1439 (
            .O(N__12611),
            .I(\eeprom.n4734 ));
    InMux I__1438 (
            .O(N__12608),
            .I(N__12602));
    CascadeMux I__1437 (
            .O(N__12607),
            .I(N__12595));
    InMux I__1436 (
            .O(N__12606),
            .I(N__12590));
    InMux I__1435 (
            .O(N__12605),
            .I(N__12590));
    LocalMux I__1434 (
            .O(N__12602),
            .I(N__12587));
    InMux I__1433 (
            .O(N__12601),
            .I(N__12578));
    InMux I__1432 (
            .O(N__12600),
            .I(N__12578));
    InMux I__1431 (
            .O(N__12599),
            .I(N__12578));
    InMux I__1430 (
            .O(N__12598),
            .I(N__12578));
    InMux I__1429 (
            .O(N__12595),
            .I(N__12575));
    LocalMux I__1428 (
            .O(N__12590),
            .I(\eeprom.n1256 ));
    Odrv4 I__1427 (
            .O(N__12587),
            .I(\eeprom.n1256 ));
    LocalMux I__1426 (
            .O(N__12578),
            .I(\eeprom.n1256 ));
    LocalMux I__1425 (
            .O(N__12575),
            .I(\eeprom.n1256 ));
    InMux I__1424 (
            .O(N__12566),
            .I(bfn_4_19_0_));
    InMux I__1423 (
            .O(N__12563),
            .I(\eeprom.n3517 ));
    InMux I__1422 (
            .O(N__12560),
            .I(\eeprom.n3518 ));
    InMux I__1421 (
            .O(N__12557),
            .I(\eeprom.n3519 ));
    InMux I__1420 (
            .O(N__12554),
            .I(\eeprom.n3520 ));
    InMux I__1419 (
            .O(N__12551),
            .I(\eeprom.n3521 ));
    InMux I__1418 (
            .O(N__12548),
            .I(\eeprom.n3522 ));
    InMux I__1417 (
            .O(N__12545),
            .I(N__12542));
    LocalMux I__1416 (
            .O(N__12542),
            .I(\eeprom.n2381 ));
    InMux I__1415 (
            .O(N__12539),
            .I(N__12536));
    LocalMux I__1414 (
            .O(N__12536),
            .I(\eeprom.n2384 ));
    CascadeMux I__1413 (
            .O(N__12533),
            .I(N__12530));
    InMux I__1412 (
            .O(N__12530),
            .I(N__12527));
    LocalMux I__1411 (
            .O(N__12527),
            .I(\eeprom.n2378 ));
    InMux I__1410 (
            .O(N__12524),
            .I(N__12521));
    LocalMux I__1409 (
            .O(N__12521),
            .I(\eeprom.n4733 ));
    InMux I__1408 (
            .O(N__12518),
            .I(N__12515));
    LocalMux I__1407 (
            .O(N__12515),
            .I(\eeprom.n1340 ));
    InMux I__1406 (
            .O(N__12512),
            .I(N__12508));
    InMux I__1405 (
            .O(N__12511),
            .I(N__12504));
    LocalMux I__1404 (
            .O(N__12508),
            .I(N__12501));
    InMux I__1403 (
            .O(N__12507),
            .I(N__12498));
    LocalMux I__1402 (
            .O(N__12504),
            .I(\eeprom.n1138 ));
    Odrv4 I__1401 (
            .O(N__12501),
            .I(\eeprom.n1138 ));
    LocalMux I__1400 (
            .O(N__12498),
            .I(\eeprom.n1138 ));
    CascadeMux I__1399 (
            .O(N__12491),
            .I(\eeprom.n1915_cascade_ ));
    CascadeMux I__1398 (
            .O(N__12488),
            .I(N__12484));
    InMux I__1397 (
            .O(N__12487),
            .I(N__12481));
    InMux I__1396 (
            .O(N__12484),
            .I(N__12478));
    LocalMux I__1395 (
            .O(N__12481),
            .I(\eeprom.n1135 ));
    LocalMux I__1394 (
            .O(N__12478),
            .I(\eeprom.n1135 ));
    CascadeMux I__1393 (
            .O(N__12473),
            .I(N__12467));
    CascadeMux I__1392 (
            .O(N__12472),
            .I(N__12463));
    CascadeMux I__1391 (
            .O(N__12471),
            .I(N__12460));
    InMux I__1390 (
            .O(N__12470),
            .I(N__12456));
    InMux I__1389 (
            .O(N__12467),
            .I(N__12453));
    InMux I__1388 (
            .O(N__12466),
            .I(N__12450));
    InMux I__1387 (
            .O(N__12463),
            .I(N__12443));
    InMux I__1386 (
            .O(N__12460),
            .I(N__12443));
    InMux I__1385 (
            .O(N__12459),
            .I(N__12443));
    LocalMux I__1384 (
            .O(N__12456),
            .I(\eeprom.n4405 ));
    LocalMux I__1383 (
            .O(N__12453),
            .I(\eeprom.n4405 ));
    LocalMux I__1382 (
            .O(N__12450),
            .I(\eeprom.n4405 ));
    LocalMux I__1381 (
            .O(N__12443),
            .I(\eeprom.n4405 ));
    InMux I__1380 (
            .O(N__12434),
            .I(N__12431));
    LocalMux I__1379 (
            .O(N__12431),
            .I(\eeprom.n1337 ));
    CascadeMux I__1378 (
            .O(N__12428),
            .I(N__12425));
    InMux I__1377 (
            .O(N__12425),
            .I(N__12422));
    LocalMux I__1376 (
            .O(N__12422),
            .I(N__12419));
    Span4Mux_v I__1375 (
            .O(N__12419),
            .I(N__12416));
    Span4Mux_v I__1374 (
            .O(N__12416),
            .I(N__12413));
    Odrv4 I__1373 (
            .O(N__12413),
            .I(\eeprom.n12_adj_411 ));
    InMux I__1372 (
            .O(N__12410),
            .I(N__12407));
    LocalMux I__1371 (
            .O(N__12407),
            .I(N__12404));
    Span12Mux_h I__1370 (
            .O(N__12404),
            .I(N__12401));
    Odrv12 I__1369 (
            .O(N__12401),
            .I(\eeprom.n25_adj_471 ));
    InMux I__1368 (
            .O(N__12398),
            .I(N__12394));
    InMux I__1367 (
            .O(N__12397),
            .I(N__12390));
    LocalMux I__1366 (
            .O(N__12394),
            .I(N__12387));
    InMux I__1365 (
            .O(N__12393),
            .I(N__12384));
    LocalMux I__1364 (
            .O(N__12390),
            .I(\eeprom.delay_counter_8 ));
    Odrv4 I__1363 (
            .O(N__12387),
            .I(\eeprom.delay_counter_8 ));
    LocalMux I__1362 (
            .O(N__12384),
            .I(\eeprom.delay_counter_8 ));
    InMux I__1361 (
            .O(N__12377),
            .I(\eeprom.n3554 ));
    InMux I__1360 (
            .O(N__12374),
            .I(\eeprom.n3555 ));
    InMux I__1359 (
            .O(N__12371),
            .I(\eeprom.n3556 ));
    InMux I__1358 (
            .O(N__12368),
            .I(\eeprom.n3557 ));
    InMux I__1357 (
            .O(N__12365),
            .I(bfn_3_24_0_));
    InMux I__1356 (
            .O(N__12362),
            .I(\eeprom.n3559 ));
    InMux I__1355 (
            .O(N__12359),
            .I(\eeprom.n3560 ));
    InMux I__1354 (
            .O(N__12356),
            .I(\eeprom.n3561 ));
    InMux I__1353 (
            .O(N__12353),
            .I(N__12350));
    LocalMux I__1352 (
            .O(N__12350),
            .I(N__12347));
    Odrv4 I__1351 (
            .O(N__12347),
            .I(\eeprom.n2386 ));
    InMux I__1350 (
            .O(N__12344),
            .I(N__12341));
    LocalMux I__1349 (
            .O(N__12341),
            .I(\eeprom.n19_adj_428 ));
    InMux I__1348 (
            .O(N__12338),
            .I(N__12335));
    LocalMux I__1347 (
            .O(N__12335),
            .I(N__12331));
    InMux I__1346 (
            .O(N__12334),
            .I(N__12327));
    Span4Mux_v I__1345 (
            .O(N__12331),
            .I(N__12324));
    InMux I__1344 (
            .O(N__12330),
            .I(N__12321));
    LocalMux I__1343 (
            .O(N__12327),
            .I(\eeprom.delay_counter_18 ));
    Odrv4 I__1342 (
            .O(N__12324),
            .I(\eeprom.delay_counter_18 ));
    LocalMux I__1341 (
            .O(N__12321),
            .I(\eeprom.delay_counter_18 ));
    InMux I__1340 (
            .O(N__12314),
            .I(N__12311));
    LocalMux I__1339 (
            .O(N__12311),
            .I(\eeprom.n15_adj_414 ));
    InMux I__1338 (
            .O(N__12308),
            .I(N__12303));
    InMux I__1337 (
            .O(N__12307),
            .I(N__12300));
    InMux I__1336 (
            .O(N__12306),
            .I(N__12297));
    LocalMux I__1335 (
            .O(N__12303),
            .I(N__12292));
    LocalMux I__1334 (
            .O(N__12300),
            .I(N__12292));
    LocalMux I__1333 (
            .O(N__12297),
            .I(\eeprom.delay_counter_23 ));
    Odrv4 I__1332 (
            .O(N__12292),
            .I(\eeprom.delay_counter_23 ));
    InMux I__1331 (
            .O(N__12287),
            .I(N__12284));
    LocalMux I__1330 (
            .O(N__12284),
            .I(\eeprom.n10 ));
    InMux I__1329 (
            .O(N__12281),
            .I(N__12278));
    LocalMux I__1328 (
            .O(N__12278),
            .I(\eeprom.n18_adj_426 ));
    InMux I__1327 (
            .O(N__12275),
            .I(N__12272));
    LocalMux I__1326 (
            .O(N__12272),
            .I(N__12268));
    InMux I__1325 (
            .O(N__12271),
            .I(N__12264));
    Span12Mux_v I__1324 (
            .O(N__12268),
            .I(N__12261));
    InMux I__1323 (
            .O(N__12267),
            .I(N__12258));
    LocalMux I__1322 (
            .O(N__12264),
            .I(\eeprom.delay_counter_15 ));
    Odrv12 I__1321 (
            .O(N__12261),
            .I(\eeprom.delay_counter_15 ));
    LocalMux I__1320 (
            .O(N__12258),
            .I(\eeprom.delay_counter_15 ));
    InMux I__1319 (
            .O(N__12251),
            .I(bfn_3_23_0_));
    InMux I__1318 (
            .O(N__12248),
            .I(\eeprom.n3551 ));
    InMux I__1317 (
            .O(N__12245),
            .I(\eeprom.n3552 ));
    CascadeMux I__1316 (
            .O(N__12242),
            .I(N__12239));
    InMux I__1315 (
            .O(N__12239),
            .I(N__12236));
    LocalMux I__1314 (
            .O(N__12236),
            .I(\eeprom.n2383 ));
    InMux I__1313 (
            .O(N__12233),
            .I(\eeprom.n3553 ));
    CascadeMux I__1312 (
            .O(N__12230),
            .I(N__12225));
    InMux I__1311 (
            .O(N__12229),
            .I(N__12222));
    InMux I__1310 (
            .O(N__12228),
            .I(N__12219));
    InMux I__1309 (
            .O(N__12225),
            .I(N__12216));
    LocalMux I__1308 (
            .O(N__12222),
            .I(\eeprom.delay_counter_26 ));
    LocalMux I__1307 (
            .O(N__12219),
            .I(\eeprom.delay_counter_26 ));
    LocalMux I__1306 (
            .O(N__12216),
            .I(\eeprom.delay_counter_26 ));
    CascadeMux I__1305 (
            .O(N__12209),
            .I(N__12206));
    InMux I__1304 (
            .O(N__12206),
            .I(N__12202));
    InMux I__1303 (
            .O(N__12205),
            .I(N__12199));
    LocalMux I__1302 (
            .O(N__12202),
            .I(N__12194));
    LocalMux I__1301 (
            .O(N__12199),
            .I(N__12194));
    Span4Mux_v I__1300 (
            .O(N__12194),
            .I(N__12191));
    Odrv4 I__1299 (
            .O(N__12191),
            .I(\eeprom.n7 ));
    CascadeMux I__1298 (
            .O(N__12188),
            .I(N__12184));
    InMux I__1297 (
            .O(N__12187),
            .I(N__12181));
    InMux I__1296 (
            .O(N__12184),
            .I(N__12178));
    LocalMux I__1295 (
            .O(N__12181),
            .I(N__12175));
    LocalMux I__1294 (
            .O(N__12178),
            .I(N__12172));
    Odrv4 I__1293 (
            .O(N__12175),
            .I(\eeprom.n1140 ));
    Odrv4 I__1292 (
            .O(N__12172),
            .I(\eeprom.n1140 ));
    InMux I__1291 (
            .O(N__12167),
            .I(N__12162));
    InMux I__1290 (
            .O(N__12166),
            .I(N__12159));
    InMux I__1289 (
            .O(N__12165),
            .I(N__12156));
    LocalMux I__1288 (
            .O(N__12162),
            .I(\eeprom.delay_counter_29 ));
    LocalMux I__1287 (
            .O(N__12159),
            .I(\eeprom.delay_counter_29 ));
    LocalMux I__1286 (
            .O(N__12156),
            .I(\eeprom.delay_counter_29 ));
    InMux I__1285 (
            .O(N__12149),
            .I(N__12146));
    LocalMux I__1284 (
            .O(N__12146),
            .I(N__12143));
    Span4Mux_h I__1283 (
            .O(N__12143),
            .I(N__12140));
    Odrv4 I__1282 (
            .O(N__12140),
            .I(\eeprom.n4 ));
    CascadeMux I__1281 (
            .O(N__12137),
            .I(N__12134));
    InMux I__1280 (
            .O(N__12134),
            .I(N__12131));
    LocalMux I__1279 (
            .O(N__12131),
            .I(N__12127));
    InMux I__1278 (
            .O(N__12130),
            .I(N__12124));
    Odrv4 I__1277 (
            .O(N__12127),
            .I(\eeprom.n1137 ));
    LocalMux I__1276 (
            .O(N__12124),
            .I(\eeprom.n1137 ));
    InMux I__1275 (
            .O(N__12119),
            .I(N__12116));
    LocalMux I__1274 (
            .O(N__12116),
            .I(N__12113));
    Odrv4 I__1273 (
            .O(N__12113),
            .I(\eeprom.n1339 ));
    CascadeMux I__1272 (
            .O(N__12110),
            .I(\eeprom.n1137_cascade_ ));
    InMux I__1271 (
            .O(N__12107),
            .I(N__12104));
    LocalMux I__1270 (
            .O(N__12104),
            .I(N__12101));
    Span4Mux_h I__1269 (
            .O(N__12101),
            .I(N__12098));
    Odrv4 I__1268 (
            .O(N__12098),
            .I(\eeprom.n24_adj_467 ));
    InMux I__1267 (
            .O(N__12095),
            .I(N__12091));
    InMux I__1266 (
            .O(N__12094),
            .I(N__12087));
    LocalMux I__1265 (
            .O(N__12091),
            .I(N__12084));
    InMux I__1264 (
            .O(N__12090),
            .I(N__12081));
    LocalMux I__1263 (
            .O(N__12087),
            .I(\eeprom.delay_counter_9 ));
    Odrv4 I__1262 (
            .O(N__12084),
            .I(\eeprom.delay_counter_9 ));
    LocalMux I__1261 (
            .O(N__12081),
            .I(\eeprom.delay_counter_9 ));
    InMux I__1260 (
            .O(N__12074),
            .I(N__12071));
    LocalMux I__1259 (
            .O(N__12071),
            .I(\eeprom.n33_adj_483 ));
    CascadeMux I__1258 (
            .O(N__12068),
            .I(N__12065));
    InMux I__1257 (
            .O(N__12065),
            .I(N__12062));
    LocalMux I__1256 (
            .O(N__12062),
            .I(N__12059));
    Odrv4 I__1255 (
            .O(N__12059),
            .I(\eeprom.n13_adj_412 ));
    CascadeMux I__1254 (
            .O(N__12056),
            .I(N__12053));
    InMux I__1253 (
            .O(N__12053),
            .I(N__12050));
    LocalMux I__1252 (
            .O(N__12050),
            .I(N__12047));
    Odrv4 I__1251 (
            .O(N__12047),
            .I(\eeprom.n10_adj_409 ));
    InMux I__1250 (
            .O(N__12044),
            .I(N__12040));
    InMux I__1249 (
            .O(N__12043),
            .I(N__12037));
    LocalMux I__1248 (
            .O(N__12040),
            .I(N__12034));
    LocalMux I__1247 (
            .O(N__12037),
            .I(N__12031));
    Span4Mux_v I__1246 (
            .O(N__12034),
            .I(N__12028));
    Span4Mux_v I__1245 (
            .O(N__12031),
            .I(N__12025));
    Odrv4 I__1244 (
            .O(N__12028),
            .I(\eeprom.n2_adj_395 ));
    Odrv4 I__1243 (
            .O(N__12025),
            .I(\eeprom.n2_adj_395 ));
    CascadeMux I__1242 (
            .O(N__12020),
            .I(\eeprom.n4399_cascade_ ));
    InMux I__1241 (
            .O(N__12017),
            .I(N__12014));
    LocalMux I__1240 (
            .O(N__12014),
            .I(N__12011));
    Odrv4 I__1239 (
            .O(N__12011),
            .I(\eeprom.n1343 ));
    CascadeMux I__1238 (
            .O(N__12008),
            .I(N__12005));
    InMux I__1237 (
            .O(N__12005),
            .I(N__12001));
    InMux I__1236 (
            .O(N__12004),
            .I(N__11998));
    LocalMux I__1235 (
            .O(N__12001),
            .I(N__11995));
    LocalMux I__1234 (
            .O(N__11998),
            .I(\eeprom.n1141 ));
    Odrv4 I__1233 (
            .O(N__11995),
            .I(\eeprom.n1141 ));
    CascadeMux I__1232 (
            .O(N__11990),
            .I(\eeprom.n4405_cascade_ ));
    InMux I__1231 (
            .O(N__11987),
            .I(N__11984));
    LocalMux I__1230 (
            .O(N__11984),
            .I(N__11979));
    InMux I__1229 (
            .O(N__11983),
            .I(N__11976));
    InMux I__1228 (
            .O(N__11982),
            .I(N__11973));
    Span4Mux_v I__1227 (
            .O(N__11979),
            .I(N__11970));
    LocalMux I__1226 (
            .O(N__11976),
            .I(N__11967));
    LocalMux I__1225 (
            .O(N__11973),
            .I(\eeprom.delay_counter_28 ));
    Odrv4 I__1224 (
            .O(N__11970),
            .I(\eeprom.delay_counter_28 ));
    Odrv4 I__1223 (
            .O(N__11967),
            .I(\eeprom.delay_counter_28 ));
    InMux I__1222 (
            .O(N__11960),
            .I(N__11957));
    LocalMux I__1221 (
            .O(N__11957),
            .I(N__11954));
    Span4Mux_v I__1220 (
            .O(N__11954),
            .I(N__11951));
    Odrv4 I__1219 (
            .O(N__11951),
            .I(\eeprom.n5 ));
    InMux I__1218 (
            .O(N__11948),
            .I(N__11945));
    LocalMux I__1217 (
            .O(N__11945),
            .I(N__11942));
    Odrv4 I__1216 (
            .O(N__11942),
            .I(\eeprom.n1342 ));
    CascadeMux I__1215 (
            .O(N__11939),
            .I(N__11936));
    InMux I__1214 (
            .O(N__11936),
            .I(N__11930));
    InMux I__1213 (
            .O(N__11935),
            .I(N__11930));
    LocalMux I__1212 (
            .O(N__11930),
            .I(N__11927));
    Span4Mux_v I__1211 (
            .O(N__11927),
            .I(N__11924));
    Odrv4 I__1210 (
            .O(N__11924),
            .I(\eeprom.n6_adj_402 ));
    InMux I__1209 (
            .O(N__11921),
            .I(N__11916));
    InMux I__1208 (
            .O(N__11920),
            .I(N__11913));
    InMux I__1207 (
            .O(N__11919),
            .I(N__11910));
    LocalMux I__1206 (
            .O(N__11916),
            .I(\eeprom.delay_counter_27 ));
    LocalMux I__1205 (
            .O(N__11913),
            .I(\eeprom.delay_counter_27 ));
    LocalMux I__1204 (
            .O(N__11910),
            .I(\eeprom.delay_counter_27 ));
    InMux I__1203 (
            .O(N__11903),
            .I(N__11899));
    InMux I__1202 (
            .O(N__11902),
            .I(N__11896));
    LocalMux I__1201 (
            .O(N__11899),
            .I(N__11893));
    LocalMux I__1200 (
            .O(N__11896),
            .I(\eeprom.n1139 ));
    Odrv4 I__1199 (
            .O(N__11893),
            .I(\eeprom.n1139 ));
    InMux I__1198 (
            .O(N__11888),
            .I(N__11885));
    LocalMux I__1197 (
            .O(N__11885),
            .I(N__11882));
    Odrv4 I__1196 (
            .O(N__11882),
            .I(\eeprom.n25 ));
    CascadeMux I__1195 (
            .O(N__11879),
            .I(N__11876));
    InMux I__1194 (
            .O(N__11876),
            .I(N__11873));
    LocalMux I__1193 (
            .O(N__11873),
            .I(N__11870));
    Span4Mux_h I__1192 (
            .O(N__11870),
            .I(N__11867));
    Odrv4 I__1191 (
            .O(N__11867),
            .I(\eeprom.n9 ));
    CascadeMux I__1190 (
            .O(N__11864),
            .I(N__11859));
    InMux I__1189 (
            .O(N__11863),
            .I(N__11856));
    InMux I__1188 (
            .O(N__11862),
            .I(N__11851));
    InMux I__1187 (
            .O(N__11859),
            .I(N__11851));
    LocalMux I__1186 (
            .O(N__11856),
            .I(\eeprom.delay_counter_24 ));
    LocalMux I__1185 (
            .O(N__11851),
            .I(\eeprom.delay_counter_24 ));
    CascadeMux I__1184 (
            .O(N__11846),
            .I(N__11843));
    InMux I__1183 (
            .O(N__11843),
            .I(N__11840));
    LocalMux I__1182 (
            .O(N__11840),
            .I(N__11837));
    Span4Mux_v I__1181 (
            .O(N__11837),
            .I(N__11834));
    Odrv4 I__1180 (
            .O(N__11834),
            .I(\eeprom.n9_adj_408 ));
    CascadeMux I__1179 (
            .O(N__11831),
            .I(N__11828));
    InMux I__1178 (
            .O(N__11828),
            .I(N__11825));
    LocalMux I__1177 (
            .O(N__11825),
            .I(\eeprom.n32 ));
    InMux I__1176 (
            .O(N__11822),
            .I(N__11819));
    LocalMux I__1175 (
            .O(N__11819),
            .I(N__11816));
    Odrv4 I__1174 (
            .O(N__11816),
            .I(\eeprom.n26 ));
    InMux I__1173 (
            .O(N__11813),
            .I(N__11809));
    InMux I__1172 (
            .O(N__11812),
            .I(N__11805));
    LocalMux I__1171 (
            .O(N__11809),
            .I(N__11802));
    InMux I__1170 (
            .O(N__11808),
            .I(N__11799));
    LocalMux I__1169 (
            .O(N__11805),
            .I(\eeprom.delay_counter_30 ));
    Odrv4 I__1168 (
            .O(N__11802),
            .I(\eeprom.delay_counter_30 ));
    LocalMux I__1167 (
            .O(N__11799),
            .I(\eeprom.delay_counter_30 ));
    InMux I__1166 (
            .O(N__11792),
            .I(N__11789));
    LocalMux I__1165 (
            .O(N__11789),
            .I(N__11786));
    Span4Mux_v I__1164 (
            .O(N__11786),
            .I(N__11783));
    Odrv4 I__1163 (
            .O(N__11783),
            .I(\eeprom.n3 ));
    InMux I__1162 (
            .O(N__11780),
            .I(N__11777));
    LocalMux I__1161 (
            .O(N__11777),
            .I(\eeprom.n1341 ));
    CascadeMux I__1160 (
            .O(N__11774),
            .I(\eeprom.n1256_cascade_ ));
    CascadeMux I__1159 (
            .O(N__11771),
            .I(N__11768));
    InMux I__1158 (
            .O(N__11768),
            .I(N__11765));
    LocalMux I__1157 (
            .O(N__11765),
            .I(N__11762));
    Span4Mux_v I__1156 (
            .O(N__11762),
            .I(N__11759));
    Odrv4 I__1155 (
            .O(N__11759),
            .I(\eeprom.n5_adj_400 ));
    CascadeMux I__1154 (
            .O(N__11756),
            .I(N__11753));
    InMux I__1153 (
            .O(N__11753),
            .I(N__11750));
    LocalMux I__1152 (
            .O(N__11750),
            .I(N__11747));
    Span4Mux_v I__1151 (
            .O(N__11747),
            .I(N__11744));
    Odrv4 I__1150 (
            .O(N__11744),
            .I(\eeprom.n15_adj_415 ));
    InMux I__1149 (
            .O(N__11741),
            .I(N__11738));
    LocalMux I__1148 (
            .O(N__11738),
            .I(N__11735));
    Odrv4 I__1147 (
            .O(N__11735),
            .I(\eeprom.n33 ));
    CascadeMux I__1146 (
            .O(N__11732),
            .I(N__11728));
    InMux I__1145 (
            .O(N__11731),
            .I(N__11724));
    InMux I__1144 (
            .O(N__11728),
            .I(N__11721));
    InMux I__1143 (
            .O(N__11727),
            .I(N__11718));
    LocalMux I__1142 (
            .O(N__11724),
            .I(\eeprom.delay_counter_25 ));
    LocalMux I__1141 (
            .O(N__11721),
            .I(\eeprom.delay_counter_25 ));
    LocalMux I__1140 (
            .O(N__11718),
            .I(\eeprom.delay_counter_25 ));
    InMux I__1139 (
            .O(N__11711),
            .I(N__11708));
    LocalMux I__1138 (
            .O(N__11708),
            .I(N__11705));
    Span4Mux_v I__1137 (
            .O(N__11705),
            .I(N__11702));
    Odrv4 I__1136 (
            .O(N__11702),
            .I(\eeprom.n8 ));
    CascadeMux I__1135 (
            .O(N__11699),
            .I(\eeprom.n1141_cascade_ ));
    CascadeMux I__1134 (
            .O(N__11696),
            .I(N__11693));
    InMux I__1133 (
            .O(N__11693),
            .I(N__11690));
    LocalMux I__1132 (
            .O(N__11690),
            .I(N__11687));
    Odrv4 I__1131 (
            .O(N__11687),
            .I(\eeprom.n11_adj_410 ));
    InMux I__1130 (
            .O(N__11684),
            .I(bfn_3_17_0_));
    InMux I__1129 (
            .O(N__11681),
            .I(\eeprom.n3448 ));
    InMux I__1128 (
            .O(N__11678),
            .I(\eeprom.n3449 ));
    InMux I__1127 (
            .O(N__11675),
            .I(\eeprom.n3450 ));
    InMux I__1126 (
            .O(N__11672),
            .I(\eeprom.n3451 ));
    InMux I__1125 (
            .O(N__11669),
            .I(\eeprom.n3452 ));
    InMux I__1124 (
            .O(N__11666),
            .I(\eeprom.n3453 ));
    CascadeMux I__1123 (
            .O(N__11663),
            .I(N__11660));
    InMux I__1122 (
            .O(N__11660),
            .I(N__11657));
    LocalMux I__1121 (
            .O(N__11657),
            .I(N__11654));
    Span4Mux_v I__1120 (
            .O(N__11654),
            .I(N__11651));
    Odrv4 I__1119 (
            .O(N__11651),
            .I(\eeprom.n30_adj_458 ));
    InMux I__1118 (
            .O(N__11648),
            .I(bfn_2_24_0_));
    CascadeMux I__1117 (
            .O(N__11645),
            .I(N__11642));
    InMux I__1116 (
            .O(N__11642),
            .I(N__11639));
    LocalMux I__1115 (
            .O(N__11639),
            .I(N__11636));
    Span4Mux_v I__1114 (
            .O(N__11636),
            .I(N__11633));
    Odrv4 I__1113 (
            .O(N__11633),
            .I(\eeprom.n8_adj_407 ));
    InMux I__1112 (
            .O(N__11630),
            .I(\eeprom.n3810 ));
    CascadeMux I__1111 (
            .O(N__11627),
            .I(N__11624));
    InMux I__1110 (
            .O(N__11624),
            .I(N__11621));
    LocalMux I__1109 (
            .O(N__11621),
            .I(N__11618));
    Span4Mux_v I__1108 (
            .O(N__11618),
            .I(N__11615));
    Odrv4 I__1107 (
            .O(N__11615),
            .I(\eeprom.n7_adj_405 ));
    InMux I__1106 (
            .O(N__11612),
            .I(\eeprom.n3811 ));
    CascadeMux I__1105 (
            .O(N__11609),
            .I(N__11606));
    InMux I__1104 (
            .O(N__11606),
            .I(N__11603));
    LocalMux I__1103 (
            .O(N__11603),
            .I(N__11600));
    Span4Mux_v I__1102 (
            .O(N__11600),
            .I(N__11597));
    Odrv4 I__1101 (
            .O(N__11597),
            .I(\eeprom.n6_adj_403 ));
    InMux I__1100 (
            .O(N__11594),
            .I(\eeprom.n3812 ));
    InMux I__1099 (
            .O(N__11591),
            .I(\eeprom.n3813 ));
    CascadeMux I__1098 (
            .O(N__11588),
            .I(N__11585));
    InMux I__1097 (
            .O(N__11585),
            .I(N__11582));
    LocalMux I__1096 (
            .O(N__11582),
            .I(N__11579));
    Span4Mux_v I__1095 (
            .O(N__11579),
            .I(N__11576));
    Odrv4 I__1094 (
            .O(N__11576),
            .I(\eeprom.n4_adj_397 ));
    InMux I__1093 (
            .O(N__11573),
            .I(\eeprom.n3814 ));
    CascadeMux I__1092 (
            .O(N__11570),
            .I(N__11567));
    InMux I__1091 (
            .O(N__11567),
            .I(N__11564));
    LocalMux I__1090 (
            .O(N__11564),
            .I(N__11561));
    Span4Mux_v I__1089 (
            .O(N__11561),
            .I(N__11558));
    Odrv4 I__1088 (
            .O(N__11558),
            .I(\eeprom.n3_adj_396 ));
    InMux I__1087 (
            .O(N__11555),
            .I(\eeprom.n3815 ));
    InMux I__1086 (
            .O(N__11552),
            .I(\eeprom.n3816 ));
    InMux I__1085 (
            .O(N__11549),
            .I(N__11546));
    LocalMux I__1084 (
            .O(N__11546),
            .I(N__11543));
    Odrv12 I__1083 (
            .O(N__11543),
            .I(\eeprom.n14 ));
    InMux I__1082 (
            .O(N__11540),
            .I(N__11537));
    LocalMux I__1081 (
            .O(N__11537),
            .I(N__11532));
    InMux I__1080 (
            .O(N__11536),
            .I(N__11529));
    InMux I__1079 (
            .O(N__11535),
            .I(N__11526));
    Span4Mux_v I__1078 (
            .O(N__11532),
            .I(N__11521));
    LocalMux I__1077 (
            .O(N__11529),
            .I(N__11521));
    LocalMux I__1076 (
            .O(N__11526),
            .I(\eeprom.delay_counter_19 ));
    Odrv4 I__1075 (
            .O(N__11521),
            .I(\eeprom.delay_counter_19 ));
    InMux I__1074 (
            .O(N__11516),
            .I(\eeprom.n3800 ));
    InMux I__1073 (
            .O(N__11513),
            .I(N__11510));
    LocalMux I__1072 (
            .O(N__11510),
            .I(\eeprom.n17_adj_425 ));
    InMux I__1071 (
            .O(N__11507),
            .I(N__11504));
    LocalMux I__1070 (
            .O(N__11504),
            .I(\eeprom.n17 ));
    InMux I__1069 (
            .O(N__11501),
            .I(bfn_2_23_0_));
    CascadeMux I__1068 (
            .O(N__11498),
            .I(N__11495));
    InMux I__1067 (
            .O(N__11495),
            .I(N__11492));
    LocalMux I__1066 (
            .O(N__11492),
            .I(\eeprom.n16_adj_424 ));
    InMux I__1065 (
            .O(N__11489),
            .I(\eeprom.n3802 ));
    InMux I__1064 (
            .O(N__11486),
            .I(\eeprom.n3803 ));
    CascadeMux I__1063 (
            .O(N__11483),
            .I(N__11480));
    InMux I__1062 (
            .O(N__11480),
            .I(N__11477));
    LocalMux I__1061 (
            .O(N__11477),
            .I(\eeprom.n14_adj_413 ));
    InMux I__1060 (
            .O(N__11474),
            .I(\eeprom.n3804 ));
    InMux I__1059 (
            .O(N__11471),
            .I(\eeprom.n3805 ));
    InMux I__1058 (
            .O(N__11468),
            .I(\eeprom.n3806 ));
    InMux I__1057 (
            .O(N__11465),
            .I(\eeprom.n3807 ));
    InMux I__1056 (
            .O(N__11462),
            .I(\eeprom.n3808 ));
    InMux I__1055 (
            .O(N__11459),
            .I(\eeprom.n3792 ));
    InMux I__1054 (
            .O(N__11456),
            .I(bfn_2_22_0_));
    CascadeMux I__1053 (
            .O(N__11453),
            .I(N__11450));
    InMux I__1052 (
            .O(N__11450),
            .I(N__11447));
    LocalMux I__1051 (
            .O(N__11447),
            .I(N__11444));
    Span4Mux_v I__1050 (
            .O(N__11444),
            .I(N__11441));
    Odrv4 I__1049 (
            .O(N__11441),
            .I(\eeprom.n24_adj_463 ));
    InMux I__1048 (
            .O(N__11438),
            .I(\eeprom.n3794 ));
    CascadeMux I__1047 (
            .O(N__11435),
            .I(N__11432));
    InMux I__1046 (
            .O(N__11432),
            .I(N__11429));
    LocalMux I__1045 (
            .O(N__11429),
            .I(N__11426));
    Span4Mux_v I__1044 (
            .O(N__11426),
            .I(N__11423));
    Odrv4 I__1043 (
            .O(N__11423),
            .I(\eeprom.n23 ));
    InMux I__1042 (
            .O(N__11420),
            .I(\eeprom.n3795 ));
    CascadeMux I__1041 (
            .O(N__11417),
            .I(N__11414));
    InMux I__1040 (
            .O(N__11414),
            .I(N__11411));
    LocalMux I__1039 (
            .O(N__11411),
            .I(N__11408));
    Span4Mux_v I__1038 (
            .O(N__11408),
            .I(N__11405));
    Odrv4 I__1037 (
            .O(N__11405),
            .I(\eeprom.n22_adj_448 ));
    InMux I__1036 (
            .O(N__11402),
            .I(N__11399));
    LocalMux I__1035 (
            .O(N__11399),
            .I(N__11396));
    Sp12to4 I__1034 (
            .O(N__11396),
            .I(N__11393));
    Odrv12 I__1033 (
            .O(N__11393),
            .I(\eeprom.n22_adj_447 ));
    InMux I__1032 (
            .O(N__11390),
            .I(\eeprom.n3796 ));
    CascadeMux I__1031 (
            .O(N__11387),
            .I(N__11384));
    InMux I__1030 (
            .O(N__11384),
            .I(N__11381));
    LocalMux I__1029 (
            .O(N__11381),
            .I(N__11378));
    Span4Mux_v I__1028 (
            .O(N__11378),
            .I(N__11375));
    Odrv4 I__1027 (
            .O(N__11375),
            .I(\eeprom.n21_adj_440 ));
    InMux I__1026 (
            .O(N__11372),
            .I(\eeprom.n3797 ));
    CascadeMux I__1025 (
            .O(N__11369),
            .I(N__11366));
    InMux I__1024 (
            .O(N__11366),
            .I(N__11363));
    LocalMux I__1023 (
            .O(N__11363),
            .I(\eeprom.n20_adj_431 ));
    InMux I__1022 (
            .O(N__11360),
            .I(N__11357));
    LocalMux I__1021 (
            .O(N__11357),
            .I(N__11354));
    Span4Mux_s1_h I__1020 (
            .O(N__11354),
            .I(N__11351));
    Odrv4 I__1019 (
            .O(N__11351),
            .I(\eeprom.n20_adj_430 ));
    InMux I__1018 (
            .O(N__11348),
            .I(\eeprom.n3798 ));
    InMux I__1017 (
            .O(N__11345),
            .I(\eeprom.n3799 ));
    CascadeMux I__1016 (
            .O(N__11342),
            .I(N__11339));
    InMux I__1015 (
            .O(N__11339),
            .I(N__11336));
    LocalMux I__1014 (
            .O(N__11336),
            .I(N__11333));
    Span4Mux_v I__1013 (
            .O(N__11333),
            .I(N__11330));
    Odrv4 I__1012 (
            .O(N__11330),
            .I(\eeprom.n18_adj_427 ));
    InMux I__1011 (
            .O(N__11327),
            .I(\eeprom.n3483 ));
    InMux I__1010 (
            .O(N__11324),
            .I(\eeprom.n3484 ));
    InMux I__1009 (
            .O(N__11321),
            .I(bfn_2_21_0_));
    InMux I__1008 (
            .O(N__11318),
            .I(\eeprom.n3786 ));
    CascadeMux I__1007 (
            .O(N__11315),
            .I(N__11312));
    InMux I__1006 (
            .O(N__11312),
            .I(N__11309));
    LocalMux I__1005 (
            .O(N__11309),
            .I(N__11306));
    Odrv4 I__1004 (
            .O(N__11306),
            .I(\eeprom.n31_adj_457 ));
    InMux I__1003 (
            .O(N__11303),
            .I(\eeprom.n3787 ));
    InMux I__1002 (
            .O(N__11300),
            .I(\eeprom.n3788 ));
    InMux I__1001 (
            .O(N__11297),
            .I(\eeprom.n3789 ));
    CascadeMux I__1000 (
            .O(N__11294),
            .I(N__11291));
    InMux I__999 (
            .O(N__11291),
            .I(N__11288));
    LocalMux I__998 (
            .O(N__11288),
            .I(N__11285));
    Odrv4 I__997 (
            .O(N__11285),
            .I(\eeprom.n28_adj_461 ));
    InMux I__996 (
            .O(N__11282),
            .I(\eeprom.n3790 ));
    CascadeMux I__995 (
            .O(N__11279),
            .I(N__11276));
    InMux I__994 (
            .O(N__11276),
            .I(N__11273));
    LocalMux I__993 (
            .O(N__11273),
            .I(N__11270));
    Span4Mux_v I__992 (
            .O(N__11270),
            .I(N__11267));
    Odrv4 I__991 (
            .O(N__11267),
            .I(\eeprom.n27_adj_462 ));
    InMux I__990 (
            .O(N__11264),
            .I(\eeprom.n3791 ));
    InMux I__989 (
            .O(N__11261),
            .I(\eeprom.n3474 ));
    InMux I__988 (
            .O(N__11258),
            .I(\eeprom.n3475 ));
    InMux I__987 (
            .O(N__11255),
            .I(\eeprom.n3476 ));
    InMux I__986 (
            .O(N__11252),
            .I(bfn_2_20_0_));
    InMux I__985 (
            .O(N__11249),
            .I(\eeprom.n3478 ));
    InMux I__984 (
            .O(N__11246),
            .I(\eeprom.n3479 ));
    InMux I__983 (
            .O(N__11243),
            .I(\eeprom.n3480 ));
    InMux I__982 (
            .O(N__11240),
            .I(\eeprom.n3481 ));
    InMux I__981 (
            .O(N__11237),
            .I(\eeprom.n3482 ));
    InMux I__980 (
            .O(N__11234),
            .I(\eeprom.n3465 ));
    InMux I__979 (
            .O(N__11231),
            .I(N__11227));
    InMux I__978 (
            .O(N__11230),
            .I(N__11223));
    LocalMux I__977 (
            .O(N__11227),
            .I(N__11220));
    InMux I__976 (
            .O(N__11226),
            .I(N__11217));
    LocalMux I__975 (
            .O(N__11223),
            .I(N__11212));
    Span4Mux_v I__974 (
            .O(N__11220),
            .I(N__11212));
    LocalMux I__973 (
            .O(N__11217),
            .I(\eeprom.delay_counter_13 ));
    Odrv4 I__972 (
            .O(N__11212),
            .I(\eeprom.delay_counter_13 ));
    InMux I__971 (
            .O(N__11207),
            .I(\eeprom.n3466 ));
    InMux I__970 (
            .O(N__11204),
            .I(\eeprom.n3467 ));
    InMux I__969 (
            .O(N__11201),
            .I(\eeprom.n3468 ));
    InMux I__968 (
            .O(N__11198),
            .I(N__11192));
    InMux I__967 (
            .O(N__11197),
            .I(N__11192));
    LocalMux I__966 (
            .O(N__11192),
            .I(N__11188));
    InMux I__965 (
            .O(N__11191),
            .I(N__11185));
    Span4Mux_v I__964 (
            .O(N__11188),
            .I(N__11182));
    LocalMux I__963 (
            .O(N__11185),
            .I(\eeprom.delay_counter_16 ));
    Odrv4 I__962 (
            .O(N__11182),
            .I(\eeprom.delay_counter_16 ));
    InMux I__961 (
            .O(N__11177),
            .I(bfn_2_19_0_));
    InMux I__960 (
            .O(N__11174),
            .I(\eeprom.n3470 ));
    InMux I__959 (
            .O(N__11171),
            .I(\eeprom.n3471 ));
    InMux I__958 (
            .O(N__11168),
            .I(\eeprom.n3472 ));
    InMux I__957 (
            .O(N__11165),
            .I(\eeprom.n3473 ));
    InMux I__956 (
            .O(N__11162),
            .I(\eeprom.n3456 ));
    InMux I__955 (
            .O(N__11159),
            .I(\eeprom.n3457 ));
    InMux I__954 (
            .O(N__11156),
            .I(\eeprom.n3458 ));
    InMux I__953 (
            .O(N__11153),
            .I(\eeprom.n3459 ));
    InMux I__952 (
            .O(N__11150),
            .I(\eeprom.n3460 ));
    InMux I__951 (
            .O(N__11147),
            .I(bfn_2_18_0_));
    InMux I__950 (
            .O(N__11144),
            .I(\eeprom.n3462 ));
    InMux I__949 (
            .O(N__11141),
            .I(\eeprom.n3463 ));
    InMux I__948 (
            .O(N__11138),
            .I(N__11133));
    InMux I__947 (
            .O(N__11137),
            .I(N__11128));
    InMux I__946 (
            .O(N__11136),
            .I(N__11128));
    LocalMux I__945 (
            .O(N__11133),
            .I(\eeprom.delay_counter_11 ));
    LocalMux I__944 (
            .O(N__11128),
            .I(\eeprom.delay_counter_11 ));
    InMux I__943 (
            .O(N__11123),
            .I(\eeprom.n3464 ));
    InMux I__942 (
            .O(N__11120),
            .I(bfn_2_17_0_));
    InMux I__941 (
            .O(N__11117),
            .I(\eeprom.n3454 ));
    InMux I__940 (
            .O(N__11114),
            .I(\eeprom.n3455 ));
    IoInMux I__939 (
            .O(N__11111),
            .I(N__11108));
    LocalMux I__938 (
            .O(N__11108),
            .I(N__11105));
    IoSpan4Mux I__937 (
            .O(N__11105),
            .I(N__11102));
    IoSpan4Mux I__936 (
            .O(N__11102),
            .I(N__11099));
    IoSpan4Mux I__935 (
            .O(N__11099),
            .I(N__11096));
    Odrv4 I__934 (
            .O(N__11096),
            .I(CLK_pad_gb_input));
    defparam IN_MUX_bfv_2_21_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_21_0_ (
            .carryinitin(),
            .carryinitout(bfn_2_21_0_));
    defparam IN_MUX_bfv_2_22_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_22_0_ (
            .carryinitin(\eeprom.n3793 ),
            .carryinitout(bfn_2_22_0_));
    defparam IN_MUX_bfv_2_23_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_23_0_ (
            .carryinitin(\eeprom.n3801 ),
            .carryinitout(bfn_2_23_0_));
    defparam IN_MUX_bfv_2_24_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_24_0_ (
            .carryinitin(\eeprom.n3809 ),
            .carryinitout(bfn_2_24_0_));
    defparam IN_MUX_bfv_15_20_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_20_0_ (
            .carryinitin(),
            .carryinitout(bfn_15_20_0_));
    defparam IN_MUX_bfv_15_21_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_21_0_ (
            .carryinitin(\eeprom.n3779 ),
            .carryinitout(bfn_15_21_0_));
    defparam IN_MUX_bfv_16_17_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_17_0_ (
            .carryinitin(),
            .carryinitout(bfn_16_17_0_));
    defparam IN_MUX_bfv_16_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_18_0_ (
            .carryinitin(\eeprom.n3756 ),
            .carryinitout(bfn_16_18_0_));
    defparam IN_MUX_bfv_16_19_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_19_0_ (
            .carryinitin(\eeprom.n3764 ),
            .carryinitout(bfn_16_19_0_));
    defparam IN_MUX_bfv_14_17_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_17_0_ (
            .carryinitin(),
            .carryinitout(bfn_14_17_0_));
    defparam IN_MUX_bfv_14_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_18_0_ (
            .carryinitin(\eeprom.n3734 ),
            .carryinitout(bfn_14_18_0_));
    defparam IN_MUX_bfv_14_19_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_19_0_ (
            .carryinitin(\eeprom.n3742 ),
            .carryinitout(bfn_14_19_0_));
    defparam IN_MUX_bfv_9_17_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_17_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_17_0_));
    defparam IN_MUX_bfv_9_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_18_0_ (
            .carryinitin(\eeprom.n3713 ),
            .carryinitout(bfn_9_18_0_));
    defparam IN_MUX_bfv_9_19_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_19_0_ (
            .carryinitin(\eeprom.n3721 ),
            .carryinitout(bfn_9_19_0_));
    defparam IN_MUX_bfv_9_20_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_20_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_20_0_));
    defparam IN_MUX_bfv_9_21_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_21_0_ (
            .carryinitin(\eeprom.n3693 ),
            .carryinitout(bfn_9_21_0_));
    defparam IN_MUX_bfv_9_22_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_22_0_ (
            .carryinitin(\eeprom.n3701 ),
            .carryinitout(bfn_9_22_0_));
    defparam IN_MUX_bfv_12_22_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_22_0_ (
            .carryinitin(),
            .carryinitout(bfn_12_22_0_));
    defparam IN_MUX_bfv_12_23_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_23_0_ (
            .carryinitin(\eeprom.n3674 ),
            .carryinitout(bfn_12_23_0_));
    defparam IN_MUX_bfv_12_24_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_24_0_ (
            .carryinitin(\eeprom.n3682 ),
            .carryinitout(bfn_12_24_0_));
    defparam IN_MUX_bfv_16_23_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_23_0_ (
            .carryinitin(),
            .carryinitout(bfn_16_23_0_));
    defparam IN_MUX_bfv_16_24_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_24_0_ (
            .carryinitin(\eeprom.n3656 ),
            .carryinitout(bfn_16_24_0_));
    defparam IN_MUX_bfv_16_25_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_25_0_ (
            .carryinitin(\eeprom.n3664 ),
            .carryinitout(bfn_16_25_0_));
    defparam IN_MUX_bfv_11_21_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_21_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_21_0_));
    defparam IN_MUX_bfv_11_22_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_22_0_ (
            .carryinitin(\eeprom.n3639 ),
            .carryinitout(bfn_11_22_0_));
    defparam IN_MUX_bfv_11_23_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_23_0_ (
            .carryinitin(\eeprom.n3647 ),
            .carryinitout(bfn_11_23_0_));
    defparam IN_MUX_bfv_9_23_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_23_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_23_0_));
    defparam IN_MUX_bfv_9_24_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_24_0_ (
            .carryinitin(\eeprom.n3623 ),
            .carryinitout(bfn_9_24_0_));
    defparam IN_MUX_bfv_9_25_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_25_0_ (
            .carryinitin(\eeprom.n3631 ),
            .carryinitout(bfn_9_25_0_));
    defparam IN_MUX_bfv_7_21_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_21_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_21_0_));
    defparam IN_MUX_bfv_7_22_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_22_0_ (
            .carryinitin(\eeprom.n3608 ),
            .carryinitout(bfn_7_22_0_));
    defparam IN_MUX_bfv_6_18_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_18_0_ (
            .carryinitin(),
            .carryinitout(bfn_6_18_0_));
    defparam IN_MUX_bfv_6_19_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_19_0_ (
            .carryinitin(\eeprom.n3594 ),
            .carryinitout(bfn_6_19_0_));
    defparam IN_MUX_bfv_6_21_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_21_0_ (
            .carryinitin(),
            .carryinitout(bfn_6_21_0_));
    defparam IN_MUX_bfv_6_22_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_22_0_ (
            .carryinitin(\eeprom.n3581 ),
            .carryinitout(bfn_6_22_0_));
    defparam IN_MUX_bfv_4_25_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_25_0_ (
            .carryinitin(),
            .carryinitout(bfn_4_25_0_));
    defparam IN_MUX_bfv_4_26_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_26_0_ (
            .carryinitin(\eeprom.n3569 ),
            .carryinitout(bfn_4_26_0_));
    defparam IN_MUX_bfv_3_23_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_23_0_ (
            .carryinitin(),
            .carryinitout(bfn_3_23_0_));
    defparam IN_MUX_bfv_3_24_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_24_0_ (
            .carryinitin(\eeprom.n3558 ),
            .carryinitout(bfn_3_24_0_));
    defparam IN_MUX_bfv_6_26_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_26_0_ (
            .carryinitin(),
            .carryinitout(bfn_6_26_0_));
    defparam IN_MUX_bfv_6_27_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_27_0_ (
            .carryinitin(\eeprom.n3548 ),
            .carryinitout(bfn_6_27_0_));
    defparam IN_MUX_bfv_5_27_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_27_0_ (
            .carryinitin(),
            .carryinitout(bfn_5_27_0_));
    defparam IN_MUX_bfv_5_28_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_28_0_ (
            .carryinitin(\eeprom.n3539 ),
            .carryinitout(bfn_5_28_0_));
    defparam IN_MUX_bfv_5_22_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_22_0_ (
            .carryinitin(),
            .carryinitout(bfn_5_22_0_));
    defparam IN_MUX_bfv_5_23_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_23_0_ (
            .carryinitin(\eeprom.n3531 ),
            .carryinitout(bfn_5_23_0_));
    defparam IN_MUX_bfv_4_19_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_19_0_ (
            .carryinitin(),
            .carryinitout(bfn_4_19_0_));
    defparam IN_MUX_bfv_2_17_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_17_0_ (
            .carryinitin(),
            .carryinitout(bfn_2_17_0_));
    defparam IN_MUX_bfv_2_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_18_0_ (
            .carryinitin(\eeprom.n3461 ),
            .carryinitout(bfn_2_18_0_));
    defparam IN_MUX_bfv_2_19_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_19_0_ (
            .carryinitin(\eeprom.n3469 ),
            .carryinitout(bfn_2_19_0_));
    defparam IN_MUX_bfv_2_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_20_0_ (
            .carryinitin(\eeprom.n3477 ),
            .carryinitout(bfn_2_20_0_));
    defparam IN_MUX_bfv_16_20_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_20_0_ (
            .carryinitin(),
            .carryinitout(bfn_16_20_0_));
    defparam IN_MUX_bfv_3_17_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_17_0_ (
            .carryinitin(),
            .carryinitout(bfn_3_17_0_));
    defparam IN_MUX_bfv_5_29_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_29_0_ (
            .carryinitin(),
            .carryinitout(bfn_5_29_0_));
    defparam IN_MUX_bfv_5_30_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_30_0_ (
            .carryinitin(n3492),
            .carryinitout(bfn_5_30_0_));
    defparam IN_MUX_bfv_5_31_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_31_0_ (
            .carryinitin(n3500),
            .carryinitout(bfn_5_31_0_));
    defparam IN_MUX_bfv_5_32_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_32_0_ (
            .carryinitin(n3508),
            .carryinitout(bfn_5_32_0_));
    ICE_GB CLK_pad_gb (
            .USERSIGNALTOGLOBALBUFFER(N__11111),
            .GLOBALBUFFEROUTPUT(CLK_N));
    VCC VCC (
            .Y(VCCG0));
    GND GND (
            .Y(GNDG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i10_1_lut_LC_1_17_1 .C_ON=1'b0;
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i10_1_lut_LC_1_17_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i10_1_lut_LC_1_17_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \eeprom.rem_4_unary_minus_2_inv_0_i10_1_lut_LC_1_17_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12090),
            .lcout(\eeprom.n24_adj_463 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i7_1_lut_LC_1_17_3 .C_ON=1'b0;
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i7_1_lut_LC_1_17_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i7_1_lut_LC_1_17_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \eeprom.rem_4_unary_minus_2_inv_0_i7_1_lut_LC_1_17_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23595),
            .lcout(\eeprom.n27_adj_462 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i11_1_lut_LC_1_17_5 .C_ON=1'b0;
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i11_1_lut_LC_1_17_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i11_1_lut_LC_1_17_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \eeprom.rem_4_unary_minus_2_inv_0_i11_1_lut_LC_1_17_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13470),
            .lcout(\eeprom.n23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_mux_3_i12_3_lut_LC_1_17_6 .C_ON=1'b0;
    defparam \eeprom.rem_4_mux_3_i12_3_lut_LC_1_17_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_mux_3_i12_3_lut_LC_1_17_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \eeprom.rem_4_mux_3_i12_3_lut_LC_1_17_6  (
            .in0(N__11137),
            .in1(N__11402),
            .in2(_gnd_net_),
            .in3(N__22970),
            .lcout(\eeprom.n3219 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i12_1_lut_LC_1_17_7 .C_ON=1'b0;
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i12_1_lut_LC_1_17_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i12_1_lut_LC_1_17_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \eeprom.rem_4_unary_minus_2_inv_0_i12_1_lut_LC_1_17_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11136),
            .lcout(\eeprom.n22_adj_448 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i16_1_lut_LC_1_18_2 .C_ON=1'b0;
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i16_1_lut_LC_1_18_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i16_1_lut_LC_1_18_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \eeprom.rem_4_unary_minus_2_inv_0_i16_1_lut_LC_1_18_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12267),
            .lcout(\eeprom.n18_adj_427 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i13_1_lut_LC_1_19_0 .C_ON=1'b0;
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i13_1_lut_LC_1_19_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i13_1_lut_LC_1_19_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \eeprom.rem_4_unary_minus_2_inv_0_i13_1_lut_LC_1_19_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14910),
            .lcout(\eeprom.n21_adj_440 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i26_1_lut_LC_1_19_1 .C_ON=1'b0;
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i26_1_lut_LC_1_19_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i26_1_lut_LC_1_19_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \eeprom.rem_4_unary_minus_2_inv_0_i26_1_lut_LC_1_19_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11727),
            .lcout(\eeprom.n8_adj_407 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i27_1_lut_LC_1_19_2 .C_ON=1'b0;
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i27_1_lut_LC_1_19_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i27_1_lut_LC_1_19_2 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \eeprom.rem_4_unary_minus_2_inv_0_i27_1_lut_LC_1_19_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__12230),
            .in3(_gnd_net_),
            .lcout(\eeprom.n7_adj_405 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i28_1_lut_LC_1_19_3 .C_ON=1'b0;
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i28_1_lut_LC_1_19_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i28_1_lut_LC_1_19_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \eeprom.rem_4_unary_minus_2_inv_0_i28_1_lut_LC_1_19_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11919),
            .lcout(\eeprom.n6_adj_403 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i30_1_lut_LC_1_19_4 .C_ON=1'b0;
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i30_1_lut_LC_1_19_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i30_1_lut_LC_1_19_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \eeprom.rem_4_unary_minus_2_inv_0_i30_1_lut_LC_1_19_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12165),
            .lcout(\eeprom.n4_adj_397 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i31_1_lut_LC_1_19_5 .C_ON=1'b0;
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i31_1_lut_LC_1_19_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i31_1_lut_LC_1_19_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \eeprom.rem_4_unary_minus_2_inv_0_i31_1_lut_LC_1_19_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11808),
            .lcout(\eeprom.n3_adj_396 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i3_1_lut_LC_1_19_6 .C_ON=1'b0;
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i3_1_lut_LC_1_19_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i3_1_lut_LC_1_19_6 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \eeprom.rem_4_unary_minus_2_inv_0_i3_1_lut_LC_1_19_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__23838),
            .in3(_gnd_net_),
            .lcout(\eeprom.n31_adj_457 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i6_1_lut_LC_1_19_7 .C_ON=1'b0;
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i6_1_lut_LC_1_19_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i6_1_lut_LC_1_19_7 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \eeprom.rem_4_unary_minus_2_inv_0_i6_1_lut_LC_1_19_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__23658),
            .in3(_gnd_net_),
            .lcout(\eeprom.n28_adj_461 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_mux_3_i14_3_lut_LC_1_20_2 .C_ON=1'b0;
    defparam \eeprom.rem_4_mux_3_i14_3_lut_LC_1_20_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_mux_3_i14_3_lut_LC_1_20_2 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \eeprom.rem_4_mux_3_i14_3_lut_LC_1_20_2  (
            .in0(N__11360),
            .in1(N__22888),
            .in2(_gnd_net_),
            .in3(N__11230),
            .lcout(\eeprom.n3019 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i14_1_lut_LC_1_22_1 .C_ON=1'b0;
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i14_1_lut_LC_1_22_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i14_1_lut_LC_1_22_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \eeprom.rem_4_unary_minus_2_inv_0_i14_1_lut_LC_1_22_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11231),
            .lcout(\eeprom.n20_adj_431 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_mux_3_i17_3_lut_LC_1_22_2 .C_ON=1'b0;
    defparam \eeprom.rem_4_mux_3_i17_3_lut_LC_1_22_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_mux_3_i17_3_lut_LC_1_22_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \eeprom.rem_4_mux_3_i17_3_lut_LC_1_22_2  (
            .in0(N__11198),
            .in1(N__11507),
            .in2(_gnd_net_),
            .in3(N__22938),
            .lcout(\eeprom.n2719 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i17_1_lut_LC_1_22_3 .C_ON=1'b0;
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i17_1_lut_LC_1_22_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i17_1_lut_LC_1_22_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \eeprom.rem_4_unary_minus_2_inv_0_i17_1_lut_LC_1_22_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11197),
            .lcout(\eeprom.n17_adj_425 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i18_1_lut_LC_1_22_5 .C_ON=1'b0;
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i18_1_lut_LC_1_22_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i18_1_lut_LC_1_22_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \eeprom.rem_4_unary_minus_2_inv_0_i18_1_lut_LC_1_22_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12661),
            .lcout(\eeprom.n16_adj_424 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i20_1_lut_LC_1_22_7 .C_ON=1'b0;
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i20_1_lut_LC_1_22_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i20_1_lut_LC_1_22_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \eeprom.rem_4_unary_minus_2_inv_0_i20_1_lut_LC_1_22_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11536),
            .lcout(\eeprom.n14_adj_413 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.delay_counter_288__i0_LC_2_17_0 .C_ON=1'b1;
    defparam \eeprom.delay_counter_288__i0_LC_2_17_0 .SEQ_MODE=4'b1000;
    defparam \eeprom.delay_counter_288__i0_LC_2_17_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.delay_counter_288__i0_LC_2_17_0  (
            .in0(_gnd_net_),
            .in1(N__23481),
            .in2(_gnd_net_),
            .in3(N__11120),
            .lcout(\eeprom.delay_counter_0 ),
            .ltout(),
            .carryin(bfn_2_17_0_),
            .carryout(\eeprom.n3454 ),
            .clk(N__24342),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.delay_counter_288__i1_LC_2_17_1 .C_ON=1'b1;
    defparam \eeprom.delay_counter_288__i1_LC_2_17_1 .SEQ_MODE=4'b1000;
    defparam \eeprom.delay_counter_288__i1_LC_2_17_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.delay_counter_288__i1_LC_2_17_1  (
            .in0(_gnd_net_),
            .in1(N__23891),
            .in2(_gnd_net_),
            .in3(N__11117),
            .lcout(\eeprom.delay_counter_1 ),
            .ltout(),
            .carryin(\eeprom.n3454 ),
            .carryout(\eeprom.n3455 ),
            .clk(N__24342),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.delay_counter_288__i2_LC_2_17_2 .C_ON=1'b1;
    defparam \eeprom.delay_counter_288__i2_LC_2_17_2 .SEQ_MODE=4'b1000;
    defparam \eeprom.delay_counter_288__i2_LC_2_17_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.delay_counter_288__i2_LC_2_17_2  (
            .in0(_gnd_net_),
            .in1(N__23828),
            .in2(_gnd_net_),
            .in3(N__11114),
            .lcout(\eeprom.delay_counter_2 ),
            .ltout(),
            .carryin(\eeprom.n3455 ),
            .carryout(\eeprom.n3456 ),
            .clk(N__24342),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.delay_counter_288__i3_LC_2_17_3 .C_ON=1'b1;
    defparam \eeprom.delay_counter_288__i3_LC_2_17_3 .SEQ_MODE=4'b1000;
    defparam \eeprom.delay_counter_288__i3_LC_2_17_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.delay_counter_288__i3_LC_2_17_3  (
            .in0(_gnd_net_),
            .in1(N__23772),
            .in2(_gnd_net_),
            .in3(N__11162),
            .lcout(\eeprom.delay_counter_3 ),
            .ltout(),
            .carryin(\eeprom.n3456 ),
            .carryout(\eeprom.n3457 ),
            .clk(N__24342),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.delay_counter_288__i4_LC_2_17_4 .C_ON=1'b1;
    defparam \eeprom.delay_counter_288__i4_LC_2_17_4 .SEQ_MODE=4'b1000;
    defparam \eeprom.delay_counter_288__i4_LC_2_17_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.delay_counter_288__i4_LC_2_17_4  (
            .in0(_gnd_net_),
            .in1(N__23703),
            .in2(_gnd_net_),
            .in3(N__11159),
            .lcout(\eeprom.delay_counter_4 ),
            .ltout(),
            .carryin(\eeprom.n3457 ),
            .carryout(\eeprom.n3458 ),
            .clk(N__24342),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.delay_counter_288__i5_LC_2_17_5 .C_ON=1'b1;
    defparam \eeprom.delay_counter_288__i5_LC_2_17_5 .SEQ_MODE=4'b1000;
    defparam \eeprom.delay_counter_288__i5_LC_2_17_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.delay_counter_288__i5_LC_2_17_5  (
            .in0(_gnd_net_),
            .in1(N__23649),
            .in2(_gnd_net_),
            .in3(N__11156),
            .lcout(\eeprom.delay_counter_5 ),
            .ltout(),
            .carryin(\eeprom.n3458 ),
            .carryout(\eeprom.n3459 ),
            .clk(N__24342),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.delay_counter_288__i6_LC_2_17_6 .C_ON=1'b1;
    defparam \eeprom.delay_counter_288__i6_LC_2_17_6 .SEQ_MODE=4'b1000;
    defparam \eeprom.delay_counter_288__i6_LC_2_17_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.delay_counter_288__i6_LC_2_17_6  (
            .in0(_gnd_net_),
            .in1(N__23599),
            .in2(_gnd_net_),
            .in3(N__11153),
            .lcout(\eeprom.delay_counter_6 ),
            .ltout(),
            .carryin(\eeprom.n3459 ),
            .carryout(\eeprom.n3460 ),
            .clk(N__24342),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.delay_counter_288__i7_LC_2_17_7 .C_ON=1'b1;
    defparam \eeprom.delay_counter_288__i7_LC_2_17_7 .SEQ_MODE=4'b1000;
    defparam \eeprom.delay_counter_288__i7_LC_2_17_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.delay_counter_288__i7_LC_2_17_7  (
            .in0(_gnd_net_),
            .in1(N__12832),
            .in2(_gnd_net_),
            .in3(N__11150),
            .lcout(\eeprom.delay_counter_7 ),
            .ltout(),
            .carryin(\eeprom.n3460 ),
            .carryout(\eeprom.n3461 ),
            .clk(N__24342),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.delay_counter_288__i8_LC_2_18_0 .C_ON=1'b1;
    defparam \eeprom.delay_counter_288__i8_LC_2_18_0 .SEQ_MODE=4'b1000;
    defparam \eeprom.delay_counter_288__i8_LC_2_18_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.delay_counter_288__i8_LC_2_18_0  (
            .in0(_gnd_net_),
            .in1(N__12397),
            .in2(_gnd_net_),
            .in3(N__11147),
            .lcout(\eeprom.delay_counter_8 ),
            .ltout(),
            .carryin(bfn_2_18_0_),
            .carryout(\eeprom.n3462 ),
            .clk(N__24343),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.delay_counter_288__i9_LC_2_18_1 .C_ON=1'b1;
    defparam \eeprom.delay_counter_288__i9_LC_2_18_1 .SEQ_MODE=4'b1000;
    defparam \eeprom.delay_counter_288__i9_LC_2_18_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.delay_counter_288__i9_LC_2_18_1  (
            .in0(_gnd_net_),
            .in1(N__12094),
            .in2(_gnd_net_),
            .in3(N__11144),
            .lcout(\eeprom.delay_counter_9 ),
            .ltout(),
            .carryin(\eeprom.n3462 ),
            .carryout(\eeprom.n3463 ),
            .clk(N__24343),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.delay_counter_288__i10_LC_2_18_2 .C_ON=1'b1;
    defparam \eeprom.delay_counter_288__i10_LC_2_18_2 .SEQ_MODE=4'b1000;
    defparam \eeprom.delay_counter_288__i10_LC_2_18_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.delay_counter_288__i10_LC_2_18_2  (
            .in0(_gnd_net_),
            .in1(N__13474),
            .in2(_gnd_net_),
            .in3(N__11141),
            .lcout(\eeprom.delay_counter_10 ),
            .ltout(),
            .carryin(\eeprom.n3463 ),
            .carryout(\eeprom.n3464 ),
            .clk(N__24343),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.delay_counter_288__i11_LC_2_18_3 .C_ON=1'b1;
    defparam \eeprom.delay_counter_288__i11_LC_2_18_3 .SEQ_MODE=4'b1000;
    defparam \eeprom.delay_counter_288__i11_LC_2_18_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.delay_counter_288__i11_LC_2_18_3  (
            .in0(_gnd_net_),
            .in1(N__11138),
            .in2(_gnd_net_),
            .in3(N__11123),
            .lcout(\eeprom.delay_counter_11 ),
            .ltout(),
            .carryin(\eeprom.n3464 ),
            .carryout(\eeprom.n3465 ),
            .clk(N__24343),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.delay_counter_288__i12_LC_2_18_4 .C_ON=1'b1;
    defparam \eeprom.delay_counter_288__i12_LC_2_18_4 .SEQ_MODE=4'b1000;
    defparam \eeprom.delay_counter_288__i12_LC_2_18_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.delay_counter_288__i12_LC_2_18_4  (
            .in0(_gnd_net_),
            .in1(N__14914),
            .in2(_gnd_net_),
            .in3(N__11234),
            .lcout(\eeprom.delay_counter_12 ),
            .ltout(),
            .carryin(\eeprom.n3465 ),
            .carryout(\eeprom.n3466 ),
            .clk(N__24343),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.delay_counter_288__i13_LC_2_18_5 .C_ON=1'b1;
    defparam \eeprom.delay_counter_288__i13_LC_2_18_5 .SEQ_MODE=4'b1000;
    defparam \eeprom.delay_counter_288__i13_LC_2_18_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.delay_counter_288__i13_LC_2_18_5  (
            .in0(_gnd_net_),
            .in1(N__11226),
            .in2(_gnd_net_),
            .in3(N__11207),
            .lcout(\eeprom.delay_counter_13 ),
            .ltout(),
            .carryin(\eeprom.n3466 ),
            .carryout(\eeprom.n3467 ),
            .clk(N__24343),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.delay_counter_288__i14_LC_2_18_6 .C_ON=1'b1;
    defparam \eeprom.delay_counter_288__i14_LC_2_18_6 .SEQ_MODE=4'b1000;
    defparam \eeprom.delay_counter_288__i14_LC_2_18_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.delay_counter_288__i14_LC_2_18_6  (
            .in0(_gnd_net_),
            .in1(N__13584),
            .in2(_gnd_net_),
            .in3(N__11204),
            .lcout(\eeprom.delay_counter_14 ),
            .ltout(),
            .carryin(\eeprom.n3467 ),
            .carryout(\eeprom.n3468 ),
            .clk(N__24343),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.delay_counter_288__i15_LC_2_18_7 .C_ON=1'b1;
    defparam \eeprom.delay_counter_288__i15_LC_2_18_7 .SEQ_MODE=4'b1000;
    defparam \eeprom.delay_counter_288__i15_LC_2_18_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.delay_counter_288__i15_LC_2_18_7  (
            .in0(_gnd_net_),
            .in1(N__12271),
            .in2(_gnd_net_),
            .in3(N__11201),
            .lcout(\eeprom.delay_counter_15 ),
            .ltout(),
            .carryin(\eeprom.n3468 ),
            .carryout(\eeprom.n3469 ),
            .clk(N__24343),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.delay_counter_288__i16_LC_2_19_0 .C_ON=1'b1;
    defparam \eeprom.delay_counter_288__i16_LC_2_19_0 .SEQ_MODE=4'b1000;
    defparam \eeprom.delay_counter_288__i16_LC_2_19_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.delay_counter_288__i16_LC_2_19_0  (
            .in0(_gnd_net_),
            .in1(N__11191),
            .in2(_gnd_net_),
            .in3(N__11177),
            .lcout(\eeprom.delay_counter_16 ),
            .ltout(),
            .carryin(bfn_2_19_0_),
            .carryout(\eeprom.n3470 ),
            .clk(N__24344),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.delay_counter_288__i17_LC_2_19_1 .C_ON=1'b1;
    defparam \eeprom.delay_counter_288__i17_LC_2_19_1 .SEQ_MODE=4'b1000;
    defparam \eeprom.delay_counter_288__i17_LC_2_19_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.delay_counter_288__i17_LC_2_19_1  (
            .in0(_gnd_net_),
            .in1(N__12660),
            .in2(_gnd_net_),
            .in3(N__11174),
            .lcout(\eeprom.delay_counter_17 ),
            .ltout(),
            .carryin(\eeprom.n3470 ),
            .carryout(\eeprom.n3471 ),
            .clk(N__24344),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.delay_counter_288__i18_LC_2_19_2 .C_ON=1'b1;
    defparam \eeprom.delay_counter_288__i18_LC_2_19_2 .SEQ_MODE=4'b1000;
    defparam \eeprom.delay_counter_288__i18_LC_2_19_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.delay_counter_288__i18_LC_2_19_2  (
            .in0(_gnd_net_),
            .in1(N__12334),
            .in2(_gnd_net_),
            .in3(N__11171),
            .lcout(\eeprom.delay_counter_18 ),
            .ltout(),
            .carryin(\eeprom.n3471 ),
            .carryout(\eeprom.n3472 ),
            .clk(N__24344),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.delay_counter_288__i19_LC_2_19_3 .C_ON=1'b1;
    defparam \eeprom.delay_counter_288__i19_LC_2_19_3 .SEQ_MODE=4'b1000;
    defparam \eeprom.delay_counter_288__i19_LC_2_19_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.delay_counter_288__i19_LC_2_19_3  (
            .in0(_gnd_net_),
            .in1(N__11535),
            .in2(_gnd_net_),
            .in3(N__11168),
            .lcout(\eeprom.delay_counter_19 ),
            .ltout(),
            .carryin(\eeprom.n3472 ),
            .carryout(\eeprom.n3473 ),
            .clk(N__24344),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.delay_counter_288__i20_LC_2_19_4 .C_ON=1'b1;
    defparam \eeprom.delay_counter_288__i20_LC_2_19_4 .SEQ_MODE=4'b1000;
    defparam \eeprom.delay_counter_288__i20_LC_2_19_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.delay_counter_288__i20_LC_2_19_4  (
            .in0(_gnd_net_),
            .in1(N__13050),
            .in2(_gnd_net_),
            .in3(N__11165),
            .lcout(\eeprom.delay_counter_20 ),
            .ltout(),
            .carryin(\eeprom.n3473 ),
            .carryout(\eeprom.n3474 ),
            .clk(N__24344),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.delay_counter_288__i21_LC_2_19_5 .C_ON=1'b1;
    defparam \eeprom.delay_counter_288__i21_LC_2_19_5 .SEQ_MODE=4'b1000;
    defparam \eeprom.delay_counter_288__i21_LC_2_19_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.delay_counter_288__i21_LC_2_19_5  (
            .in0(_gnd_net_),
            .in1(N__15609),
            .in2(_gnd_net_),
            .in3(N__11261),
            .lcout(\eeprom.delay_counter_21 ),
            .ltout(),
            .carryin(\eeprom.n3474 ),
            .carryout(\eeprom.n3475 ),
            .clk(N__24344),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.delay_counter_288__i22_LC_2_19_6 .C_ON=1'b1;
    defparam \eeprom.delay_counter_288__i22_LC_2_19_6 .SEQ_MODE=4'b1000;
    defparam \eeprom.delay_counter_288__i22_LC_2_19_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.delay_counter_288__i22_LC_2_19_6  (
            .in0(_gnd_net_),
            .in1(N__14178),
            .in2(_gnd_net_),
            .in3(N__11258),
            .lcout(\eeprom.delay_counter_22 ),
            .ltout(),
            .carryin(\eeprom.n3475 ),
            .carryout(\eeprom.n3476 ),
            .clk(N__24344),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.delay_counter_288__i23_LC_2_19_7 .C_ON=1'b1;
    defparam \eeprom.delay_counter_288__i23_LC_2_19_7 .SEQ_MODE=4'b1000;
    defparam \eeprom.delay_counter_288__i23_LC_2_19_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.delay_counter_288__i23_LC_2_19_7  (
            .in0(_gnd_net_),
            .in1(N__12306),
            .in2(_gnd_net_),
            .in3(N__11255),
            .lcout(\eeprom.delay_counter_23 ),
            .ltout(),
            .carryin(\eeprom.n3476 ),
            .carryout(\eeprom.n3477 ),
            .clk(N__24344),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.delay_counter_288__i24_LC_2_20_0 .C_ON=1'b1;
    defparam \eeprom.delay_counter_288__i24_LC_2_20_0 .SEQ_MODE=4'b1000;
    defparam \eeprom.delay_counter_288__i24_LC_2_20_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.delay_counter_288__i24_LC_2_20_0  (
            .in0(_gnd_net_),
            .in1(N__11863),
            .in2(_gnd_net_),
            .in3(N__11252),
            .lcout(\eeprom.delay_counter_24 ),
            .ltout(),
            .carryin(bfn_2_20_0_),
            .carryout(\eeprom.n3478 ),
            .clk(N__24345),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.delay_counter_288__i25_LC_2_20_1 .C_ON=1'b1;
    defparam \eeprom.delay_counter_288__i25_LC_2_20_1 .SEQ_MODE=4'b1000;
    defparam \eeprom.delay_counter_288__i25_LC_2_20_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.delay_counter_288__i25_LC_2_20_1  (
            .in0(_gnd_net_),
            .in1(N__11731),
            .in2(_gnd_net_),
            .in3(N__11249),
            .lcout(\eeprom.delay_counter_25 ),
            .ltout(),
            .carryin(\eeprom.n3478 ),
            .carryout(\eeprom.n3479 ),
            .clk(N__24345),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.delay_counter_288__i26_LC_2_20_2 .C_ON=1'b1;
    defparam \eeprom.delay_counter_288__i26_LC_2_20_2 .SEQ_MODE=4'b1000;
    defparam \eeprom.delay_counter_288__i26_LC_2_20_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.delay_counter_288__i26_LC_2_20_2  (
            .in0(_gnd_net_),
            .in1(N__12229),
            .in2(_gnd_net_),
            .in3(N__11246),
            .lcout(\eeprom.delay_counter_26 ),
            .ltout(),
            .carryin(\eeprom.n3479 ),
            .carryout(\eeprom.n3480 ),
            .clk(N__24345),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.delay_counter_288__i27_LC_2_20_3 .C_ON=1'b1;
    defparam \eeprom.delay_counter_288__i27_LC_2_20_3 .SEQ_MODE=4'b1000;
    defparam \eeprom.delay_counter_288__i27_LC_2_20_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.delay_counter_288__i27_LC_2_20_3  (
            .in0(_gnd_net_),
            .in1(N__11921),
            .in2(_gnd_net_),
            .in3(N__11243),
            .lcout(\eeprom.delay_counter_27 ),
            .ltout(),
            .carryin(\eeprom.n3480 ),
            .carryout(\eeprom.n3481 ),
            .clk(N__24345),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.delay_counter_288__i28_LC_2_20_4 .C_ON=1'b1;
    defparam \eeprom.delay_counter_288__i28_LC_2_20_4 .SEQ_MODE=4'b1000;
    defparam \eeprom.delay_counter_288__i28_LC_2_20_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.delay_counter_288__i28_LC_2_20_4  (
            .in0(_gnd_net_),
            .in1(N__11982),
            .in2(_gnd_net_),
            .in3(N__11240),
            .lcout(\eeprom.delay_counter_28 ),
            .ltout(),
            .carryin(\eeprom.n3481 ),
            .carryout(\eeprom.n3482 ),
            .clk(N__24345),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.delay_counter_288__i29_LC_2_20_5 .C_ON=1'b1;
    defparam \eeprom.delay_counter_288__i29_LC_2_20_5 .SEQ_MODE=4'b1000;
    defparam \eeprom.delay_counter_288__i29_LC_2_20_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.delay_counter_288__i29_LC_2_20_5  (
            .in0(_gnd_net_),
            .in1(N__12167),
            .in2(_gnd_net_),
            .in3(N__11237),
            .lcout(\eeprom.delay_counter_29 ),
            .ltout(),
            .carryin(\eeprom.n3482 ),
            .carryout(\eeprom.n3483 ),
            .clk(N__24345),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.delay_counter_288__i30_LC_2_20_6 .C_ON=1'b1;
    defparam \eeprom.delay_counter_288__i30_LC_2_20_6 .SEQ_MODE=4'b1000;
    defparam \eeprom.delay_counter_288__i30_LC_2_20_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.delay_counter_288__i30_LC_2_20_6  (
            .in0(_gnd_net_),
            .in1(N__11812),
            .in2(_gnd_net_),
            .in3(N__11327),
            .lcout(\eeprom.delay_counter_30 ),
            .ltout(),
            .carryin(\eeprom.n3483 ),
            .carryout(\eeprom.n3484 ),
            .clk(N__24345),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.delay_counter_288__i31_LC_2_20_7 .C_ON=1'b0;
    defparam \eeprom.delay_counter_288__i31_LC_2_20_7 .SEQ_MODE=4'b1000;
    defparam \eeprom.delay_counter_288__i31_LC_2_20_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.delay_counter_288__i31_LC_2_20_7  (
            .in0(_gnd_net_),
            .in1(N__22906),
            .in2(_gnd_net_),
            .in3(N__11324),
            .lcout(\eeprom.delay_counter_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24345),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_unary_minus_2_add_3_2_lut_LC_2_21_0 .C_ON=1'b1;
    defparam \eeprom.rem_4_unary_minus_2_add_3_2_lut_LC_2_21_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_unary_minus_2_add_3_2_lut_LC_2_21_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_unary_minus_2_add_3_2_lut_LC_2_21_0  (
            .in0(_gnd_net_),
            .in1(N__11741),
            .in2(_gnd_net_),
            .in3(N__11321),
            .lcout(\eeprom.n33_adj_483 ),
            .ltout(),
            .carryin(bfn_2_21_0_),
            .carryout(\eeprom.n3786 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_unary_minus_2_add_3_3_lut_LC_2_21_1 .C_ON=1'b1;
    defparam \eeprom.rem_4_unary_minus_2_add_3_3_lut_LC_2_21_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_unary_minus_2_add_3_3_lut_LC_2_21_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_unary_minus_2_add_3_3_lut_LC_2_21_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__11831),
            .in3(N__11318),
            .lcout(\eeprom.n32_adj_480 ),
            .ltout(),
            .carryin(\eeprom.n3786 ),
            .carryout(\eeprom.n3787 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_unary_minus_2_add_3_4_lut_LC_2_21_2 .C_ON=1'b1;
    defparam \eeprom.rem_4_unary_minus_2_add_3_4_lut_LC_2_21_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_unary_minus_2_add_3_4_lut_LC_2_21_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_unary_minus_2_add_3_4_lut_LC_2_21_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__11315),
            .in3(N__11303),
            .lcout(\eeprom.n31_adj_476 ),
            .ltout(),
            .carryin(\eeprom.n3787 ),
            .carryout(\eeprom.n3788 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_unary_minus_2_add_3_5_lut_LC_2_21_3 .C_ON=1'b1;
    defparam \eeprom.rem_4_unary_minus_2_add_3_5_lut_LC_2_21_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_unary_minus_2_add_3_5_lut_LC_2_21_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_unary_minus_2_add_3_5_lut_LC_2_21_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__11663),
            .in3(N__11300),
            .lcout(\eeprom.n30 ),
            .ltout(),
            .carryin(\eeprom.n3788 ),
            .carryout(\eeprom.n3789 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_unary_minus_2_add_3_6_lut_LC_2_21_4 .C_ON=1'b1;
    defparam \eeprom.rem_4_unary_minus_2_add_3_6_lut_LC_2_21_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_unary_minus_2_add_3_6_lut_LC_2_21_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_unary_minus_2_add_3_6_lut_LC_2_21_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__14894),
            .in3(N__11297),
            .lcout(\eeprom.n29 ),
            .ltout(),
            .carryin(\eeprom.n3789 ),
            .carryout(\eeprom.n3790 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_unary_minus_2_add_3_7_lut_LC_2_21_5 .C_ON=1'b1;
    defparam \eeprom.rem_4_unary_minus_2_add_3_7_lut_LC_2_21_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_unary_minus_2_add_3_7_lut_LC_2_21_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_unary_minus_2_add_3_7_lut_LC_2_21_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__11294),
            .in3(N__11282),
            .lcout(\eeprom.n28 ),
            .ltout(),
            .carryin(\eeprom.n3790 ),
            .carryout(\eeprom.n3791 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_unary_minus_2_add_3_8_lut_LC_2_21_6 .C_ON=1'b1;
    defparam \eeprom.rem_4_unary_minus_2_add_3_8_lut_LC_2_21_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_unary_minus_2_add_3_8_lut_LC_2_21_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_unary_minus_2_add_3_8_lut_LC_2_21_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__11279),
            .in3(N__11264),
            .lcout(\eeprom.n27 ),
            .ltout(),
            .carryin(\eeprom.n3791 ),
            .carryout(\eeprom.n3792 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_unary_minus_2_add_3_9_lut_LC_2_21_7 .C_ON=1'b1;
    defparam \eeprom.rem_4_unary_minus_2_add_3_9_lut_LC_2_21_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_unary_minus_2_add_3_9_lut_LC_2_21_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_unary_minus_2_add_3_9_lut_LC_2_21_7  (
            .in0(_gnd_net_),
            .in1(N__11822),
            .in2(_gnd_net_),
            .in3(N__11459),
            .lcout(\eeprom.n26_adj_469 ),
            .ltout(),
            .carryin(\eeprom.n3792 ),
            .carryout(\eeprom.n3793 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_unary_minus_2_add_3_10_lut_LC_2_22_0 .C_ON=1'b1;
    defparam \eeprom.rem_4_unary_minus_2_add_3_10_lut_LC_2_22_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_unary_minus_2_add_3_10_lut_LC_2_22_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_unary_minus_2_add_3_10_lut_LC_2_22_0  (
            .in0(_gnd_net_),
            .in1(N__11888),
            .in2(_gnd_net_),
            .in3(N__11456),
            .lcout(\eeprom.n25_adj_471 ),
            .ltout(),
            .carryin(bfn_2_22_0_),
            .carryout(\eeprom.n3794 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_unary_minus_2_add_3_11_lut_LC_2_22_1 .C_ON=1'b1;
    defparam \eeprom.rem_4_unary_minus_2_add_3_11_lut_LC_2_22_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_unary_minus_2_add_3_11_lut_LC_2_22_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_unary_minus_2_add_3_11_lut_LC_2_22_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__11453),
            .in3(N__11438),
            .lcout(\eeprom.n24_adj_467 ),
            .ltout(),
            .carryin(\eeprom.n3794 ),
            .carryout(\eeprom.n3795 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_unary_minus_2_add_3_12_lut_LC_2_22_2 .C_ON=1'b1;
    defparam \eeprom.rem_4_unary_minus_2_add_3_12_lut_LC_2_22_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_unary_minus_2_add_3_12_lut_LC_2_22_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_unary_minus_2_add_3_12_lut_LC_2_22_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__11435),
            .in3(N__11420),
            .lcout(\eeprom.n23_adj_464 ),
            .ltout(),
            .carryin(\eeprom.n3795 ),
            .carryout(\eeprom.n3796 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_unary_minus_2_add_3_13_lut_LC_2_22_3 .C_ON=1'b1;
    defparam \eeprom.rem_4_unary_minus_2_add_3_13_lut_LC_2_22_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_unary_minus_2_add_3_13_lut_LC_2_22_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_unary_minus_2_add_3_13_lut_LC_2_22_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__11417),
            .in3(N__11390),
            .lcout(\eeprom.n22_adj_447 ),
            .ltout(),
            .carryin(\eeprom.n3796 ),
            .carryout(\eeprom.n3797 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_unary_minus_2_add_3_14_lut_LC_2_22_4 .C_ON=1'b1;
    defparam \eeprom.rem_4_unary_minus_2_add_3_14_lut_LC_2_22_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_unary_minus_2_add_3_14_lut_LC_2_22_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_unary_minus_2_add_3_14_lut_LC_2_22_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__11387),
            .in3(N__11372),
            .lcout(\eeprom.n21 ),
            .ltout(),
            .carryin(\eeprom.n3797 ),
            .carryout(\eeprom.n3798 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_unary_minus_2_add_3_15_lut_LC_2_22_5 .C_ON=1'b1;
    defparam \eeprom.rem_4_unary_minus_2_add_3_15_lut_LC_2_22_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_unary_minus_2_add_3_15_lut_LC_2_22_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_unary_minus_2_add_3_15_lut_LC_2_22_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__11369),
            .in3(N__11348),
            .lcout(\eeprom.n20_adj_430 ),
            .ltout(),
            .carryin(\eeprom.n3798 ),
            .carryout(\eeprom.n3799 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_unary_minus_2_add_3_16_lut_LC_2_22_6 .C_ON=1'b1;
    defparam \eeprom.rem_4_unary_minus_2_add_3_16_lut_LC_2_22_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_unary_minus_2_add_3_16_lut_LC_2_22_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_unary_minus_2_add_3_16_lut_LC_2_22_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__13562),
            .in3(N__11345),
            .lcout(\eeprom.n19_adj_428 ),
            .ltout(),
            .carryin(\eeprom.n3799 ),
            .carryout(\eeprom.n3800 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_unary_minus_2_add_3_17_lut_LC_2_22_7 .C_ON=1'b1;
    defparam \eeprom.rem_4_unary_minus_2_add_3_17_lut_LC_2_22_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_unary_minus_2_add_3_17_lut_LC_2_22_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_unary_minus_2_add_3_17_lut_LC_2_22_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__11342),
            .in3(N__11516),
            .lcout(\eeprom.n18_adj_426 ),
            .ltout(),
            .carryin(\eeprom.n3800 ),
            .carryout(\eeprom.n3801 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_unary_minus_2_add_3_18_lut_LC_2_23_0 .C_ON=1'b1;
    defparam \eeprom.rem_4_unary_minus_2_add_3_18_lut_LC_2_23_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_unary_minus_2_add_3_18_lut_LC_2_23_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_unary_minus_2_add_3_18_lut_LC_2_23_0  (
            .in0(_gnd_net_),
            .in1(N__11513),
            .in2(_gnd_net_),
            .in3(N__11501),
            .lcout(\eeprom.n17 ),
            .ltout(),
            .carryin(bfn_2_23_0_),
            .carryout(\eeprom.n3802 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_unary_minus_2_add_3_19_lut_LC_2_23_1 .C_ON=1'b1;
    defparam \eeprom.rem_4_unary_minus_2_add_3_19_lut_LC_2_23_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_unary_minus_2_add_3_19_lut_LC_2_23_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_unary_minus_2_add_3_19_lut_LC_2_23_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__11498),
            .in3(N__11489),
            .lcout(\eeprom.n16_adj_377 ),
            .ltout(),
            .carryin(\eeprom.n3802 ),
            .carryout(\eeprom.n3803 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_unary_minus_2_add_3_20_lut_LC_2_23_2 .C_ON=1'b1;
    defparam \eeprom.rem_4_unary_minus_2_add_3_20_lut_LC_2_23_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_unary_minus_2_add_3_20_lut_LC_2_23_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_unary_minus_2_add_3_20_lut_LC_2_23_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__11756),
            .in3(N__11486),
            .lcout(\eeprom.n15_adj_414 ),
            .ltout(),
            .carryin(\eeprom.n3803 ),
            .carryout(\eeprom.n3804 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_unary_minus_2_add_3_21_lut_LC_2_23_3 .C_ON=1'b1;
    defparam \eeprom.rem_4_unary_minus_2_add_3_21_lut_LC_2_23_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_unary_minus_2_add_3_21_lut_LC_2_23_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_unary_minus_2_add_3_21_lut_LC_2_23_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__11483),
            .in3(N__11474),
            .lcout(\eeprom.n14 ),
            .ltout(),
            .carryin(\eeprom.n3804 ),
            .carryout(\eeprom.n3805 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_unary_minus_2_add_3_22_lut_LC_2_23_4 .C_ON=1'b1;
    defparam \eeprom.rem_4_unary_minus_2_add_3_22_lut_LC_2_23_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_unary_minus_2_add_3_22_lut_LC_2_23_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_unary_minus_2_add_3_22_lut_LC_2_23_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__12068),
            .in3(N__11471),
            .lcout(\eeprom.n13 ),
            .ltout(),
            .carryin(\eeprom.n3805 ),
            .carryout(\eeprom.n3806 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_unary_minus_2_add_3_23_lut_LC_2_23_5 .C_ON=1'b1;
    defparam \eeprom.rem_4_unary_minus_2_add_3_23_lut_LC_2_23_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_unary_minus_2_add_3_23_lut_LC_2_23_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_unary_minus_2_add_3_23_lut_LC_2_23_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__12428),
            .in3(N__11468),
            .lcout(\eeprom.n12_adj_351 ),
            .ltout(),
            .carryin(\eeprom.n3806 ),
            .carryout(\eeprom.n3807 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_unary_minus_2_add_3_24_lut_LC_2_23_6 .C_ON=1'b1;
    defparam \eeprom.rem_4_unary_minus_2_add_3_24_lut_LC_2_23_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_unary_minus_2_add_3_24_lut_LC_2_23_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_unary_minus_2_add_3_24_lut_LC_2_23_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__11696),
            .in3(N__11465),
            .lcout(\eeprom.n11 ),
            .ltout(),
            .carryin(\eeprom.n3807 ),
            .carryout(\eeprom.n3808 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_unary_minus_2_add_3_25_lut_LC_2_23_7 .C_ON=1'b1;
    defparam \eeprom.rem_4_unary_minus_2_add_3_25_lut_LC_2_23_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_unary_minus_2_add_3_25_lut_LC_2_23_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_unary_minus_2_add_3_25_lut_LC_2_23_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__12056),
            .in3(N__11462),
            .lcout(\eeprom.n10 ),
            .ltout(),
            .carryin(\eeprom.n3808 ),
            .carryout(\eeprom.n3809 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_unary_minus_2_add_3_26_lut_LC_2_24_0 .C_ON=1'b1;
    defparam \eeprom.rem_4_unary_minus_2_add_3_26_lut_LC_2_24_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_unary_minus_2_add_3_26_lut_LC_2_24_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_unary_minus_2_add_3_26_lut_LC_2_24_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__11846),
            .in3(N__11648),
            .lcout(\eeprom.n9 ),
            .ltout(),
            .carryin(bfn_2_24_0_),
            .carryout(\eeprom.n3810 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_unary_minus_2_add_3_27_lut_LC_2_24_1 .C_ON=1'b1;
    defparam \eeprom.rem_4_unary_minus_2_add_3_27_lut_LC_2_24_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_unary_minus_2_add_3_27_lut_LC_2_24_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_unary_minus_2_add_3_27_lut_LC_2_24_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__11645),
            .in3(N__11630),
            .lcout(\eeprom.n8 ),
            .ltout(),
            .carryin(\eeprom.n3810 ),
            .carryout(\eeprom.n3811 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_unary_minus_2_add_3_28_lut_LC_2_24_2 .C_ON=1'b1;
    defparam \eeprom.rem_4_unary_minus_2_add_3_28_lut_LC_2_24_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_unary_minus_2_add_3_28_lut_LC_2_24_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_unary_minus_2_add_3_28_lut_LC_2_24_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__11627),
            .in3(N__11612),
            .lcout(\eeprom.n7 ),
            .ltout(),
            .carryin(\eeprom.n3811 ),
            .carryout(\eeprom.n3812 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_unary_minus_2_add_3_29_lut_LC_2_24_3 .C_ON=1'b1;
    defparam \eeprom.rem_4_unary_minus_2_add_3_29_lut_LC_2_24_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_unary_minus_2_add_3_29_lut_LC_2_24_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_unary_minus_2_add_3_29_lut_LC_2_24_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__11609),
            .in3(N__11594),
            .lcout(\eeprom.n6_adj_402 ),
            .ltout(),
            .carryin(\eeprom.n3812 ),
            .carryout(\eeprom.n3813 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_unary_minus_2_add_3_30_lut_LC_2_24_4 .C_ON=1'b1;
    defparam \eeprom.rem_4_unary_minus_2_add_3_30_lut_LC_2_24_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_unary_minus_2_add_3_30_lut_LC_2_24_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_unary_minus_2_add_3_30_lut_LC_2_24_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__11771),
            .in3(N__11591),
            .lcout(\eeprom.n5 ),
            .ltout(),
            .carryin(\eeprom.n3813 ),
            .carryout(\eeprom.n3814 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_unary_minus_2_add_3_31_lut_LC_2_24_5 .C_ON=1'b1;
    defparam \eeprom.rem_4_unary_minus_2_add_3_31_lut_LC_2_24_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_unary_minus_2_add_3_31_lut_LC_2_24_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_unary_minus_2_add_3_31_lut_LC_2_24_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__11588),
            .in3(N__11573),
            .lcout(\eeprom.n4 ),
            .ltout(),
            .carryin(\eeprom.n3814 ),
            .carryout(\eeprom.n3815 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_unary_minus_2_add_3_32_lut_LC_2_24_6 .C_ON=1'b1;
    defparam \eeprom.rem_4_unary_minus_2_add_3_32_lut_LC_2_24_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_unary_minus_2_add_3_32_lut_LC_2_24_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_unary_minus_2_add_3_32_lut_LC_2_24_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__11570),
            .in3(N__11555),
            .lcout(\eeprom.n3 ),
            .ltout(),
            .carryin(\eeprom.n3815 ),
            .carryout(\eeprom.n3816 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_unary_minus_2_add_3_33_lut_LC_2_24_7 .C_ON=1'b0;
    defparam \eeprom.rem_4_unary_minus_2_add_3_33_lut_LC_2_24_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_unary_minus_2_add_3_33_lut_LC_2_24_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_unary_minus_2_add_3_33_lut_LC_2_24_7  (
            .in0(_gnd_net_),
            .in1(N__24004),
            .in2(_gnd_net_),
            .in3(N__11552),
            .lcout(\eeprom.n2_adj_395 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_mux_3_i20_3_lut_LC_2_25_6 .C_ON=1'b0;
    defparam \eeprom.rem_4_mux_3_i20_3_lut_LC_2_25_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_mux_3_i20_3_lut_LC_2_25_6 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \eeprom.rem_4_mux_3_i20_3_lut_LC_2_25_6  (
            .in0(N__11549),
            .in1(N__22969),
            .in2(_gnd_net_),
            .in3(N__11540),
            .lcout(\eeprom.n2419 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i23_1_lut_LC_2_26_3 .C_ON=1'b0;
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i23_1_lut_LC_2_26_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i23_1_lut_LC_2_26_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \eeprom.rem_4_unary_minus_2_inv_0_i23_1_lut_LC_2_26_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14185),
            .lcout(\eeprom.n11_adj_410 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.add_937_2_lut_LC_3_17_0 .C_ON=1'b1;
    defparam \eeprom.add_937_2_lut_LC_3_17_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.add_937_2_lut_LC_3_17_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.add_937_2_lut_LC_3_17_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__12008),
            .in3(N__11684),
            .lcout(\eeprom.n1343 ),
            .ltout(),
            .carryin(bfn_3_17_0_),
            .carryout(\eeprom.n3448 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.add_937_3_lut_LC_3_17_1 .C_ON=1'b1;
    defparam \eeprom.add_937_3_lut_LC_3_17_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.add_937_3_lut_LC_3_17_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.add_937_3_lut_LC_3_17_1  (
            .in0(_gnd_net_),
            .in1(N__27731),
            .in2(N__12188),
            .in3(N__11681),
            .lcout(\eeprom.n1342 ),
            .ltout(),
            .carryin(\eeprom.n3448 ),
            .carryout(\eeprom.n3449 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.add_937_4_lut_LC_3_17_2 .C_ON=1'b1;
    defparam \eeprom.add_937_4_lut_LC_3_17_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.add_937_4_lut_LC_3_17_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.add_937_4_lut_LC_3_17_2  (
            .in0(_gnd_net_),
            .in1(N__11903),
            .in2(_gnd_net_),
            .in3(N__11678),
            .lcout(\eeprom.n1341 ),
            .ltout(),
            .carryin(\eeprom.n3449 ),
            .carryout(\eeprom.n3450 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.add_937_5_lut_LC_3_17_3 .C_ON=1'b1;
    defparam \eeprom.add_937_5_lut_LC_3_17_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.add_937_5_lut_LC_3_17_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.add_937_5_lut_LC_3_17_3  (
            .in0(_gnd_net_),
            .in1(N__12512),
            .in2(_gnd_net_),
            .in3(N__11675),
            .lcout(\eeprom.n1340 ),
            .ltout(),
            .carryin(\eeprom.n3450 ),
            .carryout(\eeprom.n3451 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.add_937_6_lut_LC_3_17_4 .C_ON=1'b1;
    defparam \eeprom.add_937_6_lut_LC_3_17_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.add_937_6_lut_LC_3_17_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.add_937_6_lut_LC_3_17_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__12137),
            .in3(N__11672),
            .lcout(\eeprom.n1339 ),
            .ltout(),
            .carryin(\eeprom.n3451 ),
            .carryout(\eeprom.n3452 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.add_937_7_lut_LC_3_17_5 .C_ON=1'b1;
    defparam \eeprom.add_937_7_lut_LC_3_17_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.add_937_7_lut_LC_3_17_5 .LUT_INIT=16'b1110101110111110;
    LogicCell40 \eeprom.add_937_7_lut_LC_3_17_5  (
            .in0(N__12524),
            .in1(_gnd_net_),
            .in2(N__12607),
            .in3(N__11669),
            .lcout(\eeprom.n4734 ),
            .ltout(),
            .carryin(\eeprom.n3452 ),
            .carryout(\eeprom.n3453 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.add_937_8_lut_LC_3_17_6 .C_ON=1'b0;
    defparam \eeprom.add_937_8_lut_LC_3_17_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.add_937_8_lut_LC_3_17_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.add_937_8_lut_LC_3_17_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__12488),
            .in3(N__11666),
            .lcout(\eeprom.n1337 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i4_1_lut_LC_3_18_0 .C_ON=1'b0;
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i4_1_lut_LC_3_18_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i4_1_lut_LC_3_18_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \eeprom.rem_4_unary_minus_2_inv_0_i4_1_lut_LC_3_18_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23768),
            .lcout(\eeprom.n30_adj_458 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i520_2_lut_LC_3_18_1 .C_ON=1'b0;
    defparam \eeprom.i520_2_lut_LC_3_18_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.i520_2_lut_LC_3_18_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \eeprom.i520_2_lut_LC_3_18_1  (
            .in0(_gnd_net_),
            .in1(N__22955),
            .in2(_gnd_net_),
            .in3(N__12044),
            .lcout(\eeprom.n1135 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i8_1_lut_LC_3_18_2 .C_ON=1'b0;
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i8_1_lut_LC_3_18_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i8_1_lut_LC_3_18_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \eeprom.rem_4_unary_minus_2_inv_0_i8_1_lut_LC_3_18_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12828),
            .lcout(\eeprom.n26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_mux_3_i31_3_lut_LC_3_18_3 .C_ON=1'b0;
    defparam \eeprom.rem_4_mux_3_i31_3_lut_LC_3_18_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_mux_3_i31_3_lut_LC_3_18_3 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \eeprom.rem_4_mux_3_i31_3_lut_LC_3_18_3  (
            .in0(N__11813),
            .in1(N__22954),
            .in2(_gnd_net_),
            .in3(N__11792),
            .lcout(\eeprom.n1256 ),
            .ltout(\eeprom.n1256_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1224_3_lut_4_lut_LC_3_18_4 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1224_3_lut_4_lut_LC_3_18_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1224_3_lut_4_lut_LC_3_18_4 .LUT_INIT=16'b1010110011001100;
    LogicCell40 \eeprom.rem_4_i1224_3_lut_4_lut_LC_3_18_4  (
            .in0(N__11780),
            .in1(N__11902),
            .in2(N__11774),
            .in3(N__12466),
            .lcout(\eeprom.n1916 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i29_1_lut_LC_3_18_5 .C_ON=1'b0;
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i29_1_lut_LC_3_18_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i29_1_lut_LC_3_18_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \eeprom.rem_4_unary_minus_2_inv_0_i29_1_lut_LC_3_18_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11983),
            .lcout(\eeprom.n5_adj_400 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i19_1_lut_LC_3_18_6 .C_ON=1'b0;
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i19_1_lut_LC_3_18_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i19_1_lut_LC_3_18_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \eeprom.rem_4_unary_minus_2_inv_0_i19_1_lut_LC_3_18_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12330),
            .lcout(\eeprom.n15_adj_415 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i1_1_lut_LC_3_18_7 .C_ON=1'b0;
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i1_1_lut_LC_3_18_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i1_1_lut_LC_3_18_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \eeprom.rem_4_unary_minus_2_inv_0_i1_1_lut_LC_3_18_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23475),
            .lcout(\eeprom.n33 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_mux_3_i26_3_lut_LC_3_19_0 .C_ON=1'b0;
    defparam \eeprom.rem_4_mux_3_i26_3_lut_LC_3_19_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_mux_3_i26_3_lut_LC_3_19_0 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \eeprom.rem_4_mux_3_i26_3_lut_LC_3_19_0  (
            .in0(_gnd_net_),
            .in1(N__22852),
            .in2(N__11732),
            .in3(N__11711),
            .lcout(\eeprom.n1141 ),
            .ltout(\eeprom.n1141_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i1_4_lut_adj_48_LC_3_19_1 .C_ON=1'b0;
    defparam \eeprom.i1_4_lut_adj_48_LC_3_19_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.i1_4_lut_adj_48_LC_3_19_1 .LUT_INIT=16'b1000100010000000;
    LogicCell40 \eeprom.i1_4_lut_adj_48_LC_3_19_1  (
            .in0(N__22853),
            .in1(N__11935),
            .in2(N__11699),
            .in3(N__12205),
            .lcout(),
            .ltout(\eeprom.n4399_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i1_4_lut_adj_49_LC_3_19_2 .C_ON=1'b0;
    defparam \eeprom.i1_4_lut_adj_49_LC_3_19_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.i1_4_lut_adj_49_LC_3_19_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \eeprom.i1_4_lut_adj_49_LC_3_19_2  (
            .in0(N__12043),
            .in1(N__12507),
            .in2(N__12020),
            .in3(N__12130),
            .lcout(\eeprom.n4405 ),
            .ltout(\eeprom.n4405_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1226_3_lut_4_lut_LC_3_19_3 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1226_3_lut_4_lut_LC_3_19_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1226_3_lut_4_lut_LC_3_19_3 .LUT_INIT=16'b1010110011001100;
    LogicCell40 \eeprom.rem_4_i1226_3_lut_4_lut_LC_3_19_3  (
            .in0(N__12017),
            .in1(N__12004),
            .in2(N__11990),
            .in3(N__12605),
            .lcout(\eeprom.n1918 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_mux_3_i29_3_lut_LC_3_19_4 .C_ON=1'b0;
    defparam \eeprom.rem_4_mux_3_i29_3_lut_LC_3_19_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_mux_3_i29_3_lut_LC_3_19_4 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \eeprom.rem_4_mux_3_i29_3_lut_LC_3_19_4  (
            .in0(N__11987),
            .in1(N__22851),
            .in2(_gnd_net_),
            .in3(N__11960),
            .lcout(\eeprom.n1138 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1225_3_lut_4_lut_LC_3_19_5 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1225_3_lut_4_lut_LC_3_19_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1225_3_lut_4_lut_LC_3_19_5 .LUT_INIT=16'b1110101000101010;
    LogicCell40 \eeprom.rem_4_i1225_3_lut_4_lut_LC_3_19_5  (
            .in0(N__12187),
            .in1(N__12606),
            .in2(N__12473),
            .in3(N__11948),
            .lcout(\eeprom.n1917 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_mux_3_i28_3_lut_LC_3_19_6 .C_ON=1'b0;
    defparam \eeprom.rem_4_mux_3_i28_3_lut_LC_3_19_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_mux_3_i28_3_lut_LC_3_19_6 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \eeprom.rem_4_mux_3_i28_3_lut_LC_3_19_6  (
            .in0(_gnd_net_),
            .in1(N__22854),
            .in2(N__11939),
            .in3(N__11920),
            .lcout(\eeprom.n1139 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i9_1_lut_LC_3_19_7 .C_ON=1'b0;
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i9_1_lut_LC_3_19_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i9_1_lut_LC_3_19_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \eeprom.rem_4_unary_minus_2_inv_0_i9_1_lut_LC_3_19_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12393),
            .lcout(\eeprom.n25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_mux_3_i25_3_lut_LC_3_20_0 .C_ON=1'b0;
    defparam \eeprom.rem_4_mux_3_i25_3_lut_LC_3_20_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_mux_3_i25_3_lut_LC_3_20_0 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \eeprom.rem_4_mux_3_i25_3_lut_LC_3_20_0  (
            .in0(_gnd_net_),
            .in1(N__22849),
            .in2(N__11879),
            .in3(N__11862),
            .lcout(\eeprom.n1919 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i25_1_lut_LC_3_20_1 .C_ON=1'b0;
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i25_1_lut_LC_3_20_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i25_1_lut_LC_3_20_1 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \eeprom.rem_4_unary_minus_2_inv_0_i25_1_lut_LC_3_20_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__11864),
            .in3(_gnd_net_),
            .lcout(\eeprom.n9_adj_408 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i2_1_lut_LC_3_20_3 .C_ON=1'b0;
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i2_1_lut_LC_3_20_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i2_1_lut_LC_3_20_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \eeprom.rem_4_unary_minus_2_inv_0_i2_1_lut_LC_3_20_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23901),
            .lcout(\eeprom.n32 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_mux_3_i27_3_lut_LC_3_20_4 .C_ON=1'b0;
    defparam \eeprom.rem_4_mux_3_i27_3_lut_LC_3_20_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_mux_3_i27_3_lut_LC_3_20_4 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \eeprom.rem_4_mux_3_i27_3_lut_LC_3_20_4  (
            .in0(N__12228),
            .in1(_gnd_net_),
            .in2(N__12209),
            .in3(N__22848),
            .lcout(\eeprom.n1140 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_mux_3_i30_3_lut_LC_3_20_5 .C_ON=1'b0;
    defparam \eeprom.rem_4_mux_3_i30_3_lut_LC_3_20_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_mux_3_i30_3_lut_LC_3_20_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \eeprom.rem_4_mux_3_i30_3_lut_LC_3_20_5  (
            .in0(N__22847),
            .in1(N__12166),
            .in2(_gnd_net_),
            .in3(N__12149),
            .lcout(\eeprom.n1137 ),
            .ltout(\eeprom.n1137_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i4030_3_lut_4_lut_LC_3_20_6 .C_ON=1'b0;
    defparam \eeprom.i4030_3_lut_4_lut_LC_3_20_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.i4030_3_lut_4_lut_LC_3_20_6 .LUT_INIT=16'b1101100011110000;
    LogicCell40 \eeprom.i4030_3_lut_4_lut_LC_3_20_6  (
            .in0(N__12608),
            .in1(N__12119),
            .in2(N__12110),
            .in3(N__12470),
            .lcout(\eeprom.n1914 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_mux_3_i10_3_lut_LC_3_20_7 .C_ON=1'b0;
    defparam \eeprom.rem_4_mux_3_i10_3_lut_LC_3_20_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_mux_3_i10_3_lut_LC_3_20_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \eeprom.rem_4_mux_3_i10_3_lut_LC_3_20_7  (
            .in0(N__22850),
            .in1(N__12107),
            .in2(_gnd_net_),
            .in3(N__12095),
            .lcout(\eeprom.n3419 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_mux_3_i1_3_lut_LC_3_21_0 .C_ON=1'b0;
    defparam \eeprom.rem_4_mux_3_i1_3_lut_LC_3_21_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_mux_3_i1_3_lut_LC_3_21_0 .LUT_INIT=16'b0100010001110111;
    LogicCell40 \eeprom.rem_4_mux_3_i1_3_lut_LC_3_21_0  (
            .in0(N__12074),
            .in1(N__22846),
            .in2(_gnd_net_),
            .in3(N__23488),
            .lcout(\eeprom.n1166 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i21_1_lut_LC_3_21_1 .C_ON=1'b0;
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i21_1_lut_LC_3_21_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i21_1_lut_LC_3_21_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \eeprom.rem_4_unary_minus_2_inv_0_i21_1_lut_LC_3_21_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13051),
            .lcout(\eeprom.n13_adj_412 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i32_1_lut_LC_3_21_2 .C_ON=1'b0;
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i32_1_lut_LC_3_21_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i32_1_lut_LC_3_21_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \eeprom.rem_4_unary_minus_2_inv_0_i32_1_lut_LC_3_21_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22845),
            .lcout(\eeprom.n2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i24_1_lut_LC_3_21_7 .C_ON=1'b0;
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i24_1_lut_LC_3_21_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i24_1_lut_LC_3_21_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \eeprom.rem_4_unary_minus_2_inv_0_i24_1_lut_LC_3_21_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12307),
            .lcout(\eeprom.n10_adj_409 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_mux_3_i15_3_lut_LC_3_22_0 .C_ON=1'b0;
    defparam \eeprom.rem_4_mux_3_i15_3_lut_LC_3_22_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_mux_3_i15_3_lut_LC_3_22_0 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \eeprom.rem_4_mux_3_i15_3_lut_LC_3_22_0  (
            .in0(N__12344),
            .in1(N__22923),
            .in2(_gnd_net_),
            .in3(N__13589),
            .lcout(\eeprom.n2919 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i4037_3_lut_LC_3_22_2 .C_ON=1'b0;
    defparam \eeprom.i4037_3_lut_LC_3_22_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.i4037_3_lut_LC_3_22_2 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \eeprom.i4037_3_lut_LC_3_22_2  (
            .in0(_gnd_net_),
            .in1(N__15793),
            .in2(N__12242),
            .in3(N__13100),
            .lcout(\eeprom.n2415 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_mux_3_i19_3_lut_LC_3_22_5 .C_ON=1'b0;
    defparam \eeprom.rem_4_mux_3_i19_3_lut_LC_3_22_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_mux_3_i19_3_lut_LC_3_22_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \eeprom.rem_4_mux_3_i19_3_lut_LC_3_22_5  (
            .in0(N__22921),
            .in1(N__12338),
            .in2(_gnd_net_),
            .in3(N__12314),
            .lcout(\eeprom.n2519 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_mux_3_i24_3_lut_LC_3_22_6 .C_ON=1'b0;
    defparam \eeprom.rem_4_mux_3_i24_3_lut_LC_3_22_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_mux_3_i24_3_lut_LC_3_22_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \eeprom.rem_4_mux_3_i24_3_lut_LC_3_22_6  (
            .in0(N__12308),
            .in1(N__12287),
            .in2(_gnd_net_),
            .in3(N__22920),
            .lcout(\eeprom.n2019 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_mux_3_i16_3_lut_LC_3_22_7 .C_ON=1'b0;
    defparam \eeprom.rem_4_mux_3_i16_3_lut_LC_3_22_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_mux_3_i16_3_lut_LC_3_22_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \eeprom.rem_4_mux_3_i16_3_lut_LC_3_22_7  (
            .in0(N__22922),
            .in1(N__12281),
            .in2(_gnd_net_),
            .in3(N__12275),
            .lcout(\eeprom.n2819 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1553_2_lut_LC_3_23_0 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1553_2_lut_LC_3_23_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1553_2_lut_LC_3_23_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1553_2_lut_LC_3_23_0  (
            .in0(_gnd_net_),
            .in1(N__14004),
            .in2(_gnd_net_),
            .in3(N__12251),
            .lcout(\eeprom.n2386 ),
            .ltout(),
            .carryin(bfn_3_23_0_),
            .carryout(\eeprom.n3551 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1553_3_lut_LC_3_23_1 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1553_3_lut_LC_3_23_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1553_3_lut_LC_3_23_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1553_3_lut_LC_3_23_1  (
            .in0(_gnd_net_),
            .in1(N__27582),
            .in2(N__15584),
            .in3(N__12248),
            .lcout(\eeprom.n2385 ),
            .ltout(),
            .carryin(\eeprom.n3551 ),
            .carryout(\eeprom.n3552 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1553_4_lut_LC_3_23_2 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1553_4_lut_LC_3_23_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1553_4_lut_LC_3_23_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1553_4_lut_LC_3_23_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__15728),
            .in3(N__12245),
            .lcout(\eeprom.n2384 ),
            .ltout(),
            .carryin(\eeprom.n3552 ),
            .carryout(\eeprom.n3553 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1553_5_lut_LC_3_23_3 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1553_5_lut_LC_3_23_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1553_5_lut_LC_3_23_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1553_5_lut_LC_3_23_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__15794),
            .in3(N__12233),
            .lcout(\eeprom.n2383 ),
            .ltout(),
            .carryin(\eeprom.n3553 ),
            .carryout(\eeprom.n3554 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1553_6_lut_LC_3_23_4 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1553_6_lut_LC_3_23_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1553_6_lut_LC_3_23_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1553_6_lut_LC_3_23_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__14159),
            .in3(N__12377),
            .lcout(\eeprom.n2382 ),
            .ltout(),
            .carryin(\eeprom.n3554 ),
            .carryout(\eeprom.n3555 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1553_7_lut_LC_3_23_5 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1553_7_lut_LC_3_23_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1553_7_lut_LC_3_23_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1553_7_lut_LC_3_23_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__15830),
            .in3(N__12374),
            .lcout(\eeprom.n2381 ),
            .ltout(),
            .carryin(\eeprom.n3555 ),
            .carryout(\eeprom.n3556 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1553_8_lut_LC_3_23_6 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1553_8_lut_LC_3_23_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1553_8_lut_LC_3_23_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1553_8_lut_LC_3_23_6  (
            .in0(_gnd_net_),
            .in1(N__14228),
            .in2(_gnd_net_),
            .in3(N__12371),
            .lcout(\eeprom.n2380 ),
            .ltout(),
            .carryin(\eeprom.n3556 ),
            .carryout(\eeprom.n3557 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1553_9_lut_LC_3_23_7 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1553_9_lut_LC_3_23_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1553_9_lut_LC_3_23_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1553_9_lut_LC_3_23_7  (
            .in0(_gnd_net_),
            .in1(N__13172),
            .in2(N__27784),
            .in3(N__12368),
            .lcout(\eeprom.n2379 ),
            .ltout(),
            .carryin(\eeprom.n3557 ),
            .carryout(\eeprom.n3558 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1553_10_lut_LC_3_24_0 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1553_10_lut_LC_3_24_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1553_10_lut_LC_3_24_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1553_10_lut_LC_3_24_0  (
            .in0(_gnd_net_),
            .in1(N__27732),
            .in2(N__14129),
            .in3(N__12365),
            .lcout(\eeprom.n2378 ),
            .ltout(),
            .carryin(bfn_3_24_0_),
            .carryout(\eeprom.n3559 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1553_11_lut_LC_3_24_1 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1553_11_lut_LC_3_24_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1553_11_lut_LC_3_24_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1553_11_lut_LC_3_24_1  (
            .in0(_gnd_net_),
            .in1(N__13979),
            .in2(N__27783),
            .in3(N__12362),
            .lcout(\eeprom.n2377 ),
            .ltout(),
            .carryin(\eeprom.n3559 ),
            .carryout(\eeprom.n3560 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1553_12_lut_LC_3_24_2 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1553_12_lut_LC_3_24_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1553_12_lut_LC_3_24_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1553_12_lut_LC_3_24_2  (
            .in0(_gnd_net_),
            .in1(N__14036),
            .in2(N__27785),
            .in3(N__12359),
            .lcout(\eeprom.n2376 ),
            .ltout(),
            .carryin(\eeprom.n3560 ),
            .carryout(\eeprom.n3561 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1553_13_lut_LC_3_24_3 .C_ON=1'b0;
    defparam \eeprom.rem_4_add_1553_13_lut_LC_3_24_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1553_13_lut_LC_3_24_3 .LUT_INIT=16'b1001000001100000;
    LogicCell40 \eeprom.rem_4_add_1553_13_lut_LC_3_24_3  (
            .in0(N__16523),
            .in1(N__27742),
            .in2(N__13115),
            .in3(N__12356),
            .lcout(\eeprom.n2407 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1566_3_lut_LC_3_24_5 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1566_3_lut_LC_3_24_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1566_3_lut_LC_3_24_5 .LUT_INIT=16'b1111101000001010;
    LogicCell40 \eeprom.rem_4_i1566_3_lut_LC_3_24_5  (
            .in0(N__14012),
            .in1(_gnd_net_),
            .in2(N__13114),
            .in3(N__12353),
            .lcout(\eeprom.n2418 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i4035_3_lut_LC_3_24_6 .C_ON=1'b0;
    defparam \eeprom.i4035_3_lut_LC_3_24_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.i4035_3_lut_LC_3_24_6 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \eeprom.i4035_3_lut_LC_3_24_6  (
            .in0(_gnd_net_),
            .in1(N__12545),
            .in2(N__15829),
            .in3(N__13090),
            .lcout(\eeprom.n2413 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1564_3_lut_LC_3_24_7 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1564_3_lut_LC_3_24_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1564_3_lut_LC_3_24_7 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \eeprom.rem_4_i1564_3_lut_LC_3_24_7  (
            .in0(_gnd_net_),
            .in1(N__12539),
            .in2(N__13113),
            .in3(N__15727),
            .lcout(\eeprom.n2416 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1558_3_lut_LC_3_25_5 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1558_3_lut_LC_3_25_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1558_3_lut_LC_3_25_5 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \eeprom.rem_4_i1558_3_lut_LC_3_25_5  (
            .in0(_gnd_net_),
            .in1(N__14127),
            .in2(N__12533),
            .in3(N__13118),
            .lcout(\eeprom.n2410 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i3948_1_lut_LC_4_18_0 .C_ON=1'b0;
    defparam \eeprom.i3948_1_lut_LC_4_18_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.i3948_1_lut_LC_4_18_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \eeprom.i3948_1_lut_LC_4_18_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12459),
            .lcout(\eeprom.n4733 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1223_3_lut_4_lut_LC_4_18_1 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1223_3_lut_4_lut_LC_4_18_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1223_3_lut_4_lut_LC_4_18_1 .LUT_INIT=16'b1011111110000000;
    LogicCell40 \eeprom.rem_4_i1223_3_lut_4_lut_LC_4_18_1  (
            .in0(N__12518),
            .in1(N__12598),
            .in2(N__12471),
            .in3(N__12511),
            .lcout(\eeprom.n1915 ),
            .ltout(\eeprom.n1915_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i1_2_lut_3_lut_LC_4_18_2 .C_ON=1'b0;
    defparam \eeprom.i1_2_lut_3_lut_LC_4_18_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.i1_2_lut_3_lut_LC_4_18_2 .LUT_INIT=16'b1010000000000000;
    LogicCell40 \eeprom.i1_2_lut_3_lut_LC_4_18_2  (
            .in0(N__12599),
            .in1(_gnd_net_),
            .in2(N__12491),
            .in3(N__12616),
            .lcout(\eeprom.n4437 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1220_3_lut_4_lut_LC_4_18_3 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1220_3_lut_4_lut_LC_4_18_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1220_3_lut_4_lut_LC_4_18_3 .LUT_INIT=16'b1110101000101010;
    LogicCell40 \eeprom.rem_4_i1220_3_lut_4_lut_LC_4_18_3  (
            .in0(N__12487),
            .in1(N__12600),
            .in2(N__12472),
            .in3(N__12434),
            .lcout(\eeprom.n1912 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i22_1_lut_LC_4_18_4 .C_ON=1'b0;
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i22_1_lut_LC_4_18_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i22_1_lut_LC_4_18_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \eeprom.rem_4_unary_minus_2_inv_0_i22_1_lut_LC_4_18_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15616),
            .lcout(\eeprom.n12_adj_411 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_mux_3_i9_3_lut_LC_4_18_5 .C_ON=1'b0;
    defparam \eeprom.rem_4_mux_3_i9_3_lut_LC_4_18_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_mux_3_i9_3_lut_LC_4_18_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \eeprom.rem_4_mux_3_i9_3_lut_LC_4_18_5  (
            .in0(N__22957),
            .in1(N__12410),
            .in2(_gnd_net_),
            .in3(N__12398),
            .lcout(\eeprom.n3519_adj_379 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_mux_3_i18_3_lut_LC_4_18_6 .C_ON=1'b0;
    defparam \eeprom.rem_4_mux_3_i18_3_lut_LC_4_18_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_mux_3_i18_3_lut_LC_4_18_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \eeprom.rem_4_mux_3_i18_3_lut_LC_4_18_6  (
            .in0(N__12665),
            .in1(N__12635),
            .in2(_gnd_net_),
            .in3(N__22956),
            .lcout(\eeprom.n2619 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i3950_2_lut_LC_4_18_7 .C_ON=1'b0;
    defparam \eeprom.i3950_2_lut_LC_4_18_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.i3950_2_lut_LC_4_18_7 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \eeprom.i3950_2_lut_LC_4_18_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__12620),
            .in3(N__12601),
            .lcout(\eeprom.n1913 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1285_2_lut_LC_4_19_0 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1285_2_lut_LC_4_19_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1285_2_lut_LC_4_19_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1285_2_lut_LC_4_19_0  (
            .in0(_gnd_net_),
            .in1(N__12975),
            .in2(_gnd_net_),
            .in3(N__12566),
            .lcout(\eeprom.n1986 ),
            .ltout(),
            .carryin(bfn_4_19_0_),
            .carryout(\eeprom.n3517 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1285_3_lut_LC_4_19_1 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1285_3_lut_LC_4_19_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1285_3_lut_LC_4_19_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1285_3_lut_LC_4_19_1  (
            .in0(_gnd_net_),
            .in1(N__27730),
            .in2(N__12767),
            .in3(N__12563),
            .lcout(\eeprom.n1985 ),
            .ltout(),
            .carryin(\eeprom.n3517 ),
            .carryout(\eeprom.n3518 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1285_4_lut_LC_4_19_2 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1285_4_lut_LC_4_19_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1285_4_lut_LC_4_19_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1285_4_lut_LC_4_19_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__12794),
            .in3(N__12560),
            .lcout(\eeprom.n1984 ),
            .ltout(),
            .carryin(\eeprom.n3518 ),
            .carryout(\eeprom.n3519 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1285_5_lut_LC_4_19_3 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1285_5_lut_LC_4_19_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1285_5_lut_LC_4_19_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1285_5_lut_LC_4_19_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__12727),
            .in3(N__12557),
            .lcout(\eeprom.n1983 ),
            .ltout(),
            .carryin(\eeprom.n3519 ),
            .carryout(\eeprom.n3520 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1285_6_lut_LC_4_19_4 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1285_6_lut_LC_4_19_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1285_6_lut_LC_4_19_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1285_6_lut_LC_4_19_4  (
            .in0(_gnd_net_),
            .in1(N__13009),
            .in2(_gnd_net_),
            .in3(N__12554),
            .lcout(\eeprom.n1982 ),
            .ltout(),
            .carryin(\eeprom.n3520 ),
            .carryout(\eeprom.n3521 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1285_7_lut_LC_4_19_5 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1285_7_lut_LC_4_19_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1285_7_lut_LC_4_19_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1285_7_lut_LC_4_19_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__12686),
            .in3(N__12551),
            .lcout(\eeprom.n1981 ),
            .ltout(),
            .carryin(\eeprom.n3521 ),
            .carryout(\eeprom.n3522 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1285_8_lut_LC_4_19_6 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1285_8_lut_LC_4_19_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1285_8_lut_LC_4_19_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1285_8_lut_LC_4_19_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__12946),
            .in3(N__12548),
            .lcout(\eeprom.n1980 ),
            .ltout(),
            .carryin(\eeprom.n3522 ),
            .carryout(\eeprom.n3523 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1285_9_lut_LC_4_19_7 .C_ON=1'b0;
    defparam \eeprom.rem_4_add_1285_9_lut_LC_4_19_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1285_9_lut_LC_4_19_7 .LUT_INIT=16'b1001000001100000;
    LogicCell40 \eeprom.rem_4_add_1285_9_lut_LC_4_19_7  (
            .in0(N__27383),
            .in1(N__12742),
            .in2(N__12929),
            .in3(N__12851),
            .lcout(\eeprom.n2011 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_mux_3_i8_3_lut_LC_4_20_0 .C_ON=1'b0;
    defparam \eeprom.rem_4_mux_3_i8_3_lut_LC_4_20_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_mux_3_i8_3_lut_LC_4_20_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \eeprom.rem_4_mux_3_i8_3_lut_LC_4_20_0  (
            .in0(N__22943),
            .in1(N__12848),
            .in2(_gnd_net_),
            .in3(N__12836),
            .lcout(\eeprom.n3619_adj_352 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1292_3_lut_LC_4_20_1 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1292_3_lut_LC_4_20_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1292_3_lut_LC_4_20_1 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \eeprom.rem_4_i1292_3_lut_LC_4_20_1  (
            .in0(N__12793),
            .in1(_gnd_net_),
            .in2(N__12812),
            .in3(N__12911),
            .lcout(\eeprom.n2016 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1293_3_lut_LC_4_20_2 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1293_3_lut_LC_4_20_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1293_3_lut_LC_4_20_2 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \eeprom.rem_4_i1293_3_lut_LC_4_20_2  (
            .in0(N__12803),
            .in1(_gnd_net_),
            .in2(N__12926),
            .in3(N__12766),
            .lcout(\eeprom.n2017 ),
            .ltout(\eeprom.n2017_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i1_3_lut_adj_68_LC_4_20_3 .C_ON=1'b0;
    defparam \eeprom.i1_3_lut_adj_68_LC_4_20_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.i1_3_lut_adj_68_LC_4_20_3 .LUT_INIT=16'b1100000000000000;
    LogicCell40 \eeprom.i1_3_lut_adj_68_LC_4_20_3  (
            .in0(_gnd_net_),
            .in1(N__13632),
            .in2(N__12797),
            .in3(N__13743),
            .lcout(\eeprom.n4415 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i1_4_lut_adj_65_LC_4_20_5 .C_ON=1'b0;
    defparam \eeprom.i1_4_lut_adj_65_LC_4_20_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.i1_4_lut_adj_65_LC_4_20_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \eeprom.i1_4_lut_adj_65_LC_4_20_5  (
            .in0(N__12792),
            .in1(N__12681),
            .in2(N__12728),
            .in3(N__12776),
            .lcout(),
            .ltout(\eeprom.n4441_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i3028_4_lut_LC_4_20_6 .C_ON=1'b0;
    defparam \eeprom.i3028_4_lut_LC_4_20_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.i3028_4_lut_LC_4_20_6 .LUT_INIT=16'b1111111111100000;
    LogicCell40 \eeprom.i3028_4_lut_LC_4_20_6  (
            .in0(N__12765),
            .in1(N__12976),
            .in2(N__12746),
            .in3(N__12743),
            .lcout(\eeprom.n1945 ),
            .ltout(\eeprom.n1945_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1291_3_lut_LC_4_20_7 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1291_3_lut_LC_4_20_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1291_3_lut_LC_4_20_7 .LUT_INIT=16'b1111101000001010;
    LogicCell40 \eeprom.rem_4_i1291_3_lut_LC_4_20_7  (
            .in0(N__12726),
            .in1(_gnd_net_),
            .in2(N__12704),
            .in3(N__12701),
            .lcout(\eeprom.n2015 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i4031_3_lut_LC_4_21_0 .C_ON=1'b0;
    defparam \eeprom.i4031_3_lut_LC_4_21_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.i4031_3_lut_LC_4_21_0 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \eeprom.i4031_3_lut_LC_4_21_0  (
            .in0(_gnd_net_),
            .in1(N__12695),
            .in2(N__12928),
            .in3(N__12685),
            .lcout(\eeprom.n2013 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1290_3_lut_LC_4_21_1 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1290_3_lut_LC_4_21_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1290_3_lut_LC_4_21_1 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \eeprom.rem_4_i1290_3_lut_LC_4_21_1  (
            .in0(_gnd_net_),
            .in1(N__13013),
            .in2(N__12998),
            .in3(N__12916),
            .lcout(\eeprom.n2014 ),
            .ltout(\eeprom.n2014_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i1_4_lut_adj_70_LC_4_21_2 .C_ON=1'b0;
    defparam \eeprom.i1_4_lut_adj_70_LC_4_21_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.i1_4_lut_adj_70_LC_4_21_2 .LUT_INIT=16'b1110000000000000;
    LogicCell40 \eeprom.i1_4_lut_adj_70_LC_4_21_2  (
            .in0(N__14064),
            .in1(N__13674),
            .in2(N__12986),
            .in3(N__12983),
            .lcout(\eeprom.n4419 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1294_3_lut_LC_4_21_3 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1294_3_lut_LC_4_21_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1294_3_lut_LC_4_21_3 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \eeprom.rem_4_i1294_3_lut_LC_4_21_3  (
            .in0(_gnd_net_),
            .in1(N__12977),
            .in2(N__12959),
            .in3(N__12915),
            .lcout(\eeprom.n2018 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i3_4_lut_adj_80_LC_4_21_5 .C_ON=1'b0;
    defparam \eeprom.i3_4_lut_adj_80_LC_4_21_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.i3_4_lut_adj_80_LC_4_21_5 .LUT_INIT=16'b1111111011110000;
    LogicCell40 \eeprom.i3_4_lut_adj_80_LC_4_21_5  (
            .in0(N__15180),
            .in1(N__15144),
            .in2(N__15370),
            .in3(N__12869),
            .lcout(\eeprom.n11_adj_473 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1288_3_lut_LC_4_21_6 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1288_3_lut_LC_4_21_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1288_3_lut_LC_4_21_6 .LUT_INIT=16'b1111101000001010;
    LogicCell40 \eeprom.rem_4_i1288_3_lut_LC_4_21_6  (
            .in0(N__12947),
            .in1(_gnd_net_),
            .in2(N__12927),
            .in3(N__12887),
            .lcout(\eeprom.n2012 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i1_4_lut_adj_71_LC_4_22_0 .C_ON=1'b0;
    defparam \eeprom.i1_4_lut_adj_71_LC_4_22_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.i1_4_lut_adj_71_LC_4_22_0 .LUT_INIT=16'b1111111011101110;
    LogicCell40 \eeprom.i1_4_lut_adj_71_LC_4_22_0  (
            .in0(N__13843),
            .in1(N__13792),
            .in2(N__13885),
            .in3(N__12878),
            .lcout(\eeprom.n2044 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i1_2_lut_adj_78_LC_4_22_1 .C_ON=1'b0;
    defparam \eeprom.i1_2_lut_adj_78_LC_4_22_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.i1_2_lut_adj_78_LC_4_22_1 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \eeprom.i1_2_lut_adj_78_LC_4_22_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__15006),
            .in3(N__15537),
            .lcout(),
            .ltout(\eeprom.n4575_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i1_4_lut_adj_79_LC_4_22_2 .C_ON=1'b0;
    defparam \eeprom.i1_4_lut_adj_79_LC_4_22_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.i1_4_lut_adj_79_LC_4_22_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \eeprom.i1_4_lut_adj_79_LC_4_22_2  (
            .in0(N__15096),
            .in1(N__15051),
            .in2(N__12872),
            .in3(N__14958),
            .lcout(\eeprom.n4579 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_mux_3_i21_3_lut_LC_4_22_4 .C_ON=1'b0;
    defparam \eeprom.rem_4_mux_3_i21_3_lut_LC_4_22_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_mux_3_i21_3_lut_LC_4_22_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \eeprom.rem_4_mux_3_i21_3_lut_LC_4_22_4  (
            .in0(N__12863),
            .in1(N__13055),
            .in2(_gnd_net_),
            .in3(N__22959),
            .lcout(\eeprom.n2319 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1632_3_lut_LC_4_22_5 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1632_3_lut_LC_4_22_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1632_3_lut_LC_4_22_5 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \eeprom.rem_4_i1632_3_lut_LC_4_22_5  (
            .in0(_gnd_net_),
            .in1(N__13324),
            .in2(N__13304),
            .in3(N__15961),
            .lcout(\eeprom.n2516 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1630_3_lut_LC_4_22_7 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1630_3_lut_LC_4_22_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1630_3_lut_LC_4_22_7 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \eeprom.rem_4_i1630_3_lut_LC_4_22_7  (
            .in0(_gnd_net_),
            .in1(N__13254),
            .in2(N__13232),
            .in3(N__15960),
            .lcout(\eeprom.n2514 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i1_3_lut_adj_74_LC_4_23_0 .C_ON=1'b0;
    defparam \eeprom.i1_3_lut_adj_74_LC_4_23_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.i1_3_lut_adj_74_LC_4_23_0 .LUT_INIT=16'b1100000000000000;
    LogicCell40 \eeprom.i1_3_lut_adj_74_LC_4_23_0  (
            .in0(_gnd_net_),
            .in1(N__13320),
            .in2(N__13288),
            .in3(N__13209),
            .lcout(),
            .ltout(\eeprom.n4479_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i1_4_lut_adj_75_LC_4_23_1 .C_ON=1'b0;
    defparam \eeprom.i1_4_lut_adj_75_LC_4_23_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.i1_4_lut_adj_75_LC_4_23_1 .LUT_INIT=16'b1110000000000000;
    LogicCell40 \eeprom.i1_4_lut_adj_75_LC_4_23_1  (
            .in0(N__13720),
            .in1(N__13359),
            .in2(N__13031),
            .in3(N__13028),
            .lcout(\eeprom.n4133 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i1_2_lut_adj_73_LC_4_23_2 .C_ON=1'b0;
    defparam \eeprom.i1_2_lut_adj_73_LC_4_23_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.i1_2_lut_adj_73_LC_4_23_2 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \eeprom.i1_2_lut_adj_73_LC_4_23_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__13255),
            .in3(N__16083),
            .lcout(\eeprom.n4477 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i5_4_lut_LC_4_23_3 .C_ON=1'b0;
    defparam \eeprom.i5_4_lut_LC_4_23_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.i5_4_lut_LC_4_23_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \eeprom.i5_4_lut_LC_4_23_3  (
            .in0(N__13171),
            .in1(N__13730),
            .in2(N__14128),
            .in3(N__13985),
            .lcout(\eeprom.n2341 ),
            .ltout(\eeprom.n2341_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1565_3_lut_LC_4_23_4 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1565_3_lut_LC_4_23_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1565_3_lut_LC_4_23_4 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \eeprom.rem_4_i1565_3_lut_LC_4_23_4  (
            .in0(N__13022),
            .in1(_gnd_net_),
            .in2(N__13016),
            .in3(N__15583),
            .lcout(\eeprom.n2417 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1629_3_lut_LC_4_23_5 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1629_3_lut_LC_4_23_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1629_3_lut_LC_4_23_5 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \eeprom.rem_4_i1629_3_lut_LC_4_23_5  (
            .in0(_gnd_net_),
            .in1(N__13196),
            .in2(N__13216),
            .in3(N__15931),
            .lcout(\eeprom.n2513 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1631_3_lut_LC_4_23_6 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1631_3_lut_LC_4_23_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1631_3_lut_LC_4_23_6 .LUT_INIT=16'b1111101000001010;
    LogicCell40 \eeprom.rem_4_i1631_3_lut_LC_4_23_6  (
            .in0(N__13284),
            .in1(_gnd_net_),
            .in2(N__15959),
            .in3(N__13268),
            .lcout(\eeprom.n2515 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1633_3_lut_LC_4_23_7 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1633_3_lut_LC_4_23_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1633_3_lut_LC_4_23_7 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \eeprom.rem_4_i1633_3_lut_LC_4_23_7  (
            .in0(_gnd_net_),
            .in1(N__13360),
            .in2(N__13343),
            .in3(N__15935),
            .lcout(\eeprom.n2517 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1556_3_lut_LC_4_24_0 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1556_3_lut_LC_4_24_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1556_3_lut_LC_4_24_0 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \eeprom.rem_4_i1556_3_lut_LC_4_24_0  (
            .in0(_gnd_net_),
            .in1(N__13178),
            .in2(N__13117),
            .in3(N__14034),
            .lcout(\eeprom.n2408 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1492_3_lut_LC_4_24_1 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1492_3_lut_LC_4_24_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1492_3_lut_LC_4_24_1 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \eeprom.rem_4_i1492_3_lut_LC_4_24_1  (
            .in0(_gnd_net_),
            .in1(N__16115),
            .in2(N__16727),
            .in3(N__16603),
            .lcout(\eeprom.n2312 ),
            .ltout(\eeprom.n2312_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1559_3_lut_LC_4_24_2 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1559_3_lut_LC_4_24_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1559_3_lut_LC_4_24_2 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \eeprom.rem_4_i1559_3_lut_LC_4_24_2  (
            .in0(N__13102),
            .in1(_gnd_net_),
            .in2(N__13160),
            .in3(N__13157),
            .lcout(\eeprom.n2411 ),
            .ltout(\eeprom.n2411_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i5_4_lut_adj_76_LC_4_24_3 .C_ON=1'b0;
    defparam \eeprom.i5_4_lut_adj_76_LC_4_24_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.i5_4_lut_adj_76_LC_4_24_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \eeprom.i5_4_lut_adj_76_LC_4_24_3  (
            .in0(N__13375),
            .in1(N__13413),
            .in2(N__13151),
            .in3(N__13148),
            .lcout(),
            .ltout(\eeprom.n12_adj_472_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i6_4_lut_adj_77_LC_4_24_4 .C_ON=1'b0;
    defparam \eeprom.i6_4_lut_adj_77_LC_4_24_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.i6_4_lut_adj_77_LC_4_24_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \eeprom.i6_4_lut_adj_77_LC_4_24_4  (
            .in0(N__16014),
            .in1(N__13429),
            .in2(N__13142),
            .in3(N__15685),
            .lcout(\eeprom.n2440 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1562_3_lut_LC_4_24_5 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1562_3_lut_LC_4_24_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1562_3_lut_LC_4_24_5 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \eeprom.rem_4_i1562_3_lut_LC_4_24_5  (
            .in0(_gnd_net_),
            .in1(N__13139),
            .in2(N__14155),
            .in3(N__13101),
            .lcout(\eeprom.n2414 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1557_3_lut_LC_4_24_6 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1557_3_lut_LC_4_24_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1557_3_lut_LC_4_24_6 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \eeprom.rem_4_i1557_3_lut_LC_4_24_6  (
            .in0(_gnd_net_),
            .in1(N__13133),
            .in2(N__13116),
            .in3(N__13978),
            .lcout(\eeprom.n2409 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1560_3_lut_LC_4_24_7 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1560_3_lut_LC_4_24_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1560_3_lut_LC_4_24_7 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \eeprom.rem_4_i1560_3_lut_LC_4_24_7  (
            .in0(_gnd_net_),
            .in1(N__14224),
            .in2(N__13127),
            .in3(N__13103),
            .lcout(\eeprom.n2412 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1620_2_lut_LC_4_25_0 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1620_2_lut_LC_4_25_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1620_2_lut_LC_4_25_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1620_2_lut_LC_4_25_0  (
            .in0(_gnd_net_),
            .in1(N__13719),
            .in2(_gnd_net_),
            .in3(N__13364),
            .lcout(\eeprom.n2486 ),
            .ltout(),
            .carryin(bfn_4_25_0_),
            .carryout(\eeprom.n3562 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1620_3_lut_LC_4_25_1 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1620_3_lut_LC_4_25_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1620_3_lut_LC_4_25_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1620_3_lut_LC_4_25_1  (
            .in0(_gnd_net_),
            .in1(N__27371),
            .in2(N__13361),
            .in3(N__13331),
            .lcout(\eeprom.n2485 ),
            .ltout(),
            .carryin(\eeprom.n3562 ),
            .carryout(\eeprom.n3563 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1620_4_lut_LC_4_25_2 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1620_4_lut_LC_4_25_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1620_4_lut_LC_4_25_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1620_4_lut_LC_4_25_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__13328),
            .in3(N__13292),
            .lcout(\eeprom.n2484 ),
            .ltout(),
            .carryin(\eeprom.n3563 ),
            .carryout(\eeprom.n3564 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1620_5_lut_LC_4_25_3 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1620_5_lut_LC_4_25_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1620_5_lut_LC_4_25_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1620_5_lut_LC_4_25_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__13289),
            .in3(N__13259),
            .lcout(\eeprom.n2483 ),
            .ltout(),
            .carryin(\eeprom.n3564 ),
            .carryout(\eeprom.n3565 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1620_6_lut_LC_4_25_4 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1620_6_lut_LC_4_25_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1620_6_lut_LC_4_25_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1620_6_lut_LC_4_25_4  (
            .in0(_gnd_net_),
            .in1(N__13256),
            .in2(_gnd_net_),
            .in3(N__13220),
            .lcout(\eeprom.n2482 ),
            .ltout(),
            .carryin(\eeprom.n3565 ),
            .carryout(\eeprom.n3566 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1620_7_lut_LC_4_25_5 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1620_7_lut_LC_4_25_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1620_7_lut_LC_4_25_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1620_7_lut_LC_4_25_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__13217),
            .in3(N__13187),
            .lcout(\eeprom.n2481 ),
            .ltout(),
            .carryin(\eeprom.n3566 ),
            .carryout(\eeprom.n3567 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1620_8_lut_LC_4_25_6 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1620_8_lut_LC_4_25_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1620_8_lut_LC_4_25_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1620_8_lut_LC_4_25_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__16090),
            .in3(N__13184),
            .lcout(\eeprom.n2480 ),
            .ltout(),
            .carryin(\eeprom.n3567 ),
            .carryout(\eeprom.n3568 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1620_9_lut_LC_4_25_7 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1620_9_lut_LC_4_25_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1620_9_lut_LC_4_25_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1620_9_lut_LC_4_25_7  (
            .in0(_gnd_net_),
            .in1(N__15684),
            .in2(N__27581),
            .in3(N__13181),
            .lcout(\eeprom.n2479 ),
            .ltout(),
            .carryin(\eeprom.n3568 ),
            .carryout(\eeprom.n3569 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1620_10_lut_LC_4_26_0 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1620_10_lut_LC_4_26_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1620_10_lut_LC_4_26_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1620_10_lut_LC_4_26_0  (
            .in0(_gnd_net_),
            .in1(N__13531),
            .in2(N__27744),
            .in3(N__13445),
            .lcout(\eeprom.n2478 ),
            .ltout(),
            .carryin(bfn_4_26_0_),
            .carryout(\eeprom.n3570 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1620_11_lut_LC_4_26_1 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1620_11_lut_LC_4_26_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1620_11_lut_LC_4_26_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1620_11_lut_LC_4_26_1  (
            .in0(_gnd_net_),
            .in1(N__13414),
            .in2(N__27746),
            .in3(N__13442),
            .lcout(\eeprom.n2477 ),
            .ltout(),
            .carryin(\eeprom.n3570 ),
            .carryout(\eeprom.n3571 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1620_12_lut_LC_4_26_2 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1620_12_lut_LC_4_26_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1620_12_lut_LC_4_26_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1620_12_lut_LC_4_26_2  (
            .in0(_gnd_net_),
            .in1(N__13381),
            .in2(N__27745),
            .in3(N__13439),
            .lcout(\eeprom.n2476 ),
            .ltout(),
            .carryin(\eeprom.n3571 ),
            .carryout(\eeprom.n3572 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1620_13_lut_LC_4_26_3 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1620_13_lut_LC_4_26_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1620_13_lut_LC_4_26_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1620_13_lut_LC_4_26_3  (
            .in0(_gnd_net_),
            .in1(N__16021),
            .in2(N__27747),
            .in3(N__13436),
            .lcout(\eeprom.n2475 ),
            .ltout(),
            .carryin(\eeprom.n3572 ),
            .carryout(\eeprom.n3573 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1620_14_lut_LC_4_26_4 .C_ON=1'b0;
    defparam \eeprom.rem_4_add_1620_14_lut_LC_4_26_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1620_14_lut_LC_4_26_4 .LUT_INIT=16'b1001000001100000;
    LogicCell40 \eeprom.rem_4_add_1620_14_lut_LC_4_26_4  (
            .in0(N__27620),
            .in1(N__13433),
            .in2(N__15977),
            .in3(N__13418),
            .lcout(\eeprom.n2506 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1625_3_lut_LC_4_26_5 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1625_3_lut_LC_4_26_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1625_3_lut_LC_4_26_5 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \eeprom.rem_4_i1625_3_lut_LC_4_26_5  (
            .in0(_gnd_net_),
            .in1(N__13415),
            .in2(N__13400),
            .in3(N__15963),
            .lcout(\eeprom.n2509 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1624_3_lut_LC_4_26_7 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1624_3_lut_LC_4_26_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1624_3_lut_LC_4_26_7 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \eeprom.rem_4_i1624_3_lut_LC_4_26_7  (
            .in0(_gnd_net_),
            .in1(N__13391),
            .in2(N__13385),
            .in3(N__15962),
            .lcout(\eeprom.n2508 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i3982_4_lut_LC_4_31_0.C_ON=1'b0;
    defparam i3982_4_lut_LC_4_31_0.SEQ_MODE=4'b0000;
    defparam i3982_4_lut_LC_4_31_0.LUT_INIT=16'b1111110111100000;
    LogicCell40 i3982_4_lut_LC_4_31_0 (
            .in0(N__14783),
            .in1(N__14744),
            .in2(N__14804),
            .in3(N__14764),
            .lcout(n4826),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i3981_4_lut_LC_4_31_3.C_ON=1'b0;
    defparam i3981_4_lut_LC_4_31_3.SEQ_MODE=4'b0000;
    defparam i3981_4_lut_LC_4_31_3.LUT_INIT=16'b1101110101000000;
    LogicCell40 i3981_4_lut_LC_4_31_3 (
            .in0(N__14743),
            .in1(N__14782),
            .in2(N__14765),
            .in3(N__14800),
            .lcout(),
            .ltout(n4825_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i3983_3_lut_LC_4_31_4.C_ON=1'b0;
    defparam i3983_3_lut_LC_4_31_4.SEQ_MODE=4'b0000;
    defparam i3983_3_lut_LC_4_31_4.LUT_INIT=16'b0011001100001111;
    LogicCell40 i3983_3_lut_LC_4_31_4 (
            .in0(_gnd_net_),
            .in1(N__13505),
            .in2(N__13499),
            .in3(N__14723),
            .lcout(LED_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_mux_3_i11_3_lut_LC_5_18_2 .C_ON=1'b0;
    defparam \eeprom.rem_4_mux_3_i11_3_lut_LC_5_18_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_mux_3_i11_3_lut_LC_5_18_2 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \eeprom.rem_4_mux_3_i11_3_lut_LC_5_18_2  (
            .in0(N__13487),
            .in1(N__22958),
            .in2(_gnd_net_),
            .in3(N__13475),
            .lcout(\eeprom.n3319 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1700_3_lut_LC_5_19_0 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1700_3_lut_LC_5_19_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1700_3_lut_LC_5_19_0 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \eeprom.rem_4_i1700_3_lut_LC_5_19_0  (
            .in0(_gnd_net_),
            .in1(N__15080),
            .in2(N__15518),
            .in3(N__15112),
            .lcout(\eeprom.n2616 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1699_3_lut_LC_5_19_1 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1699_3_lut_LC_5_19_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1699_3_lut_LC_5_19_1 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \eeprom.rem_4_i1699_3_lut_LC_5_19_1  (
            .in0(_gnd_net_),
            .in1(N__15504),
            .in2(N__15035),
            .in3(N__15067),
            .lcout(\eeprom.n2615 ),
            .ltout(\eeprom.n2615_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i1_2_lut_adj_83_LC_5_19_2 .C_ON=1'b0;
    defparam \eeprom.i1_2_lut_adj_83_LC_5_19_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.i1_2_lut_adj_83_LC_5_19_2 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \eeprom.i1_2_lut_adj_83_LC_5_19_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__13454),
            .in3(N__16413),
            .lcout(),
            .ltout(\eeprom.n4497_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i1_4_lut_adj_84_LC_5_19_3 .C_ON=1'b0;
    defparam \eeprom.i1_4_lut_adj_84_LC_5_19_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.i1_4_lut_adj_84_LC_5_19_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \eeprom.i1_4_lut_adj_84_LC_5_19_3  (
            .in0(N__16884),
            .in1(N__16842),
            .in2(N__13451),
            .in3(N__16908),
            .lcout(),
            .ltout(\eeprom.n4501_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i3_4_lut_adj_86_LC_5_19_4 .C_ON=1'b0;
    defparam \eeprom.i3_4_lut_adj_86_LC_5_19_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.i3_4_lut_adj_86_LC_5_19_4 .LUT_INIT=16'b1111110011101100;
    LogicCell40 \eeprom.i3_4_lut_adj_86_LC_5_19_4  (
            .in0(N__16762),
            .in1(N__14874),
            .in2(N__13448),
            .in3(N__16809),
            .lcout(\eeprom.n12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1701_3_lut_LC_5_19_5 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1701_3_lut_LC_5_19_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1701_3_lut_LC_5_19_5 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \eeprom.rem_4_i1701_3_lut_LC_5_19_5  (
            .in0(_gnd_net_),
            .in1(N__15125),
            .in2(N__15152),
            .in3(N__15500),
            .lcout(\eeprom.n2617 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1698_3_lut_LC_5_20_0 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1698_3_lut_LC_5_20_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1698_3_lut_LC_5_20_0 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \eeprom.rem_4_i1698_3_lut_LC_5_20_0  (
            .in0(_gnd_net_),
            .in1(N__14981),
            .in2(N__15020),
            .in3(N__15505),
            .lcout(\eeprom.n2614 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1693_3_lut_LC_5_20_1 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1693_3_lut_LC_5_20_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1693_3_lut_LC_5_20_1 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \eeprom.rem_4_i1693_3_lut_LC_5_20_1  (
            .in0(_gnd_net_),
            .in1(N__15347),
            .in2(N__15519),
            .in3(N__15369),
            .lcout(\eeprom.n2609 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i5_4_lut_adj_81_LC_5_20_3 .C_ON=1'b0;
    defparam \eeprom.i5_4_lut_adj_81_LC_5_20_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.i5_4_lut_adj_81_LC_5_20_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \eeprom.i5_4_lut_adj_81_LC_5_20_3  (
            .in0(N__15327),
            .in1(N__15223),
            .in2(N__15276),
            .in3(N__15899),
            .lcout(),
            .ltout(\eeprom.n13_adj_474_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i7_4_lut_adj_82_LC_5_20_4 .C_ON=1'b0;
    defparam \eeprom.i7_4_lut_adj_82_LC_5_20_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.i7_4_lut_adj_82_LC_5_20_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \eeprom.i7_4_lut_adj_82_LC_5_20_4  (
            .in0(N__15653),
            .in1(N__16050),
            .in2(N__13601),
            .in3(N__13598),
            .lcout(\eeprom.n2539 ),
            .ltout(\eeprom.n2539_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1697_3_lut_LC_5_20_5 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1697_3_lut_LC_5_20_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1697_3_lut_LC_5_20_5 .LUT_INIT=16'b1111110000001100;
    LogicCell40 \eeprom.rem_4_i1697_3_lut_LC_5_20_5  (
            .in0(_gnd_net_),
            .in1(N__14968),
            .in2(N__13592),
            .in3(N__15398),
            .lcout(\eeprom.n2613 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i15_1_lut_LC_5_20_6 .C_ON=1'b0;
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i15_1_lut_LC_5_20_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i15_1_lut_LC_5_20_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \eeprom.rem_4_unary_minus_2_inv_0_i15_1_lut_LC_5_20_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13585),
            .lcout(\eeprom.n19_adj_429 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_mux_3_i4_3_lut_LC_5_21_0 .C_ON=1'b0;
    defparam \eeprom.rem_4_mux_3_i4_3_lut_LC_5_21_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_mux_3_i4_3_lut_LC_5_21_0 .LUT_INIT=16'b0010011100100111;
    LogicCell40 \eeprom.rem_4_mux_3_i4_3_lut_LC_5_21_0  (
            .in0(N__22983),
            .in1(N__13547),
            .in2(N__23788),
            .in3(_gnd_net_),
            .lcout(\eeprom.n3722_adj_433 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1358_3_lut_LC_5_21_1 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1358_3_lut_LC_5_21_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1358_3_lut_LC_5_21_1 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \eeprom.rem_4_i1358_3_lut_LC_5_21_1  (
            .in0(_gnd_net_),
            .in1(N__13636),
            .in2(N__13616),
            .in3(N__13935),
            .lcout(\eeprom.n2114 ),
            .ltout(\eeprom.n2114_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i1_3_lut_LC_5_21_2 .C_ON=1'b0;
    defparam \eeprom.i1_3_lut_LC_5_21_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.i1_3_lut_LC_5_21_2 .LUT_INIT=16'b1100000000000000;
    LogicCell40 \eeprom.i1_3_lut_LC_5_21_2  (
            .in0(_gnd_net_),
            .in1(N__14262),
            .in2(N__13538),
            .in3(N__14295),
            .lcout(\eeprom.n4463 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1356_3_lut_LC_5_21_3 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1356_3_lut_LC_5_21_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1356_3_lut_LC_5_21_3 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \eeprom.rem_4_i1356_3_lut_LC_5_21_3  (
            .in0(_gnd_net_),
            .in1(N__13884),
            .in2(N__13862),
            .in3(N__13936),
            .lcout(\eeprom.n2112 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1626_3_lut_LC_5_21_4 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1626_3_lut_LC_5_21_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1626_3_lut_LC_5_21_4 .LUT_INIT=16'b1111110000001100;
    LogicCell40 \eeprom.rem_4_i1626_3_lut_LC_5_21_4  (
            .in0(_gnd_net_),
            .in1(N__13535),
            .in2(N__15983),
            .in3(N__13517),
            .lcout(\eeprom.n2510 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1361_3_lut_LC_5_21_5 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1361_3_lut_LC_5_21_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1361_3_lut_LC_5_21_5 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \eeprom.rem_4_i1361_3_lut_LC_5_21_5  (
            .in0(_gnd_net_),
            .in1(N__13678),
            .in2(N__13658),
            .in3(N__13931),
            .lcout(\eeprom.n2117 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1360_3_lut_LC_5_21_6 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1360_3_lut_LC_5_21_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1360_3_lut_LC_5_21_6 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \eeprom.rem_4_i1360_3_lut_LC_5_21_6  (
            .in0(_gnd_net_),
            .in1(N__13897),
            .in2(N__13949),
            .in3(N__15858),
            .lcout(\eeprom.n2116 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1634_3_lut_LC_5_21_7 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1634_3_lut_LC_5_21_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1634_3_lut_LC_5_21_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \eeprom.rem_4_i1634_3_lut_LC_5_21_7  (
            .in0(N__13724),
            .in1(N__13694),
            .in2(_gnd_net_),
            .in3(N__15978),
            .lcout(\eeprom.n2518 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1352_2_lut_LC_5_22_0 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1352_2_lut_LC_5_22_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1352_2_lut_LC_5_22_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1352_2_lut_LC_5_22_0  (
            .in0(_gnd_net_),
            .in1(N__14068),
            .in2(_gnd_net_),
            .in3(N__13682),
            .lcout(\eeprom.n2086 ),
            .ltout(),
            .carryin(bfn_5_22_0_),
            .carryout(\eeprom.n3524 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1352_3_lut_LC_5_22_1 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1352_3_lut_LC_5_22_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1352_3_lut_LC_5_22_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1352_3_lut_LC_5_22_1  (
            .in0(_gnd_net_),
            .in1(N__27181),
            .in2(N__13679),
            .in3(N__13649),
            .lcout(\eeprom.n2085 ),
            .ltout(),
            .carryin(\eeprom.n3524 ),
            .carryout(\eeprom.n3525 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1352_4_lut_LC_5_22_2 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1352_4_lut_LC_5_22_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1352_4_lut_LC_5_22_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1352_4_lut_LC_5_22_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__15868),
            .in3(N__13646),
            .lcout(\eeprom.n2084 ),
            .ltout(),
            .carryin(\eeprom.n3525 ),
            .carryout(\eeprom.n3526 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1352_5_lut_LC_5_22_3 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1352_5_lut_LC_5_22_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1352_5_lut_LC_5_22_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1352_5_lut_LC_5_22_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__13756),
            .in3(N__13643),
            .lcout(\eeprom.n2083 ),
            .ltout(),
            .carryin(\eeprom.n3526 ),
            .carryout(\eeprom.n3527 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1352_6_lut_LC_5_22_4 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1352_6_lut_LC_5_22_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1352_6_lut_LC_5_22_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1352_6_lut_LC_5_22_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__13640),
            .in3(N__13607),
            .lcout(\eeprom.n2082 ),
            .ltout(),
            .carryin(\eeprom.n3527 ),
            .carryout(\eeprom.n3528 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1352_7_lut_LC_5_22_5 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1352_7_lut_LC_5_22_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1352_7_lut_LC_5_22_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1352_7_lut_LC_5_22_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__13813),
            .in3(N__13604),
            .lcout(\eeprom.n2081 ),
            .ltout(),
            .carryin(\eeprom.n3528 ),
            .carryout(\eeprom.n3529 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1352_8_lut_LC_5_22_6 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1352_8_lut_LC_5_22_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1352_8_lut_LC_5_22_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1352_8_lut_LC_5_22_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__13886),
            .in3(N__13853),
            .lcout(\eeprom.n2080 ),
            .ltout(),
            .carryin(\eeprom.n3529 ),
            .carryout(\eeprom.n3530 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1352_9_lut_LC_5_22_7 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1352_9_lut_LC_5_22_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1352_9_lut_LC_5_22_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1352_9_lut_LC_5_22_7  (
            .in0(_gnd_net_),
            .in1(N__13791),
            .in2(N__27729),
            .in3(N__13850),
            .lcout(\eeprom.n2079 ),
            .ltout(),
            .carryin(\eeprom.n3530 ),
            .carryout(\eeprom.n3531 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1352_10_lut_LC_5_23_0 .C_ON=1'b0;
    defparam \eeprom.rem_4_add_1352_10_lut_LC_5_23_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1352_10_lut_LC_5_23_0 .LUT_INIT=16'b1001000001100000;
    LogicCell40 \eeprom.rem_4_add_1352_10_lut_LC_5_23_0  (
            .in0(N__27629),
            .in1(N__13847),
            .in2(N__13950),
            .in3(N__13826),
            .lcout(\eeprom.n2110 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1357_3_lut_LC_5_23_1 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1357_3_lut_LC_5_23_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1357_3_lut_LC_5_23_1 .LUT_INIT=16'b1010101011110000;
    LogicCell40 \eeprom.rem_4_i1357_3_lut_LC_5_23_1  (
            .in0(N__13823),
            .in1(_gnd_net_),
            .in2(N__13817),
            .in3(N__13937),
            .lcout(\eeprom.n2113 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1355_3_lut_LC_5_23_2 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1355_3_lut_LC_5_23_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1355_3_lut_LC_5_23_2 .LUT_INIT=16'b1100101011001010;
    LogicCell40 \eeprom.rem_4_i1355_3_lut_LC_5_23_2  (
            .in0(N__13796),
            .in1(N__13772),
            .in2(N__13951),
            .in3(_gnd_net_),
            .lcout(\eeprom.n2111 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i1_2_lut_LC_5_23_4 .C_ON=1'b0;
    defparam \eeprom.i1_2_lut_LC_5_23_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.i1_2_lut_LC_5_23_4 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \eeprom.i1_2_lut_LC_5_23_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__14556),
            .in3(N__16386),
            .lcout(\eeprom.n4461 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1359_3_lut_LC_5_23_5 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1359_3_lut_LC_5_23_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1359_3_lut_LC_5_23_5 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \eeprom.rem_4_i1359_3_lut_LC_5_23_5  (
            .in0(_gnd_net_),
            .in1(N__13766),
            .in2(N__13760),
            .in3(N__13938),
            .lcout(\eeprom.n2115 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i1_2_lut_adj_72_LC_5_23_6 .C_ON=1'b0;
    defparam \eeprom.i1_2_lut_adj_72_LC_5_23_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.i1_2_lut_adj_72_LC_5_23_6 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \eeprom.i1_2_lut_adj_72_LC_5_23_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__14035),
            .in3(N__16522),
            .lcout(\eeprom.n7_adj_470 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1362_3_lut_LC_5_23_7 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1362_3_lut_LC_5_23_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1362_3_lut_LC_5_23_7 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \eeprom.rem_4_i1362_3_lut_LC_5_23_7  (
            .in0(N__14072),
            .in1(_gnd_net_),
            .in2(N__14045),
            .in3(N__13939),
            .lcout(\eeprom.n2118 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1489_3_lut_LC_5_24_0 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1489_3_lut_LC_5_24_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1489_3_lut_LC_5_24_0 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \eeprom.rem_4_i1489_3_lut_LC_5_24_0  (
            .in0(_gnd_net_),
            .in1(N__16616),
            .in2(N__16636),
            .in3(N__16601),
            .lcout(\eeprom.n2309 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i1_4_lut_adj_50_LC_5_24_2 .C_ON=1'b0;
    defparam \eeprom.i1_4_lut_adj_50_LC_5_24_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.i1_4_lut_adj_50_LC_5_24_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \eeprom.i1_4_lut_adj_50_LC_5_24_2  (
            .in0(N__15780),
            .in1(N__15717),
            .in2(N__15819),
            .in3(N__14207),
            .lcout(),
            .ltout(\eeprom.n4509_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i2_4_lut_LC_5_24_3 .C_ON=1'b0;
    defparam \eeprom.i2_4_lut_LC_5_24_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.i2_4_lut_LC_5_24_3 .LUT_INIT=16'b1111111111100000;
    LogicCell40 \eeprom.i2_4_lut_LC_5_24_3  (
            .in0(N__14011),
            .in1(N__15579),
            .in2(N__13988),
            .in3(N__13974),
            .lcout(\eeprom.n8_adj_468 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1490_3_lut_LC_5_24_4 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1490_3_lut_LC_5_24_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1490_3_lut_LC_5_24_4 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \eeprom.rem_4_i1490_3_lut_LC_5_24_4  (
            .in0(_gnd_net_),
            .in1(N__16602),
            .in2(N__16655),
            .in3(N__16675),
            .lcout(\eeprom.n2310 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i1_2_lut_adj_25_LC_5_24_5 .C_ON=1'b0;
    defparam \eeprom.i1_2_lut_adj_25_LC_5_24_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.i1_2_lut_adj_25_LC_5_24_5 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \eeprom.i1_2_lut_adj_25_LC_5_24_5  (
            .in0(_gnd_net_),
            .in1(N__16629),
            .in2(_gnd_net_),
            .in3(N__16547),
            .lcout(),
            .ltout(\eeprom.n6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i4_4_lut_LC_5_24_6 .C_ON=1'b0;
    defparam \eeprom.i4_4_lut_LC_5_24_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.i4_4_lut_LC_5_24_6 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \eeprom.i4_4_lut_LC_5_24_6  (
            .in0(N__16708),
            .in1(N__16674),
            .in2(N__13958),
            .in3(N__15698),
            .lcout(\eeprom.n2242 ),
            .ltout(\eeprom.n2242_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i4028_3_lut_LC_5_24_7 .C_ON=1'b0;
    defparam \eeprom.i4028_3_lut_LC_5_24_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.i4028_3_lut_LC_5_24_7 .LUT_INIT=16'b1111111111111100;
    LogicCell40 \eeprom.i4028_3_lut_LC_5_24_7  (
            .in0(_gnd_net_),
            .in1(N__16369),
            .in2(N__13955),
            .in3(N__13952),
            .lcout(\eeprom.n4872 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1360_rep_36_3_lut_LC_5_25_0 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1360_rep_36_3_lut_LC_5_25_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1360_rep_36_3_lut_LC_5_25_0 .LUT_INIT=16'b1111110000001100;
    LogicCell40 \eeprom.rem_4_i1360_rep_36_3_lut_LC_5_25_0  (
            .in0(_gnd_net_),
            .in1(N__13901),
            .in2(N__16365),
            .in3(N__14249),
            .lcout(\eeprom.n4801 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1426_3_lut_LC_5_25_1 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1426_3_lut_LC_5_25_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1426_3_lut_LC_5_25_1 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \eeprom.rem_4_i1426_3_lut_LC_5_25_1  (
            .in0(_gnd_net_),
            .in1(N__14531),
            .in2(N__14561),
            .in3(N__16339),
            .lcout(\eeprom.n2214 ),
            .ltout(\eeprom.n2214_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1493_3_lut_LC_5_25_2 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1493_3_lut_LC_5_25_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1493_3_lut_LC_5_25_2 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \eeprom.rem_4_i1493_3_lut_LC_5_25_2  (
            .in0(N__16592),
            .in1(_gnd_net_),
            .in2(N__14231),
            .in3(N__16124),
            .lcout(\eeprom.n2313 ),
            .ltout(\eeprom.n2313_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i1_2_lut_adj_46_LC_5_25_3 .C_ON=1'b0;
    defparam \eeprom.i1_2_lut_adj_46_LC_5_25_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.i1_2_lut_adj_46_LC_5_25_3 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \eeprom.i1_2_lut_adj_46_LC_5_25_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__14210),
            .in3(N__14145),
            .lcout(\eeprom.n4505 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_mux_3_i23_3_lut_LC_5_25_4 .C_ON=1'b0;
    defparam \eeprom.rem_4_mux_3_i23_3_lut_LC_5_25_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_mux_3_i23_3_lut_LC_5_25_4 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \eeprom.rem_4_mux_3_i23_3_lut_LC_5_25_4  (
            .in0(N__14201),
            .in1(N__22978),
            .in2(_gnd_net_),
            .in3(N__14189),
            .lcout(\eeprom.n2119 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1495_3_lut_LC_5_25_5 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1495_3_lut_LC_5_25_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1495_3_lut_LC_5_25_5 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \eeprom.rem_4_i1495_3_lut_LC_5_25_5  (
            .in0(_gnd_net_),
            .in1(N__16203),
            .in2(N__16181),
            .in3(N__16591),
            .lcout(\eeprom.n2315 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1422_3_lut_LC_5_25_6 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1422_3_lut_LC_5_25_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1422_3_lut_LC_5_25_6 .LUT_INIT=16'b1010110010101100;
    LogicCell40 \eeprom.rem_4_i1422_3_lut_LC_5_25_6  (
            .in0(N__14414),
            .in1(N__14440),
            .in2(N__16364),
            .in3(_gnd_net_),
            .lcout(\eeprom.n2210 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1491_3_lut_LC_5_25_7 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1491_3_lut_LC_5_25_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1491_3_lut_LC_5_25_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \eeprom.rem_4_i1491_3_lut_LC_5_25_7  (
            .in0(N__16685),
            .in1(N__16707),
            .in2(_gnd_net_),
            .in3(N__16593),
            .lcout(\eeprom.n2311 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i1_4_lut_LC_5_26_0 .C_ON=1'b0;
    defparam \eeprom.i1_4_lut_LC_5_26_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.i1_4_lut_LC_5_26_0 .LUT_INIT=16'b1110000000000000;
    LogicCell40 \eeprom.i1_4_lut_LC_5_26_0  (
            .in0(N__14343),
            .in1(N__15750),
            .in2(N__14096),
            .in3(N__14084),
            .lcout(),
            .ltout(\eeprom.n4225_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i3_4_lut_LC_5_26_1 .C_ON=1'b0;
    defparam \eeprom.i3_4_lut_LC_5_26_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.i3_4_lut_LC_5_26_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \eeprom.i3_4_lut_LC_5_26_1  (
            .in0(N__14436),
            .in1(N__14478),
            .in2(N__14075),
            .in3(N__14398),
            .lcout(\eeprom.n2143 ),
            .ltout(\eeprom.n2143_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i4033_3_lut_LC_5_26_2 .C_ON=1'b0;
    defparam \eeprom.i4033_3_lut_LC_5_26_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.i4033_3_lut_LC_5_26_2 .LUT_INIT=16'b1111101000001010;
    LogicCell40 \eeprom.i4033_3_lut_LC_5_26_2  (
            .in0(N__14272),
            .in1(_gnd_net_),
            .in2(N__14351),
            .in3(N__14245),
            .lcout(\eeprom.n2215 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1425_3_lut_LC_5_26_3 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1425_3_lut_LC_5_26_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1425_3_lut_LC_5_26_3 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \eeprom.rem_4_i1425_3_lut_LC_5_26_3  (
            .in0(N__14492),
            .in1(_gnd_net_),
            .in2(N__16367),
            .in3(N__14519),
            .lcout(\eeprom.n2213 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1428_3_lut_LC_5_26_4 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1428_3_lut_LC_5_26_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1428_3_lut_LC_5_26_4 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \eeprom.rem_4_i1428_3_lut_LC_5_26_4  (
            .in0(_gnd_net_),
            .in1(N__14282),
            .in2(N__14315),
            .in3(N__16346),
            .lcout(\eeprom.n2216 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1423_3_lut_LC_5_26_5 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1423_3_lut_LC_5_26_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1423_3_lut_LC_5_26_5 .LUT_INIT=16'b1110010011100100;
    LogicCell40 \eeprom.rem_4_i1423_3_lut_LC_5_26_5  (
            .in0(N__16353),
            .in1(N__14479),
            .in2(N__14456),
            .in3(_gnd_net_),
            .lcout(\eeprom.n2211 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1429_rep_30_3_lut_LC_5_26_7 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1429_rep_30_3_lut_LC_5_26_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1429_rep_30_3_lut_LC_5_26_7 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \eeprom.rem_4_i1429_rep_30_3_lut_LC_5_26_7  (
            .in0(_gnd_net_),
            .in1(N__14324),
            .in2(N__16366),
            .in3(N__14344),
            .lcout(\eeprom.n2217 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1419_2_lut_LC_5_27_0 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1419_2_lut_LC_5_27_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1419_2_lut_LC_5_27_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1419_2_lut_LC_5_27_0  (
            .in0(_gnd_net_),
            .in1(N__15752),
            .in2(_gnd_net_),
            .in3(N__14348),
            .lcout(\eeprom.n2186 ),
            .ltout(),
            .carryin(bfn_5_27_0_),
            .carryout(\eeprom.n3532 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1419_3_lut_LC_5_27_1 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1419_3_lut_LC_5_27_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1419_3_lut_LC_5_27_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1419_3_lut_LC_5_27_1  (
            .in0(_gnd_net_),
            .in1(N__27627),
            .in2(N__14345),
            .in3(N__14318),
            .lcout(\eeprom.n2185 ),
            .ltout(),
            .carryin(\eeprom.n3532 ),
            .carryout(\eeprom.n3533 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1419_4_lut_LC_5_27_2 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1419_4_lut_LC_5_27_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1419_4_lut_LC_5_27_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1419_4_lut_LC_5_27_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__14314),
            .in3(N__14276),
            .lcout(\eeprom.n2184 ),
            .ltout(),
            .carryin(\eeprom.n3533 ),
            .carryout(\eeprom.n3534 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1419_5_lut_LC_5_27_3 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1419_5_lut_LC_5_27_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1419_5_lut_LC_5_27_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1419_5_lut_LC_5_27_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__14273),
            .in3(N__14234),
            .lcout(\eeprom.n2183 ),
            .ltout(),
            .carryin(\eeprom.n3534 ),
            .carryout(\eeprom.n3535 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1419_6_lut_LC_5_27_4 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1419_6_lut_LC_5_27_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1419_6_lut_LC_5_27_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1419_6_lut_LC_5_27_4  (
            .in0(_gnd_net_),
            .in1(N__14557),
            .in2(_gnd_net_),
            .in3(N__14522),
            .lcout(\eeprom.n2182 ),
            .ltout(),
            .carryin(\eeprom.n3535 ),
            .carryout(\eeprom.n3536 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1419_7_lut_LC_5_27_5 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1419_7_lut_LC_5_27_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1419_7_lut_LC_5_27_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1419_7_lut_LC_5_27_5  (
            .in0(_gnd_net_),
            .in1(N__14515),
            .in2(_gnd_net_),
            .in3(N__14486),
            .lcout(\eeprom.n2181 ),
            .ltout(),
            .carryin(\eeprom.n3536 ),
            .carryout(\eeprom.n3537 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1419_8_lut_LC_5_27_6 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1419_8_lut_LC_5_27_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1419_8_lut_LC_5_27_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1419_8_lut_LC_5_27_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__16397),
            .in3(N__14483),
            .lcout(\eeprom.n2180 ),
            .ltout(),
            .carryin(\eeprom.n3537 ),
            .carryout(\eeprom.n3538 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1419_9_lut_LC_5_27_7 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1419_9_lut_LC_5_27_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1419_9_lut_LC_5_27_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1419_9_lut_LC_5_27_7  (
            .in0(_gnd_net_),
            .in1(N__27628),
            .in2(N__14480),
            .in3(N__14447),
            .lcout(\eeprom.n2179 ),
            .ltout(),
            .carryin(\eeprom.n3538 ),
            .carryout(\eeprom.n3539 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1419_10_lut_LC_5_28_0 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1419_10_lut_LC_5_28_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1419_10_lut_LC_5_28_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1419_10_lut_LC_5_28_0  (
            .in0(_gnd_net_),
            .in1(N__27612),
            .in2(N__14444),
            .in3(N__14405),
            .lcout(\eeprom.n2178 ),
            .ltout(),
            .carryin(bfn_5_28_0_),
            .carryout(\eeprom.n3540 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1419_11_lut_LC_5_28_1 .C_ON=1'b0;
    defparam \eeprom.rem_4_add_1419_11_lut_LC_5_28_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1419_11_lut_LC_5_28_1 .LUT_INIT=16'b1001000001100000;
    LogicCell40 \eeprom.rem_4_add_1419_11_lut_LC_5_28_1  (
            .in0(N__27613),
            .in1(N__14402),
            .in2(N__16370),
            .in3(N__14381),
            .lcout(\eeprom.n2209 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_287__i0_LC_5_29_0.C_ON=1'b1;
    defparam blink_counter_287__i0_LC_5_29_0.SEQ_MODE=4'b1000;
    defparam blink_counter_287__i0_LC_5_29_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_287__i0_LC_5_29_0 (
            .in0(_gnd_net_),
            .in1(N__14378),
            .in2(_gnd_net_),
            .in3(N__14372),
            .lcout(n26),
            .ltout(),
            .carryin(bfn_5_29_0_),
            .carryout(n3485),
            .clk(N__24346),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_287__i1_LC_5_29_1.C_ON=1'b1;
    defparam blink_counter_287__i1_LC_5_29_1.SEQ_MODE=4'b1000;
    defparam blink_counter_287__i1_LC_5_29_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_287__i1_LC_5_29_1 (
            .in0(_gnd_net_),
            .in1(N__14369),
            .in2(_gnd_net_),
            .in3(N__14363),
            .lcout(n25),
            .ltout(),
            .carryin(n3485),
            .carryout(n3486),
            .clk(N__24346),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_287__i2_LC_5_29_2.C_ON=1'b1;
    defparam blink_counter_287__i2_LC_5_29_2.SEQ_MODE=4'b1000;
    defparam blink_counter_287__i2_LC_5_29_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_287__i2_LC_5_29_2 (
            .in0(_gnd_net_),
            .in1(N__14360),
            .in2(_gnd_net_),
            .in3(N__14354),
            .lcout(n24),
            .ltout(),
            .carryin(n3486),
            .carryout(n3487),
            .clk(N__24346),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_287__i3_LC_5_29_3.C_ON=1'b1;
    defparam blink_counter_287__i3_LC_5_29_3.SEQ_MODE=4'b1000;
    defparam blink_counter_287__i3_LC_5_29_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_287__i3_LC_5_29_3 (
            .in0(_gnd_net_),
            .in1(N__14633),
            .in2(_gnd_net_),
            .in3(N__14627),
            .lcout(n23),
            .ltout(),
            .carryin(n3487),
            .carryout(n3488),
            .clk(N__24346),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_287__i4_LC_5_29_4.C_ON=1'b1;
    defparam blink_counter_287__i4_LC_5_29_4.SEQ_MODE=4'b1000;
    defparam blink_counter_287__i4_LC_5_29_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_287__i4_LC_5_29_4 (
            .in0(_gnd_net_),
            .in1(N__14624),
            .in2(_gnd_net_),
            .in3(N__14618),
            .lcout(n22),
            .ltout(),
            .carryin(n3488),
            .carryout(n3489),
            .clk(N__24346),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_287__i5_LC_5_29_5.C_ON=1'b1;
    defparam blink_counter_287__i5_LC_5_29_5.SEQ_MODE=4'b1000;
    defparam blink_counter_287__i5_LC_5_29_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_287__i5_LC_5_29_5 (
            .in0(_gnd_net_),
            .in1(N__14615),
            .in2(_gnd_net_),
            .in3(N__14609),
            .lcout(n21),
            .ltout(),
            .carryin(n3489),
            .carryout(n3490),
            .clk(N__24346),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_287__i6_LC_5_29_6.C_ON=1'b1;
    defparam blink_counter_287__i6_LC_5_29_6.SEQ_MODE=4'b1000;
    defparam blink_counter_287__i6_LC_5_29_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_287__i6_LC_5_29_6 (
            .in0(_gnd_net_),
            .in1(N__14606),
            .in2(_gnd_net_),
            .in3(N__14600),
            .lcout(n20),
            .ltout(),
            .carryin(n3490),
            .carryout(n3491),
            .clk(N__24346),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_287__i7_LC_5_29_7.C_ON=1'b1;
    defparam blink_counter_287__i7_LC_5_29_7.SEQ_MODE=4'b1000;
    defparam blink_counter_287__i7_LC_5_29_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_287__i7_LC_5_29_7 (
            .in0(_gnd_net_),
            .in1(N__14597),
            .in2(_gnd_net_),
            .in3(N__14591),
            .lcout(n19),
            .ltout(),
            .carryin(n3491),
            .carryout(n3492),
            .clk(N__24346),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_287__i8_LC_5_30_0.C_ON=1'b1;
    defparam blink_counter_287__i8_LC_5_30_0.SEQ_MODE=4'b1000;
    defparam blink_counter_287__i8_LC_5_30_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_287__i8_LC_5_30_0 (
            .in0(_gnd_net_),
            .in1(N__14588),
            .in2(_gnd_net_),
            .in3(N__14582),
            .lcout(n18),
            .ltout(),
            .carryin(bfn_5_30_0_),
            .carryout(n3493),
            .clk(N__24347),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_287__i9_LC_5_30_1.C_ON=1'b1;
    defparam blink_counter_287__i9_LC_5_30_1.SEQ_MODE=4'b1000;
    defparam blink_counter_287__i9_LC_5_30_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_287__i9_LC_5_30_1 (
            .in0(_gnd_net_),
            .in1(N__14579),
            .in2(_gnd_net_),
            .in3(N__14573),
            .lcout(n17),
            .ltout(),
            .carryin(n3493),
            .carryout(n3494),
            .clk(N__24347),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_287__i10_LC_5_30_2.C_ON=1'b1;
    defparam blink_counter_287__i10_LC_5_30_2.SEQ_MODE=4'b1000;
    defparam blink_counter_287__i10_LC_5_30_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_287__i10_LC_5_30_2 (
            .in0(_gnd_net_),
            .in1(N__14570),
            .in2(_gnd_net_),
            .in3(N__14564),
            .lcout(n16),
            .ltout(),
            .carryin(n3494),
            .carryout(n3495),
            .clk(N__24347),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_287__i11_LC_5_30_3.C_ON=1'b1;
    defparam blink_counter_287__i11_LC_5_30_3.SEQ_MODE=4'b1000;
    defparam blink_counter_287__i11_LC_5_30_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_287__i11_LC_5_30_3 (
            .in0(_gnd_net_),
            .in1(N__14705),
            .in2(_gnd_net_),
            .in3(N__14699),
            .lcout(n15),
            .ltout(),
            .carryin(n3495),
            .carryout(n3496),
            .clk(N__24347),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_287__i12_LC_5_30_4.C_ON=1'b1;
    defparam blink_counter_287__i12_LC_5_30_4.SEQ_MODE=4'b1000;
    defparam blink_counter_287__i12_LC_5_30_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_287__i12_LC_5_30_4 (
            .in0(_gnd_net_),
            .in1(N__14696),
            .in2(_gnd_net_),
            .in3(N__14690),
            .lcout(n14),
            .ltout(),
            .carryin(n3496),
            .carryout(n3497),
            .clk(N__24347),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_287__i13_LC_5_30_5.C_ON=1'b1;
    defparam blink_counter_287__i13_LC_5_30_5.SEQ_MODE=4'b1000;
    defparam blink_counter_287__i13_LC_5_30_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_287__i13_LC_5_30_5 (
            .in0(_gnd_net_),
            .in1(N__14687),
            .in2(_gnd_net_),
            .in3(N__14681),
            .lcout(n13),
            .ltout(),
            .carryin(n3497),
            .carryout(n3498),
            .clk(N__24347),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_287__i14_LC_5_30_6.C_ON=1'b1;
    defparam blink_counter_287__i14_LC_5_30_6.SEQ_MODE=4'b1000;
    defparam blink_counter_287__i14_LC_5_30_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_287__i14_LC_5_30_6 (
            .in0(_gnd_net_),
            .in1(N__14678),
            .in2(_gnd_net_),
            .in3(N__14672),
            .lcout(n12),
            .ltout(),
            .carryin(n3498),
            .carryout(n3499),
            .clk(N__24347),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_287__i15_LC_5_30_7.C_ON=1'b1;
    defparam blink_counter_287__i15_LC_5_30_7.SEQ_MODE=4'b1000;
    defparam blink_counter_287__i15_LC_5_30_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_287__i15_LC_5_30_7 (
            .in0(_gnd_net_),
            .in1(N__14669),
            .in2(_gnd_net_),
            .in3(N__14663),
            .lcout(n11),
            .ltout(),
            .carryin(n3499),
            .carryout(n3500),
            .clk(N__24347),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_287__i16_LC_5_31_0.C_ON=1'b1;
    defparam blink_counter_287__i16_LC_5_31_0.SEQ_MODE=4'b1000;
    defparam blink_counter_287__i16_LC_5_31_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_287__i16_LC_5_31_0 (
            .in0(_gnd_net_),
            .in1(N__14660),
            .in2(_gnd_net_),
            .in3(N__14654),
            .lcout(n10),
            .ltout(),
            .carryin(bfn_5_31_0_),
            .carryout(n3501),
            .clk(N__24348),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_287__i17_LC_5_31_1.C_ON=1'b1;
    defparam blink_counter_287__i17_LC_5_31_1.SEQ_MODE=4'b1000;
    defparam blink_counter_287__i17_LC_5_31_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_287__i17_LC_5_31_1 (
            .in0(_gnd_net_),
            .in1(N__14651),
            .in2(_gnd_net_),
            .in3(N__14645),
            .lcout(n9),
            .ltout(),
            .carryin(n3501),
            .carryout(n3502),
            .clk(N__24348),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_287__i18_LC_5_31_2.C_ON=1'b1;
    defparam blink_counter_287__i18_LC_5_31_2.SEQ_MODE=4'b1000;
    defparam blink_counter_287__i18_LC_5_31_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_287__i18_LC_5_31_2 (
            .in0(_gnd_net_),
            .in1(N__14642),
            .in2(_gnd_net_),
            .in3(N__14636),
            .lcout(n8),
            .ltout(),
            .carryin(n3502),
            .carryout(n3503),
            .clk(N__24348),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_287__i19_LC_5_31_3.C_ON=1'b1;
    defparam blink_counter_287__i19_LC_5_31_3.SEQ_MODE=4'b1000;
    defparam blink_counter_287__i19_LC_5_31_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_287__i19_LC_5_31_3 (
            .in0(_gnd_net_),
            .in1(N__14822),
            .in2(_gnd_net_),
            .in3(N__14816),
            .lcout(n7),
            .ltout(),
            .carryin(n3503),
            .carryout(n3504),
            .clk(N__24348),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_287__i20_LC_5_31_4.C_ON=1'b1;
    defparam blink_counter_287__i20_LC_5_31_4.SEQ_MODE=4'b1000;
    defparam blink_counter_287__i20_LC_5_31_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_287__i20_LC_5_31_4 (
            .in0(_gnd_net_),
            .in1(N__14813),
            .in2(_gnd_net_),
            .in3(N__14807),
            .lcout(n6),
            .ltout(),
            .carryin(n3504),
            .carryout(n3505),
            .clk(N__24348),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_287__i21_LC_5_31_5.C_ON=1'b1;
    defparam blink_counter_287__i21_LC_5_31_5.SEQ_MODE=4'b1000;
    defparam blink_counter_287__i21_LC_5_31_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_287__i21_LC_5_31_5 (
            .in0(_gnd_net_),
            .in1(N__14799),
            .in2(_gnd_net_),
            .in3(N__14786),
            .lcout(blink_counter_21),
            .ltout(),
            .carryin(n3505),
            .carryout(n3506),
            .clk(N__24348),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_287__i22_LC_5_31_6.C_ON=1'b1;
    defparam blink_counter_287__i22_LC_5_31_6.SEQ_MODE=4'b1000;
    defparam blink_counter_287__i22_LC_5_31_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_287__i22_LC_5_31_6 (
            .in0(_gnd_net_),
            .in1(N__14781),
            .in2(_gnd_net_),
            .in3(N__14768),
            .lcout(blink_counter_22),
            .ltout(),
            .carryin(n3506),
            .carryout(n3507),
            .clk(N__24348),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_287__i23_LC_5_31_7.C_ON=1'b1;
    defparam blink_counter_287__i23_LC_5_31_7.SEQ_MODE=4'b1000;
    defparam blink_counter_287__i23_LC_5_31_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_287__i23_LC_5_31_7 (
            .in0(_gnd_net_),
            .in1(N__14760),
            .in2(_gnd_net_),
            .in3(N__14747),
            .lcout(blink_counter_23),
            .ltout(),
            .carryin(n3507),
            .carryout(n3508),
            .clk(N__24348),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_287__i24_LC_5_32_0.C_ON=1'b1;
    defparam blink_counter_287__i24_LC_5_32_0.SEQ_MODE=4'b1000;
    defparam blink_counter_287__i24_LC_5_32_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_287__i24_LC_5_32_0 (
            .in0(_gnd_net_),
            .in1(N__14742),
            .in2(_gnd_net_),
            .in3(N__14729),
            .lcout(blink_counter_24),
            .ltout(),
            .carryin(bfn_5_32_0_),
            .carryout(n3509),
            .clk(N__24350),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_287__i25_LC_5_32_1.C_ON=1'b0;
    defparam blink_counter_287__i25_LC_5_32_1.SEQ_MODE=4'b1000;
    defparam blink_counter_287__i25_LC_5_32_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_287__i25_LC_5_32_1 (
            .in0(_gnd_net_),
            .in1(N__14722),
            .in2(_gnd_net_),
            .in3(N__14726),
            .lcout(blink_counter_25),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24350),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1754_2_lut_LC_6_18_0 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1754_2_lut_LC_6_18_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1754_2_lut_LC_6_18_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1754_2_lut_LC_6_18_0  (
            .in0(_gnd_net_),
            .in1(N__16761),
            .in2(_gnd_net_),
            .in3(N__14711),
            .lcout(\eeprom.n2686 ),
            .ltout(),
            .carryin(bfn_6_18_0_),
            .carryout(\eeprom.n3587 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1754_3_lut_LC_6_18_1 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1754_3_lut_LC_6_18_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1754_3_lut_LC_6_18_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1754_3_lut_LC_6_18_1  (
            .in0(_gnd_net_),
            .in1(N__27779),
            .in2(N__16811),
            .in3(N__14708),
            .lcout(\eeprom.n2685 ),
            .ltout(),
            .carryin(\eeprom.n3587 ),
            .carryout(\eeprom.n3588 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1754_4_lut_LC_6_18_2 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1754_4_lut_LC_6_18_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1754_4_lut_LC_6_18_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1754_4_lut_LC_6_18_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__16891),
            .in3(N__14849),
            .lcout(\eeprom.n2684 ),
            .ltout(),
            .carryin(\eeprom.n3588 ),
            .carryout(\eeprom.n3589 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1754_5_lut_LC_6_18_3 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1754_5_lut_LC_6_18_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1754_5_lut_LC_6_18_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1754_5_lut_LC_6_18_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__16915),
            .in3(N__14846),
            .lcout(\eeprom.n2683 ),
            .ltout(),
            .carryin(\eeprom.n3589 ),
            .carryout(\eeprom.n3590 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1754_6_lut_LC_6_18_4 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1754_6_lut_LC_6_18_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1754_6_lut_LC_6_18_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1754_6_lut_LC_6_18_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__17002),
            .in3(N__14843),
            .lcout(\eeprom.n2682 ),
            .ltout(),
            .carryin(\eeprom.n3590 ),
            .carryout(\eeprom.n3591 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1754_7_lut_LC_6_18_5 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1754_7_lut_LC_6_18_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1754_7_lut_LC_6_18_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1754_7_lut_LC_6_18_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__16855),
            .in3(N__14840),
            .lcout(\eeprom.n2681 ),
            .ltout(),
            .carryin(\eeprom.n3591 ),
            .carryout(\eeprom.n3592 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1754_8_lut_LC_6_18_6 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1754_8_lut_LC_6_18_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1754_8_lut_LC_6_18_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1754_8_lut_LC_6_18_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__16426),
            .in3(N__14837),
            .lcout(\eeprom.n2680 ),
            .ltout(),
            .carryin(\eeprom.n3592 ),
            .carryout(\eeprom.n3593 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1754_9_lut_LC_6_18_7 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1754_9_lut_LC_6_18_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1754_9_lut_LC_6_18_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1754_9_lut_LC_6_18_7  (
            .in0(_gnd_net_),
            .in1(N__27780),
            .in2(N__16498),
            .in3(N__14834),
            .lcout(\eeprom.n2679 ),
            .ltout(),
            .carryin(\eeprom.n3593 ),
            .carryout(\eeprom.n3594 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1754_10_lut_LC_6_19_0 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1754_10_lut_LC_6_19_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1754_10_lut_LC_6_19_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1754_10_lut_LC_6_19_0  (
            .in0(_gnd_net_),
            .in1(N__27756),
            .in2(N__15419),
            .in3(N__14831),
            .lcout(\eeprom.n2678 ),
            .ltout(),
            .carryin(bfn_6_19_0_),
            .carryout(\eeprom.n3595 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1754_11_lut_LC_6_19_1 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1754_11_lut_LC_6_19_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1754_11_lut_LC_6_19_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1754_11_lut_LC_6_19_1  (
            .in0(_gnd_net_),
            .in1(N__17254),
            .in2(N__27786),
            .in3(N__14828),
            .lcout(\eeprom.n2677 ),
            .ltout(),
            .carryin(\eeprom.n3595 ),
            .carryout(\eeprom.n3596 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1754_12_lut_LC_6_19_2 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1754_12_lut_LC_6_19_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1754_12_lut_LC_6_19_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1754_12_lut_LC_6_19_2  (
            .in0(_gnd_net_),
            .in1(N__27760),
            .in2(N__14879),
            .in3(N__14825),
            .lcout(\eeprom.n2676 ),
            .ltout(),
            .carryin(\eeprom.n3596 ),
            .carryout(\eeprom.n3597 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1754_13_lut_LC_6_19_3 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1754_13_lut_LC_6_19_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1754_13_lut_LC_6_19_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1754_13_lut_LC_6_19_3  (
            .in0(_gnd_net_),
            .in1(N__27748),
            .in2(N__16985),
            .in3(N__14942),
            .lcout(\eeprom.n2675 ),
            .ltout(),
            .carryin(\eeprom.n3597 ),
            .carryout(\eeprom.n3598 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1754_14_lut_LC_6_19_4 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1754_14_lut_LC_6_19_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1754_14_lut_LC_6_19_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1754_14_lut_LC_6_19_4  (
            .in0(_gnd_net_),
            .in1(N__27761),
            .in2(N__16958),
            .in3(N__14939),
            .lcout(\eeprom.n2674 ),
            .ltout(),
            .carryin(\eeprom.n3598 ),
            .carryout(\eeprom.n3599 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1754_15_lut_LC_6_19_5 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1754_15_lut_LC_6_19_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1754_15_lut_LC_6_19_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1754_15_lut_LC_6_19_5  (
            .in0(_gnd_net_),
            .in1(N__16456),
            .in2(N__27787),
            .in3(N__14936),
            .lcout(\eeprom.n2673 ),
            .ltout(),
            .carryin(\eeprom.n3599 ),
            .carryout(\eeprom.n3600 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1754_16_lut_LC_6_19_6 .C_ON=1'b0;
    defparam \eeprom.rem_4_add_1754_16_lut_LC_6_19_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1754_16_lut_LC_6_19_6 .LUT_INIT=16'b1000010001001000;
    LogicCell40 \eeprom.rem_4_add_1754_16_lut_LC_6_19_6  (
            .in0(N__27749),
            .in1(N__17213),
            .in2(N__15437),
            .in3(N__14933),
            .lcout(\eeprom.n2704 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1702_3_lut_LC_6_19_7 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1702_3_lut_LC_6_19_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1702_3_lut_LC_6_19_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \eeprom.rem_4_i1702_3_lut_LC_6_19_7  (
            .in0(N__15164),
            .in1(N__15191),
            .in2(_gnd_net_),
            .in3(N__15499),
            .lcout(\eeprom.n2618 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_mux_3_i13_3_lut_LC_6_20_0 .C_ON=1'b0;
    defparam \eeprom.rem_4_mux_3_i13_3_lut_LC_6_20_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_mux_3_i13_3_lut_LC_6_20_0 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \eeprom.rem_4_mux_3_i13_3_lut_LC_6_20_0  (
            .in0(N__14930),
            .in1(N__22942),
            .in2(_gnd_net_),
            .in3(N__14918),
            .lcout(\eeprom.n3119 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i5_1_lut_LC_6_20_2 .C_ON=1'b0;
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i5_1_lut_LC_6_20_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i5_1_lut_LC_6_20_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \eeprom.rem_4_unary_minus_2_inv_0_i5_1_lut_LC_6_20_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23710),
            .lcout(\eeprom.n29_adj_460 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1760_3_lut_LC_6_20_3 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1760_3_lut_LC_6_20_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1760_3_lut_LC_6_20_3 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \eeprom.rem_4_i1760_3_lut_LC_6_20_3  (
            .in0(_gnd_net_),
            .in1(N__14878),
            .in2(N__14858),
            .in3(N__17212),
            .lcout(\eeprom.n2708 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1695_3_lut_LC_6_20_4 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1695_3_lut_LC_6_20_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1695_3_lut_LC_6_20_4 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \eeprom.rem_4_i1695_3_lut_LC_6_20_4  (
            .in0(N__16052),
            .in1(_gnd_net_),
            .in2(N__15386),
            .in3(N__15494),
            .lcout(\eeprom.n2611 ),
            .ltout(\eeprom.n2611_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1762_3_lut_LC_6_20_5 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1762_3_lut_LC_6_20_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1762_3_lut_LC_6_20_5 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \eeprom.rem_4_i1762_3_lut_LC_6_20_5  (
            .in0(_gnd_net_),
            .in1(N__15200),
            .in2(N__15194),
            .in3(N__17211),
            .lcout(\eeprom.n2710 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1691_3_lut_LC_6_20_6 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1691_3_lut_LC_6_20_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1691_3_lut_LC_6_20_6 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \eeprom.rem_4_i1691_3_lut_LC_6_20_6  (
            .in0(_gnd_net_),
            .in1(N__15284),
            .in2(N__15242),
            .in3(N__15498),
            .lcout(\eeprom.n2607 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1692_3_lut_LC_6_20_7 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1692_3_lut_LC_6_20_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1692_3_lut_LC_6_20_7 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \eeprom.rem_4_i1692_3_lut_LC_6_20_7  (
            .in0(_gnd_net_),
            .in1(N__15296),
            .in2(N__15517),
            .in3(N__15335),
            .lcout(\eeprom.n2608 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1687_2_lut_LC_6_21_0 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1687_2_lut_LC_6_21_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1687_2_lut_LC_6_21_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1687_2_lut_LC_6_21_0  (
            .in0(_gnd_net_),
            .in1(N__15187),
            .in2(_gnd_net_),
            .in3(N__15155),
            .lcout(\eeprom.n2586 ),
            .ltout(),
            .carryin(bfn_6_21_0_),
            .carryout(\eeprom.n3574 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1687_3_lut_LC_6_21_1 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1687_3_lut_LC_6_21_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1687_3_lut_LC_6_21_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1687_3_lut_LC_6_21_1  (
            .in0(_gnd_net_),
            .in1(N__27754),
            .in2(N__15148),
            .in3(N__15116),
            .lcout(\eeprom.n2585 ),
            .ltout(),
            .carryin(\eeprom.n3574 ),
            .carryout(\eeprom.n3575 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1687_4_lut_LC_6_21_2 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1687_4_lut_LC_6_21_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1687_4_lut_LC_6_21_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1687_4_lut_LC_6_21_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__15113),
            .in3(N__15071),
            .lcout(\eeprom.n2584 ),
            .ltout(),
            .carryin(\eeprom.n3575 ),
            .carryout(\eeprom.n3576 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1687_5_lut_LC_6_21_3 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1687_5_lut_LC_6_21_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1687_5_lut_LC_6_21_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1687_5_lut_LC_6_21_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__15068),
            .in3(N__15023),
            .lcout(\eeprom.n2583 ),
            .ltout(),
            .carryin(\eeprom.n3576 ),
            .carryout(\eeprom.n3577 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1687_6_lut_LC_6_21_4 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1687_6_lut_LC_6_21_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1687_6_lut_LC_6_21_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1687_6_lut_LC_6_21_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__15019),
            .in3(N__14975),
            .lcout(\eeprom.n2582 ),
            .ltout(),
            .carryin(\eeprom.n3577 ),
            .carryout(\eeprom.n3578 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1687_7_lut_LC_6_21_5 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1687_7_lut_LC_6_21_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1687_7_lut_LC_6_21_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1687_7_lut_LC_6_21_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__14972),
            .in3(N__15392),
            .lcout(\eeprom.n2581 ),
            .ltout(),
            .carryin(\eeprom.n3578 ),
            .carryout(\eeprom.n3579 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1687_8_lut_LC_6_21_6 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1687_8_lut_LC_6_21_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1687_8_lut_LC_6_21_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1687_8_lut_LC_6_21_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__15551),
            .in3(N__15389),
            .lcout(\eeprom.n2580 ),
            .ltout(),
            .carryin(\eeprom.n3579 ),
            .carryout(\eeprom.n3580 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1687_9_lut_LC_6_21_7 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1687_9_lut_LC_6_21_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1687_9_lut_LC_6_21_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1687_9_lut_LC_6_21_7  (
            .in0(_gnd_net_),
            .in1(N__27755),
            .in2(N__16051),
            .in3(N__15377),
            .lcout(\eeprom.n2579 ),
            .ltout(),
            .carryin(\eeprom.n3580 ),
            .carryout(\eeprom.n3581 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1687_10_lut_LC_6_22_0 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1687_10_lut_LC_6_22_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1687_10_lut_LC_6_22_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1687_10_lut_LC_6_22_0  (
            .in0(_gnd_net_),
            .in1(N__27179),
            .in2(N__15652),
            .in3(N__15374),
            .lcout(\eeprom.n2578 ),
            .ltout(),
            .carryin(bfn_6_22_0_),
            .carryout(\eeprom.n3582 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1687_11_lut_LC_6_22_1 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1687_11_lut_LC_6_22_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1687_11_lut_LC_6_22_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1687_11_lut_LC_6_22_1  (
            .in0(_gnd_net_),
            .in1(N__27648),
            .in2(N__15371),
            .in3(N__15338),
            .lcout(\eeprom.n2577 ),
            .ltout(),
            .carryin(\eeprom.n3582 ),
            .carryout(\eeprom.n3583 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1687_12_lut_LC_6_22_2 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1687_12_lut_LC_6_22_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1687_12_lut_LC_6_22_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1687_12_lut_LC_6_22_2  (
            .in0(_gnd_net_),
            .in1(N__27180),
            .in2(N__15334),
            .in3(N__15287),
            .lcout(\eeprom.n2576 ),
            .ltout(),
            .carryin(\eeprom.n3583 ),
            .carryout(\eeprom.n3584 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1687_13_lut_LC_6_22_3 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1687_13_lut_LC_6_22_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1687_13_lut_LC_6_22_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1687_13_lut_LC_6_22_3  (
            .in0(_gnd_net_),
            .in1(N__27649),
            .in2(N__15283),
            .in3(N__15230),
            .lcout(\eeprom.n2575 ),
            .ltout(),
            .carryin(\eeprom.n3584 ),
            .carryout(\eeprom.n3585 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1687_14_lut_LC_6_22_4 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1687_14_lut_LC_6_22_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1687_14_lut_LC_6_22_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1687_14_lut_LC_6_22_4  (
            .in0(_gnd_net_),
            .in1(N__15897),
            .in2(N__27753),
            .in3(N__15227),
            .lcout(\eeprom.n2574 ),
            .ltout(),
            .carryin(\eeprom.n3585 ),
            .carryout(\eeprom.n3586 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1687_15_lut_LC_6_22_5 .C_ON=1'b0;
    defparam \eeprom.rem_4_add_1687_15_lut_LC_6_22_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1687_15_lut_LC_6_22_5 .LUT_INIT=16'b1001000001100000;
    LogicCell40 \eeprom.rem_4_add_1687_15_lut_LC_6_22_5  (
            .in0(N__15224),
            .in1(N__27653),
            .in2(N__15520),
            .in3(N__15203),
            .lcout(\eeprom.n2605 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1627_3_lut_LC_6_22_6 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1627_3_lut_LC_6_22_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1627_3_lut_LC_6_22_6 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \eeprom.rem_4_i1627_3_lut_LC_6_22_6  (
            .in0(_gnd_net_),
            .in1(N__15692),
            .in2(N__15668),
            .in3(N__15982),
            .lcout(\eeprom.n2511 ),
            .ltout(\eeprom.n2511_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1694_3_lut_LC_6_22_7 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1694_3_lut_LC_6_22_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1694_3_lut_LC_6_22_7 .LUT_INIT=16'b1101100011011000;
    LogicCell40 \eeprom.rem_4_i1694_3_lut_LC_6_22_7  (
            .in0(N__15512),
            .in1(N__15635),
            .in2(N__15629),
            .in3(_gnd_net_),
            .lcout(\eeprom.n2610 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_mux_3_i22_3_lut_LC_6_23_2 .C_ON=1'b0;
    defparam \eeprom.rem_4_mux_3_i22_3_lut_LC_6_23_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_mux_3_i22_3_lut_LC_6_23_2 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \eeprom.rem_4_mux_3_i22_3_lut_LC_6_23_2  (
            .in0(N__15626),
            .in1(N__22979),
            .in2(_gnd_net_),
            .in3(N__15617),
            .lcout(\eeprom.n2219 ),
            .ltout(\eeprom.n2219_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1498_3_lut_LC_6_23_3 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1498_3_lut_LC_6_23_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1498_3_lut_LC_6_23_3 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \eeprom.rem_4_i1498_3_lut_LC_6_23_3  (
            .in0(_gnd_net_),
            .in1(N__16274),
            .in2(N__15587),
            .in3(N__16600),
            .lcout(\eeprom.n2318 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1696_3_lut_LC_6_23_4 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1696_3_lut_LC_6_23_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1696_3_lut_LC_6_23_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \eeprom.rem_4_i1696_3_lut_LC_6_23_4  (
            .in0(N__15560),
            .in1(N__15547),
            .in2(_gnd_net_),
            .in3(N__15513),
            .lcout(\eeprom.n2612 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1690_3_lut_LC_6_23_5 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1690_3_lut_LC_6_23_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1690_3_lut_LC_6_23_5 .LUT_INIT=16'b1111110000001100;
    LogicCell40 \eeprom.rem_4_i1690_3_lut_LC_6_23_5  (
            .in0(_gnd_net_),
            .in1(N__15898),
            .in2(N__15521),
            .in3(N__15446),
            .lcout(\eeprom.n2606 ),
            .ltout(\eeprom.n2606_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i1_2_lut_adj_85_LC_6_23_6 .C_ON=1'b0;
    defparam \eeprom.i1_2_lut_adj_85_LC_6_23_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.i1_2_lut_adj_85_LC_6_23_6 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \eeprom.i1_2_lut_adj_85_LC_6_23_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__15440),
            .in3(N__15430),
            .lcout(),
            .ltout(\eeprom.n10_adj_475_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i7_4_lut_adj_87_LC_6_23_7 .C_ON=1'b0;
    defparam \eeprom.i7_4_lut_adj_87_LC_6_23_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.i7_4_lut_adj_87_LC_6_23_7 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \eeprom.i7_4_lut_adj_87_LC_6_23_7  (
            .in0(N__17247),
            .in1(N__15418),
            .in2(N__15401),
            .in3(N__16485),
            .lcout(\eeprom.n16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1628_3_lut_LC_6_24_1 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1628_3_lut_LC_6_24_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1628_3_lut_LC_6_24_1 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \eeprom.rem_4_i1628_3_lut_LC_6_24_1  (
            .in0(_gnd_net_),
            .in1(N__16091),
            .in2(N__16067),
            .in3(N__15973),
            .lcout(\eeprom.n2512 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1623_3_lut_LC_6_24_5 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1623_3_lut_LC_6_24_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1623_3_lut_LC_6_24_5 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \eeprom.rem_4_i1623_3_lut_LC_6_24_5  (
            .in0(_gnd_net_),
            .in1(N__16022),
            .in2(N__15998),
            .in3(N__15972),
            .lcout(\eeprom.n2507 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1427_rep_34_3_lut_LC_6_24_6 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1427_rep_34_3_lut_LC_6_24_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1427_rep_34_3_lut_LC_6_24_6 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \eeprom.rem_4_i1427_rep_34_3_lut_LC_6_24_6  (
            .in0(_gnd_net_),
            .in1(N__15875),
            .in2(N__16154),
            .in3(N__16597),
            .lcout(),
            .ltout(\eeprom.n4799_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1494_3_lut_LC_6_24_7 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1494_3_lut_LC_6_24_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1494_3_lut_LC_6_24_7 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \eeprom.rem_4_i1494_3_lut_LC_6_24_7  (
            .in0(N__15869),
            .in1(_gnd_net_),
            .in2(N__15839),
            .in3(N__15836),
            .lcout(\eeprom.n2314 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i4036_3_lut_LC_6_25_1 .C_ON=1'b0;
    defparam \eeprom.i4036_3_lut_LC_6_25_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.i4036_3_lut_LC_6_25_1 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \eeprom.i4036_3_lut_LC_6_25_1  (
            .in0(_gnd_net_),
            .in1(N__16214),
            .in2(N__16238),
            .in3(N__16599),
            .lcout(\eeprom.n2316 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1430_3_lut_LC_6_25_2 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1430_3_lut_LC_6_25_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1430_3_lut_LC_6_25_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \eeprom.rem_4_i1430_3_lut_LC_6_25_2  (
            .in0(N__15761),
            .in1(N__15751),
            .in2(_gnd_net_),
            .in3(N__16354),
            .lcout(\eeprom.n2218 ),
            .ltout(\eeprom.n2218_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1497_3_lut_LC_6_25_3 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1497_3_lut_LC_6_25_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1497_3_lut_LC_6_25_3 .LUT_INIT=16'b1010101011110000;
    LogicCell40 \eeprom.rem_4_i1497_3_lut_LC_6_25_3  (
            .in0(N__16247),
            .in1(_gnd_net_),
            .in2(N__15731),
            .in3(N__16598),
            .lcout(\eeprom.n2317 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i1_4_lut_adj_24_LC_6_25_5 .C_ON=1'b0;
    defparam \eeprom.i1_4_lut_adj_24_LC_6_25_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.i1_4_lut_adj_24_LC_6_25_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \eeprom.i1_4_lut_adj_24_LC_6_25_5  (
            .in0(N__16165),
            .in1(N__16135),
            .in2(N__16204),
            .in3(N__16230),
            .lcout(),
            .ltout(\eeprom.n4447_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i1_4_lut_adj_26_LC_6_25_6 .C_ON=1'b0;
    defparam \eeprom.i1_4_lut_adj_26_LC_6_25_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.i1_4_lut_adj_26_LC_6_25_6 .LUT_INIT=16'b1100000010000000;
    LogicCell40 \eeprom.i1_4_lut_adj_26_LC_6_25_6  (
            .in0(N__16289),
            .in1(N__16107),
            .in2(N__15701),
            .in3(N__16258),
            .lcout(\eeprom.n4218 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1424_3_lut_LC_6_25_7 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1424_3_lut_LC_6_25_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1424_3_lut_LC_6_25_7 .LUT_INIT=16'b1111110000001100;
    LogicCell40 \eeprom.rem_4_i1424_3_lut_LC_6_25_7  (
            .in0(_gnd_net_),
            .in1(N__16396),
            .in2(N__16368),
            .in3(N__16298),
            .lcout(\eeprom.n2212 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1486_2_lut_LC_6_26_0 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1486_2_lut_LC_6_26_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1486_2_lut_LC_6_26_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1486_2_lut_LC_6_26_0  (
            .in0(_gnd_net_),
            .in1(N__16288),
            .in2(_gnd_net_),
            .in3(N__16265),
            .lcout(\eeprom.n2286 ),
            .ltout(),
            .carryin(bfn_6_26_0_),
            .carryout(\eeprom.n3541 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1486_3_lut_LC_6_26_1 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1486_3_lut_LC_6_26_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1486_3_lut_LC_6_26_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1486_3_lut_LC_6_26_1  (
            .in0(_gnd_net_),
            .in1(N__27421),
            .in2(N__16262),
            .in3(N__16241),
            .lcout(\eeprom.n2285 ),
            .ltout(),
            .carryin(\eeprom.n3541 ),
            .carryout(\eeprom.n3542 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1486_4_lut_LC_6_26_2 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1486_4_lut_LC_6_26_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1486_4_lut_LC_6_26_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1486_4_lut_LC_6_26_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__16237),
            .in3(N__16208),
            .lcout(\eeprom.n2284 ),
            .ltout(),
            .carryin(\eeprom.n3542 ),
            .carryout(\eeprom.n3543 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1486_5_lut_LC_6_26_3 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1486_5_lut_LC_6_26_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1486_5_lut_LC_6_26_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1486_5_lut_LC_6_26_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__16205),
            .in3(N__16172),
            .lcout(\eeprom.n2283 ),
            .ltout(),
            .carryin(\eeprom.n3543 ),
            .carryout(\eeprom.n3544 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1486_6_lut_LC_6_26_4 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1486_6_lut_LC_6_26_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1486_6_lut_LC_6_26_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1486_6_lut_LC_6_26_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__16169),
            .in3(N__16142),
            .lcout(\eeprom.n2282 ),
            .ltout(),
            .carryin(\eeprom.n3544 ),
            .carryout(\eeprom.n3545 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1486_7_lut_LC_6_26_5 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1486_7_lut_LC_6_26_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1486_7_lut_LC_6_26_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1486_7_lut_LC_6_26_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__16139),
            .in3(N__16118),
            .lcout(\eeprom.n2281 ),
            .ltout(),
            .carryin(\eeprom.n3545 ),
            .carryout(\eeprom.n3546 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1486_8_lut_LC_6_26_6 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1486_8_lut_LC_6_26_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1486_8_lut_LC_6_26_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1486_8_lut_LC_6_26_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__16114),
            .in3(N__16712),
            .lcout(\eeprom.n2280 ),
            .ltout(),
            .carryin(\eeprom.n3546 ),
            .carryout(\eeprom.n3547 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1486_9_lut_LC_6_26_7 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1486_9_lut_LC_6_26_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1486_9_lut_LC_6_26_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1486_9_lut_LC_6_26_7  (
            .in0(_gnd_net_),
            .in1(N__27422),
            .in2(N__16709),
            .in3(N__16679),
            .lcout(\eeprom.n2279 ),
            .ltout(),
            .carryin(\eeprom.n3547 ),
            .carryout(\eeprom.n3548 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1486_10_lut_LC_6_27_0 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1486_10_lut_LC_6_27_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1486_10_lut_LC_6_27_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1486_10_lut_LC_6_27_0  (
            .in0(_gnd_net_),
            .in1(N__27607),
            .in2(N__16676),
            .in3(N__16640),
            .lcout(\eeprom.n2278 ),
            .ltout(),
            .carryin(bfn_6_27_0_),
            .carryout(\eeprom.n3549 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1486_11_lut_LC_6_27_1 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1486_11_lut_LC_6_27_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1486_11_lut_LC_6_27_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1486_11_lut_LC_6_27_1  (
            .in0(_gnd_net_),
            .in1(N__16637),
            .in2(N__27743),
            .in3(N__16607),
            .lcout(\eeprom.n2277 ),
            .ltout(),
            .carryin(\eeprom.n3549 ),
            .carryout(\eeprom.n3550 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1486_12_lut_LC_6_27_2 .C_ON=1'b0;
    defparam \eeprom.rem_4_add_1486_12_lut_LC_6_27_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1486_12_lut_LC_6_27_2 .LUT_INIT=16'b1000010001001000;
    LogicCell40 \eeprom.rem_4_add_1486_12_lut_LC_6_27_2  (
            .in0(N__27611),
            .in1(N__16604),
            .in2(N__16546),
            .in3(N__16526),
            .lcout(\eeprom.n2308 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1763_3_lut_LC_7_17_3 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1763_3_lut_LC_7_17_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1763_3_lut_LC_7_17_3 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \eeprom.rem_4_i1763_3_lut_LC_7_17_3  (
            .in0(_gnd_net_),
            .in1(N__16499),
            .in2(N__16469),
            .in3(N__17222),
            .lcout(\eeprom.n2711 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1757_3_lut_LC_7_18_0 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1757_3_lut_LC_7_18_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1757_3_lut_LC_7_18_0 .LUT_INIT=16'b1111101000001010;
    LogicCell40 \eeprom.rem_4_i1757_3_lut_LC_7_18_0  (
            .in0(N__16460),
            .in1(_gnd_net_),
            .in2(N__17220),
            .in3(N__16439),
            .lcout(\eeprom.n2705 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1764_3_lut_LC_7_18_1 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1764_3_lut_LC_7_18_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1764_3_lut_LC_7_18_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \eeprom.rem_4_i1764_3_lut_LC_7_18_1  (
            .in0(N__16433),
            .in1(N__16427),
            .in2(_gnd_net_),
            .in3(N__17210),
            .lcout(\eeprom.n2712 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1765_3_lut_LC_7_18_2 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1765_3_lut_LC_7_18_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1765_3_lut_LC_7_18_2 .LUT_INIT=16'b1111110000001100;
    LogicCell40 \eeprom.rem_4_i1765_3_lut_LC_7_18_2  (
            .in0(_gnd_net_),
            .in1(N__16856),
            .in2(N__17221),
            .in3(N__16826),
            .lcout(\eeprom.n2713 ),
            .ltout(\eeprom.n2713_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i1_2_lut_adj_29_LC_7_18_3 .C_ON=1'b0;
    defparam \eeprom.i1_2_lut_adj_29_LC_7_18_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.i1_2_lut_adj_29_LC_7_18_3 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \eeprom.i1_2_lut_adj_29_LC_7_18_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__16820),
            .in3(N__17376),
            .lcout(),
            .ltout(\eeprom.n4695_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i1_4_lut_adj_30_LC_7_18_4 .C_ON=1'b0;
    defparam \eeprom.i1_4_lut_adj_30_LC_7_18_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.i1_4_lut_adj_30_LC_7_18_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \eeprom.i1_4_lut_adj_30_LC_7_18_4  (
            .in0(N__17046),
            .in1(N__17430),
            .in2(N__16817),
            .in3(N__17319),
            .lcout(\eeprom.n4699 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i6_4_lut_LC_7_18_5 .C_ON=1'b0;
    defparam \eeprom.i6_4_lut_LC_7_18_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.i6_4_lut_LC_7_18_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \eeprom.i6_4_lut_LC_7_18_5  (
            .in0(N__18132),
            .in1(N__17706),
            .in2(N__17518),
            .in3(N__18459),
            .lcout(),
            .ltout(\eeprom.n16_adj_416_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i8_3_lut_LC_7_18_6 .C_ON=1'b0;
    defparam \eeprom.i8_3_lut_LC_7_18_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.i8_3_lut_LC_7_18_6 .LUT_INIT=16'b1111111111111100;
    LogicCell40 \eeprom.i8_3_lut_LC_7_18_6  (
            .in0(_gnd_net_),
            .in1(N__18504),
            .in2(N__16814),
            .in3(N__17487),
            .lcout(\eeprom.n18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1769_3_lut_LC_7_18_7 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1769_3_lut_LC_7_18_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1769_3_lut_LC_7_18_7 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \eeprom.rem_4_i1769_3_lut_LC_7_18_7  (
            .in0(_gnd_net_),
            .in1(N__16810),
            .in2(N__16790),
            .in3(N__17203),
            .lcout(\eeprom.n2717 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1758_3_lut_LC_7_19_0 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1758_3_lut_LC_7_19_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1758_3_lut_LC_7_19_0 .LUT_INIT=16'b1010110010101100;
    LogicCell40 \eeprom.rem_4_i1758_3_lut_LC_7_19_0  (
            .in0(N__16781),
            .in1(N__16953),
            .in2(N__17219),
            .in3(_gnd_net_),
            .lcout(\eeprom.n2706 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1770_3_lut_LC_7_19_1 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1770_3_lut_LC_7_19_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1770_3_lut_LC_7_19_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \eeprom.rem_4_i1770_3_lut_LC_7_19_1  (
            .in0(N__16775),
            .in1(N__16763),
            .in2(_gnd_net_),
            .in3(N__17194),
            .lcout(\eeprom.n2718 ),
            .ltout(\eeprom.n2718_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i3_4_lut_adj_31_LC_7_19_2 .C_ON=1'b0;
    defparam \eeprom.i3_4_lut_adj_31_LC_7_19_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.i3_4_lut_adj_31_LC_7_19_2 .LUT_INIT=16'b1111111011001100;
    LogicCell40 \eeprom.i3_4_lut_adj_31_LC_7_19_2  (
            .in0(N__17126),
            .in1(N__18369),
            .in2(N__16736),
            .in3(N__16733),
            .lcout(\eeprom.n13_adj_417 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1759_3_lut_LC_7_19_3 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1759_3_lut_LC_7_19_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1759_3_lut_LC_7_19_3 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \eeprom.rem_4_i1759_3_lut_LC_7_19_3  (
            .in0(N__16981),
            .in1(_gnd_net_),
            .in2(N__17018),
            .in3(N__17202),
            .lcout(\eeprom.n2707 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1766_3_lut_LC_7_19_4 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1766_3_lut_LC_7_19_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1766_3_lut_LC_7_19_4 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \eeprom.rem_4_i1766_3_lut_LC_7_19_4  (
            .in0(_gnd_net_),
            .in1(N__17009),
            .in2(N__17218),
            .in3(N__17003),
            .lcout(\eeprom.n2714 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i8_4_lut_LC_7_19_5 .C_ON=1'b0;
    defparam \eeprom.i8_4_lut_LC_7_19_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.i8_4_lut_LC_7_19_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \eeprom.i8_4_lut_LC_7_19_5  (
            .in0(N__16980),
            .in1(N__16967),
            .in2(N__16957),
            .in3(N__16937),
            .lcout(\eeprom.n2638 ),
            .ltout(\eeprom.n2638_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1767_3_lut_LC_7_19_6 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1767_3_lut_LC_7_19_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1767_3_lut_LC_7_19_6 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \eeprom.rem_4_i1767_3_lut_LC_7_19_6  (
            .in0(N__16925),
            .in1(_gnd_net_),
            .in2(N__16919),
            .in3(N__16916),
            .lcout(\eeprom.n2715 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1768_3_lut_LC_7_19_7 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1768_3_lut_LC_7_19_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1768_3_lut_LC_7_19_7 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \eeprom.rem_4_i1768_3_lut_LC_7_19_7  (
            .in0(_gnd_net_),
            .in1(N__16892),
            .in2(N__16868),
            .in3(N__17198),
            .lcout(\eeprom.n2716 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1837_3_lut_LC_7_20_0 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1837_3_lut_LC_7_20_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1837_3_lut_LC_7_20_0 .LUT_INIT=16'b1010110010101100;
    LogicCell40 \eeprom.rem_4_i1837_3_lut_LC_7_20_0  (
            .in0(N__17066),
            .in1(N__17080),
            .in2(N__18313),
            .in3(_gnd_net_),
            .lcout(\eeprom.n2817 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1838_3_lut_LC_7_20_1 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1838_3_lut_LC_7_20_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1838_3_lut_LC_7_20_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \eeprom.rem_4_i1838_3_lut_LC_7_20_1  (
            .in0(N__17122),
            .in1(N__17093),
            .in2(_gnd_net_),
            .in3(N__18278),
            .lcout(\eeprom.n2818 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1835_3_lut_LC_7_20_2 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1835_3_lut_LC_7_20_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1835_3_lut_LC_7_20_2 .LUT_INIT=16'b1111110000001100;
    LogicCell40 \eeprom.rem_4_i1835_3_lut_LC_7_20_2  (
            .in0(_gnd_net_),
            .in1(N__17050),
            .in2(N__18314),
            .in3(N__17030),
            .lcout(\eeprom.n2815 ),
            .ltout(\eeprom.n2815_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i1_2_lut_adj_32_LC_7_20_3 .C_ON=1'b0;
    defparam \eeprom.i1_2_lut_adj_32_LC_7_20_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.i1_2_lut_adj_32_LC_7_20_3 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \eeprom.i1_2_lut_adj_32_LC_7_20_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__16859),
            .in3(N__19615),
            .lcout(\eeprom.n4529 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_mux_3_i6_3_lut_LC_7_20_4 .C_ON=1'b0;
    defparam \eeprom.rem_4_mux_3_i6_3_lut_LC_7_20_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_mux_3_i6_3_lut_LC_7_20_4 .LUT_INIT=16'b0010001001110111;
    LogicCell40 \eeprom.rem_4_mux_3_i6_3_lut_LC_7_20_4  (
            .in0(N__22990),
            .in1(N__17273),
            .in2(_gnd_net_),
            .in3(N__23665),
            .lcout(\eeprom.n3720_adj_435 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1761_3_lut_LC_7_20_5 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1761_3_lut_LC_7_20_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1761_3_lut_LC_7_20_5 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \eeprom.rem_4_i1761_3_lut_LC_7_20_5  (
            .in0(_gnd_net_),
            .in1(N__17258),
            .in2(N__17231),
            .in3(N__17217),
            .lcout(\eeprom.n2709 ),
            .ltout(\eeprom.n2709_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i9_4_lut_LC_7_20_6 .C_ON=1'b0;
    defparam \eeprom.i9_4_lut_LC_7_20_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.i9_4_lut_LC_7_20_6 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \eeprom.i9_4_lut_LC_7_20_6  (
            .in0(N__17458),
            .in1(N__17147),
            .in2(N__17138),
            .in3(N__17135),
            .lcout(\eeprom.n2737 ),
            .ltout(\eeprom.n2737_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1833_3_lut_LC_7_20_7 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1833_3_lut_LC_7_20_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1833_3_lut_LC_7_20_7 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \eeprom.rem_4_i1833_3_lut_LC_7_20_7  (
            .in0(N__17303),
            .in1(_gnd_net_),
            .in2(N__17129),
            .in3(N__17323),
            .lcout(\eeprom.n2813 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1821_2_lut_LC_7_21_0 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1821_2_lut_LC_7_21_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1821_2_lut_LC_7_21_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1821_2_lut_LC_7_21_0  (
            .in0(_gnd_net_),
            .in1(N__17121),
            .in2(_gnd_net_),
            .in3(N__17087),
            .lcout(\eeprom.n2786 ),
            .ltout(),
            .carryin(bfn_7_21_0_),
            .carryout(\eeprom.n3601 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1821_3_lut_LC_7_21_1 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1821_3_lut_LC_7_21_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1821_3_lut_LC_7_21_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1821_3_lut_LC_7_21_1  (
            .in0(_gnd_net_),
            .in1(N__27589),
            .in2(N__17084),
            .in3(N__17060),
            .lcout(\eeprom.n2785 ),
            .ltout(),
            .carryin(\eeprom.n3601 ),
            .carryout(\eeprom.n3602 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1821_4_lut_LC_7_21_2 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1821_4_lut_LC_7_21_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1821_4_lut_LC_7_21_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1821_4_lut_LC_7_21_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__17437),
            .in3(N__17057),
            .lcout(\eeprom.n2784 ),
            .ltout(),
            .carryin(\eeprom.n3602 ),
            .carryout(\eeprom.n3603 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1821_5_lut_LC_7_21_3 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1821_5_lut_LC_7_21_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1821_5_lut_LC_7_21_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1821_5_lut_LC_7_21_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__17054),
            .in3(N__17024),
            .lcout(\eeprom.n2783 ),
            .ltout(),
            .carryin(\eeprom.n3603 ),
            .carryout(\eeprom.n3604 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1821_6_lut_LC_7_21_4 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1821_6_lut_LC_7_21_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1821_6_lut_LC_7_21_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1821_6_lut_LC_7_21_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__17389),
            .in3(N__17021),
            .lcout(\eeprom.n2782 ),
            .ltout(),
            .carryin(\eeprom.n3604 ),
            .carryout(\eeprom.n3605 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1821_7_lut_LC_7_21_5 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1821_7_lut_LC_7_21_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1821_7_lut_LC_7_21_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1821_7_lut_LC_7_21_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__17327),
            .in3(N__17297),
            .lcout(\eeprom.n2781 ),
            .ltout(),
            .carryin(\eeprom.n3605 ),
            .carryout(\eeprom.n3606 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1821_8_lut_LC_7_21_6 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1821_8_lut_LC_7_21_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1821_8_lut_LC_7_21_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1821_8_lut_LC_7_21_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__17362),
            .in3(N__17294),
            .lcout(\eeprom.n2780 ),
            .ltout(),
            .carryin(\eeprom.n3606 ),
            .carryout(\eeprom.n3607 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1821_9_lut_LC_7_21_7 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1821_9_lut_LC_7_21_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1821_9_lut_LC_7_21_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1821_9_lut_LC_7_21_7  (
            .in0(_gnd_net_),
            .in1(N__27590),
            .in2(N__18511),
            .in3(N__17291),
            .lcout(\eeprom.n2779 ),
            .ltout(),
            .carryin(\eeprom.n3607 ),
            .carryout(\eeprom.n3608 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1821_10_lut_LC_7_22_0 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1821_10_lut_LC_7_22_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1821_10_lut_LC_7_22_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1821_10_lut_LC_7_22_0  (
            .in0(_gnd_net_),
            .in1(N__17457),
            .in2(N__27381),
            .in3(N__17288),
            .lcout(\eeprom.n2778 ),
            .ltout(),
            .carryin(bfn_7_22_0_),
            .carryout(\eeprom.n3609 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1821_11_lut_LC_7_22_1 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1821_11_lut_LC_7_22_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1821_11_lut_LC_7_22_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1821_11_lut_LC_7_22_1  (
            .in0(_gnd_net_),
            .in1(N__27174),
            .in2(N__17492),
            .in3(N__17285),
            .lcout(\eeprom.n2777 ),
            .ltout(),
            .carryin(\eeprom.n3609 ),
            .carryout(\eeprom.n3610 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1821_12_lut_LC_7_22_2 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1821_12_lut_LC_7_22_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1821_12_lut_LC_7_22_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1821_12_lut_LC_7_22_2  (
            .in0(_gnd_net_),
            .in1(N__27642),
            .in2(N__17680),
            .in3(N__17282),
            .lcout(\eeprom.n2776 ),
            .ltout(),
            .carryin(\eeprom.n3610 ),
            .carryout(\eeprom.n3611 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1821_13_lut_LC_7_22_3 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1821_13_lut_LC_7_22_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1821_13_lut_LC_7_22_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1821_13_lut_LC_7_22_3  (
            .in0(_gnd_net_),
            .in1(N__27175),
            .in2(N__18382),
            .in3(N__17279),
            .lcout(\eeprom.n2775 ),
            .ltout(),
            .carryin(\eeprom.n3611 ),
            .carryout(\eeprom.n3612 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1821_14_lut_LC_7_22_4 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1821_14_lut_LC_7_22_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1821_14_lut_LC_7_22_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1821_14_lut_LC_7_22_4  (
            .in0(_gnd_net_),
            .in1(N__27643),
            .in2(N__18472),
            .in3(N__17276),
            .lcout(\eeprom.n2774 ),
            .ltout(),
            .carryin(\eeprom.n3612 ),
            .carryout(\eeprom.n3613 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1821_15_lut_LC_7_22_5 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1821_15_lut_LC_7_22_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1821_15_lut_LC_7_22_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1821_15_lut_LC_7_22_5  (
            .in0(_gnd_net_),
            .in1(N__17713),
            .in2(N__27752),
            .in3(N__17528),
            .lcout(\eeprom.n2773 ),
            .ltout(),
            .carryin(\eeprom.n3613 ),
            .carryout(\eeprom.n3614 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1821_16_lut_LC_7_22_6 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1821_16_lut_LC_7_22_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1821_16_lut_LC_7_22_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1821_16_lut_LC_7_22_6  (
            .in0(_gnd_net_),
            .in1(N__18139),
            .in2(N__27382),
            .in3(N__17525),
            .lcout(\eeprom.n2772 ),
            .ltout(),
            .carryin(\eeprom.n3614 ),
            .carryout(\eeprom.n3615 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1821_17_lut_LC_7_22_7 .C_ON=1'b0;
    defparam \eeprom.rem_4_add_1821_17_lut_LC_7_22_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1821_17_lut_LC_7_22_7 .LUT_INIT=16'b1000010001001000;
    LogicCell40 \eeprom.rem_4_add_1821_17_lut_LC_7_22_7  (
            .in0(N__27647),
            .in1(N__18326),
            .in2(N__17522),
            .in3(N__17501),
            .lcout(\eeprom.n2803 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1829_3_lut_LC_7_23_0 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1829_3_lut_LC_7_23_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1829_3_lut_LC_7_23_0 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \eeprom.rem_4_i1829_3_lut_LC_7_23_0  (
            .in0(_gnd_net_),
            .in1(N__17498),
            .in2(N__18339),
            .in3(N__17491),
            .lcout(\eeprom.n2809 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1830_3_lut_LC_7_23_2 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1830_3_lut_LC_7_23_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1830_3_lut_LC_7_23_2 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \eeprom.rem_4_i1830_3_lut_LC_7_23_2  (
            .in0(N__17465),
            .in1(_gnd_net_),
            .in2(N__18338),
            .in3(N__17459),
            .lcout(\eeprom.n2810 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1836_3_lut_LC_7_23_3 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1836_3_lut_LC_7_23_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1836_3_lut_LC_7_23_3 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \eeprom.rem_4_i1836_3_lut_LC_7_23_3  (
            .in0(_gnd_net_),
            .in1(N__17438),
            .in2(N__17411),
            .in3(N__18315),
            .lcout(\eeprom.n2816 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1834_3_lut_LC_7_23_4 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1834_3_lut_LC_7_23_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1834_3_lut_LC_7_23_4 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \eeprom.rem_4_i1834_3_lut_LC_7_23_4  (
            .in0(_gnd_net_),
            .in1(N__17399),
            .in2(N__18337),
            .in3(N__17390),
            .lcout(\eeprom.n2814 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1832_3_lut_LC_7_23_5 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1832_3_lut_LC_7_23_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1832_3_lut_LC_7_23_5 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \eeprom.rem_4_i1832_3_lut_LC_7_23_5  (
            .in0(_gnd_net_),
            .in1(N__17363),
            .in2(N__17342),
            .in3(N__18319),
            .lcout(\eeprom.n2812 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2223_2_lut_LC_9_17_0 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2223_2_lut_LC_9_17_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2223_2_lut_LC_9_17_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2223_2_lut_LC_9_17_0  (
            .in0(_gnd_net_),
            .in1(N__20274),
            .in2(_gnd_net_),
            .in3(N__17330),
            .lcout(\eeprom.n3386 ),
            .ltout(),
            .carryin(bfn_9_17_0_),
            .carryout(\eeprom.n3706 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2223_3_lut_LC_9_17_1 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2223_3_lut_LC_9_17_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2223_3_lut_LC_9_17_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2223_3_lut_LC_9_17_1  (
            .in0(_gnd_net_),
            .in1(N__27727),
            .in2(N__18809),
            .in3(N__17555),
            .lcout(\eeprom.n3385 ),
            .ltout(),
            .carryin(\eeprom.n3706 ),
            .carryout(\eeprom.n3707 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2223_4_lut_LC_9_17_2 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2223_4_lut_LC_9_17_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2223_4_lut_LC_9_17_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2223_4_lut_LC_9_17_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__19064),
            .in3(N__17552),
            .lcout(\eeprom.n3384 ),
            .ltout(),
            .carryin(\eeprom.n3707 ),
            .carryout(\eeprom.n3708 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2223_5_lut_LC_9_17_3 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2223_5_lut_LC_9_17_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2223_5_lut_LC_9_17_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2223_5_lut_LC_9_17_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__20249),
            .in3(N__17549),
            .lcout(\eeprom.n3383 ),
            .ltout(),
            .carryin(\eeprom.n3708 ),
            .carryout(\eeprom.n3709 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2223_6_lut_LC_9_17_4 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2223_6_lut_LC_9_17_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2223_6_lut_LC_9_17_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2223_6_lut_LC_9_17_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__19787),
            .in3(N__17546),
            .lcout(\eeprom.n3382 ),
            .ltout(),
            .carryin(\eeprom.n3709 ),
            .carryout(\eeprom.n3710 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2223_7_lut_LC_9_17_5 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2223_7_lut_LC_9_17_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2223_7_lut_LC_9_17_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2223_7_lut_LC_9_17_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__20206),
            .in3(N__17543),
            .lcout(\eeprom.n3381 ),
            .ltout(),
            .carryin(\eeprom.n3710 ),
            .carryout(\eeprom.n3711 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2223_8_lut_LC_9_17_6 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2223_8_lut_LC_9_17_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2223_8_lut_LC_9_17_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2223_8_lut_LC_9_17_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__20353),
            .in3(N__17540),
            .lcout(\eeprom.n3380 ),
            .ltout(),
            .carryin(\eeprom.n3711 ),
            .carryout(\eeprom.n3712 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2223_9_lut_LC_9_17_7 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2223_9_lut_LC_9_17_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2223_9_lut_LC_9_17_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2223_9_lut_LC_9_17_7  (
            .in0(_gnd_net_),
            .in1(N__27728),
            .in2(N__17950),
            .in3(N__17537),
            .lcout(\eeprom.n3379 ),
            .ltout(),
            .carryin(\eeprom.n3712 ),
            .carryout(\eeprom.n3713 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2223_10_lut_LC_9_18_0 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2223_10_lut_LC_9_18_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2223_10_lut_LC_9_18_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2223_10_lut_LC_9_18_0  (
            .in0(_gnd_net_),
            .in1(N__27769),
            .in2(N__20155),
            .in3(N__17534),
            .lcout(\eeprom.n3378 ),
            .ltout(),
            .carryin(bfn_9_18_0_),
            .carryout(\eeprom.n3714 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2223_11_lut_LC_9_18_1 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2223_11_lut_LC_9_18_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2223_11_lut_LC_9_18_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2223_11_lut_LC_9_18_1  (
            .in0(_gnd_net_),
            .in1(N__20385),
            .in2(N__27788),
            .in3(N__17531),
            .lcout(\eeprom.n3377 ),
            .ltout(),
            .carryin(\eeprom.n3714 ),
            .carryout(\eeprom.n3715 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2223_12_lut_LC_9_18_2 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2223_12_lut_LC_9_18_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2223_12_lut_LC_9_18_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2223_12_lut_LC_9_18_2  (
            .in0(_gnd_net_),
            .in1(N__27773),
            .in2(N__18910),
            .in3(N__17582),
            .lcout(\eeprom.n3376 ),
            .ltout(),
            .carryin(\eeprom.n3715 ),
            .carryout(\eeprom.n3716 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2223_13_lut_LC_9_18_3 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2223_13_lut_LC_9_18_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2223_13_lut_LC_9_18_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2223_13_lut_LC_9_18_3  (
            .in0(_gnd_net_),
            .in1(N__27776),
            .in2(N__19021),
            .in3(N__17579),
            .lcout(\eeprom.n3375 ),
            .ltout(),
            .carryin(\eeprom.n3716 ),
            .carryout(\eeprom.n3717 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2223_14_lut_LC_9_18_4 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2223_14_lut_LC_9_18_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2223_14_lut_LC_9_18_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2223_14_lut_LC_9_18_4  (
            .in0(_gnd_net_),
            .in1(N__27774),
            .in2(N__17915),
            .in3(N__17576),
            .lcout(\eeprom.n3374 ),
            .ltout(),
            .carryin(\eeprom.n3717 ),
            .carryout(\eeprom.n3718 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2223_15_lut_LC_9_18_5 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2223_15_lut_LC_9_18_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2223_15_lut_LC_9_18_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2223_15_lut_LC_9_18_5  (
            .in0(_gnd_net_),
            .in1(N__27777),
            .in2(N__18980),
            .in3(N__17573),
            .lcout(\eeprom.n3373 ),
            .ltout(),
            .carryin(\eeprom.n3718 ),
            .carryout(\eeprom.n3719 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2223_16_lut_LC_9_18_6 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2223_16_lut_LC_9_18_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2223_16_lut_LC_9_18_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2223_16_lut_LC_9_18_6  (
            .in0(_gnd_net_),
            .in1(N__27775),
            .in2(N__18947),
            .in3(N__17570),
            .lcout(\eeprom.n3372 ),
            .ltout(),
            .carryin(\eeprom.n3719 ),
            .carryout(\eeprom.n3720 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2223_17_lut_LC_9_18_7 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2223_17_lut_LC_9_18_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2223_17_lut_LC_9_18_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2223_17_lut_LC_9_18_7  (
            .in0(_gnd_net_),
            .in1(N__27778),
            .in2(N__18782),
            .in3(N__17567),
            .lcout(\eeprom.n3371 ),
            .ltout(),
            .carryin(\eeprom.n3720 ),
            .carryout(\eeprom.n3721 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2223_18_lut_LC_9_19_0 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2223_18_lut_LC_9_19_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2223_18_lut_LC_9_19_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2223_18_lut_LC_9_19_0  (
            .in0(_gnd_net_),
            .in1(N__27560),
            .in2(N__20693),
            .in3(N__17564),
            .lcout(\eeprom.n3370 ),
            .ltout(),
            .carryin(bfn_9_19_0_),
            .carryout(\eeprom.n3722 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2223_19_lut_LC_9_19_1 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2223_19_lut_LC_9_19_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2223_19_lut_LC_9_19_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2223_19_lut_LC_9_19_1  (
            .in0(_gnd_net_),
            .in1(N__18756),
            .in2(N__27725),
            .in3(N__17561),
            .lcout(\eeprom.n3369 ),
            .ltout(),
            .carryin(\eeprom.n3722 ),
            .carryout(\eeprom.n3723 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2223_20_lut_LC_9_19_2 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2223_20_lut_LC_9_19_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2223_20_lut_LC_9_19_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2223_20_lut_LC_9_19_2  (
            .in0(_gnd_net_),
            .in1(N__19309),
            .in2(N__27726),
            .in3(N__17558),
            .lcout(\eeprom.n3368 ),
            .ltout(),
            .carryin(\eeprom.n3723 ),
            .carryout(\eeprom.n3724 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2223_21_lut_LC_9_19_3 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2223_21_lut_LC_9_19_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2223_21_lut_LC_9_19_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2223_21_lut_LC_9_19_3  (
            .in0(_gnd_net_),
            .in1(N__27569),
            .in2(N__19360),
            .in3(N__17615),
            .lcout(\eeprom.n3367 ),
            .ltout(),
            .carryin(\eeprom.n3724 ),
            .carryout(\eeprom.n3725 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2223_22_lut_LC_9_19_4 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2223_22_lut_LC_9_19_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2223_22_lut_LC_9_19_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2223_22_lut_LC_9_19_4  (
            .in0(_gnd_net_),
            .in1(N__27564),
            .in2(N__20647),
            .in3(N__17612),
            .lcout(\eeprom.n3366 ),
            .ltout(),
            .carryin(\eeprom.n3725 ),
            .carryout(\eeprom.n3726 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2223_23_lut_LC_9_19_5 .C_ON=1'b0;
    defparam \eeprom.rem_4_add_2223_23_lut_LC_9_19_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2223_23_lut_LC_9_19_5 .LUT_INIT=16'b1001000001100000;
    LogicCell40 \eeprom.rem_4_add_2223_23_lut_LC_9_19_5  (
            .in0(N__27565),
            .in1(N__19336),
            .in2(N__20615),
            .in3(N__17609),
            .lcout(\eeprom.n3397 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2173_3_lut_LC_9_19_6 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2173_3_lut_LC_9_19_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2173_3_lut_LC_9_19_6 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \eeprom.rem_4_i2173_3_lut_LC_9_19_6  (
            .in0(_gnd_net_),
            .in1(N__20804),
            .in2(N__17591),
            .in3(N__19211),
            .lcout(\eeprom.n3313 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2156_2_lut_LC_9_20_0 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2156_2_lut_LC_9_20_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2156_2_lut_LC_9_20_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2156_2_lut_LC_9_20_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__19445),
            .in3(N__17606),
            .lcout(\eeprom.n3286 ),
            .ltout(),
            .carryin(bfn_9_20_0_),
            .carryout(\eeprom.n3686 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2156_3_lut_LC_9_20_1 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2156_3_lut_LC_9_20_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2156_3_lut_LC_9_20_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2156_3_lut_LC_9_20_1  (
            .in0(_gnd_net_),
            .in1(N__27556),
            .in2(N__19399),
            .in3(N__17603),
            .lcout(\eeprom.n3285 ),
            .ltout(),
            .carryin(\eeprom.n3686 ),
            .carryout(\eeprom.n3687 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2156_4_lut_LC_9_20_2 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2156_4_lut_LC_9_20_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2156_4_lut_LC_9_20_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2156_4_lut_LC_9_20_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__20426),
            .in3(N__17600),
            .lcout(\eeprom.n3284 ),
            .ltout(),
            .carryin(\eeprom.n3687 ),
            .carryout(\eeprom.n3688 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2156_5_lut_LC_9_20_3 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2156_5_lut_LC_9_20_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2156_5_lut_LC_9_20_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2156_5_lut_LC_9_20_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__20482),
            .in3(N__17597),
            .lcout(\eeprom.n3283 ),
            .ltout(),
            .carryin(\eeprom.n3688 ),
            .carryout(\eeprom.n3689 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2156_6_lut_LC_9_20_4 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2156_6_lut_LC_9_20_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2156_6_lut_LC_9_20_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2156_6_lut_LC_9_20_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__19519),
            .in3(N__17594),
            .lcout(\eeprom.n3282 ),
            .ltout(),
            .carryin(\eeprom.n3689 ),
            .carryout(\eeprom.n3690 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2156_7_lut_LC_9_20_5 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2156_7_lut_LC_9_20_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2156_7_lut_LC_9_20_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2156_7_lut_LC_9_20_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__20803),
            .in3(N__17645),
            .lcout(\eeprom.n3281 ),
            .ltout(),
            .carryin(\eeprom.n3690 ),
            .carryout(\eeprom.n3691 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2156_8_lut_LC_9_20_6 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2156_8_lut_LC_9_20_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2156_8_lut_LC_9_20_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2156_8_lut_LC_9_20_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__19550),
            .in3(N__17642),
            .lcout(\eeprom.n3280 ),
            .ltout(),
            .carryin(\eeprom.n3691 ),
            .carryout(\eeprom.n3692 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2156_9_lut_LC_9_20_7 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2156_9_lut_LC_9_20_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2156_9_lut_LC_9_20_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2156_9_lut_LC_9_20_7  (
            .in0(_gnd_net_),
            .in1(N__19112),
            .in2(N__27724),
            .in3(N__17639),
            .lcout(\eeprom.n3279 ),
            .ltout(),
            .carryin(\eeprom.n3692 ),
            .carryout(\eeprom.n3693 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2156_10_lut_LC_9_21_0 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2156_10_lut_LC_9_21_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2156_10_lut_LC_9_21_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2156_10_lut_LC_9_21_0  (
            .in0(_gnd_net_),
            .in1(N__27670),
            .in2(N__21264),
            .in3(N__17636),
            .lcout(\eeprom.n3278 ),
            .ltout(),
            .carryin(bfn_9_21_0_),
            .carryout(\eeprom.n3694 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2156_11_lut_LC_9_21_1 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2156_11_lut_LC_9_21_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2156_11_lut_LC_9_21_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2156_11_lut_LC_9_21_1  (
            .in0(_gnd_net_),
            .in1(N__19139),
            .in2(N__27765),
            .in3(N__17633),
            .lcout(\eeprom.n3277 ),
            .ltout(),
            .carryin(\eeprom.n3694 ),
            .carryout(\eeprom.n3695 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2156_12_lut_LC_9_21_2 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2156_12_lut_LC_9_21_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2156_12_lut_LC_9_21_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2156_12_lut_LC_9_21_2  (
            .in0(_gnd_net_),
            .in1(N__18035),
            .in2(N__27721),
            .in3(N__17630),
            .lcout(\eeprom.n3276 ),
            .ltout(),
            .carryin(\eeprom.n3695 ),
            .carryout(\eeprom.n3696 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2156_13_lut_LC_9_21_3 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2156_13_lut_LC_9_21_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2156_13_lut_LC_9_21_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2156_13_lut_LC_9_21_3  (
            .in0(_gnd_net_),
            .in1(N__19090),
            .in2(N__27766),
            .in3(N__17627),
            .lcout(\eeprom.n3275 ),
            .ltout(),
            .carryin(\eeprom.n3696 ),
            .carryout(\eeprom.n3697 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2156_14_lut_LC_9_21_4 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2156_14_lut_LC_9_21_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2156_14_lut_LC_9_21_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2156_14_lut_LC_9_21_4  (
            .in0(_gnd_net_),
            .in1(N__21559),
            .in2(N__27722),
            .in3(N__17624),
            .lcout(\eeprom.n3274 ),
            .ltout(),
            .carryin(\eeprom.n3697 ),
            .carryout(\eeprom.n3698 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2156_15_lut_LC_9_21_5 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2156_15_lut_LC_9_21_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2156_15_lut_LC_9_21_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2156_15_lut_LC_9_21_5  (
            .in0(_gnd_net_),
            .in1(N__20830),
            .in2(N__27767),
            .in3(N__17621),
            .lcout(\eeprom.n3273 ),
            .ltout(),
            .carryin(\eeprom.n3698 ),
            .carryout(\eeprom.n3699 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2156_16_lut_LC_9_21_6 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2156_16_lut_LC_9_21_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2156_16_lut_LC_9_21_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2156_16_lut_LC_9_21_6  (
            .in0(_gnd_net_),
            .in1(N__21676),
            .in2(N__27723),
            .in3(N__17618),
            .lcout(\eeprom.n3272 ),
            .ltout(),
            .carryin(\eeprom.n3699 ),
            .carryout(\eeprom.n3700 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2156_17_lut_LC_9_21_7 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2156_17_lut_LC_9_21_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2156_17_lut_LC_9_21_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2156_17_lut_LC_9_21_7  (
            .in0(_gnd_net_),
            .in1(N__21306),
            .in2(N__27768),
            .in3(N__17735),
            .lcout(\eeprom.n3271 ),
            .ltout(),
            .carryin(\eeprom.n3700 ),
            .carryout(\eeprom.n3701 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2156_18_lut_LC_9_22_0 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2156_18_lut_LC_9_22_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2156_18_lut_LC_9_22_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2156_18_lut_LC_9_22_0  (
            .in0(_gnd_net_),
            .in1(N__20449),
            .in2(N__27750),
            .in3(N__17732),
            .lcout(\eeprom.n3270 ),
            .ltout(),
            .carryin(bfn_9_22_0_),
            .carryout(\eeprom.n3702 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2156_19_lut_LC_9_22_1 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2156_19_lut_LC_9_22_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2156_19_lut_LC_9_22_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2156_19_lut_LC_9_22_1  (
            .in0(_gnd_net_),
            .in1(N__21925),
            .in2(N__27333),
            .in3(N__17729),
            .lcout(\eeprom.n3269 ),
            .ltout(),
            .carryin(\eeprom.n3702 ),
            .carryout(\eeprom.n3703 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2156_20_lut_LC_9_22_2 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2156_20_lut_LC_9_22_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2156_20_lut_LC_9_22_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2156_20_lut_LC_9_22_2  (
            .in0(_gnd_net_),
            .in1(N__21580),
            .in2(N__27751),
            .in3(N__17726),
            .lcout(\eeprom.n3268 ),
            .ltout(),
            .carryin(\eeprom.n3703 ),
            .carryout(\eeprom.n3704 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2156_21_lut_LC_9_22_3 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2156_21_lut_LC_9_22_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2156_21_lut_LC_9_22_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2156_21_lut_LC_9_22_3  (
            .in0(_gnd_net_),
            .in1(N__21889),
            .in2(N__27334),
            .in3(N__17723),
            .lcout(\eeprom.n3267 ),
            .ltout(),
            .carryin(\eeprom.n3704 ),
            .carryout(\eeprom.n3705 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2156_22_lut_LC_9_22_4 .C_ON=1'b0;
    defparam \eeprom.rem_4_add_2156_22_lut_LC_9_22_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2156_22_lut_LC_9_22_4 .LUT_INIT=16'b1001000001100000;
    LogicCell40 \eeprom.rem_4_add_2156_22_lut_LC_9_22_4  (
            .in0(N__27641),
            .in1(N__21650),
            .in2(N__19268),
            .in3(N__17720),
            .lcout(\eeprom.n3298 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1825_3_lut_LC_9_22_6 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1825_3_lut_LC_9_22_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1825_3_lut_LC_9_22_6 .LUT_INIT=16'b1111110000001100;
    LogicCell40 \eeprom.rem_4_i1825_3_lut_LC_9_22_6  (
            .in0(_gnd_net_),
            .in1(N__17717),
            .in2(N__18340),
            .in3(N__17690),
            .lcout(\eeprom.n2805 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1828_3_lut_LC_9_22_7 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1828_3_lut_LC_9_22_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1828_3_lut_LC_9_22_7 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \eeprom.rem_4_i1828_3_lut_LC_9_22_7  (
            .in0(_gnd_net_),
            .in1(N__17681),
            .in2(N__17657),
            .in3(N__18327),
            .lcout(\eeprom.n2808 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1888_2_lut_LC_9_23_0 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1888_2_lut_LC_9_23_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1888_2_lut_LC_9_23_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1888_2_lut_LC_9_23_0  (
            .in0(_gnd_net_),
            .in1(N__18693),
            .in2(_gnd_net_),
            .in3(N__17765),
            .lcout(\eeprom.n2886 ),
            .ltout(),
            .carryin(bfn_9_23_0_),
            .carryout(\eeprom.n3616 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1888_3_lut_LC_9_23_1 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1888_3_lut_LC_9_23_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1888_3_lut_LC_9_23_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1888_3_lut_LC_9_23_1  (
            .in0(_gnd_net_),
            .in1(N__27459),
            .in2(N__18550),
            .in3(N__17762),
            .lcout(\eeprom.n2885 ),
            .ltout(),
            .carryin(\eeprom.n3616 ),
            .carryout(\eeprom.n3617 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1888_4_lut_LC_9_23_2 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1888_4_lut_LC_9_23_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1888_4_lut_LC_9_23_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1888_4_lut_LC_9_23_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__20131),
            .in3(N__17759),
            .lcout(\eeprom.n2884 ),
            .ltout(),
            .carryin(\eeprom.n3617 ),
            .carryout(\eeprom.n3618 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1888_5_lut_LC_9_23_3 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1888_5_lut_LC_9_23_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1888_5_lut_LC_9_23_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1888_5_lut_LC_9_23_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__18654),
            .in3(N__17756),
            .lcout(\eeprom.n2883 ),
            .ltout(),
            .carryin(\eeprom.n3618 ),
            .carryout(\eeprom.n3619 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1888_6_lut_LC_9_23_4 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1888_6_lut_LC_9_23_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1888_6_lut_LC_9_23_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1888_6_lut_LC_9_23_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__18202),
            .in3(N__17753),
            .lcout(\eeprom.n2882 ),
            .ltout(),
            .carryin(\eeprom.n3619 ),
            .carryout(\eeprom.n3620 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1888_7_lut_LC_9_23_5 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1888_7_lut_LC_9_23_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1888_7_lut_LC_9_23_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1888_7_lut_LC_9_23_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__18719),
            .in3(N__17750),
            .lcout(\eeprom.n2881 ),
            .ltout(),
            .carryin(\eeprom.n3620 ),
            .carryout(\eeprom.n3621 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1888_8_lut_LC_9_23_6 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1888_8_lut_LC_9_23_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1888_8_lut_LC_9_23_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1888_8_lut_LC_9_23_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__19633),
            .in3(N__17747),
            .lcout(\eeprom.n2880 ),
            .ltout(),
            .carryin(\eeprom.n3621 ),
            .carryout(\eeprom.n3622 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1888_9_lut_LC_9_23_7 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1888_9_lut_LC_9_23_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1888_9_lut_LC_9_23_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1888_9_lut_LC_9_23_7  (
            .in0(_gnd_net_),
            .in1(N__19668),
            .in2(N__27546),
            .in3(N__17744),
            .lcout(\eeprom.n2879 ),
            .ltout(),
            .carryin(\eeprom.n3622 ),
            .carryout(\eeprom.n3623 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1888_10_lut_LC_9_24_0 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1888_10_lut_LC_9_24_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1888_10_lut_LC_9_24_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1888_10_lut_LC_9_24_0  (
            .in0(_gnd_net_),
            .in1(N__27411),
            .in2(N__19996),
            .in3(N__17741),
            .lcout(\eeprom.n2878 ),
            .ltout(),
            .carryin(bfn_9_24_0_),
            .carryout(\eeprom.n3624 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1888_11_lut_LC_9_24_1 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1888_11_lut_LC_9_24_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1888_11_lut_LC_9_24_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1888_11_lut_LC_9_24_1  (
            .in0(_gnd_net_),
            .in1(N__20071),
            .in2(N__27604),
            .in3(N__17738),
            .lcout(\eeprom.n2877 ),
            .ltout(),
            .carryin(\eeprom.n3624 ),
            .carryout(\eeprom.n3625 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1888_12_lut_LC_9_24_2 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1888_12_lut_LC_9_24_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1888_12_lut_LC_9_24_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1888_12_lut_LC_9_24_2  (
            .in0(_gnd_net_),
            .in1(N__18621),
            .in2(N__27586),
            .in3(N__17801),
            .lcout(\eeprom.n2876 ),
            .ltout(),
            .carryin(\eeprom.n3625 ),
            .carryout(\eeprom.n3626 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1888_13_lut_LC_9_24_3 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1888_13_lut_LC_9_24_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1888_13_lut_LC_9_24_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1888_13_lut_LC_9_24_3  (
            .in0(_gnd_net_),
            .in1(N__18862),
            .in2(N__27605),
            .in3(N__17798),
            .lcout(\eeprom.n2875 ),
            .ltout(),
            .carryin(\eeprom.n3626 ),
            .carryout(\eeprom.n3627 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1888_14_lut_LC_9_24_4 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1888_14_lut_LC_9_24_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1888_14_lut_LC_9_24_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1888_14_lut_LC_9_24_4  (
            .in0(_gnd_net_),
            .in1(N__18251),
            .in2(N__27587),
            .in3(N__17795),
            .lcout(\eeprom.n2874 ),
            .ltout(),
            .carryin(\eeprom.n3627 ),
            .carryout(\eeprom.n3628 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1888_15_lut_LC_9_24_5 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1888_15_lut_LC_9_24_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1888_15_lut_LC_9_24_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1888_15_lut_LC_9_24_5  (
            .in0(_gnd_net_),
            .in1(N__27393),
            .in2(N__18433),
            .in3(N__17792),
            .lcout(\eeprom.n2873 ),
            .ltout(),
            .carryin(\eeprom.n3628 ),
            .carryout(\eeprom.n3629 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1888_16_lut_LC_9_24_6 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1888_16_lut_LC_9_24_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1888_16_lut_LC_9_24_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1888_16_lut_LC_9_24_6  (
            .in0(_gnd_net_),
            .in1(N__18409),
            .in2(N__27588),
            .in3(N__17789),
            .lcout(\eeprom.n2872 ),
            .ltout(),
            .carryin(\eeprom.n3629 ),
            .carryout(\eeprom.n3630 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1888_17_lut_LC_9_24_7 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1888_17_lut_LC_9_24_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1888_17_lut_LC_9_24_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1888_17_lut_LC_9_24_7  (
            .in0(_gnd_net_),
            .in1(N__18587),
            .in2(N__27606),
            .in3(N__17786),
            .lcout(\eeprom.n2871 ),
            .ltout(),
            .carryin(\eeprom.n3630 ),
            .carryout(\eeprom.n3631 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1888_18_lut_LC_9_25_0 .C_ON=1'b0;
    defparam \eeprom.rem_4_add_1888_18_lut_LC_9_25_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1888_18_lut_LC_9_25_0 .LUT_INIT=16'b1000010001001000;
    LogicCell40 \eeprom.rem_4_add_1888_18_lut_LC_9_25_0  (
            .in0(N__27410),
            .in1(N__19959),
            .in2(N__18101),
            .in3(N__17783),
            .lcout(\eeprom.n2902 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1893_3_lut_LC_9_25_1 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1893_3_lut_LC_9_25_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1893_3_lut_LC_9_25_1 .LUT_INIT=16'b1111110000001100;
    LogicCell40 \eeprom.rem_4_i1893_3_lut_LC_9_25_1  (
            .in0(_gnd_net_),
            .in1(N__18434),
            .in2(N__19967),
            .in3(N__17780),
            .lcout(\eeprom.n2905 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1892_3_lut_LC_9_25_2 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1892_3_lut_LC_9_25_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1892_3_lut_LC_9_25_2 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \eeprom.rem_4_i1892_3_lut_LC_9_25_2  (
            .in0(_gnd_net_),
            .in1(N__18410),
            .in2(N__17774),
            .in3(N__19963),
            .lcout(\eeprom.n2904 ),
            .ltout(\eeprom.n2904_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i7_4_lut_adj_37_LC_9_25_3 .C_ON=1'b0;
    defparam \eeprom.i7_4_lut_adj_37_LC_9_25_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.i7_4_lut_adj_37_LC_9_25_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \eeprom.i7_4_lut_adj_37_LC_9_25_3  (
            .in0(N__19703),
            .in1(N__19747),
            .in2(N__17870),
            .in3(N__21481),
            .lcout(\eeprom.n19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2178_3_lut_LC_10_17_0 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2178_3_lut_LC_10_17_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2178_3_lut_LC_10_17_0 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \eeprom.rem_4_i2178_3_lut_LC_10_17_0  (
            .in0(N__19431),
            .in1(_gnd_net_),
            .in2(N__17867),
            .in3(N__19239),
            .lcout(\eeprom.n3318 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2177_3_lut_LC_10_17_2 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2177_3_lut_LC_10_17_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2177_3_lut_LC_10_17_2 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \eeprom.rem_4_i2177_3_lut_LC_10_17_2  (
            .in0(_gnd_net_),
            .in1(N__17852),
            .in2(N__19403),
            .in3(N__19240),
            .lcout(\eeprom.n3317 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2231_3_lut_LC_10_17_4 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2231_3_lut_LC_10_17_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2231_3_lut_LC_10_17_4 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \eeprom.rem_4_i2231_3_lut_LC_10_17_4  (
            .in0(_gnd_net_),
            .in1(N__18781),
            .in2(N__17843),
            .in3(N__20596),
            .lcout(\eeprom.n3403 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2174_3_lut_LC_10_17_5 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2174_3_lut_LC_10_17_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2174_3_lut_LC_10_17_5 .LUT_INIT=16'b1111110000001100;
    LogicCell40 \eeprom.rem_4_i2174_3_lut_LC_10_17_5  (
            .in0(_gnd_net_),
            .in1(N__19520),
            .in2(N__19262),
            .in3(N__17834),
            .lcout(\eeprom.n3314 ),
            .ltout(\eeprom.n3314_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i1_3_lut_adj_96_LC_10_17_6 .C_ON=1'b0;
    defparam \eeprom.i1_3_lut_adj_96_LC_10_17_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.i1_3_lut_adj_96_LC_10_17_6 .LUT_INIT=16'b1100000000000000;
    LogicCell40 \eeprom.i1_3_lut_adj_96_LC_10_17_6  (
            .in0(_gnd_net_),
            .in1(N__19062),
            .in2(N__17825),
            .in3(N__20248),
            .lcout(\eeprom.n4721 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2164_3_lut_LC_10_18_0 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2164_3_lut_LC_10_18_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2164_3_lut_LC_10_18_0 .LUT_INIT=16'b1111110000001100;
    LogicCell40 \eeprom.rem_4_i2164_3_lut_LC_10_18_0  (
            .in0(_gnd_net_),
            .in1(N__21680),
            .in2(N__19256),
            .in3(N__17822),
            .lcout(\eeprom.n3304 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i12_4_lut_adj_98_LC_10_18_1 .C_ON=1'b0;
    defparam \eeprom.i12_4_lut_adj_98_LC_10_18_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.i12_4_lut_adj_98_LC_10_18_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \eeprom.i12_4_lut_adj_98_LC_10_18_1  (
            .in0(N__17914),
            .in1(N__19017),
            .in2(N__17951),
            .in3(N__18906),
            .lcout(\eeprom.n28_adj_484 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2166_3_lut_LC_10_18_2 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2166_3_lut_LC_10_18_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2166_3_lut_LC_10_18_2 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \eeprom.rem_4_i2166_3_lut_LC_10_18_2  (
            .in0(N__17810),
            .in1(_gnd_net_),
            .in2(N__19257),
            .in3(N__21563),
            .lcout(\eeprom.n3306 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2165_3_lut_LC_10_18_3 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2165_3_lut_LC_10_18_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2165_3_lut_LC_10_18_3 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \eeprom.rem_4_i2165_3_lut_LC_10_18_3  (
            .in0(_gnd_net_),
            .in1(N__17969),
            .in2(N__20840),
            .in3(N__19224),
            .lcout(\eeprom.n3305 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2172_3_lut_LC_10_18_4 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2172_3_lut_LC_10_18_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2172_3_lut_LC_10_18_4 .LUT_INIT=16'b1010110010101100;
    LogicCell40 \eeprom.rem_4_i2172_3_lut_LC_10_18_4  (
            .in0(N__17960),
            .in1(N__19549),
            .in2(N__19254),
            .in3(_gnd_net_),
            .lcout(\eeprom.n3312 ),
            .ltout(\eeprom.n3312_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2239_3_lut_LC_10_18_5 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2239_3_lut_LC_10_18_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2239_3_lut_LC_10_18_5 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \eeprom.rem_4_i2239_3_lut_LC_10_18_5  (
            .in0(_gnd_net_),
            .in1(N__17933),
            .in2(N__17927),
            .in3(N__20607),
            .lcout(\eeprom.n3411 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2167_3_lut_LC_10_18_6 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2167_3_lut_LC_10_18_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2167_3_lut_LC_10_18_6 .LUT_INIT=16'b1111110000001100;
    LogicCell40 \eeprom.rem_4_i2167_3_lut_LC_10_18_6  (
            .in0(_gnd_net_),
            .in1(N__19094),
            .in2(N__19255),
            .in3(N__17924),
            .lcout(\eeprom.n3307 ),
            .ltout(\eeprom.n3307_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2234_3_lut_LC_10_18_7 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2234_3_lut_LC_10_18_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2234_3_lut_LC_10_18_7 .LUT_INIT=16'b1010101011110000;
    LogicCell40 \eeprom.rem_4_i2234_3_lut_LC_10_18_7  (
            .in0(N__17900),
            .in1(_gnd_net_),
            .in2(N__17894),
            .in3(N__20606),
            .lcout(\eeprom.n3406 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i13_4_lut_adj_94_LC_10_19_0 .C_ON=1'b0;
    defparam \eeprom.i13_4_lut_adj_94_LC_10_19_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.i13_4_lut_adj_94_LC_10_19_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \eeprom.i13_4_lut_adj_94_LC_10_19_0  (
            .in0(N__19110),
            .in1(N__18033),
            .in2(N__19073),
            .in3(N__19373),
            .lcout(),
            .ltout(\eeprom.n28_adj_482_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i14_4_lut_LC_10_19_1 .C_ON=1'b0;
    defparam \eeprom.i14_4_lut_LC_10_19_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.i14_4_lut_LC_10_19_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \eeprom.i14_4_lut_LC_10_19_1  (
            .in0(N__21533),
            .in1(N__21265),
            .in2(N__17891),
            .in3(N__21632),
            .lcout(\eeprom.n3232 ),
            .ltout(\eeprom.n3232_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2170_3_lut_LC_10_19_2 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2170_3_lut_LC_10_19_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2170_3_lut_LC_10_19_2 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \eeprom.rem_4_i2170_3_lut_LC_10_19_2  (
            .in0(N__17888),
            .in1(_gnd_net_),
            .in2(N__17879),
            .in3(N__21269),
            .lcout(\eeprom.n3310 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2227_3_lut_LC_10_19_3 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2227_3_lut_LC_10_19_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2227_3_lut_LC_10_19_3 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \eeprom.rem_4_i2227_3_lut_LC_10_19_3  (
            .in0(_gnd_net_),
            .in1(N__17876),
            .in2(N__19361),
            .in3(N__20578),
            .lcout(\eeprom.n3399 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2168_3_lut_LC_10_19_4 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2168_3_lut_LC_10_19_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2168_3_lut_LC_10_19_4 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \eeprom.rem_4_i2168_3_lut_LC_10_19_4  (
            .in0(_gnd_net_),
            .in1(N__18074),
            .in2(N__19258),
            .in3(N__18034),
            .lcout(\eeprom.n3308 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2171_3_lut_LC_10_19_5 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2171_3_lut_LC_10_19_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2171_3_lut_LC_10_19_5 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \eeprom.rem_4_i2171_3_lut_LC_10_19_5  (
            .in0(_gnd_net_),
            .in1(N__19111),
            .in2(N__18065),
            .in3(N__19225),
            .lcout(\eeprom.n3311 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2163_3_lut_LC_10_19_6 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2163_3_lut_LC_10_19_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2163_3_lut_LC_10_19_6 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \eeprom.rem_4_i2163_3_lut_LC_10_19_6  (
            .in0(N__18056),
            .in1(_gnd_net_),
            .in2(N__19259),
            .in3(N__21311),
            .lcout(\eeprom.n3303 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2169_rep_54_3_lut_LC_10_19_7 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2169_rep_54_3_lut_LC_10_19_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2169_rep_54_3_lut_LC_10_19_7 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \eeprom.rem_4_i2169_rep_54_3_lut_LC_10_19_7  (
            .in0(_gnd_net_),
            .in1(N__19135),
            .in2(N__18047),
            .in3(N__19226),
            .lcout(\eeprom.n3309 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2101_3_lut_LC_10_20_0 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2101_3_lut_LC_10_20_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2101_3_lut_LC_10_20_0 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \eeprom.rem_4_i2101_3_lut_LC_10_20_0  (
            .in0(_gnd_net_),
            .in1(N__24215),
            .in2(N__20873),
            .in3(N__21793),
            .lcout(\eeprom.n3209 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2229_3_lut_LC_10_20_1 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2229_3_lut_LC_10_20_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2229_3_lut_LC_10_20_1 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \eeprom.rem_4_i2229_3_lut_LC_10_20_1  (
            .in0(_gnd_net_),
            .in1(N__18020),
            .in2(N__20611),
            .in3(N__18757),
            .lcout(\eeprom.n3401 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_mux_3_i7_3_lut_LC_10_20_3 .C_ON=1'b0;
    defparam \eeprom.rem_4_mux_3_i7_3_lut_LC_10_20_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_mux_3_i7_3_lut_LC_10_20_3 .LUT_INIT=16'b0100010001110111;
    LogicCell40 \eeprom.rem_4_mux_3_i7_3_lut_LC_10_20_3  (
            .in0(N__18014),
            .in1(N__22950),
            .in2(_gnd_net_),
            .in3(N__23611),
            .lcout(\eeprom.n3719_adj_436 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2160_3_lut_LC_10_20_4 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2160_3_lut_LC_10_20_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2160_3_lut_LC_10_20_4 .LUT_INIT=16'b1111110000001100;
    LogicCell40 \eeprom.rem_4_i2160_3_lut_LC_10_20_4  (
            .in0(_gnd_net_),
            .in1(N__21584),
            .in2(N__19260),
            .in3(N__17996),
            .lcout(\eeprom.n3300 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_mux_3_i2_3_lut_LC_10_20_5 .C_ON=1'b0;
    defparam \eeprom.rem_4_mux_3_i2_3_lut_LC_10_20_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_mux_3_i2_3_lut_LC_10_20_5 .LUT_INIT=16'b0100010001110111;
    LogicCell40 \eeprom.rem_4_mux_3_i2_3_lut_LC_10_20_5  (
            .in0(N__17987),
            .in1(N__22949),
            .in2(_gnd_net_),
            .in3(N__23908),
            .lcout(\eeprom.n3724_adj_335 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2161_3_lut_LC_10_20_6 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2161_3_lut_LC_10_20_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2161_3_lut_LC_10_20_6 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \eeprom.rem_4_i2161_3_lut_LC_10_20_6  (
            .in0(_gnd_net_),
            .in1(N__18212),
            .in2(N__19261),
            .in3(N__21926),
            .lcout(\eeprom.n3301 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1902_3_lut_LC_10_21_0 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1902_3_lut_LC_10_21_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1902_3_lut_LC_10_21_0 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \eeprom.rem_4_i1902_3_lut_LC_10_21_0  (
            .in0(_gnd_net_),
            .in1(N__18203),
            .in2(N__18179),
            .in3(N__19954),
            .lcout(\eeprom.n2914 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2110_3_lut_LC_10_21_1 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2110_3_lut_LC_10_21_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2110_3_lut_LC_10_21_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \eeprom.rem_4_i2110_3_lut_LC_10_21_1  (
            .in0(N__20767),
            .in1(N__20726),
            .in2(_gnd_net_),
            .in3(N__21789),
            .lcout(\eeprom.n3218 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1906_3_lut_LC_10_21_3 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1906_3_lut_LC_10_21_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1906_3_lut_LC_10_21_3 .LUT_INIT=16'b1111101000001010;
    LogicCell40 \eeprom.rem_4_i1906_3_lut_LC_10_21_3  (
            .in0(N__18698),
            .in1(_gnd_net_),
            .in2(N__19966),
            .in3(N__18167),
            .lcout(\eeprom.n2918 ),
            .ltout(\eeprom.n2918_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1973_3_lut_LC_10_21_4 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1973_3_lut_LC_10_21_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1973_3_lut_LC_10_21_4 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \eeprom.rem_4_i1973_3_lut_LC_10_21_4  (
            .in0(_gnd_net_),
            .in1(N__19466),
            .in2(N__18155),
            .in3(N__24735),
            .lcout(\eeprom.n3017 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2100_3_lut_LC_10_21_5 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2100_3_lut_LC_10_21_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2100_3_lut_LC_10_21_5 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \eeprom.rem_4_i2100_3_lut_LC_10_21_5  (
            .in0(_gnd_net_),
            .in1(N__24248),
            .in2(N__21053),
            .in3(N__21790),
            .lcout(\eeprom.n3208 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2159_3_lut_LC_10_21_7 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2159_3_lut_LC_10_21_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2159_3_lut_LC_10_21_7 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \eeprom.rem_4_i2159_3_lut_LC_10_21_7  (
            .in0(_gnd_net_),
            .in1(N__21890),
            .in2(N__18152),
            .in3(N__19267),
            .lcout(\eeprom.n3299 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1824_3_lut_LC_10_22_0 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1824_3_lut_LC_10_22_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1824_3_lut_LC_10_22_0 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \eeprom.rem_4_i1824_3_lut_LC_10_22_0  (
            .in0(_gnd_net_),
            .in1(N__18143),
            .in2(N__18116),
            .in3(N__18336),
            .lcout(\eeprom.n2804 ),
            .ltout(\eeprom.n2804_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i9_4_lut_adj_34_LC_10_22_1 .C_ON=1'b0;
    defparam \eeprom.i9_4_lut_adj_34_LC_10_22_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.i9_4_lut_adj_34_LC_10_22_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \eeprom.i9_4_lut_adj_34_LC_10_22_1  (
            .in0(N__18094),
            .in1(N__19983),
            .in2(N__18077),
            .in3(N__18389),
            .lcout(\eeprom.n20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2162_3_lut_LC_10_22_2 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2162_3_lut_LC_10_22_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2162_3_lut_LC_10_22_2 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \eeprom.rem_4_i2162_3_lut_LC_10_22_2  (
            .in0(_gnd_net_),
            .in1(N__18521),
            .in2(N__20453),
            .in3(N__19266),
            .lcout(\eeprom.n3302 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1831_3_lut_LC_10_22_3 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1831_3_lut_LC_10_22_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1831_3_lut_LC_10_22_3 .LUT_INIT=16'b1111110000001100;
    LogicCell40 \eeprom.rem_4_i1831_3_lut_LC_10_22_3  (
            .in0(_gnd_net_),
            .in1(N__18515),
            .in2(N__18341),
            .in3(N__18485),
            .lcout(\eeprom.n2811 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1826_3_lut_LC_10_22_4 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1826_3_lut_LC_10_22_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1826_3_lut_LC_10_22_4 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \eeprom.rem_4_i1826_3_lut_LC_10_22_4  (
            .in0(_gnd_net_),
            .in1(N__18473),
            .in2(N__18446),
            .in3(N__18332),
            .lcout(\eeprom.n2806 ),
            .ltout(\eeprom.n2806_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i7_4_lut_LC_10_22_5 .C_ON=1'b0;
    defparam \eeprom.i7_4_lut_LC_10_22_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.i7_4_lut_LC_10_22_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \eeprom.i7_4_lut_LC_10_22_5  (
            .in0(N__18247),
            .in1(N__18855),
            .in2(N__18413),
            .in3(N__18402),
            .lcout(\eeprom.n18_adj_418 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1827_3_lut_LC_10_22_6 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1827_3_lut_LC_10_22_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1827_3_lut_LC_10_22_6 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \eeprom.rem_4_i1827_3_lut_LC_10_22_6  (
            .in0(_gnd_net_),
            .in1(N__18383),
            .in2(N__18353),
            .in3(N__18331),
            .lcout(\eeprom.n2807 ),
            .ltout(\eeprom.n2807_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1894_3_lut_LC_10_22_7 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1894_3_lut_LC_10_22_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1894_3_lut_LC_10_22_7 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \eeprom.rem_4_i1894_3_lut_LC_10_22_7  (
            .in0(_gnd_net_),
            .in1(N__18236),
            .in2(N__18227),
            .in3(N__19935),
            .lcout(\eeprom.n2906 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1901_3_lut_LC_10_23_0 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1901_3_lut_LC_10_23_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1901_3_lut_LC_10_23_0 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \eeprom.rem_4_i1901_3_lut_LC_10_23_0  (
            .in0(_gnd_net_),
            .in1(N__18718),
            .in2(N__18224),
            .in3(N__19930),
            .lcout(\eeprom.n2913 ),
            .ltout(\eeprom.n2913_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i1_2_lut_adj_27_LC_10_23_1 .C_ON=1'b0;
    defparam \eeprom.i1_2_lut_adj_27_LC_10_23_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.i1_2_lut_adj_27_LC_10_23_1 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \eeprom.i1_2_lut_adj_27_LC_10_23_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__18215),
            .in3(N__19869),
            .lcout(\eeprom.n4703 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i1_4_lut_adj_33_LC_10_23_2 .C_ON=1'b0;
    defparam \eeprom.i1_4_lut_adj_33_LC_10_23_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.i1_4_lut_adj_33_LC_10_23_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \eeprom.i1_4_lut_adj_33_LC_10_23_2  (
            .in0(N__18731),
            .in1(N__18655),
            .in2(N__20132),
            .in3(N__18717),
            .lcout(),
            .ltout(\eeprom.n4533_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i4_4_lut_adj_35_LC_10_23_3 .C_ON=1'b0;
    defparam \eeprom.i4_4_lut_adj_35_LC_10_23_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.i4_4_lut_adj_35_LC_10_23_3 .LUT_INIT=16'b1111111111100000;
    LogicCell40 \eeprom.i4_4_lut_adj_35_LC_10_23_3  (
            .in0(N__18546),
            .in1(N__18694),
            .in2(N__18668),
            .in3(N__18622),
            .lcout(),
            .ltout(\eeprom.n15_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i10_4_lut_LC_10_23_4 .C_ON=1'b0;
    defparam \eeprom.i10_4_lut_LC_10_23_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.i10_4_lut_LC_10_23_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \eeprom.i10_4_lut_LC_10_23_4  (
            .in0(N__20070),
            .in1(N__18665),
            .in2(N__18659),
            .in3(N__19669),
            .lcout(\eeprom.n2836 ),
            .ltout(\eeprom.n2836_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1903_3_lut_LC_10_23_5 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1903_3_lut_LC_10_23_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1903_3_lut_LC_10_23_5 .LUT_INIT=16'b1111101000001010;
    LogicCell40 \eeprom.rem_4_i1903_3_lut_LC_10_23_5  (
            .in0(N__18656),
            .in1(_gnd_net_),
            .in2(N__18632),
            .in3(N__18629),
            .lcout(\eeprom.n2915 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1896_3_lut_LC_10_23_6 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1896_3_lut_LC_10_23_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1896_3_lut_LC_10_23_6 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \eeprom.rem_4_i1896_3_lut_LC_10_23_6  (
            .in0(N__18623),
            .in1(_gnd_net_),
            .in2(N__18596),
            .in3(N__19934),
            .lcout(\eeprom.n2908 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1891_3_lut_LC_10_23_7 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1891_3_lut_LC_10_23_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1891_3_lut_LC_10_23_7 .LUT_INIT=16'b1111110000001100;
    LogicCell40 \eeprom.rem_4_i1891_3_lut_LC_10_23_7  (
            .in0(_gnd_net_),
            .in1(N__18586),
            .in2(N__19958),
            .in3(N__18572),
            .lcout(\eeprom.n2903 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i10_4_lut_adj_38_LC_10_24_0 .C_ON=1'b0;
    defparam \eeprom.i10_4_lut_adj_38_LC_10_24_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.i10_4_lut_adj_38_LC_10_24_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \eeprom.i10_4_lut_adj_38_LC_10_24_0  (
            .in0(N__23178),
            .in1(N__18566),
            .in2(N__22125),
            .in3(N__18875),
            .lcout(),
            .ltout(\eeprom.n22_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i11_4_lut_LC_10_24_1 .C_ON=1'b0;
    defparam \eeprom.i11_4_lut_LC_10_24_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.i11_4_lut_LC_10_24_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \eeprom.i11_4_lut_LC_10_24_1  (
            .in0(N__20022),
            .in1(N__19842),
            .in2(N__18560),
            .in3(N__20042),
            .lcout(\eeprom.n2935 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1905_3_lut_LC_10_24_2 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1905_3_lut_LC_10_24_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1905_3_lut_LC_10_24_2 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \eeprom.rem_4_i1905_3_lut_LC_10_24_2  (
            .in0(_gnd_net_),
            .in1(N__18557),
            .in2(N__18551),
            .in3(N__19948),
            .lcout(\eeprom.n2917 ),
            .ltout(\eeprom.n2917_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i1_4_lut_adj_28_LC_10_24_3 .C_ON=1'b0;
    defparam \eeprom.i1_4_lut_adj_28_LC_10_24_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.i1_4_lut_adj_28_LC_10_24_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \eeprom.i1_4_lut_adj_28_LC_10_24_3  (
            .in0(N__21831),
            .in1(N__18887),
            .in2(N__18881),
            .in3(N__22080),
            .lcout(),
            .ltout(\eeprom.n4707_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i3_4_lut_adj_36_LC_10_24_4 .C_ON=1'b0;
    defparam \eeprom.i3_4_lut_adj_36_LC_10_24_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.i3_4_lut_adj_36_LC_10_24_4 .LUT_INIT=16'b1111101011101010;
    LogicCell40 \eeprom.i3_4_lut_adj_36_LC_10_24_4  (
            .in0(N__19733),
            .in1(N__24825),
            .in2(N__18878),
            .in3(N__19483),
            .lcout(\eeprom.n15_adj_419 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1895_3_lut_LC_10_24_5 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1895_3_lut_LC_10_24_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1895_3_lut_LC_10_24_5 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \eeprom.rem_4_i1895_3_lut_LC_10_24_5  (
            .in0(_gnd_net_),
            .in1(N__18869),
            .in2(N__19965),
            .in3(N__18863),
            .lcout(\eeprom.n2907 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2245_3_lut_LC_11_17_1 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2245_3_lut_LC_11_17_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2245_3_lut_LC_11_17_1 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \eeprom.rem_4_i2245_3_lut_LC_11_17_1  (
            .in0(_gnd_net_),
            .in1(N__18805),
            .in2(N__18839),
            .in3(N__20580),
            .lcout(\eeprom.n3417 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2175_3_lut_LC_11_17_3 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2175_3_lut_LC_11_17_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2175_3_lut_LC_11_17_3 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \eeprom.rem_4_i2175_3_lut_LC_11_17_3  (
            .in0(_gnd_net_),
            .in1(N__20483),
            .in2(N__18827),
            .in3(N__19253),
            .lcout(\eeprom.n3315 ),
            .ltout(\eeprom.n3315_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i1_2_lut_adj_95_LC_11_17_4 .C_ON=1'b0;
    defparam \eeprom.i1_2_lut_adj_95_LC_11_17_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.i1_2_lut_adj_95_LC_11_17_4 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \eeprom.i1_2_lut_adj_95_LC_11_17_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__18812),
            .in3(N__20354),
            .lcout(),
            .ltout(\eeprom.n4719_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i1_4_lut_adj_97_LC_11_17_5 .C_ON=1'b0;
    defparam \eeprom.i1_4_lut_adj_97_LC_11_17_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.i1_4_lut_adj_97_LC_11_17_5 .LUT_INIT=16'b1110000000000000;
    LogicCell40 \eeprom.i1_4_lut_adj_97_LC_11_17_5  (
            .in0(N__20281),
            .in1(N__18804),
            .in2(N__18791),
            .in3(N__18788),
            .lcout(),
            .ltout(\eeprom.n4151_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i10_4_lut_adj_99_LC_11_17_6 .C_ON=1'b0;
    defparam \eeprom.i10_4_lut_adj_99_LC_11_17_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.i10_4_lut_adj_99_LC_11_17_6 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \eeprom.i10_4_lut_adj_99_LC_11_17_6  (
            .in0(N__18777),
            .in1(N__20688),
            .in2(N__18761),
            .in3(N__18758),
            .lcout(\eeprom.n26_adj_485 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2244_3_lut_LC_11_17_7 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2244_3_lut_LC_11_17_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2244_3_lut_LC_11_17_7 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \eeprom.rem_4_i2244_3_lut_LC_11_17_7  (
            .in0(_gnd_net_),
            .in1(N__19063),
            .in2(N__19043),
            .in3(N__20579),
            .lcout(\eeprom.n3416 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2235_3_lut_LC_11_18_0 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2235_3_lut_LC_11_18_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2235_3_lut_LC_11_18_0 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \eeprom.rem_4_i2235_3_lut_LC_11_18_0  (
            .in0(_gnd_net_),
            .in1(N__19031),
            .in2(N__20610),
            .in3(N__19022),
            .lcout(\eeprom.n3407 ),
            .ltout(\eeprom.n3407_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i12_4_lut_adj_108_LC_11_18_1 .C_ON=1'b0;
    defparam \eeprom.i12_4_lut_adj_108_LC_11_18_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.i12_4_lut_adj_108_LC_11_18_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \eeprom.i12_4_lut_adj_108_LC_11_18_1  (
            .in0(N__22155),
            .in1(N__22297),
            .in2(N__18998),
            .in3(N__22230),
            .lcout(\eeprom.n29_adj_491 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i11_4_lut_adj_100_LC_11_18_3 .C_ON=1'b0;
    defparam \eeprom.i11_4_lut_adj_100_LC_11_18_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.i11_4_lut_adj_100_LC_11_18_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \eeprom.i11_4_lut_adj_100_LC_11_18_3  (
            .in0(N__20386),
            .in1(N__18945),
            .in2(N__18979),
            .in3(N__20151),
            .lcout(),
            .ltout(\eeprom.n27_adj_486_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i15_4_lut_LC_11_18_4 .C_ON=1'b0;
    defparam \eeprom.i15_4_lut_LC_11_18_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.i15_4_lut_LC_11_18_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \eeprom.i15_4_lut_LC_11_18_4  (
            .in0(N__19316),
            .in1(N__18995),
            .in2(N__18989),
            .in3(N__18986),
            .lcout(\eeprom.n3331 ),
            .ltout(\eeprom.n3331_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2233_3_lut_LC_11_18_5 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2233_3_lut_LC_11_18_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2233_3_lut_LC_11_18_5 .LUT_INIT=16'b1111101000001010;
    LogicCell40 \eeprom.rem_4_i2233_3_lut_LC_11_18_5  (
            .in0(N__18975),
            .in1(_gnd_net_),
            .in2(N__18959),
            .in3(N__18956),
            .lcout(\eeprom.n3405 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2232_3_lut_LC_11_18_6 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2232_3_lut_LC_11_18_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2232_3_lut_LC_11_18_6 .LUT_INIT=16'b1111101000001010;
    LogicCell40 \eeprom.rem_4_i2232_3_lut_LC_11_18_6  (
            .in0(N__18946),
            .in1(_gnd_net_),
            .in2(N__20609),
            .in3(N__18929),
            .lcout(\eeprom.n3404 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i4038_3_lut_LC_11_18_7 .C_ON=1'b0;
    defparam \eeprom.i4038_3_lut_LC_11_18_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.i4038_3_lut_LC_11_18_7 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \eeprom.i4038_3_lut_LC_11_18_7  (
            .in0(_gnd_net_),
            .in1(N__18920),
            .in2(N__18911),
            .in3(N__20588),
            .lcout(\eeprom.n3408 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i1_4_lut_adj_89_LC_11_19_0 .C_ON=1'b0;
    defparam \eeprom.i1_4_lut_adj_89_LC_11_19_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.i1_4_lut_adj_89_LC_11_19_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \eeprom.i1_4_lut_adj_89_LC_11_19_0  (
            .in0(N__20415),
            .in1(N__20469),
            .in2(N__20796),
            .in3(N__19367),
            .lcout(),
            .ltout(\eeprom.n4615_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i6_4_lut_adj_90_LC_11_19_1 .C_ON=1'b0;
    defparam \eeprom.i6_4_lut_adj_90_LC_11_19_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.i6_4_lut_adj_90_LC_11_19_1 .LUT_INIT=16'b1111110011101100;
    LogicCell40 \eeprom.i6_4_lut_adj_90_LC_11_19_1  (
            .in0(N__19438),
            .in1(N__19131),
            .in2(N__19406),
            .in3(N__19395),
            .lcout(\eeprom.n21_adj_477 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i1_2_lut_adj_88_LC_11_19_2 .C_ON=1'b0;
    defparam \eeprom.i1_2_lut_adj_88_LC_11_19_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.i1_2_lut_adj_88_LC_11_19_2 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \eeprom.i1_2_lut_adj_88_LC_11_19_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__19512),
            .in3(N__19539),
            .lcout(\eeprom.n4611 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i9_4_lut_adj_101_LC_11_19_5 .C_ON=1'b0;
    defparam \eeprom.i9_4_lut_adj_101_LC_11_19_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.i9_4_lut_adj_101_LC_11_19_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \eeprom.i9_4_lut_adj_101_LC_11_19_5  (
            .in0(N__19353),
            .in1(N__19337),
            .in2(N__19310),
            .in3(N__20643),
            .lcout(\eeprom.n25_adj_487 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2228_3_lut_LC_11_19_6 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2228_3_lut_LC_11_19_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2228_3_lut_LC_11_19_6 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \eeprom.rem_4_i2228_3_lut_LC_11_19_6  (
            .in0(_gnd_net_),
            .in1(N__19308),
            .in2(N__19292),
            .in3(N__20595),
            .lcout(\eeprom.n3400 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2176_3_lut_LC_11_19_7 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2176_3_lut_LC_11_19_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2176_3_lut_LC_11_19_7 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \eeprom.rem_4_i2176_3_lut_LC_11_19_7  (
            .in0(_gnd_net_),
            .in1(N__19280),
            .in2(N__20425),
            .in3(N__19193),
            .lcout(\eeprom.n3316 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2102_3_lut_LC_11_20_0 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2102_3_lut_LC_11_20_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2102_3_lut_LC_11_20_0 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \eeprom.rem_4_i2102_3_lut_LC_11_20_0  (
            .in0(_gnd_net_),
            .in1(N__20888),
            .in2(N__21777),
            .in3(N__24283),
            .lcout(\eeprom.n3210 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2037_3_lut_LC_11_20_1 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2037_3_lut_LC_11_20_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2037_3_lut_LC_11_20_1 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \eeprom.rem_4_i2037_3_lut_LC_11_20_1  (
            .in0(_gnd_net_),
            .in1(N__26146),
            .in2(N__26117),
            .in3(N__27911),
            .lcout(\eeprom.n3113 ),
            .ltout(\eeprom.n3113_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2104_3_lut_LC_11_20_2 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2104_3_lut_LC_11_20_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2104_3_lut_LC_11_20_2 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \eeprom.rem_4_i2104_3_lut_LC_11_20_2  (
            .in0(N__21746),
            .in1(_gnd_net_),
            .in2(N__19115),
            .in3(N__20906),
            .lcout(\eeprom.n3212 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i10_4_lut_adj_91_LC_11_20_4 .C_ON=1'b0;
    defparam \eeprom.i10_4_lut_adj_91_LC_11_20_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.i10_4_lut_adj_91_LC_11_20_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \eeprom.i10_4_lut_adj_91_LC_11_20_4  (
            .in0(N__20437),
            .in1(N__19089),
            .in2(N__20829),
            .in3(N__21310),
            .lcout(\eeprom.n25_adj_478 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2105_3_lut_LC_11_20_5 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2105_3_lut_LC_11_20_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2105_3_lut_LC_11_20_5 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \eeprom.rem_4_i2105_3_lut_LC_11_20_5  (
            .in0(_gnd_net_),
            .in1(N__21521),
            .in2(N__20939),
            .in3(N__21741),
            .lcout(\eeprom.n3213 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2040_3_lut_LC_11_20_6 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2040_3_lut_LC_11_20_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2040_3_lut_LC_11_20_6 .LUT_INIT=16'b1111110000001100;
    LogicCell40 \eeprom.rem_4_i2040_3_lut_LC_11_20_6  (
            .in0(_gnd_net_),
            .in1(N__26283),
            .in2(N__27919),
            .in3(N__26267),
            .lcout(\eeprom.n3116 ),
            .ltout(\eeprom.n3116_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2107_3_lut_LC_11_20_7 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2107_3_lut_LC_11_20_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2107_3_lut_LC_11_20_7 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \eeprom.rem_4_i2107_3_lut_LC_11_20_7  (
            .in0(_gnd_net_),
            .in1(N__20960),
            .in2(N__19523),
            .in3(N__21742),
            .lcout(\eeprom.n3215 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1955_2_lut_LC_11_21_0 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1955_2_lut_LC_11_21_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1955_2_lut_LC_11_21_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1955_2_lut_LC_11_21_0  (
            .in0(_gnd_net_),
            .in1(N__24832),
            .in2(_gnd_net_),
            .in3(N__19487),
            .lcout(\eeprom.n2986 ),
            .ltout(),
            .carryin(bfn_11_21_0_),
            .carryout(\eeprom.n3632 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1955_3_lut_LC_11_21_1 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1955_3_lut_LC_11_21_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1955_3_lut_LC_11_21_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1955_3_lut_LC_11_21_1  (
            .in0(_gnd_net_),
            .in1(N__27325),
            .in2(N__19484),
            .in3(N__19460),
            .lcout(\eeprom.n2985 ),
            .ltout(),
            .carryin(\eeprom.n3632 ),
            .carryout(\eeprom.n3633 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1955_4_lut_LC_11_21_2 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1955_4_lut_LC_11_21_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1955_4_lut_LC_11_21_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1955_4_lut_LC_11_21_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__19805),
            .in3(N__19457),
            .lcout(\eeprom.n2984 ),
            .ltout(),
            .carryin(\eeprom.n3633 ),
            .carryout(\eeprom.n3634 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1955_5_lut_LC_11_21_3 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1955_5_lut_LC_11_21_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1955_5_lut_LC_11_21_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1955_5_lut_LC_11_21_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__21844),
            .in3(N__19454),
            .lcout(\eeprom.n2983 ),
            .ltout(),
            .carryin(\eeprom.n3634 ),
            .carryout(\eeprom.n3635 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1955_6_lut_LC_11_21_4 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1955_6_lut_LC_11_21_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1955_6_lut_LC_11_21_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1955_6_lut_LC_11_21_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__19877),
            .in3(N__19451),
            .lcout(\eeprom.n2982 ),
            .ltout(),
            .carryin(\eeprom.n3635 ),
            .carryout(\eeprom.n3636 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1955_7_lut_LC_11_21_5 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1955_7_lut_LC_11_21_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1955_7_lut_LC_11_21_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1955_7_lut_LC_11_21_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__22081),
            .in3(N__19448),
            .lcout(\eeprom.n2981 ),
            .ltout(),
            .carryin(\eeprom.n3636 ),
            .carryout(\eeprom.n3637 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1955_8_lut_LC_11_21_6 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1955_8_lut_LC_11_21_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1955_8_lut_LC_11_21_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1955_8_lut_LC_11_21_6  (
            .in0(_gnd_net_),
            .in1(N__19604),
            .in2(_gnd_net_),
            .in3(N__19577),
            .lcout(\eeprom.n2980 ),
            .ltout(),
            .carryin(\eeprom.n3637 ),
            .carryout(\eeprom.n3638 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1955_9_lut_LC_11_21_7 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1955_9_lut_LC_11_21_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1955_9_lut_LC_11_21_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1955_9_lut_LC_11_21_7  (
            .in0(_gnd_net_),
            .in1(N__27326),
            .in2(N__23188),
            .in3(N__19574),
            .lcout(\eeprom.n2979 ),
            .ltout(),
            .carryin(\eeprom.n3638 ),
            .carryout(\eeprom.n3639 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1955_10_lut_LC_11_22_0 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1955_10_lut_LC_11_22_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1955_10_lut_LC_11_22_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1955_10_lut_LC_11_22_0  (
            .in0(_gnd_net_),
            .in1(N__19843),
            .in2(N__27543),
            .in3(N__19571),
            .lcout(\eeprom.n2978 ),
            .ltout(),
            .carryin(bfn_11_22_0_),
            .carryout(\eeprom.n3640 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1955_11_lut_LC_11_22_1 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1955_11_lut_LC_11_22_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1955_11_lut_LC_11_22_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1955_11_lut_LC_11_22_1  (
            .in0(_gnd_net_),
            .in1(N__27318),
            .in2(N__21080),
            .in3(N__19568),
            .lcout(\eeprom.n2977 ),
            .ltout(),
            .carryin(\eeprom.n3640 ),
            .carryout(\eeprom.n3641 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1955_12_lut_LC_11_22_2 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1955_12_lut_LC_11_22_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1955_12_lut_LC_11_22_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1955_12_lut_LC_11_22_2  (
            .in0(_gnd_net_),
            .in1(N__27126),
            .in2(N__24797),
            .in3(N__19565),
            .lcout(\eeprom.n2976 ),
            .ltout(),
            .carryin(\eeprom.n3641 ),
            .carryout(\eeprom.n3642 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1955_13_lut_LC_11_22_3 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1955_13_lut_LC_11_22_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1955_13_lut_LC_11_22_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1955_13_lut_LC_11_22_3  (
            .in0(_gnd_net_),
            .in1(N__20023),
            .in2(N__27330),
            .in3(N__19562),
            .lcout(\eeprom.n2975 ),
            .ltout(),
            .carryin(\eeprom.n3642 ),
            .carryout(\eeprom.n3643 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1955_14_lut_LC_11_22_4 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1955_14_lut_LC_11_22_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1955_14_lut_LC_11_22_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1955_14_lut_LC_11_22_4  (
            .in0(_gnd_net_),
            .in1(N__22126),
            .in2(N__27544),
            .in3(N__19559),
            .lcout(\eeprom.n2974 ),
            .ltout(),
            .carryin(\eeprom.n3643 ),
            .carryout(\eeprom.n3644 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1955_15_lut_LC_11_22_5 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1955_15_lut_LC_11_22_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1955_15_lut_LC_11_22_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1955_15_lut_LC_11_22_5  (
            .in0(_gnd_net_),
            .in1(N__19731),
            .in2(N__27331),
            .in3(N__19556),
            .lcout(\eeprom.n2973 ),
            .ltout(),
            .carryin(\eeprom.n3644 ),
            .carryout(\eeprom.n3645 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1955_16_lut_LC_11_22_6 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1955_16_lut_LC_11_22_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1955_16_lut_LC_11_22_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1955_16_lut_LC_11_22_6  (
            .in0(_gnd_net_),
            .in1(N__21493),
            .in2(N__27545),
            .in3(N__19553),
            .lcout(\eeprom.n2972 ),
            .ltout(),
            .carryin(\eeprom.n3645 ),
            .carryout(\eeprom.n3646 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1955_17_lut_LC_11_22_7 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1955_17_lut_LC_11_22_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1955_17_lut_LC_11_22_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1955_17_lut_LC_11_22_7  (
            .in0(_gnd_net_),
            .in1(N__21106),
            .in2(N__27332),
            .in3(N__19760),
            .lcout(\eeprom.n2971 ),
            .ltout(),
            .carryin(\eeprom.n3646 ),
            .carryout(\eeprom.n3647 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1955_18_lut_LC_11_23_0 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1955_18_lut_LC_11_23_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1955_18_lut_LC_11_23_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1955_18_lut_LC_11_23_0  (
            .in0(_gnd_net_),
            .in1(N__19701),
            .in2(N__27541),
            .in3(N__19757),
            .lcout(\eeprom.n2970 ),
            .ltout(),
            .carryin(bfn_11_23_0_),
            .carryout(\eeprom.n3648 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1955_19_lut_LC_11_23_1 .C_ON=1'b0;
    defparam \eeprom.rem_4_add_1955_19_lut_LC_11_23_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1955_19_lut_LC_11_23_1 .LUT_INIT=16'b1001000001100000;
    LogicCell40 \eeprom.rem_4_add_1955_19_lut_LC_11_23_1  (
            .in0(N__19754),
            .in1(N__27310),
            .in2(N__24758),
            .in3(N__19736),
            .lcout(\eeprom.n3001 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1961_3_lut_LC_11_23_2 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1961_3_lut_LC_11_23_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1961_3_lut_LC_11_23_2 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \eeprom.rem_4_i1961_3_lut_LC_11_23_2  (
            .in0(_gnd_net_),
            .in1(N__19732),
            .in2(N__19712),
            .in3(N__24727),
            .lcout(\eeprom.n3005 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1958_3_lut_LC_11_23_3 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1958_3_lut_LC_11_23_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1958_3_lut_LC_11_23_3 .LUT_INIT=16'b1111101000001010;
    LogicCell40 \eeprom.rem_4_i1958_3_lut_LC_11_23_3  (
            .in0(N__19702),
            .in1(_gnd_net_),
            .in2(N__24757),
            .in3(N__19685),
            .lcout(\eeprom.n3002 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1899_3_lut_LC_11_23_4 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1899_3_lut_LC_11_23_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1899_3_lut_LC_11_23_4 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \eeprom.rem_4_i1899_3_lut_LC_11_23_4  (
            .in0(_gnd_net_),
            .in1(N__19679),
            .in2(N__19964),
            .in3(N__19670),
            .lcout(\eeprom.n2911 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1900_3_lut_LC_11_23_5 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1900_3_lut_LC_11_23_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1900_3_lut_LC_11_23_5 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \eeprom.rem_4_i1900_3_lut_LC_11_23_5  (
            .in0(_gnd_net_),
            .in1(N__19646),
            .in2(N__19637),
            .in3(N__19944),
            .lcout(\eeprom.n2912 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1968_3_lut_LC_11_23_6 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1968_3_lut_LC_11_23_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1968_3_lut_LC_11_23_6 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \eeprom.rem_4_i1968_3_lut_LC_11_23_6  (
            .in0(_gnd_net_),
            .in1(N__19603),
            .in2(N__19589),
            .in3(N__24728),
            .lcout(\eeprom.n3012 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1904_3_lut_LC_11_23_7 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1904_3_lut_LC_11_23_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1904_3_lut_LC_11_23_7 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \eeprom.rem_4_i1904_3_lut_LC_11_23_7  (
            .in0(N__20130),
            .in1(_gnd_net_),
            .in2(N__20096),
            .in3(N__19943),
            .lcout(\eeprom.n2916 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1897_3_lut_LC_11_24_0 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1897_3_lut_LC_11_24_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1897_3_lut_LC_11_24_0 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \eeprom.rem_4_i1897_3_lut_LC_11_24_0  (
            .in0(N__19953),
            .in1(_gnd_net_),
            .in2(N__20084),
            .in3(N__20072),
            .lcout(\eeprom.n2909 ),
            .ltout(\eeprom.n2909_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i6_2_lut_LC_11_24_1 .C_ON=1'b0;
    defparam \eeprom.i6_2_lut_LC_11_24_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.i6_2_lut_LC_11_24_1 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \eeprom.i6_2_lut_LC_11_24_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__20045),
            .in3(N__21072),
            .lcout(\eeprom.n18_adj_420 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1963_3_lut_LC_11_24_2 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1963_3_lut_LC_11_24_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1963_3_lut_LC_11_24_2 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \eeprom.rem_4_i1963_3_lut_LC_11_24_2  (
            .in0(N__24705),
            .in1(_gnd_net_),
            .in2(N__20036),
            .in3(N__20024),
            .lcout(\eeprom.n3007 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1898_3_lut_LC_11_24_3 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1898_3_lut_LC_11_24_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1898_3_lut_LC_11_24_3 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \eeprom.rem_4_i1898_3_lut_LC_11_24_3  (
            .in0(_gnd_net_),
            .in1(N__20006),
            .in2(N__19997),
            .in3(N__19952),
            .lcout(\eeprom.n2910 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1970_3_lut_LC_11_24_4 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1970_3_lut_LC_11_24_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1970_3_lut_LC_11_24_4 .LUT_INIT=16'b1111101000001010;
    LogicCell40 \eeprom.rem_4_i1970_3_lut_LC_11_24_4  (
            .in0(N__19873),
            .in1(_gnd_net_),
            .in2(N__24736),
            .in3(N__19853),
            .lcout(\eeprom.n3014 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1966_3_lut_LC_11_24_5 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1966_3_lut_LC_11_24_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1966_3_lut_LC_11_24_5 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \eeprom.rem_4_i1966_3_lut_LC_11_24_5  (
            .in0(_gnd_net_),
            .in1(N__19844),
            .in2(N__19826),
            .in3(N__24706),
            .lcout(\eeprom.n3010 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1972_3_lut_LC_11_24_7 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1972_3_lut_LC_11_24_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1972_3_lut_LC_11_24_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \eeprom.rem_4_i1972_3_lut_LC_11_24_7  (
            .in0(N__19814),
            .in1(N__19801),
            .in2(_gnd_net_),
            .in3(N__24701),
            .lcout(\eeprom.n3016 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2242_3_lut_LC_12_17_0 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2242_3_lut_LC_12_17_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2242_3_lut_LC_12_17_0 .LUT_INIT=16'b1111110000001100;
    LogicCell40 \eeprom.rem_4_i2242_3_lut_LC_12_17_0  (
            .in0(_gnd_net_),
            .in1(N__19783),
            .in2(N__20599),
            .in3(N__19769),
            .lcout(\eeprom.n3414 ),
            .ltout(\eeprom.n3414_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i1_3_lut_adj_104_LC_12_17_1 .C_ON=1'b0;
    defparam \eeprom.i1_3_lut_adj_104_LC_12_17_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.i1_3_lut_adj_104_LC_12_17_1 .LUT_INIT=16'b1100000000000000;
    LogicCell40 \eeprom.i1_3_lut_adj_104_LC_12_17_1  (
            .in0(_gnd_net_),
            .in1(N__23106),
            .in2(N__20303),
            .in3(N__23031),
            .lcout(),
            .ltout(\eeprom.n4689_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i1_4_lut_adj_105_LC_12_17_2 .C_ON=1'b0;
    defparam \eeprom.i1_4_lut_adj_105_LC_12_17_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.i1_4_lut_adj_105_LC_12_17_2 .LUT_INIT=16'b1110000000000000;
    LogicCell40 \eeprom.i1_4_lut_adj_105_LC_12_17_2  (
            .in0(N__23421),
            .in1(N__23073),
            .in2(N__20300),
            .in3(N__20177),
            .lcout(),
            .ltout(\eeprom.n4144_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i11_4_lut_adj_107_LC_12_17_3 .C_ON=1'b0;
    defparam \eeprom.i11_4_lut_adj_107_LC_12_17_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.i11_4_lut_adj_107_LC_12_17_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \eeprom.i11_4_lut_adj_107_LC_12_17_3  (
            .in0(N__23244),
            .in1(N__22674),
            .in2(N__20297),
            .in3(N__22635),
            .lcout(\eeprom.n28_adj_490 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2246_3_lut_LC_12_17_4 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2246_3_lut_LC_12_17_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2246_3_lut_LC_12_17_4 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \eeprom.rem_4_i2246_3_lut_LC_12_17_4  (
            .in0(_gnd_net_),
            .in1(N__20294),
            .in2(N__20597),
            .in3(N__20282),
            .lcout(\eeprom.n3418 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2243_3_lut_LC_12_17_5 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2243_3_lut_LC_12_17_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2243_3_lut_LC_12_17_5 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \eeprom.rem_4_i2243_3_lut_LC_12_17_5  (
            .in0(_gnd_net_),
            .in1(N__20244),
            .in2(N__20219),
            .in3(N__20557),
            .lcout(\eeprom.n3415 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2241_3_lut_LC_12_17_6 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2241_3_lut_LC_12_17_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2241_3_lut_LC_12_17_6 .LUT_INIT=16'b1111110000001100;
    LogicCell40 \eeprom.rem_4_i2241_3_lut_LC_12_17_6  (
            .in0(_gnd_net_),
            .in1(N__20207),
            .in2(N__20598),
            .in3(N__20189),
            .lcout(\eeprom.n3413 ),
            .ltout(\eeprom.n3413_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i1_2_lut_adj_103_LC_12_17_7 .C_ON=1'b0;
    defparam \eeprom.i1_2_lut_adj_103_LC_12_17_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.i1_2_lut_adj_103_LC_12_17_7 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \eeprom.i1_2_lut_adj_103_LC_12_17_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__20180),
            .in3(N__22002),
            .lcout(\eeprom.n4687 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2238_3_lut_LC_12_18_0 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2238_3_lut_LC_12_18_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2238_3_lut_LC_12_18_0 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \eeprom.rem_4_i2238_3_lut_LC_12_18_0  (
            .in0(_gnd_net_),
            .in1(N__20171),
            .in2(N__20162),
            .in3(N__20586),
            .lcout(\eeprom.n3410 ),
            .ltout(\eeprom.n3410_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2305_3_lut_LC_12_18_1 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2305_3_lut_LC_12_18_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2305_3_lut_LC_12_18_1 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \eeprom.rem_4_i2305_3_lut_LC_12_18_1  (
            .in0(_gnd_net_),
            .in1(N__22286),
            .in2(N__20399),
            .in3(N__23345),
            .lcout(\eeprom.n3509 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2373_3_lut_LC_12_18_2 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2373_3_lut_LC_12_18_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2373_3_lut_LC_12_18_2 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \eeprom.rem_4_i2373_3_lut_LC_12_18_2  (
            .in0(_gnd_net_),
            .in1(N__25013),
            .in2(N__25033),
            .in3(N__25659),
            .lcout(\eeprom.n3609_adj_445 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2301_3_lut_LC_12_18_4 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2301_3_lut_LC_12_18_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2301_3_lut_LC_12_18_4 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \eeprom.rem_4_i2301_3_lut_LC_12_18_4  (
            .in0(N__23347),
            .in1(_gnd_net_),
            .in2(N__22142),
            .in3(N__22165),
            .lcout(\eeprom.n3505 ),
            .ltout(\eeprom.n3505_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i13_4_lut_adj_117_LC_12_18_5 .C_ON=1'b0;
    defparam \eeprom.i13_4_lut_adj_117_LC_12_18_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.i13_4_lut_adj_117_LC_12_18_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \eeprom.i13_4_lut_adj_117_LC_12_18_5  (
            .in0(N__24984),
            .in1(N__25026),
            .in2(N__20396),
            .in3(N__24870),
            .lcout(\eeprom.n31_adj_496 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2237_3_lut_LC_12_18_6 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2237_3_lut_LC_12_18_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2237_3_lut_LC_12_18_6 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \eeprom.rem_4_i2237_3_lut_LC_12_18_6  (
            .in0(_gnd_net_),
            .in1(N__20393),
            .in2(N__20369),
            .in3(N__20587),
            .lcout(\eeprom.n3409 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2302_3_lut_LC_12_18_7 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2302_3_lut_LC_12_18_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2302_3_lut_LC_12_18_7 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \eeprom.rem_4_i2302_3_lut_LC_12_18_7  (
            .in0(_gnd_net_),
            .in1(N__22178),
            .in2(N__22198),
            .in3(N__23346),
            .lcout(\eeprom.n3506 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2372_3_lut_LC_12_19_1 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2372_3_lut_LC_12_19_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2372_3_lut_LC_12_19_1 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \eeprom.rem_4_i2372_3_lut_LC_12_19_1  (
            .in0(_gnd_net_),
            .in1(N__24968),
            .in2(N__24994),
            .in3(N__25678),
            .lcout(),
            .ltout(\eeprom.n3608_adj_451_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i1_4_lut_adj_54_LC_12_19_2 .C_ON=1'b0;
    defparam \eeprom.i1_4_lut_adj_54_LC_12_19_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.i1_4_lut_adj_54_LC_12_19_2 .LUT_INIT=16'b1111111011110100;
    LogicCell40 \eeprom.i1_4_lut_adj_54_LC_12_19_2  (
            .in0(N__25679),
            .in1(N__25072),
            .in2(N__20357),
            .in3(N__25052),
            .lcout(\eeprom.n4581 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2240_3_lut_LC_12_19_3 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2240_3_lut_LC_12_19_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2240_3_lut_LC_12_19_3 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \eeprom.rem_4_i2240_3_lut_LC_12_19_3  (
            .in0(_gnd_net_),
            .in1(N__20352),
            .in2(N__20321),
            .in3(N__20581),
            .lcout(\eeprom.n3412 ),
            .ltout(\eeprom.n3412_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2307_3_lut_LC_12_19_4 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2307_3_lut_LC_12_19_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2307_3_lut_LC_12_19_4 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \eeprom.rem_4_i2307_3_lut_LC_12_19_4  (
            .in0(_gnd_net_),
            .in1(N__22355),
            .in2(N__20306),
            .in3(N__23353),
            .lcout(\eeprom.n3511_adj_362 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2230_3_lut_LC_12_19_6 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2230_3_lut_LC_12_19_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2230_3_lut_LC_12_19_6 .LUT_INIT=16'b1111110000001100;
    LogicCell40 \eeprom.rem_4_i2230_3_lut_LC_12_19_6  (
            .in0(_gnd_net_),
            .in1(N__20692),
            .in2(N__20608),
            .in3(N__20666),
            .lcout(\eeprom.n3402 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2226_3_lut_LC_12_19_7 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2226_3_lut_LC_12_19_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2226_3_lut_LC_12_19_7 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \eeprom.rem_4_i2226_3_lut_LC_12_19_7  (
            .in0(_gnd_net_),
            .in1(N__20657),
            .in2(N__20648),
            .in3(N__20585),
            .lcout(\eeprom.n3398 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2296_3_lut_LC_12_20_0 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2296_3_lut_LC_12_20_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2296_3_lut_LC_12_20_0 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \eeprom.rem_4_i2296_3_lut_LC_12_20_0  (
            .in0(_gnd_net_),
            .in1(N__22544),
            .in2(N__22570),
            .in3(N__23362),
            .lcout(\eeprom.n3500 ),
            .ltout(\eeprom.n3500_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i11_4_lut_adj_118_LC_12_20_1 .C_ON=1'b0;
    defparam \eeprom.i11_4_lut_adj_118_LC_12_20_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.i11_4_lut_adj_118_LC_12_20_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \eeprom.i11_4_lut_adj_118_LC_12_20_1  (
            .in0(N__25393),
            .in1(N__25341),
            .in2(N__20486),
            .in3(N__25308),
            .lcout(\eeprom.n29_adj_497 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i10_4_lut_adj_109_LC_12_20_2 .C_ON=1'b0;
    defparam \eeprom.i10_4_lut_adj_109_LC_12_20_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.i10_4_lut_adj_109_LC_12_20_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \eeprom.i10_4_lut_adj_109_LC_12_20_2  (
            .in0(N__22563),
            .in1(N__22605),
            .in2(N__22524),
            .in3(N__22479),
            .lcout(\eeprom.n27_adj_492 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2108_3_lut_LC_12_20_3 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2108_3_lut_LC_12_20_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2108_3_lut_LC_12_20_3 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \eeprom.rem_4_i2108_3_lut_LC_12_20_3  (
            .in0(_gnd_net_),
            .in1(N__21391),
            .in2(N__20993),
            .in3(N__21772),
            .lcout(\eeprom.n3216 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2297_3_lut_LC_12_20_4 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2297_3_lut_LC_12_20_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2297_3_lut_LC_12_20_4 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \eeprom.rem_4_i2297_3_lut_LC_12_20_4  (
            .in0(_gnd_net_),
            .in1(N__22606),
            .in2(N__22592),
            .in3(N__23361),
            .lcout(\eeprom.n3501 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2095_3_lut_LC_12_20_6 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2095_3_lut_LC_12_20_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2095_3_lut_LC_12_20_6 .LUT_INIT=16'b1111101000001010;
    LogicCell40 \eeprom.rem_4_i2095_3_lut_LC_12_20_6  (
            .in0(N__21953),
            .in1(_gnd_net_),
            .in2(N__21791),
            .in3(N__21014),
            .lcout(\eeprom.n3203 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2109_3_lut_LC_12_20_7 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2109_3_lut_LC_12_20_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2109_3_lut_LC_12_20_7 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \eeprom.rem_4_i2109_3_lut_LC_12_20_7  (
            .in0(N__21458),
            .in1(_gnd_net_),
            .in2(N__20708),
            .in3(N__21771),
            .lcout(\eeprom.n3217 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i4_4_lut_adj_47_LC_12_21_0 .C_ON=1'b0;
    defparam \eeprom.i4_4_lut_adj_47_LC_12_21_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.i4_4_lut_adj_47_LC_12_21_0 .LUT_INIT=16'b1111111011001100;
    LogicCell40 \eeprom.i4_4_lut_adj_47_LC_12_21_0  (
            .in0(N__20768),
            .in1(N__21818),
            .in2(N__21454),
            .in3(N__20846),
            .lcout(),
            .ltout(\eeprom.n18_adj_432_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i12_4_lut_adj_69_LC_12_21_1 .C_ON=1'b0;
    defparam \eeprom.i12_4_lut_adj_69_LC_12_21_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.i12_4_lut_adj_69_LC_12_21_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \eeprom.i12_4_lut_adj_69_LC_12_21_1  (
            .in0(N__21952),
            .in1(N__21340),
            .in2(N__20855),
            .in3(N__22772),
            .lcout(),
            .ltout(\eeprom.n26_adj_466_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i13_4_lut_LC_12_21_2 .C_ON=1'b0;
    defparam \eeprom.i13_4_lut_LC_12_21_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.i13_4_lut_LC_12_21_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \eeprom.i13_4_lut_LC_12_21_2  (
            .in0(N__23222),
            .in1(N__21370),
            .in2(N__20852),
            .in3(N__21413),
            .lcout(\eeprom.n3133 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i1_2_lut_adj_44_LC_12_21_3 .C_ON=1'b0;
    defparam \eeprom.i1_2_lut_adj_44_LC_12_21_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.i1_2_lut_adj_44_LC_12_21_3 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \eeprom.i1_2_lut_adj_44_LC_12_21_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__21615),
            .in3(N__20917),
            .lcout(),
            .ltout(\eeprom.n4711_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i1_4_lut_adj_45_LC_12_21_4 .C_ON=1'b0;
    defparam \eeprom.i1_4_lut_adj_45_LC_12_21_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.i1_4_lut_adj_45_LC_12_21_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \eeprom.i1_4_lut_adj_45_LC_12_21_4  (
            .in0(N__21390),
            .in1(N__21510),
            .in2(N__20849),
            .in3(N__20974),
            .lcout(\eeprom.n4715 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2098_3_lut_LC_12_21_5 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2098_3_lut_LC_12_21_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2098_3_lut_LC_12_21_5 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \eeprom.rem_4_i2098_3_lut_LC_12_21_5  (
            .in0(_gnd_net_),
            .in1(N__21032),
            .in2(N__24185),
            .in3(N__21762),
            .lcout(\eeprom.n3206 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2106_3_lut_LC_12_21_7 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2106_3_lut_LC_12_21_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2106_3_lut_LC_12_21_7 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \eeprom.rem_4_i2106_3_lut_LC_12_21_7  (
            .in0(_gnd_net_),
            .in1(N__20948),
            .in2(N__21616),
            .in3(N__21761),
            .lcout(\eeprom.n3214 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2089_2_lut_LC_12_22_0 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2089_2_lut_LC_12_22_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2089_2_lut_LC_12_22_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2089_2_lut_LC_12_22_0  (
            .in0(_gnd_net_),
            .in1(N__20763),
            .in2(_gnd_net_),
            .in3(N__20711),
            .lcout(\eeprom.n3186 ),
            .ltout(),
            .carryin(bfn_12_22_0_),
            .carryout(\eeprom.n3667 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2089_3_lut_LC_12_22_1 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2089_3_lut_LC_12_22_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2089_3_lut_LC_12_22_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2089_3_lut_LC_12_22_1  (
            .in0(_gnd_net_),
            .in1(N__27311),
            .in2(N__21453),
            .in3(N__20696),
            .lcout(\eeprom.n3185 ),
            .ltout(),
            .carryin(\eeprom.n3667 ),
            .carryout(\eeprom.n3668 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2089_4_lut_LC_12_22_2 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2089_4_lut_LC_12_22_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2089_4_lut_LC_12_22_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2089_4_lut_LC_12_22_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__21392),
            .in3(N__20981),
            .lcout(\eeprom.n3184 ),
            .ltout(),
            .carryin(\eeprom.n3668 ),
            .carryout(\eeprom.n3669 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2089_5_lut_LC_12_22_3 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2089_5_lut_LC_12_22_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2089_5_lut_LC_12_22_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2089_5_lut_LC_12_22_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__20978),
            .in3(N__20951),
            .lcout(\eeprom.n3183 ),
            .ltout(),
            .carryin(\eeprom.n3669 ),
            .carryout(\eeprom.n3670 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2089_6_lut_LC_12_22_4 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2089_6_lut_LC_12_22_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2089_6_lut_LC_12_22_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2089_6_lut_LC_12_22_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__21617),
            .in3(N__20942),
            .lcout(\eeprom.n3182 ),
            .ltout(),
            .carryin(\eeprom.n3670 ),
            .carryout(\eeprom.n3671 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2089_7_lut_LC_12_22_5 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2089_7_lut_LC_12_22_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2089_7_lut_LC_12_22_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2089_7_lut_LC_12_22_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__21517),
            .in3(N__20927),
            .lcout(\eeprom.n3181 ),
            .ltout(),
            .carryin(\eeprom.n3671 ),
            .carryout(\eeprom.n3672 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2089_8_lut_LC_12_22_6 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2089_8_lut_LC_12_22_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2089_8_lut_LC_12_22_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2089_8_lut_LC_12_22_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__20924),
            .in3(N__20894),
            .lcout(\eeprom.n3180 ),
            .ltout(),
            .carryin(\eeprom.n3672 ),
            .carryout(\eeprom.n3673 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2089_9_lut_LC_12_22_7 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2089_9_lut_LC_12_22_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2089_9_lut_LC_12_22_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2089_9_lut_LC_12_22_7  (
            .in0(_gnd_net_),
            .in1(N__23220),
            .in2(N__27542),
            .in3(N__20891),
            .lcout(\eeprom.n3179 ),
            .ltout(),
            .carryin(\eeprom.n3673 ),
            .carryout(\eeprom.n3674 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2089_10_lut_LC_12_23_0 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2089_10_lut_LC_12_23_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2089_10_lut_LC_12_23_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2089_10_lut_LC_12_23_0  (
            .in0(_gnd_net_),
            .in1(N__27080),
            .in2(N__24284),
            .in3(N__20876),
            .lcout(\eeprom.n3178 ),
            .ltout(),
            .carryin(bfn_12_23_0_),
            .carryout(\eeprom.n3675 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2089_11_lut_LC_12_23_1 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2089_11_lut_LC_12_23_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2089_11_lut_LC_12_23_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2089_11_lut_LC_12_23_1  (
            .in0(_gnd_net_),
            .in1(N__24208),
            .in2(N__27302),
            .in3(N__20858),
            .lcout(\eeprom.n3177 ),
            .ltout(),
            .carryin(\eeprom.n3675 ),
            .carryout(\eeprom.n3676 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2089_12_lut_LC_12_23_2 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2089_12_lut_LC_12_23_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2089_12_lut_LC_12_23_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2089_12_lut_LC_12_23_2  (
            .in0(_gnd_net_),
            .in1(N__27084),
            .in2(N__24244),
            .in3(N__21038),
            .lcout(\eeprom.n3176 ),
            .ltout(),
            .carryin(\eeprom.n3676 ),
            .carryout(\eeprom.n3677 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2089_13_lut_LC_12_23_3 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2089_13_lut_LC_12_23_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2089_13_lut_LC_12_23_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2089_13_lut_LC_12_23_3  (
            .in0(_gnd_net_),
            .in1(N__21371),
            .in2(N__27303),
            .in3(N__21035),
            .lcout(\eeprom.n3175 ),
            .ltout(),
            .carryin(\eeprom.n3677 ),
            .carryout(\eeprom.n3678 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2089_14_lut_LC_12_23_4 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2089_14_lut_LC_12_23_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2089_14_lut_LC_12_23_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2089_14_lut_LC_12_23_4  (
            .in0(_gnd_net_),
            .in1(N__24178),
            .in2(N__27306),
            .in3(N__21023),
            .lcout(\eeprom.n3174 ),
            .ltout(),
            .carryin(\eeprom.n3678 ),
            .carryout(\eeprom.n3679 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2089_15_lut_LC_12_23_5 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2089_15_lut_LC_12_23_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2089_15_lut_LC_12_23_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2089_15_lut_LC_12_23_5  (
            .in0(_gnd_net_),
            .in1(N__21817),
            .in2(N__27304),
            .in3(N__21020),
            .lcout(\eeprom.n3173 ),
            .ltout(),
            .carryin(\eeprom.n3679 ),
            .carryout(\eeprom.n3680 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2089_16_lut_LC_12_23_6 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2089_16_lut_LC_12_23_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2089_16_lut_LC_12_23_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2089_16_lut_LC_12_23_6  (
            .in0(_gnd_net_),
            .in1(N__27091),
            .in2(N__21344),
            .in3(N__21017),
            .lcout(\eeprom.n3172 ),
            .ltout(),
            .carryin(\eeprom.n3680 ),
            .carryout(\eeprom.n3681 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2089_17_lut_LC_12_23_7 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2089_17_lut_LC_12_23_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2089_17_lut_LC_12_23_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2089_17_lut_LC_12_23_7  (
            .in0(_gnd_net_),
            .in1(N__21951),
            .in2(N__27305),
            .in3(N__21005),
            .lcout(\eeprom.n3171 ),
            .ltout(),
            .carryin(\eeprom.n3681 ),
            .carryout(\eeprom.n3682 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2089_18_lut_LC_12_24_0 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2089_18_lut_LC_12_24_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2089_18_lut_LC_12_24_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2089_18_lut_LC_12_24_0  (
            .in0(_gnd_net_),
            .in1(N__23144),
            .in2(N__27384),
            .in3(N__21002),
            .lcout(\eeprom.n3170 ),
            .ltout(),
            .carryin(bfn_12_24_0_),
            .carryout(\eeprom.n3683 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2089_19_lut_LC_12_24_1 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2089_19_lut_LC_12_24_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2089_19_lut_LC_12_24_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2089_19_lut_LC_12_24_1  (
            .in0(_gnd_net_),
            .in1(N__21427),
            .in2(N__27386),
            .in3(N__20999),
            .lcout(\eeprom.n3169 ),
            .ltout(),
            .carryin(\eeprom.n3683 ),
            .carryout(\eeprom.n3684 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2089_20_lut_LC_12_24_2 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2089_20_lut_LC_12_24_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2089_20_lut_LC_12_24_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2089_20_lut_LC_12_24_2  (
            .in0(_gnd_net_),
            .in1(N__22042),
            .in2(N__27385),
            .in3(N__20996),
            .lcout(\eeprom.n3168 ),
            .ltout(),
            .carryin(\eeprom.n3684 ),
            .carryout(\eeprom.n3685 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2089_21_lut_LC_12_24_3 .C_ON=1'b0;
    defparam \eeprom.rem_4_add_2089_21_lut_LC_12_24_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2089_21_lut_LC_12_24_3 .LUT_INIT=16'b1001000001100000;
    LogicCell40 \eeprom.rem_4_add_2089_21_lut_LC_12_24_3  (
            .in0(N__27205),
            .in1(N__27806),
            .in2(N__21792),
            .in3(N__21125),
            .lcout(\eeprom.n3199 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1959_3_lut_LC_12_24_5 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1959_3_lut_LC_12_24_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1959_3_lut_LC_12_24_5 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \eeprom.rem_4_i1959_3_lut_LC_12_24_5  (
            .in0(_gnd_net_),
            .in1(N__21122),
            .in2(N__21113),
            .in3(N__24753),
            .lcout(\eeprom.n3003 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1965_3_lut_LC_12_24_6 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1965_3_lut_LC_12_24_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1965_3_lut_LC_12_24_6 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \eeprom.rem_4_i1965_3_lut_LC_12_24_6  (
            .in0(N__21089),
            .in1(_gnd_net_),
            .in2(N__24764),
            .in3(N__21076),
            .lcout(\eeprom.n3009 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2309_3_lut_LC_13_17_0 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2309_3_lut_LC_13_17_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2309_3_lut_LC_13_17_0 .LUT_INIT=16'b1111110000001100;
    LogicCell40 \eeprom.rem_4_i2309_3_lut_LC_13_17_0  (
            .in0(_gnd_net_),
            .in1(N__21976),
            .in2(N__23363),
            .in3(N__21962),
            .lcout(\eeprom.n3513_adj_366 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2310_3_lut_LC_13_17_1 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2310_3_lut_LC_13_17_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2310_3_lut_LC_13_17_1 .LUT_INIT=16'b1010101011110000;
    LogicCell40 \eeprom.rem_4_i2310_3_lut_LC_13_17_1  (
            .in0(N__21986),
            .in1(_gnd_net_),
            .in2(N__22012),
            .in3(N__23324),
            .lcout(\eeprom.n3514_adj_368 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2308_3_lut_LC_13_17_3 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2308_3_lut_LC_13_17_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2308_3_lut_LC_13_17_3 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \eeprom.rem_4_i2308_3_lut_LC_13_17_3  (
            .in0(_gnd_net_),
            .in1(N__22385),
            .in2(N__22406),
            .in3(N__23331),
            .lcout(\eeprom.n3512_adj_364 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2294_3_lut_LC_13_17_4 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2294_3_lut_LC_13_17_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2294_3_lut_LC_13_17_4 .LUT_INIT=16'b1111110000001100;
    LogicCell40 \eeprom.rem_4_i2294_3_lut_LC_13_17_4  (
            .in0(_gnd_net_),
            .in1(N__22489),
            .in2(N__23364),
            .in3(N__22457),
            .lcout(\eeprom.n3498 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2293_3_lut_LC_13_17_5 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2293_3_lut_LC_13_17_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2293_3_lut_LC_13_17_5 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \eeprom.rem_4_i2293_3_lut_LC_13_17_5  (
            .in0(_gnd_net_),
            .in1(N__22445),
            .in2(N__22418),
            .in3(N__23332),
            .lcout(\eeprom.n3497 ),
            .ltout(\eeprom.n3497_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i10_4_lut_adj_110_LC_13_17_6 .C_ON=1'b0;
    defparam \eeprom.i10_4_lut_adj_110_LC_13_17_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.i10_4_lut_adj_110_LC_13_17_6 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \eeprom.i10_4_lut_adj_110_LC_13_17_6  (
            .in0(N__25723),
            .in1(N__25240),
            .in2(N__21056),
            .in3(N__25186),
            .lcout(),
            .ltout(\eeprom.n28_adj_493_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i14_3_lut_LC_13_17_7 .C_ON=1'b0;
    defparam \eeprom.i14_3_lut_LC_13_17_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.i14_3_lut_LC_13_17_7 .LUT_INIT=16'b1111111111111100;
    LogicCell40 \eeprom.i14_3_lut_LC_13_17_7  (
            .in0(_gnd_net_),
            .in1(N__24946),
            .in2(N__21170),
            .in3(N__25113),
            .lcout(\eeprom.n32_adj_494 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i4039_3_lut_LC_13_18_0 .C_ON=1'b0;
    defparam \eeprom.i4039_3_lut_LC_13_18_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.i4039_3_lut_LC_13_18_0 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \eeprom.i4039_3_lut_LC_13_18_0  (
            .in0(_gnd_net_),
            .in1(N__22240),
            .in2(N__22214),
            .in3(N__23352),
            .lcout(\eeprom.n3507 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2300_3_lut_LC_13_18_1 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2300_3_lut_LC_13_18_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2300_3_lut_LC_13_18_1 .LUT_INIT=16'b1111110000001100;
    LogicCell40 \eeprom.rem_4_i2300_3_lut_LC_13_18_1  (
            .in0(_gnd_net_),
            .in1(N__22684),
            .in2(N__23371),
            .in3(N__22661),
            .lcout(\eeprom.n3504 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2306_3_lut_LC_13_18_2 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2306_3_lut_LC_13_18_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2306_3_lut_LC_13_18_2 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \eeprom.rem_4_i2306_3_lut_LC_13_18_2  (
            .in0(_gnd_net_),
            .in1(N__22339),
            .in2(N__22316),
            .in3(N__23348),
            .lcout(\eeprom.n3510_adj_360 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i1_2_lut_adj_102_LC_13_18_3 .C_ON=1'b0;
    defparam \eeprom.i1_2_lut_adj_102_LC_13_18_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.i1_2_lut_adj_102_LC_13_18_3 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \eeprom.i1_2_lut_adj_102_LC_13_18_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__22443),
            .in3(N__22732),
            .lcout(),
            .ltout(\eeprom.n18_adj_488_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i13_4_lut_adj_106_LC_13_18_4 .C_ON=1'b0;
    defparam \eeprom.i13_4_lut_adj_106_LC_13_18_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.i13_4_lut_adj_106_LC_13_18_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \eeprom.i13_4_lut_adj_106_LC_13_18_4  (
            .in0(N__22338),
            .in1(N__22369),
            .in2(N__21167),
            .in3(N__22269),
            .lcout(),
            .ltout(\eeprom.n30_adj_489_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i16_4_lut_LC_13_18_5 .C_ON=1'b0;
    defparam \eeprom.i16_4_lut_LC_13_18_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.i16_4_lut_LC_13_18_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \eeprom.i16_4_lut_LC_13_18_5  (
            .in0(N__21164),
            .in1(N__21155),
            .in2(N__21149),
            .in3(N__21146),
            .lcout(\eeprom.n3430 ),
            .ltout(\eeprom.n3430_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2304_3_lut_LC_13_18_6 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2304_3_lut_LC_13_18_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2304_3_lut_LC_13_18_6 .LUT_INIT=16'b1111110000001100;
    LogicCell40 \eeprom.rem_4_i2304_3_lut_LC_13_18_6  (
            .in0(_gnd_net_),
            .in1(N__22270),
            .in2(N__21137),
            .in3(N__22253),
            .lcout(\eeprom.n3508 ),
            .ltout(\eeprom.n3508_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i1_4_lut_adj_52_LC_13_18_7 .C_ON=1'b0;
    defparam \eeprom.i1_4_lut_adj_52_LC_13_18_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.i1_4_lut_adj_52_LC_13_18_7 .LUT_INIT=16'b1110111011111010;
    LogicCell40 \eeprom.i1_4_lut_adj_52_LC_13_18_7  (
            .in0(N__21134),
            .in1(N__24935),
            .in2(N__21128),
            .in3(N__25660),
            .lcout(\eeprom.n4429 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2298_3_lut_LC_13_19_0 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2298_3_lut_LC_13_19_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2298_3_lut_LC_13_19_0 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \eeprom.rem_4_i2298_3_lut_LC_13_19_0  (
            .in0(_gnd_net_),
            .in1(N__22619),
            .in2(N__23370),
            .in3(N__22645),
            .lcout(\eeprom.n3502 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i12_4_lut_adj_116_LC_13_19_1 .C_ON=1'b0;
    defparam \eeprom.i12_4_lut_adj_116_LC_13_19_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.i12_4_lut_adj_116_LC_13_19_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \eeprom.i12_4_lut_adj_116_LC_13_19_1  (
            .in0(N__25425),
            .in1(N__25071),
            .in2(N__24922),
            .in3(N__23126),
            .lcout(),
            .ltout(\eeprom.n30_adj_495_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i17_4_lut_LC_13_19_2 .C_ON=1'b0;
    defparam \eeprom.i17_4_lut_LC_13_19_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.i17_4_lut_LC_13_19_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \eeprom.i17_4_lut_LC_13_19_2  (
            .in0(N__21233),
            .in1(N__21227),
            .in2(N__21221),
            .in3(N__21218),
            .lcout(\eeprom.n3529_adj_336 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2295_3_lut_LC_13_19_3 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2295_3_lut_LC_13_19_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2295_3_lut_LC_13_19_3 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \eeprom.rem_4_i2295_3_lut_LC_13_19_3  (
            .in0(_gnd_net_),
            .in1(N__22528),
            .in2(N__22502),
            .in3(N__23341),
            .lcout(\eeprom.n3499 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2370_3_lut_LC_13_19_4 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2370_3_lut_LC_13_19_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2370_3_lut_LC_13_19_4 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \eeprom.rem_4_i2370_3_lut_LC_13_19_4  (
            .in0(_gnd_net_),
            .in1(N__24918),
            .in2(N__24902),
            .in3(N__25680),
            .lcout(),
            .ltout(\eeprom.n3606_adj_446_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i1_4_lut_adj_51_LC_13_19_5 .C_ON=1'b0;
    defparam \eeprom.i1_4_lut_adj_51_LC_13_19_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.i1_4_lut_adj_51_LC_13_19_5 .LUT_INIT=16'b1111110111111000;
    LogicCell40 \eeprom.i1_4_lut_adj_51_LC_13_19_5  (
            .in0(N__25681),
            .in1(N__25409),
            .in2(N__21209),
            .in3(N__25429),
            .lcout(),
            .ltout(\eeprom.n4451_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i1_4_lut_adj_53_LC_13_19_6 .C_ON=1'b0;
    defparam \eeprom.i1_4_lut_adj_53_LC_13_19_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.i1_4_lut_adj_53_LC_13_19_6 .LUT_INIT=16'b1111101011111100;
    LogicCell40 \eeprom.i1_4_lut_adj_53_LC_13_19_6  (
            .in0(N__25361),
            .in1(N__25394),
            .in2(N__21206),
            .in3(N__25682),
            .lcout(\eeprom.n4453 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2363_3_lut_LC_13_20_0 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2363_3_lut_LC_13_20_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2363_3_lut_LC_13_20_0 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \eeprom.rem_4_i2363_3_lut_LC_13_20_0  (
            .in0(_gnd_net_),
            .in1(N__25256),
            .in2(N__25276),
            .in3(N__25632),
            .lcout(),
            .ltout(\eeprom.n3599_adj_450_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i1_4_lut_adj_57_LC_13_20_1 .C_ON=1'b0;
    defparam \eeprom.i1_4_lut_adj_57_LC_13_20_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.i1_4_lut_adj_57_LC_13_20_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \eeprom.i1_4_lut_adj_57_LC_13_20_1  (
            .in0(N__21404),
            .in1(N__21203),
            .in2(N__21197),
            .in3(N__21194),
            .lcout(\eeprom.n4433 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_mux_3_i5_3_lut_LC_13_20_2 .C_ON=1'b0;
    defparam \eeprom.rem_4_mux_3_i5_3_lut_LC_13_20_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_mux_3_i5_3_lut_LC_13_20_2 .LUT_INIT=16'b0010001001110111;
    LogicCell40 \eeprom.rem_4_mux_3_i5_3_lut_LC_13_20_2  (
            .in0(N__22977),
            .in1(N__21185),
            .in2(_gnd_net_),
            .in3(N__23722),
            .lcout(\eeprom.n3721_adj_434 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2364_3_lut_LC_13_20_3 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2364_3_lut_LC_13_20_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2364_3_lut_LC_13_20_3 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \eeprom.rem_4_i2364_3_lut_LC_13_20_3  (
            .in0(_gnd_net_),
            .in1(N__25292),
            .in2(N__25672),
            .in3(N__25312),
            .lcout(\eeprom.n3600_adj_449 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2377_3_lut_LC_13_20_4 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2377_3_lut_LC_13_20_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2377_3_lut_LC_13_20_4 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \eeprom.rem_4_i2377_3_lut_LC_13_20_4  (
            .in0(_gnd_net_),
            .in1(N__24487),
            .in2(N__24461),
            .in3(N__25628),
            .lcout(\eeprom.n3613_adj_342 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i1_4_lut_adj_55_LC_13_20_6 .C_ON=1'b0;
    defparam \eeprom.i1_4_lut_adj_55_LC_13_20_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.i1_4_lut_adj_55_LC_13_20_6 .LUT_INIT=16'b1111101011101110;
    LogicCell40 \eeprom.i1_4_lut_adj_55_LC_13_20_6  (
            .in0(N__21398),
            .in1(N__25123),
            .in2(N__25097),
            .in3(N__25633),
            .lcout(\eeprom.n4583 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2041_3_lut_LC_13_21_0 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2041_3_lut_LC_13_21_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2041_3_lut_LC_13_21_0 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \eeprom.rem_4_i2041_3_lut_LC_13_21_0  (
            .in0(_gnd_net_),
            .in1(N__26312),
            .in2(N__27915),
            .in3(N__26339),
            .lcout(\eeprom.n3117 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2032_3_lut_LC_13_21_1 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2032_3_lut_LC_13_21_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2032_3_lut_LC_13_21_1 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \eeprom.rem_4_i2032_3_lut_LC_13_21_1  (
            .in0(_gnd_net_),
            .in1(N__26594),
            .in2(N__26561),
            .in3(N__27902),
            .lcout(\eeprom.n3108 ),
            .ltout(\eeprom.n3108_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2099_3_lut_LC_13_21_2 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2099_3_lut_LC_13_21_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2099_3_lut_LC_13_21_2 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \eeprom.rem_4_i2099_3_lut_LC_13_21_2  (
            .in0(_gnd_net_),
            .in1(N__21356),
            .in2(N__21347),
            .in3(N__21764),
            .lcout(\eeprom.n3207 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2029_3_lut_LC_13_21_3 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2029_3_lut_LC_13_21_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2029_3_lut_LC_13_21_3 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \eeprom.rem_4_i2029_3_lut_LC_13_21_3  (
            .in0(_gnd_net_),
            .in1(N__26468),
            .in2(N__26444),
            .in3(N__27903),
            .lcout(\eeprom.n3105 ),
            .ltout(\eeprom.n3105_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2096_3_lut_LC_13_21_4 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2096_3_lut_LC_13_21_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2096_3_lut_LC_13_21_4 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \eeprom.rem_4_i2096_3_lut_LC_13_21_4  (
            .in0(_gnd_net_),
            .in1(N__21326),
            .in2(N__21314),
            .in3(N__21763),
            .lcout(\eeprom.n3204 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2103_3_lut_LC_13_21_6 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2103_3_lut_LC_13_21_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2103_3_lut_LC_13_21_6 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \eeprom.rem_4_i2103_3_lut_LC_13_21_6  (
            .in0(_gnd_net_),
            .in1(N__23221),
            .in2(N__21278),
            .in3(N__21765),
            .lcout(\eeprom.n3211 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2039_3_lut_LC_13_22_0 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2039_3_lut_LC_13_22_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2039_3_lut_LC_13_22_0 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \eeprom.rem_4_i2039_3_lut_LC_13_22_0  (
            .in0(_gnd_net_),
            .in1(N__27874),
            .in2(N__26213),
            .in3(N__26245),
            .lcout(\eeprom.n3115 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2093_3_lut_LC_13_22_1 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2093_3_lut_LC_13_22_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2093_3_lut_LC_13_22_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \eeprom.rem_4_i2093_3_lut_LC_13_22_1  (
            .in0(N__21593),
            .in1(N__21428),
            .in2(_gnd_net_),
            .in3(N__21776),
            .lcout(\eeprom.n3201 ),
            .ltout(\eeprom.n3201_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i9_4_lut_adj_93_LC_13_22_2 .C_ON=1'b0;
    defparam \eeprom.i9_4_lut_adj_93_LC_13_22_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.i9_4_lut_adj_93_LC_13_22_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \eeprom.i9_4_lut_adj_93_LC_13_22_2  (
            .in0(N__21876),
            .in1(N__21552),
            .in2(N__21536),
            .in3(N__21912),
            .lcout(\eeprom.n24_adj_481 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2038_3_lut_LC_13_22_3 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2038_3_lut_LC_13_22_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2038_3_lut_LC_13_22_3 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \eeprom.rem_4_i2038_3_lut_LC_13_22_3  (
            .in0(N__26165),
            .in1(_gnd_net_),
            .in2(N__27908),
            .in3(N__26191),
            .lcout(\eeprom.n3114 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1960_3_lut_LC_13_22_5 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1960_3_lut_LC_13_22_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1960_3_lut_LC_13_22_5 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \eeprom.rem_4_i1960_3_lut_LC_13_22_5  (
            .in0(_gnd_net_),
            .in1(N__21494),
            .in2(N__21470),
            .in3(N__24763),
            .lcout(\eeprom.n3004 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2042_3_lut_LC_13_22_7 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2042_3_lut_LC_13_22_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2042_3_lut_LC_13_22_7 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \eeprom.rem_4_i2042_3_lut_LC_13_22_7  (
            .in0(_gnd_net_),
            .in1(N__26354),
            .in2(N__27907),
            .in3(N__26390),
            .lcout(\eeprom.n3118 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i8_4_lut_adj_42_LC_13_23_0 .C_ON=1'b0;
    defparam \eeprom.i8_4_lut_adj_42_LC_13_23_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.i8_4_lut_adj_42_LC_13_23_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \eeprom.i8_4_lut_adj_42_LC_13_23_0  (
            .in0(N__26418),
            .in1(N__26460),
            .in2(N__28030),
            .in3(N__28062),
            .lcout(\eeprom.n21_adj_422 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2026_3_lut_LC_13_23_1 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2026_3_lut_LC_13_23_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2026_3_lut_LC_13_23_1 .LUT_INIT=16'b1111110000001100;
    LogicCell40 \eeprom.rem_4_i2026_3_lut_LC_13_23_1  (
            .in0(_gnd_net_),
            .in1(N__28026),
            .in2(N__27910),
            .in3(N__28010),
            .lcout(\eeprom.n3102 ),
            .ltout(\eeprom.n3102_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i8_4_lut_adj_67_LC_13_23_2 .C_ON=1'b0;
    defparam \eeprom.i8_4_lut_adj_67_LC_13_23_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.i8_4_lut_adj_67_LC_13_23_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \eeprom.i8_4_lut_adj_67_LC_13_23_2  (
            .in0(N__27805),
            .in1(N__23139),
            .in2(N__21416),
            .in3(N__22038),
            .lcout(\eeprom.n22_adj_465 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2028_3_lut_LC_13_23_4 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2028_3_lut_LC_13_23_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2028_3_lut_LC_13_23_4 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \eeprom.rem_4_i2028_3_lut_LC_13_23_4  (
            .in0(N__26419),
            .in1(_gnd_net_),
            .in2(N__28091),
            .in3(N__27890),
            .lcout(\eeprom.n3104 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i7_3_lut_LC_13_23_5 .C_ON=1'b0;
    defparam \eeprom.i7_3_lut_LC_13_23_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.i7_3_lut_LC_13_23_5 .LUT_INIT=16'b1111111111111010;
    LogicCell40 \eeprom.i7_3_lut_LC_13_23_5  (
            .in0(N__26703),
            .in1(_gnd_net_),
            .in2(N__27943),
            .in3(N__27987),
            .lcout(\eeprom.n20_adj_423 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2094_3_lut_LC_13_23_6 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2094_3_lut_LC_13_23_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2094_3_lut_LC_13_23_6 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \eeprom.rem_4_i2094_3_lut_LC_13_23_6  (
            .in0(_gnd_net_),
            .in1(N__21932),
            .in2(N__21794),
            .in3(N__23140),
            .lcout(\eeprom.n3202 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2092_3_lut_LC_13_23_7 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2092_3_lut_LC_13_23_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2092_3_lut_LC_13_23_7 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \eeprom.rem_4_i2092_3_lut_LC_13_23_7  (
            .in0(_gnd_net_),
            .in1(N__21896),
            .in2(N__22043),
            .in3(N__21784),
            .lcout(\eeprom.n3200 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1971_3_lut_LC_13_24_0 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1971_3_lut_LC_13_24_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1971_3_lut_LC_13_24_0 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \eeprom.rem_4_i1971_3_lut_LC_13_24_0  (
            .in0(_gnd_net_),
            .in1(N__21860),
            .in2(N__21848),
            .in3(N__24737),
            .lcout(\eeprom.n3015 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2030_3_lut_LC_13_24_1 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2030_3_lut_LC_13_24_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2030_3_lut_LC_13_24_1 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \eeprom.rem_4_i2030_3_lut_LC_13_24_1  (
            .in0(N__27889),
            .in1(_gnd_net_),
            .in2(N__26483),
            .in3(N__26512),
            .lcout(\eeprom.n3106 ),
            .ltout(\eeprom.n3106_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2097_3_lut_LC_13_24_2 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2097_3_lut_LC_13_24_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2097_3_lut_LC_13_24_2 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \eeprom.rem_4_i2097_3_lut_LC_13_24_2  (
            .in0(_gnd_net_),
            .in1(N__21803),
            .in2(N__21797),
            .in3(N__21788),
            .lcout(\eeprom.n3205 ),
            .ltout(\eeprom.n3205_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i1_2_lut_adj_92_LC_13_24_3 .C_ON=1'b0;
    defparam \eeprom.i1_2_lut_adj_92_LC_13_24_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.i1_2_lut_adj_92_LC_13_24_3 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \eeprom.i1_2_lut_adj_92_LC_13_24_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__21653),
            .in3(N__21643),
            .lcout(\eeprom.n16_adj_479 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1962_3_lut_LC_13_24_4 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1962_3_lut_LC_13_24_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1962_3_lut_LC_13_24_4 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \eeprom.rem_4_i1962_3_lut_LC_13_24_4  (
            .in0(_gnd_net_),
            .in1(N__22127),
            .in2(N__22100),
            .in3(N__24741),
            .lcout(\eeprom.n3006 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1969_3_lut_LC_13_24_5 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1969_3_lut_LC_13_24_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1969_3_lut_LC_13_24_5 .LUT_INIT=16'b1111110000001100;
    LogicCell40 \eeprom.rem_4_i1969_3_lut_LC_13_24_5  (
            .in0(_gnd_net_),
            .in1(N__22085),
            .in2(N__24759),
            .in3(N__22055),
            .lcout(\eeprom.n3013 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2025_3_lut_LC_13_24_6 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2025_3_lut_LC_13_24_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2025_3_lut_LC_13_24_6 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \eeprom.rem_4_i2025_3_lut_LC_13_24_6  (
            .in0(_gnd_net_),
            .in1(N__27994),
            .in2(N__27965),
            .in3(N__27888),
            .lcout(\eeprom.n3101 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2290_2_lut_LC_14_17_0 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2290_2_lut_LC_14_17_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2290_2_lut_LC_14_17_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2290_2_lut_LC_14_17_0  (
            .in0(_gnd_net_),
            .in1(N__23425),
            .in2(_gnd_net_),
            .in3(N__22025),
            .lcout(\eeprom.n3486 ),
            .ltout(),
            .carryin(bfn_14_17_0_),
            .carryout(\eeprom.n3727 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2290_3_lut_LC_14_17_1 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2290_3_lut_LC_14_17_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2290_3_lut_LC_14_17_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2290_3_lut_LC_14_17_1  (
            .in0(_gnd_net_),
            .in1(N__27781),
            .in2(N__23078),
            .in3(N__22022),
            .lcout(\eeprom.n3485 ),
            .ltout(),
            .carryin(\eeprom.n3727 ),
            .carryout(\eeprom.n3728 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2290_4_lut_LC_14_17_2 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2290_4_lut_LC_14_17_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2290_4_lut_LC_14_17_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2290_4_lut_LC_14_17_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__23113),
            .in3(N__22019),
            .lcout(\eeprom.n3484_adj_406 ),
            .ltout(),
            .carryin(\eeprom.n3728 ),
            .carryout(\eeprom.n3729 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2290_5_lut_LC_14_17_3 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2290_5_lut_LC_14_17_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2290_5_lut_LC_14_17_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2290_5_lut_LC_14_17_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__23036),
            .in3(N__22016),
            .lcout(\eeprom.n3483_adj_404 ),
            .ltout(),
            .carryin(\eeprom.n3729 ),
            .carryout(\eeprom.n3730 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2290_6_lut_LC_14_17_4 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2290_6_lut_LC_14_17_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2290_6_lut_LC_14_17_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2290_6_lut_LC_14_17_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__22013),
            .in3(N__21980),
            .lcout(\eeprom.n3482_adj_401 ),
            .ltout(),
            .carryin(\eeprom.n3730 ),
            .carryout(\eeprom.n3731 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2290_7_lut_LC_14_17_5 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2290_7_lut_LC_14_17_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2290_7_lut_LC_14_17_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2290_7_lut_LC_14_17_5  (
            .in0(_gnd_net_),
            .in1(N__21977),
            .in2(_gnd_net_),
            .in3(N__21956),
            .lcout(\eeprom.n3481_adj_399 ),
            .ltout(),
            .carryin(\eeprom.n3731 ),
            .carryout(\eeprom.n3732 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2290_8_lut_LC_14_17_6 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2290_8_lut_LC_14_17_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2290_8_lut_LC_14_17_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2290_8_lut_LC_14_17_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__22405),
            .in3(N__22379),
            .lcout(\eeprom.n3480_adj_398 ),
            .ltout(),
            .carryin(\eeprom.n3732 ),
            .carryout(\eeprom.n3733 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2290_9_lut_LC_14_17_7 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2290_9_lut_LC_14_17_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2290_9_lut_LC_14_17_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2290_9_lut_LC_14_17_7  (
            .in0(_gnd_net_),
            .in1(N__27782),
            .in2(N__22376),
            .in3(N__22343),
            .lcout(\eeprom.n3479_adj_394 ),
            .ltout(),
            .carryin(\eeprom.n3733 ),
            .carryout(\eeprom.n3734 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2290_10_lut_LC_14_18_0 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2290_10_lut_LC_14_18_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2290_10_lut_LC_14_18_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2290_10_lut_LC_14_18_0  (
            .in0(_gnd_net_),
            .in1(N__27708),
            .in2(N__22340),
            .in3(N__22307),
            .lcout(\eeprom.n3478_adj_393 ),
            .ltout(),
            .carryin(bfn_14_18_0_),
            .carryout(\eeprom.n3735 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2290_11_lut_LC_14_18_1 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2290_11_lut_LC_14_18_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2290_11_lut_LC_14_18_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2290_11_lut_LC_14_18_1  (
            .in0(_gnd_net_),
            .in1(N__27712),
            .in2(N__22304),
            .in3(N__22277),
            .lcout(\eeprom.n3477_adj_392 ),
            .ltout(),
            .carryin(\eeprom.n3735 ),
            .carryout(\eeprom.n3736 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2290_12_lut_LC_14_18_2 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2290_12_lut_LC_14_18_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2290_12_lut_LC_14_18_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2290_12_lut_LC_14_18_2  (
            .in0(_gnd_net_),
            .in1(N__27709),
            .in2(N__22274),
            .in3(N__22244),
            .lcout(\eeprom.n3476_adj_391 ),
            .ltout(),
            .carryin(\eeprom.n3736 ),
            .carryout(\eeprom.n3737 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2290_13_lut_LC_14_18_3 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2290_13_lut_LC_14_18_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2290_13_lut_LC_14_18_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2290_13_lut_LC_14_18_3  (
            .in0(_gnd_net_),
            .in1(N__27713),
            .in2(N__22241),
            .in3(N__22202),
            .lcout(\eeprom.n3475_adj_390 ),
            .ltout(),
            .carryin(\eeprom.n3737 ),
            .carryout(\eeprom.n3738 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2290_14_lut_LC_14_18_4 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2290_14_lut_LC_14_18_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2290_14_lut_LC_14_18_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2290_14_lut_LC_14_18_4  (
            .in0(_gnd_net_),
            .in1(N__27710),
            .in2(N__22199),
            .in3(N__22169),
            .lcout(\eeprom.n3474_adj_389 ),
            .ltout(),
            .carryin(\eeprom.n3738 ),
            .carryout(\eeprom.n3739 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2290_15_lut_LC_14_18_5 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2290_15_lut_LC_14_18_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2290_15_lut_LC_14_18_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2290_15_lut_LC_14_18_5  (
            .in0(_gnd_net_),
            .in1(N__27714),
            .in2(N__22166),
            .in3(N__22130),
            .lcout(\eeprom.n3473_adj_388 ),
            .ltout(),
            .carryin(\eeprom.n3739 ),
            .carryout(\eeprom.n3740 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2290_16_lut_LC_14_18_6 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2290_16_lut_LC_14_18_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2290_16_lut_LC_14_18_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2290_16_lut_LC_14_18_6  (
            .in0(_gnd_net_),
            .in1(N__27711),
            .in2(N__22685),
            .in3(N__22652),
            .lcout(\eeprom.n3472_adj_387 ),
            .ltout(),
            .carryin(\eeprom.n3740 ),
            .carryout(\eeprom.n3741 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2290_17_lut_LC_14_18_7 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2290_17_lut_LC_14_18_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2290_17_lut_LC_14_18_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2290_17_lut_LC_14_18_7  (
            .in0(_gnd_net_),
            .in1(N__27715),
            .in2(N__23255),
            .in3(N__22649),
            .lcout(\eeprom.n3471_adj_386 ),
            .ltout(),
            .carryin(\eeprom.n3741 ),
            .carryout(\eeprom.n3742 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2290_18_lut_LC_14_19_0 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2290_18_lut_LC_14_19_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2290_18_lut_LC_14_19_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2290_18_lut_LC_14_19_0  (
            .in0(_gnd_net_),
            .in1(N__27509),
            .in2(N__22646),
            .in3(N__22613),
            .lcout(\eeprom.n3470_adj_385 ),
            .ltout(),
            .carryin(bfn_14_19_0_),
            .carryout(\eeprom.n3743 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2290_19_lut_LC_14_19_1 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2290_19_lut_LC_14_19_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2290_19_lut_LC_14_19_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2290_19_lut_LC_14_19_1  (
            .in0(_gnd_net_),
            .in1(N__22610),
            .in2(N__27706),
            .in3(N__22577),
            .lcout(\eeprom.n3469_adj_384 ),
            .ltout(),
            .carryin(\eeprom.n3743 ),
            .carryout(\eeprom.n3744 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2290_20_lut_LC_14_19_2 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2290_20_lut_LC_14_19_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2290_20_lut_LC_14_19_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2290_20_lut_LC_14_19_2  (
            .in0(_gnd_net_),
            .in1(N__27513),
            .in2(N__22574),
            .in3(N__22532),
            .lcout(\eeprom.n3468_adj_383 ),
            .ltout(),
            .carryin(\eeprom.n3744 ),
            .carryout(\eeprom.n3745 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2290_21_lut_LC_14_19_3 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2290_21_lut_LC_14_19_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2290_21_lut_LC_14_19_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2290_21_lut_LC_14_19_3  (
            .in0(_gnd_net_),
            .in1(N__27518),
            .in2(N__22529),
            .in3(N__22493),
            .lcout(\eeprom.n3467_adj_382 ),
            .ltout(),
            .carryin(\eeprom.n3745 ),
            .carryout(\eeprom.n3746 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2290_22_lut_LC_14_19_4 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2290_22_lut_LC_14_19_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2290_22_lut_LC_14_19_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2290_22_lut_LC_14_19_4  (
            .in0(_gnd_net_),
            .in1(N__27514),
            .in2(N__22490),
            .in3(N__22448),
            .lcout(\eeprom.n3466_adj_381 ),
            .ltout(),
            .carryin(\eeprom.n3746 ),
            .carryout(\eeprom.n3747 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2290_23_lut_LC_14_19_5 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2290_23_lut_LC_14_19_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2290_23_lut_LC_14_19_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2290_23_lut_LC_14_19_5  (
            .in0(_gnd_net_),
            .in1(N__22444),
            .in2(N__27707),
            .in3(N__22736),
            .lcout(\eeprom.n3465_adj_380 ),
            .ltout(),
            .carryin(\eeprom.n3747 ),
            .carryout(\eeprom.n3748 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2290_24_lut_LC_14_19_6 .C_ON=1'b0;
    defparam \eeprom.rem_4_add_2290_24_lut_LC_14_19_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2290_24_lut_LC_14_19_6 .LUT_INIT=16'b1001000001100000;
    LogicCell40 \eeprom.rem_4_add_2290_24_lut_LC_14_19_6  (
            .in0(N__27519),
            .in1(N__22733),
            .in2(N__23369),
            .in3(N__22712),
            .lcout(\eeprom.n3496 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i1_2_lut_adj_58_LC_14_19_7 .C_ON=1'b0;
    defparam \eeprom.i1_2_lut_adj_58_LC_14_19_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.i1_2_lut_adj_58_LC_14_19_7 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \eeprom.i1_2_lut_adj_58_LC_14_19_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__26056),
            .in3(N__25525),
            .lcout(\eeprom.n4619 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i1_4_lut_adj_56_LC_14_20_0 .C_ON=1'b0;
    defparam \eeprom.i1_4_lut_adj_56_LC_14_20_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.i1_4_lut_adj_56_LC_14_20_0 .LUT_INIT=16'b1111101011111100;
    LogicCell40 \eeprom.i1_4_lut_adj_56_LC_14_20_0  (
            .in0(N__25445),
            .in1(N__25466),
            .in2(N__22709),
            .in3(N__25663),
            .lcout(),
            .ltout(\eeprom.n31_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i1_4_lut_adj_62_LC_14_20_1 .C_ON=1'b0;
    defparam \eeprom.i1_4_lut_adj_62_LC_14_20_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.i1_4_lut_adj_62_LC_14_20_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \eeprom.i1_4_lut_adj_62_LC_14_20_1  (
            .in0(N__26014),
            .in1(N__22691),
            .in2(N__22700),
            .in3(N__22697),
            .lcout(\eeprom.n4567 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2445_3_lut_LC_14_20_2 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2445_3_lut_LC_14_20_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2445_3_lut_LC_14_20_2 .LUT_INIT=16'b0011000000111111;
    LogicCell40 \eeprom.rem_4_i2445_3_lut_LC_14_20_2  (
            .in0(_gnd_net_),
            .in1(N__25478),
            .in2(N__25832),
            .in3(N__25502),
            .lcout(\eeprom.n3713_adj_443 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2362_3_lut_LC_14_20_3 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2362_3_lut_LC_14_20_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2362_3_lut_LC_14_20_3 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \eeprom.rem_4_i2362_3_lut_LC_14_20_3  (
            .in0(N__25662),
            .in1(_gnd_net_),
            .in2(N__25217),
            .in3(N__25239),
            .lcout(\eeprom.n3598_adj_452 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2376_3_lut_LC_14_20_4 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2376_3_lut_LC_14_20_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2376_3_lut_LC_14_20_4 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \eeprom.rem_4_i2376_3_lut_LC_14_20_4  (
            .in0(_gnd_net_),
            .in1(N__25139),
            .in2(N__25175),
            .in3(N__25661),
            .lcout(\eeprom.n3612_adj_339 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2444_3_lut_LC_14_20_5 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2444_3_lut_LC_14_20_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2444_3_lut_LC_14_20_5 .LUT_INIT=16'b0000111100110011;
    LogicCell40 \eeprom.rem_4_i2444_3_lut_LC_14_20_5  (
            .in0(_gnd_net_),
            .in1(N__26055),
            .in2(N__26033),
            .in3(N__25817),
            .lcout(\eeprom.n3712_adj_444 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2360_3_lut_LC_14_20_7 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2360_3_lut_LC_14_20_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2360_3_lut_LC_14_20_7 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \eeprom.rem_4_i2360_3_lut_LC_14_20_7  (
            .in0(N__25664),
            .in1(_gnd_net_),
            .in2(N__25766),
            .in3(N__25739),
            .lcout(\eeprom.n3596_adj_454 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_mux_3_i3_3_lut_LC_14_21_1 .C_ON=1'b0;
    defparam \eeprom.rem_4_mux_3_i3_3_lut_LC_14_21_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_mux_3_i3_3_lut_LC_14_21_1 .LUT_INIT=16'b0011001101010101;
    LogicCell40 \eeprom.rem_4_mux_3_i3_3_lut_LC_14_21_1  (
            .in0(N__23845),
            .in1(N__23003),
            .in2(_gnd_net_),
            .in3(N__22991),
            .lcout(\eeprom.n3723_adj_334 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i4077_1_lut_LC_14_21_3 .C_ON=1'b0;
    defparam \eeprom.i4077_1_lut_LC_14_21_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.i4077_1_lut_LC_14_21_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \eeprom.i4077_1_lut_LC_14_21_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24091),
            .lcout(\eeprom.n4921 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i4080_1_lut_2_lut_LC_14_21_7 .C_ON=1'b0;
    defparam \eeprom.i4080_1_lut_2_lut_LC_14_21_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.i4080_1_lut_2_lut_LC_14_21_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \eeprom.i4080_1_lut_2_lut_LC_14_21_7  (
            .in0(_gnd_net_),
            .in1(N__25952),
            .in2(_gnd_net_),
            .in3(N__25833),
            .lcout(\eeprom.n4924 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i10_4_lut_adj_66_LC_14_22_5 .C_ON=1'b0;
    defparam \eeprom.i10_4_lut_adj_66_LC_14_22_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.i10_4_lut_adj_66_LC_14_22_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \eeprom.i10_4_lut_adj_66_LC_14_22_5  (
            .in0(N__24201),
            .in1(N__24231),
            .in2(N__24273),
            .in3(N__24171),
            .lcout(\eeprom.n24_adj_459 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i1_2_lut_adj_39_LC_14_23_2 .C_ON=1'b0;
    defparam \eeprom.i1_2_lut_adj_39_LC_14_23_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.i1_2_lut_adj_39_LC_14_23_2 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \eeprom.i1_2_lut_adj_39_LC_14_23_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__26092),
            .in3(N__26184),
            .lcout(),
            .ltout(\eeprom.n4559_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i1_4_lut_adj_40_LC_14_23_3 .C_ON=1'b0;
    defparam \eeprom.i1_4_lut_adj_40_LC_14_23_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.i1_4_lut_adj_40_LC_14_23_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \eeprom.i1_4_lut_adj_40_LC_14_23_3  (
            .in0(N__26244),
            .in1(N__26145),
            .in2(N__22760),
            .in3(N__26293),
            .lcout(),
            .ltout(\eeprom.n4563_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i4_4_lut_adj_41_LC_14_23_4 .C_ON=1'b0;
    defparam \eeprom.i4_4_lut_adj_41_LC_14_23_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.i4_4_lut_adj_41_LC_14_23_4 .LUT_INIT=16'b1111101011101010;
    LogicCell40 \eeprom.i4_4_lut_adj_41_LC_14_23_4  (
            .in0(N__26513),
            .in1(N__26385),
            .in2(N__22757),
            .in3(N__26331),
            .lcout(),
            .ltout(\eeprom.n17_adj_421_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i11_4_lut_adj_43_LC_14_23_5 .C_ON=1'b0;
    defparam \eeprom.i11_4_lut_adj_43_LC_14_23_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.i11_4_lut_adj_43_LC_14_23_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \eeprom.i11_4_lut_adj_43_LC_14_23_5  (
            .in0(N__22754),
            .in1(N__26539),
            .in2(N__22748),
            .in3(N__26593),
            .lcout(),
            .ltout(\eeprom.n24_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i12_4_lut_LC_14_23_6 .C_ON=1'b0;
    defparam \eeprom.i12_4_lut_LC_14_23_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.i12_4_lut_LC_14_23_6 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \eeprom.i12_4_lut_LC_14_23_6  (
            .in0(N__26667),
            .in1(N__26635),
            .in2(N__22745),
            .in3(N__22742),
            .lcout(\eeprom.n3034 ),
            .ltout(\eeprom.n3034_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2036_3_lut_LC_14_23_7 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2036_3_lut_LC_14_23_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2036_3_lut_LC_14_23_7 .LUT_INIT=16'b1111110000001100;
    LogicCell40 \eeprom.rem_4_i2036_3_lut_LC_14_23_7  (
            .in0(_gnd_net_),
            .in1(N__26088),
            .in2(N__23225),
            .in3(N__26069),
            .lcout(\eeprom.n3112 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1967_3_lut_LC_14_24_5 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1967_3_lut_LC_14_24_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1967_3_lut_LC_14_24_5 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \eeprom.rem_4_i1967_3_lut_LC_14_24_5  (
            .in0(_gnd_net_),
            .in1(N__23189),
            .in2(N__23159),
            .in3(N__24762),
            .lcout(\eeprom.n3011 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2027_3_lut_LC_14_24_7 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2027_3_lut_LC_14_24_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2027_3_lut_LC_14_24_7 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \eeprom.rem_4_i2027_3_lut_LC_14_24_7  (
            .in0(_gnd_net_),
            .in1(N__28072),
            .in2(N__28049),
            .in3(N__27887),
            .lcout(\eeprom.n3103 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i1_4_lut_adj_115_LC_15_17_0 .C_ON=1'b0;
    defparam \eeprom.i1_4_lut_adj_115_LC_15_17_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.i1_4_lut_adj_115_LC_15_17_0 .LUT_INIT=16'b1110000000000000;
    LogicCell40 \eeprom.i1_4_lut_adj_115_LC_15_17_0  (
            .in0(N__24600),
            .in1(N__24658),
            .in2(N__23435),
            .in3(N__23042),
            .lcout(\eeprom.n4137 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2312_3_lut_LC_15_17_1 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2312_3_lut_LC_15_17_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2312_3_lut_LC_15_17_1 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \eeprom.rem_4_i2312_3_lut_LC_15_17_1  (
            .in0(_gnd_net_),
            .in1(N__23114),
            .in2(N__23087),
            .in3(N__23372),
            .lcout(\eeprom.n3516_adj_372 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2380_3_lut_LC_15_17_2 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2380_3_lut_LC_15_17_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2380_3_lut_LC_15_17_2 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \eeprom.rem_4_i2380_3_lut_LC_15_17_2  (
            .in0(N__24560),
            .in1(_gnd_net_),
            .in2(N__25705),
            .in3(N__24574),
            .lcout(\eeprom.n3616_adj_345 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2313_3_lut_LC_15_17_3 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2313_3_lut_LC_15_17_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2313_3_lut_LC_15_17_3 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \eeprom.rem_4_i2313_3_lut_LC_15_17_3  (
            .in0(_gnd_net_),
            .in1(N__23077),
            .in2(N__23054),
            .in3(N__23374),
            .lcout(\eeprom.n3517_adj_374 ),
            .ltout(\eeprom.n3517_adj_374_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i1_3_lut_adj_114_LC_15_17_4 .C_ON=1'b0;
    defparam \eeprom.i1_3_lut_adj_114_LC_15_17_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.i1_3_lut_adj_114_LC_15_17_4 .LUT_INIT=16'b1100000000000000;
    LogicCell40 \eeprom.i1_3_lut_adj_114_LC_15_17_4  (
            .in0(_gnd_net_),
            .in1(N__24483),
            .in2(N__23045),
            .in3(N__24543),
            .lcout(\eeprom.n4729 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2311_3_lut_LC_15_17_5 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2311_3_lut_LC_15_17_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2311_3_lut_LC_15_17_5 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \eeprom.rem_4_i2311_3_lut_LC_15_17_5  (
            .in0(_gnd_net_),
            .in1(N__23035),
            .in2(N__23012),
            .in3(N__23373),
            .lcout(\eeprom.n3515_adj_370 ),
            .ltout(\eeprom.n3515_adj_370_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i1_2_lut_adj_111_LC_15_17_6 .C_ON=1'b0;
    defparam \eeprom.i1_2_lut_adj_111_LC_15_17_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.i1_2_lut_adj_111_LC_15_17_6 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \eeprom.i1_2_lut_adj_111_LC_15_17_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__23438),
            .in3(N__25161),
            .lcout(\eeprom.n4727 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2378_3_lut_LC_15_17_7 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2378_3_lut_LC_15_17_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2378_3_lut_LC_15_17_7 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \eeprom.rem_4_i2378_3_lut_LC_15_17_7  (
            .in0(_gnd_net_),
            .in1(N__24517),
            .in2(N__24503),
            .in3(N__25696),
            .lcout(\eeprom.n3614_adj_343 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2314_3_lut_LC_15_18_0 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2314_3_lut_LC_15_18_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2314_3_lut_LC_15_18_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \eeprom.rem_4_i2314_3_lut_LC_15_18_0  (
            .in0(N__23426),
            .in1(N__23387),
            .in2(_gnd_net_),
            .in3(N__23365),
            .lcout(\eeprom.n3518_adj_376 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2299_3_lut_LC_15_18_1 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2299_3_lut_LC_15_18_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2299_3_lut_LC_15_18_1 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \eeprom.rem_4_i2299_3_lut_LC_15_18_1  (
            .in0(_gnd_net_),
            .in1(N__23381),
            .in2(N__23375),
            .in3(N__23254),
            .lcout(\eeprom.n3503 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2369_3_lut_LC_15_18_2 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2369_3_lut_LC_15_18_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2369_3_lut_LC_15_18_2 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \eeprom.rem_4_i2369_3_lut_LC_15_18_2  (
            .in0(_gnd_net_),
            .in1(N__24857),
            .in2(N__25704),
            .in3(N__24884),
            .lcout(\eeprom.n3605_adj_453 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2379_3_lut_LC_15_18_3 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2379_3_lut_LC_15_18_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2379_3_lut_LC_15_18_3 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \eeprom.rem_4_i2379_3_lut_LC_15_18_3  (
            .in0(_gnd_net_),
            .in1(N__24527),
            .in2(N__24551),
            .in3(N__25689),
            .lcout(\eeprom.n3615_adj_344 ),
            .ltout(\eeprom.n3615_adj_344_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2446_3_lut_LC_15_18_4 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2446_3_lut_LC_15_18_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2446_3_lut_LC_15_18_4 .LUT_INIT=16'b0011001100001111;
    LogicCell40 \eeprom.rem_4_i2446_3_lut_LC_15_18_4  (
            .in0(_gnd_net_),
            .in1(N__25514),
            .in2(N__23231),
            .in3(N__25816),
            .lcout(\eeprom.n3714_adj_442 ),
            .ltout(\eeprom.n3714_adj_442_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i4071_1_lut_LC_15_18_5 .C_ON=1'b0;
    defparam \eeprom.i4071_1_lut_LC_15_18_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.i4071_1_lut_LC_15_18_5 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \eeprom.i4071_1_lut_LC_15_18_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__23228),
            .in3(_gnd_net_),
            .lcout(\eeprom.n4915 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2381_3_lut_LC_15_18_6 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2381_3_lut_LC_15_18_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2381_3_lut_LC_15_18_6 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \eeprom.rem_4_i2381_3_lut_LC_15_18_6  (
            .in0(N__24584),
            .in1(_gnd_net_),
            .in2(N__25703),
            .in3(N__24604),
            .lcout(\eeprom.n3617_adj_346 ),
            .ltout(\eeprom.n3617_adj_346_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i1_4_lut_adj_59_LC_15_18_7 .C_ON=1'b0;
    defparam \eeprom.i1_4_lut_adj_59_LC_15_18_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.i1_4_lut_adj_59_LC_15_18_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \eeprom.i1_4_lut_adj_59_LC_15_18_7  (
            .in0(N__25494),
            .in1(N__25980),
            .in2(N__23555),
            .in3(N__23552),
            .lcout(\eeprom.n4623 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i1_4_lut_adj_61_LC_15_19_0 .C_ON=1'b0;
    defparam \eeprom.i1_4_lut_adj_61_LC_15_19_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.i1_4_lut_adj_61_LC_15_19_0 .LUT_INIT=16'b1111111111100010;
    LogicCell40 \eeprom.i1_4_lut_adj_61_LC_15_19_0  (
            .in0(N__25349),
            .in1(N__25684),
            .in2(N__25328),
            .in3(N__23507),
            .lcout(),
            .ltout(\eeprom.n4427_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i1_4_lut_adj_63_LC_15_19_1 .C_ON=1'b0;
    defparam \eeprom.i1_4_lut_adj_63_LC_15_19_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.i1_4_lut_adj_63_LC_15_19_1 .LUT_INIT=16'b1111110111111000;
    LogicCell40 \eeprom.i1_4_lut_adj_63_LC_15_19_1  (
            .in0(N__25685),
            .in1(N__25775),
            .in2(N__23546),
            .in3(N__25199),
            .lcout(),
            .ltout(\eeprom.n28_adj_455_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i1_4_lut_adj_64_LC_15_19_2 .C_ON=1'b0;
    defparam \eeprom.i1_4_lut_adj_64_LC_15_19_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.i1_4_lut_adj_64_LC_15_19_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \eeprom.i1_4_lut_adj_64_LC_15_19_2  (
            .in0(N__25571),
            .in1(N__23543),
            .in2(N__23537),
            .in3(N__23534),
            .lcout(\eeprom.n3628_adj_437 ),
            .ltout(\eeprom.n3628_adj_437_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2448_3_lut_LC_15_19_3 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2448_3_lut_LC_15_19_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2448_3_lut_LC_15_19_3 .LUT_INIT=16'b0011000000111111;
    LogicCell40 \eeprom.rem_4_i2448_3_lut_LC_15_19_3  (
            .in0(_gnd_net_),
            .in1(N__25544),
            .in2(N__23528),
            .in3(N__25558),
            .lcout(\eeprom.n3716_adj_439 ),
            .ltout(\eeprom.n3716_adj_439_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i4065_1_lut_LC_15_19_4 .C_ON=1'b0;
    defparam \eeprom.i4065_1_lut_LC_15_19_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.i4065_1_lut_LC_15_19_4 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \eeprom.i4065_1_lut_LC_15_19_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__23525),
            .in3(_gnd_net_),
            .lcout(\eeprom.n4909 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2382_3_lut_LC_15_19_6 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2382_3_lut_LC_15_19_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2382_3_lut_LC_15_19_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \eeprom.rem_4_i2382_3_lut_LC_15_19_6  (
            .in0(N__24620),
            .in1(N__24654),
            .in2(_gnd_net_),
            .in3(N__25683),
            .lcout(\eeprom.n3618_adj_350 ),
            .ltout(\eeprom.n3618_adj_350_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i1_4_lut_adj_60_LC_15_19_7 .C_ON=1'b0;
    defparam \eeprom.i1_4_lut_adj_60_LC_15_19_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.i1_4_lut_adj_60_LC_15_19_7 .LUT_INIT=16'b1111111011001100;
    LogicCell40 \eeprom.i1_4_lut_adj_60_LC_15_19_7  (
            .in0(N__25876),
            .in1(N__23522),
            .in2(N__23516),
            .in3(N__23513),
            .lcout(\eeprom.n4425 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2473_2_lut_LC_15_20_0 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2473_2_lut_LC_15_20_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2473_2_lut_LC_15_20_0 .LUT_INIT=16'b1000101110111000;
    LogicCell40 \eeprom.rem_4_add_2473_2_lut_LC_15_20_0  (
            .in0(N__23501),
            .in1(N__24062),
            .in2(N__23459),
            .in3(N__23441),
            .lcout(\eeprom.number_of_bytes_7_N_68_0 ),
            .ltout(),
            .carryin(bfn_15_20_0_),
            .carryout(\eeprom.n3772 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2473_3_lut_LC_15_20_1 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2473_3_lut_LC_15_20_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2473_3_lut_LC_15_20_1 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \eeprom.rem_4_add_2473_3_lut_LC_15_20_1  (
            .in0(N__23912),
            .in1(N__23867),
            .in2(N__24075),
            .in3(N__23855),
            .lcout(\eeprom.number_of_bytes_7_N_68_1 ),
            .ltout(),
            .carryin(\eeprom.n3772 ),
            .carryout(\eeprom.n3773 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2473_4_lut_LC_15_20_2 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2473_4_lut_LC_15_20_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2473_4_lut_LC_15_20_2 .LUT_INIT=16'b1000101110111000;
    LogicCell40 \eeprom.rem_4_add_2473_4_lut_LC_15_20_2  (
            .in0(N__23852),
            .in1(N__24066),
            .in2(N__23804),
            .in3(N__23792),
            .lcout(\eeprom.number_of_bytes_7_N_68_2 ),
            .ltout(),
            .carryin(\eeprom.n3773 ),
            .carryout(\eeprom.n3774 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2473_5_lut_LC_15_20_3 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2473_5_lut_LC_15_20_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2473_5_lut_LC_15_20_3 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \eeprom.rem_4_add_2473_5_lut_LC_15_20_3  (
            .in0(N__23789),
            .in1(N__23747),
            .in2(N__24076),
            .in3(N__23729),
            .lcout(\eeprom.number_of_bytes_7_N_68_3 ),
            .ltout(),
            .carryin(\eeprom.n3774 ),
            .carryout(\eeprom.n3775 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2473_6_lut_LC_15_20_4 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2473_6_lut_LC_15_20_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2473_6_lut_LC_15_20_4 .LUT_INIT=16'b1000101110111000;
    LogicCell40 \eeprom.rem_4_add_2473_6_lut_LC_15_20_4  (
            .in0(N__23726),
            .in1(N__24070),
            .in2(N__23687),
            .in3(N__23675),
            .lcout(\eeprom.number_of_bytes_7_N_68_4 ),
            .ltout(),
            .carryin(\eeprom.n3775 ),
            .carryout(\eeprom.n3776 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2473_7_lut_LC_15_20_5 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2473_7_lut_LC_15_20_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2473_7_lut_LC_15_20_5 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \eeprom.rem_4_add_2473_7_lut_LC_15_20_5  (
            .in0(N__23672),
            .in1(N__23630),
            .in2(N__24077),
            .in3(N__23621),
            .lcout(\eeprom.number_of_bytes_7_N_68_5 ),
            .ltout(),
            .carryin(\eeprom.n3776 ),
            .carryout(\eeprom.n3777 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2473_8_lut_LC_15_20_6 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2473_8_lut_LC_15_20_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2473_8_lut_LC_15_20_6 .LUT_INIT=16'b1000101110111000;
    LogicCell40 \eeprom.rem_4_add_2473_8_lut_LC_15_20_6  (
            .in0(N__23618),
            .in1(N__24074),
            .in2(N__23579),
            .in3(N__23564),
            .lcout(\eeprom.number_of_bytes_7_N_68_6 ),
            .ltout(),
            .carryin(\eeprom.n3777 ),
            .carryout(\eeprom.n3778 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2473_9_lut_LC_15_20_7 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2473_9_lut_LC_15_20_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2473_9_lut_LC_15_20_7 .LUT_INIT=16'b1000101110111000;
    LogicCell40 \eeprom.rem_4_add_2473_9_lut_LC_15_20_7  (
            .in0(N__26396),
            .in1(N__24059),
            .in2(N__25784),
            .in3(N__23561),
            .lcout(\eeprom.number_of_bytes_7_N_68_7 ),
            .ltout(),
            .carryin(\eeprom.n3778 ),
            .carryout(\eeprom.n3779 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2473_10_lut_LC_15_21_0 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2473_10_lut_LC_15_21_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2473_10_lut_LC_15_21_0 .LUT_INIT=16'b1000101110111000;
    LogicCell40 \eeprom.rem_4_add_2473_10_lut_LC_15_21_0  (
            .in0(N__25889),
            .in1(N__24043),
            .in2(N__25901),
            .in3(N__23558),
            .lcout(\eeprom.number_of_bytes_7_N_68_8 ),
            .ltout(),
            .carryin(bfn_15_21_0_),
            .carryout(\eeprom.n3780 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2473_11_lut_LC_15_21_1 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2473_11_lut_LC_15_21_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2473_11_lut_LC_15_21_1 .LUT_INIT=16'b1000101110111000;
    LogicCell40 \eeprom.rem_4_add_2473_11_lut_LC_15_21_1  (
            .in0(N__24155),
            .in1(N__24033),
            .in2(N__24146),
            .in3(N__24134),
            .lcout(\eeprom.number_of_bytes_7_N_68_9 ),
            .ltout(),
            .carryin(\eeprom.n3780 ),
            .carryout(\eeprom.n3781 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2473_12_lut_LC_15_21_2 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2473_12_lut_LC_15_21_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2473_12_lut_LC_15_21_2 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \eeprom.rem_4_add_2473_12_lut_LC_15_21_2  (
            .in0(N__25958),
            .in1(N__25967),
            .in2(N__24060),
            .in3(N__24131),
            .lcout(\eeprom.number_of_bytes_7_N_68_10 ),
            .ltout(),
            .carryin(\eeprom.n3781 ),
            .carryout(\eeprom.n3782 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2473_13_lut_LC_15_21_3 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2473_13_lut_LC_15_21_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2473_13_lut_LC_15_21_3 .LUT_INIT=16'b1000101110111000;
    LogicCell40 \eeprom.rem_4_add_2473_13_lut_LC_15_21_3  (
            .in0(N__24128),
            .in1(N__24037),
            .in2(N__24119),
            .in3(N__24107),
            .lcout(\eeprom.number_of_bytes_7_N_68_11 ),
            .ltout(),
            .carryin(\eeprom.n3782 ),
            .carryout(\eeprom.n3783 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2473_14_lut_LC_15_21_4 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2473_14_lut_LC_15_21_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2473_14_lut_LC_15_21_4 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \eeprom.rem_4_add_2473_14_lut_LC_15_21_4  (
            .in0(N__23948),
            .in1(N__23959),
            .in2(N__24061),
            .in3(N__24104),
            .lcout(\eeprom.number_of_bytes_7_N_68_12 ),
            .ltout(),
            .carryin(\eeprom.n3783 ),
            .carryout(\eeprom.n3784 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2473_15_lut_LC_15_21_5 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2473_15_lut_LC_15_21_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2473_15_lut_LC_15_21_5 .LUT_INIT=16'b1000101110111000;
    LogicCell40 \eeprom.rem_4_add_2473_15_lut_LC_15_21_5  (
            .in0(N__24101),
            .in1(N__24041),
            .in2(N__24095),
            .in3(N__24080),
            .lcout(\eeprom.number_of_bytes_7_N_68_13 ),
            .ltout(),
            .carryin(\eeprom.n3784 ),
            .carryout(\eeprom.n3785 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2473_16_lut_LC_15_21_6 .C_ON=1'b0;
    defparam \eeprom.rem_4_add_2473_16_lut_LC_15_21_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2473_16_lut_LC_15_21_6 .LUT_INIT=16'b1000110111011000;
    LogicCell40 \eeprom.rem_4_add_2473_16_lut_LC_15_21_6  (
            .in0(N__24042),
            .in1(N__23969),
            .in2(N__25934),
            .in3(N__23963),
            .lcout(\eeprom.number_of_bytes_7_N_68_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i4074_1_lut_LC_15_21_7 .C_ON=1'b0;
    defparam \eeprom.i4074_1_lut_LC_15_21_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.i4074_1_lut_LC_15_21_7 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \eeprom.i4074_1_lut_LC_15_21_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__23960),
            .in3(_gnd_net_),
            .lcout(\eeprom.n4918 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i1_4_lut_adj_113_LC_15_22_0 .C_ON=1'b0;
    defparam \eeprom.i1_4_lut_adj_113_LC_15_22_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.i1_4_lut_adj_113_LC_15_22_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \eeprom.i1_4_lut_adj_113_LC_15_22_0  (
            .in0(N__23942),
            .in1(N__23933),
            .in2(N__23924),
            .in3(N__24290),
            .lcout(),
            .ltout(\eeprom.n4301_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i1_4_lut_adj_119_LC_15_22_1 .C_ON=1'b0;
    defparam \eeprom.i1_4_lut_adj_119_LC_15_22_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.i1_4_lut_adj_119_LC_15_22_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \eeprom.i1_4_lut_adj_119_LC_15_22_1  (
            .in0(N__24443),
            .in1(N__24434),
            .in2(N__24428),
            .in3(N__24425),
            .lcout(),
            .ltout(\eeprom.n4307_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i1_4_lut_adj_120_LC_15_22_2 .C_ON=1'b0;
    defparam \eeprom.i1_4_lut_adj_120_LC_15_22_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.i1_4_lut_adj_120_LC_15_22_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \eeprom.i1_4_lut_adj_120_LC_15_22_2  (
            .in0(N__24416),
            .in1(N__24410),
            .in2(N__24404),
            .in3(N__24401),
            .lcout(),
            .ltout(\eeprom.n4313_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.ena_12_LC_15_22_3 .C_ON=1'b0;
    defparam \eeprom.ena_12_LC_15_22_3 .SEQ_MODE=4'b1000;
    defparam \eeprom.ena_12_LC_15_22_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \eeprom.ena_12_LC_15_22_3  (
            .in0(N__24395),
            .in1(N__24389),
            .in2(N__24383),
            .in3(N__24380),
            .lcout(sda_enable),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24349),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i1_3_lut_adj_112_LC_15_22_7 .C_ON=1'b0;
    defparam \eeprom.i1_3_lut_adj_112_LC_15_22_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.i1_3_lut_adj_112_LC_15_22_7 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \eeprom.i1_3_lut_adj_112_LC_15_22_7  (
            .in0(N__24317),
            .in1(N__24308),
            .in2(_gnd_net_),
            .in3(N__24299),
            .lcout(\eeprom.n4295 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2035_3_lut_LC_15_23_0 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2035_3_lut_LC_15_23_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2035_3_lut_LC_15_23_0 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \eeprom.rem_4_i2035_3_lut_LC_15_23_0  (
            .in0(_gnd_net_),
            .in1(N__26681),
            .in2(N__27909),
            .in3(N__26704),
            .lcout(\eeprom.n3111 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2033_3_lut_LC_15_23_3 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2033_3_lut_LC_15_23_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2033_3_lut_LC_15_23_3 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \eeprom.rem_4_i2033_3_lut_LC_15_23_3  (
            .in0(_gnd_net_),
            .in1(N__26639),
            .in2(N__26606),
            .in3(N__27882),
            .lcout(\eeprom.n3109 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2034_3_lut_LC_15_23_5 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2034_3_lut_LC_15_23_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2034_3_lut_LC_15_23_5 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \eeprom.rem_4_i2034_3_lut_LC_15_23_5  (
            .in0(_gnd_net_),
            .in1(N__26671),
            .in2(N__26651),
            .in3(N__27881),
            .lcout(\eeprom.n3110 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2031_3_lut_LC_15_23_7 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2031_3_lut_LC_15_23_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2031_3_lut_LC_15_23_7 .LUT_INIT=16'b1010101011110000;
    LogicCell40 \eeprom.rem_4_i2031_3_lut_LC_15_23_7  (
            .in0(N__26522),
            .in1(_gnd_net_),
            .in2(N__26543),
            .in3(N__27886),
            .lcout(\eeprom.n3107 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1974_3_lut_LC_15_24_2 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1974_3_lut_LC_15_24_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1974_3_lut_LC_15_24_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \eeprom.rem_4_i1974_3_lut_LC_15_24_2  (
            .in0(N__24848),
            .in1(N__24836),
            .in2(_gnd_net_),
            .in3(N__24760),
            .lcout(\eeprom.n3018 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1964_3_lut_LC_15_24_6 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1964_3_lut_LC_15_24_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1964_3_lut_LC_15_24_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \eeprom.rem_4_i1964_3_lut_LC_15_24_6  (
            .in0(N__24796),
            .in1(N__24776),
            .in2(_gnd_net_),
            .in3(N__24761),
            .lcout(\eeprom.n3008 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2357_2_lut_LC_16_17_0 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2357_2_lut_LC_16_17_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2357_2_lut_LC_16_17_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2357_2_lut_LC_16_17_0  (
            .in0(_gnd_net_),
            .in1(N__24659),
            .in2(_gnd_net_),
            .in3(N__24608),
            .lcout(\eeprom.n3586_adj_378 ),
            .ltout(),
            .carryin(bfn_16_17_0_),
            .carryout(\eeprom.n3749 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2357_3_lut_LC_16_17_1 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2357_3_lut_LC_16_17_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2357_3_lut_LC_16_17_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2357_3_lut_LC_16_17_1  (
            .in0(_gnd_net_),
            .in1(N__27024),
            .in2(N__24605),
            .in3(N__24578),
            .lcout(\eeprom.n3585_adj_375 ),
            .ltout(),
            .carryin(\eeprom.n3749 ),
            .carryout(\eeprom.n3750 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2357_4_lut_LC_16_17_2 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2357_4_lut_LC_16_17_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2357_4_lut_LC_16_17_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2357_4_lut_LC_16_17_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__24575),
            .in3(N__24554),
            .lcout(\eeprom.n3584_adj_373 ),
            .ltout(),
            .carryin(\eeprom.n3750 ),
            .carryout(\eeprom.n3751 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2357_5_lut_LC_16_17_3 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2357_5_lut_LC_16_17_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2357_5_lut_LC_16_17_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2357_5_lut_LC_16_17_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__24550),
            .in3(N__24521),
            .lcout(\eeprom.n3583_adj_371 ),
            .ltout(),
            .carryin(\eeprom.n3751 ),
            .carryout(\eeprom.n3752 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2357_6_lut_LC_16_17_4 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2357_6_lut_LC_16_17_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2357_6_lut_LC_16_17_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2357_6_lut_LC_16_17_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__24518),
            .in3(N__24494),
            .lcout(\eeprom.n3582_adj_369 ),
            .ltout(),
            .carryin(\eeprom.n3752 ),
            .carryout(\eeprom.n3753 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2357_7_lut_LC_16_17_5 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2357_7_lut_LC_16_17_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2357_7_lut_LC_16_17_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2357_7_lut_LC_16_17_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__24491),
            .in3(N__24446),
            .lcout(\eeprom.n3581_adj_367 ),
            .ltout(),
            .carryin(\eeprom.n3753 ),
            .carryout(\eeprom.n3754 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2357_8_lut_LC_16_17_6 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2357_8_lut_LC_16_17_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2357_8_lut_LC_16_17_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2357_8_lut_LC_16_17_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__25174),
            .in3(N__25127),
            .lcout(\eeprom.n3580_adj_365 ),
            .ltout(),
            .carryin(\eeprom.n3754 ),
            .carryout(\eeprom.n3755 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2357_9_lut_LC_16_17_7 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2357_9_lut_LC_16_17_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2357_9_lut_LC_16_17_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2357_9_lut_LC_16_17_7  (
            .in0(_gnd_net_),
            .in1(N__27025),
            .in2(N__25124),
            .in3(N__25082),
            .lcout(\eeprom.n3579_adj_363 ),
            .ltout(),
            .carryin(\eeprom.n3755 ),
            .carryout(\eeprom.n3756 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2357_10_lut_LC_16_18_0 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2357_10_lut_LC_16_18_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2357_10_lut_LC_16_18_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2357_10_lut_LC_16_18_0  (
            .in0(_gnd_net_),
            .in1(N__27008),
            .in2(N__25079),
            .in3(N__25040),
            .lcout(\eeprom.n3578_adj_361 ),
            .ltout(),
            .carryin(bfn_16_18_0_),
            .carryout(\eeprom.n3757 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2357_11_lut_LC_16_18_1 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2357_11_lut_LC_16_18_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2357_11_lut_LC_16_18_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2357_11_lut_LC_16_18_1  (
            .in0(_gnd_net_),
            .in1(N__27016),
            .in2(N__25037),
            .in3(N__25001),
            .lcout(\eeprom.n3577_adj_359 ),
            .ltout(),
            .carryin(\eeprom.n3757 ),
            .carryout(\eeprom.n3758 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2357_12_lut_LC_16_18_2 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2357_12_lut_LC_16_18_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2357_12_lut_LC_16_18_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2357_12_lut_LC_16_18_2  (
            .in0(_gnd_net_),
            .in1(N__27009),
            .in2(N__24998),
            .in3(N__24956),
            .lcout(\eeprom.n3576_adj_358 ),
            .ltout(),
            .carryin(\eeprom.n3758 ),
            .carryout(\eeprom.n3759 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2357_13_lut_LC_16_18_3 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2357_13_lut_LC_16_18_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2357_13_lut_LC_16_18_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2357_13_lut_LC_16_18_3  (
            .in0(_gnd_net_),
            .in1(N__27017),
            .in2(N__24953),
            .in3(N__24926),
            .lcout(\eeprom.n3575_adj_357 ),
            .ltout(),
            .carryin(\eeprom.n3759 ),
            .carryout(\eeprom.n3760 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2357_14_lut_LC_16_18_4 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2357_14_lut_LC_16_18_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2357_14_lut_LC_16_18_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2357_14_lut_LC_16_18_4  (
            .in0(_gnd_net_),
            .in1(N__24923),
            .in2(N__27194),
            .in3(N__24887),
            .lcout(\eeprom.n3574_adj_356 ),
            .ltout(),
            .carryin(\eeprom.n3760 ),
            .carryout(\eeprom.n3761 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2357_15_lut_LC_16_18_5 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2357_15_lut_LC_16_18_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2357_15_lut_LC_16_18_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2357_15_lut_LC_16_18_5  (
            .in0(_gnd_net_),
            .in1(N__24883),
            .in2(N__27192),
            .in3(N__24851),
            .lcout(\eeprom.n3573_adj_355 ),
            .ltout(),
            .carryin(\eeprom.n3761 ),
            .carryout(\eeprom.n3762 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2357_16_lut_LC_16_18_6 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2357_16_lut_LC_16_18_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2357_16_lut_LC_16_18_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2357_16_lut_LC_16_18_6  (
            .in0(_gnd_net_),
            .in1(N__25462),
            .in2(N__27195),
            .in3(N__25433),
            .lcout(\eeprom.n3572_adj_354 ),
            .ltout(),
            .carryin(\eeprom.n3762 ),
            .carryout(\eeprom.n3763 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2357_17_lut_LC_16_18_7 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2357_17_lut_LC_16_18_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2357_17_lut_LC_16_18_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2357_17_lut_LC_16_18_7  (
            .in0(_gnd_net_),
            .in1(N__25430),
            .in2(N__27193),
            .in3(N__25397),
            .lcout(\eeprom.n3571_adj_353 ),
            .ltout(),
            .carryin(\eeprom.n3763 ),
            .carryout(\eeprom.n3764 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2357_18_lut_LC_16_19_0 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2357_18_lut_LC_16_19_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2357_18_lut_LC_16_19_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2357_18_lut_LC_16_19_0  (
            .in0(_gnd_net_),
            .in1(N__26988),
            .in2(N__25389),
            .in3(N__25352),
            .lcout(\eeprom.n3570_adj_349 ),
            .ltout(),
            .carryin(bfn_16_19_0_),
            .carryout(\eeprom.n3765 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2357_19_lut_LC_16_19_1 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2357_19_lut_LC_16_19_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2357_19_lut_LC_16_19_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2357_19_lut_LC_16_19_1  (
            .in0(_gnd_net_),
            .in1(N__25348),
            .in2(N__27186),
            .in3(N__25319),
            .lcout(\eeprom.n3569_adj_348 ),
            .ltout(),
            .carryin(\eeprom.n3765 ),
            .carryout(\eeprom.n3766 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2357_20_lut_LC_16_19_2 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2357_20_lut_LC_16_19_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2357_20_lut_LC_16_19_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2357_20_lut_LC_16_19_2  (
            .in0(_gnd_net_),
            .in1(N__25316),
            .in2(N__27189),
            .in3(N__25280),
            .lcout(\eeprom.n3568_adj_347 ),
            .ltout(),
            .carryin(\eeprom.n3766 ),
            .carryout(\eeprom.n3767 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2357_21_lut_LC_16_19_3 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2357_21_lut_LC_16_19_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2357_21_lut_LC_16_19_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2357_21_lut_LC_16_19_3  (
            .in0(_gnd_net_),
            .in1(N__25277),
            .in2(N__27187),
            .in3(N__25244),
            .lcout(\eeprom.n3567_adj_341 ),
            .ltout(),
            .carryin(\eeprom.n3767 ),
            .carryout(\eeprom.n3768 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2357_22_lut_LC_16_19_4 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2357_22_lut_LC_16_19_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2357_22_lut_LC_16_19_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2357_22_lut_LC_16_19_4  (
            .in0(_gnd_net_),
            .in1(N__25241),
            .in2(N__27190),
            .in3(N__25202),
            .lcout(\eeprom.n3566_adj_340 ),
            .ltout(),
            .carryin(\eeprom.n3768 ),
            .carryout(\eeprom.n3769 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2357_23_lut_LC_16_19_5 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2357_23_lut_LC_16_19_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2357_23_lut_LC_16_19_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2357_23_lut_LC_16_19_5  (
            .in0(_gnd_net_),
            .in1(N__25198),
            .in2(N__27188),
            .in3(N__25769),
            .lcout(\eeprom.n3565_adj_338 ),
            .ltout(),
            .carryin(\eeprom.n3769 ),
            .carryout(\eeprom.n3770 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2357_24_lut_LC_16_19_6 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2357_24_lut_LC_16_19_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2357_24_lut_LC_16_19_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2357_24_lut_LC_16_19_6  (
            .in0(_gnd_net_),
            .in1(N__25762),
            .in2(N__27191),
            .in3(N__25727),
            .lcout(\eeprom.n3564_adj_337 ),
            .ltout(),
            .carryin(\eeprom.n3770 ),
            .carryout(\eeprom.n3771 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2357_25_lut_LC_16_19_7 .C_ON=1'b0;
    defparam \eeprom.rem_4_add_2357_25_lut_LC_16_19_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2357_25_lut_LC_16_19_7 .LUT_INIT=16'b1001000001100000;
    LogicCell40 \eeprom.rem_4_add_2357_25_lut_LC_16_19_7  (
            .in0(N__26998),
            .in1(N__25724),
            .in2(N__25706),
            .in3(N__25574),
            .lcout(\eeprom.n4765 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.add_938_2_lut_LC_16_20_0 .C_ON=1'b1;
    defparam \eeprom.add_938_2_lut_LC_16_20_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.add_938_2_lut_LC_16_20_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.add_938_2_lut_LC_16_20_0  (
            .in0(_gnd_net_),
            .in1(N__25877),
            .in2(_gnd_net_),
            .in3(N__25565),
            .lcout(\eeprom.n1353 ),
            .ltout(),
            .carryin(bfn_16_20_0_),
            .carryout(\eeprom.n3510 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.add_938_3_lut_LC_16_20_1 .C_ON=1'b1;
    defparam \eeprom.add_938_3_lut_LC_16_20_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.add_938_3_lut_LC_16_20_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.add_938_3_lut_LC_16_20_1  (
            .in0(_gnd_net_),
            .in1(N__25912),
            .in2(N__27185),
            .in3(N__25562),
            .lcout(\eeprom.n1352 ),
            .ltout(),
            .carryin(\eeprom.n3510 ),
            .carryout(\eeprom.n3511 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.add_938_4_lut_LC_16_20_2 .C_ON=1'b1;
    defparam \eeprom.add_938_4_lut_LC_16_20_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.add_938_4_lut_LC_16_20_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.add_938_4_lut_LC_16_20_2  (
            .in0(_gnd_net_),
            .in1(N__25559),
            .in2(_gnd_net_),
            .in3(N__25538),
            .lcout(\eeprom.n1351 ),
            .ltout(),
            .carryin(\eeprom.n3511 ),
            .carryout(\eeprom.n3512 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.add_938_5_lut_LC_16_20_3 .C_ON=1'b1;
    defparam \eeprom.add_938_5_lut_LC_16_20_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.add_938_5_lut_LC_16_20_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.add_938_5_lut_LC_16_20_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__25993),
            .in3(N__25535),
            .lcout(\eeprom.n1350 ),
            .ltout(),
            .carryin(\eeprom.n3512 ),
            .carryout(\eeprom.n3513 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.add_938_6_lut_LC_16_20_4 .C_ON=1'b1;
    defparam \eeprom.add_938_6_lut_LC_16_20_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.add_938_6_lut_LC_16_20_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.add_938_6_lut_LC_16_20_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__25532),
            .in3(N__25505),
            .lcout(\eeprom.n1349 ),
            .ltout(),
            .carryin(\eeprom.n3513 ),
            .carryout(\eeprom.n3514 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.add_938_7_lut_LC_16_20_5 .C_ON=1'b1;
    defparam \eeprom.add_938_7_lut_LC_16_20_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.add_938_7_lut_LC_16_20_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.add_938_7_lut_LC_16_20_5  (
            .in0(_gnd_net_),
            .in1(N__25501),
            .in2(_gnd_net_),
            .in3(N__25469),
            .lcout(\eeprom.n1348 ),
            .ltout(),
            .carryin(\eeprom.n3514 ),
            .carryout(\eeprom.n3515 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.add_938_8_lut_LC_16_20_6 .C_ON=1'b1;
    defparam \eeprom.add_938_8_lut_LC_16_20_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.add_938_8_lut_LC_16_20_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.add_938_8_lut_LC_16_20_6  (
            .in0(_gnd_net_),
            .in1(N__26057),
            .in2(_gnd_net_),
            .in3(N__26021),
            .lcout(\eeprom.n1347 ),
            .ltout(),
            .carryin(\eeprom.n3515 ),
            .carryout(\eeprom.n3516 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.add_938_9_lut_LC_16_20_7 .C_ON=1'b0;
    defparam \eeprom.add_938_9_lut_LC_16_20_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.add_938_9_lut_LC_16_20_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \eeprom.add_938_9_lut_LC_16_20_7  (
            .in0(N__26987),
            .in1(N__26018),
            .in2(_gnd_net_),
            .in3(N__26003),
            .lcout(\eeprom.n1346 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2447_3_lut_LC_16_21_1 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2447_3_lut_LC_16_21_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2447_3_lut_LC_16_21_1 .LUT_INIT=16'b0011000000111111;
    LogicCell40 \eeprom.rem_4_i2447_3_lut_LC_16_21_1  (
            .in0(_gnd_net_),
            .in1(N__26000),
            .in2(N__25834),
            .in3(N__25994),
            .lcout(\eeprom.n3715_adj_441 ),
            .ltout(\eeprom.n3715_adj_441_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i4068_1_lut_LC_16_21_2 .C_ON=1'b0;
    defparam \eeprom.i4068_1_lut_LC_16_21_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.i4068_1_lut_LC_16_21_2 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \eeprom.i4068_1_lut_LC_16_21_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__25961),
            .in3(_gnd_net_),
            .lcout(\eeprom.n4912 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i4083_2_lut_LC_16_21_3 .C_ON=1'b0;
    defparam \eeprom.i4083_2_lut_LC_16_21_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.i4083_2_lut_LC_16_21_3 .LUT_INIT=16'b0000111111111111;
    LogicCell40 \eeprom.i4083_2_lut_LC_16_21_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__25835),
            .in3(N__25948),
            .lcout(\eeprom.n3711_adj_456 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2449_3_lut_LC_16_21_4 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2449_3_lut_LC_16_21_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2449_3_lut_LC_16_21_4 .LUT_INIT=16'b0011001100001111;
    LogicCell40 \eeprom.rem_4_i2449_3_lut_LC_16_21_4  (
            .in0(_gnd_net_),
            .in1(N__25925),
            .in2(N__25919),
            .in3(N__25825),
            .lcout(\eeprom.n3717_adj_438 ),
            .ltout(\eeprom.n3717_adj_438_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i4062_1_lut_LC_16_21_5 .C_ON=1'b0;
    defparam \eeprom.i4062_1_lut_LC_16_21_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.i4062_1_lut_LC_16_21_5 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \eeprom.i4062_1_lut_LC_16_21_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__25892),
            .in3(_gnd_net_),
            .lcout(\eeprom.n4906 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2450_rep_1_3_lut_LC_16_21_6 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2450_rep_1_3_lut_LC_16_21_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2450_rep_1_3_lut_LC_16_21_6 .LUT_INIT=16'b0101010100110011;
    LogicCell40 \eeprom.rem_4_i2450_rep_1_3_lut_LC_16_21_6  (
            .in0(N__25883),
            .in1(N__25875),
            .in2(_gnd_net_),
            .in3(N__25824),
            .lcout(\eeprom.n4766 ),
            .ltout(\eeprom.n4766_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i4059_1_lut_LC_16_21_7 .C_ON=1'b0;
    defparam \eeprom.i4059_1_lut_LC_16_21_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.i4059_1_lut_LC_16_21_7 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \eeprom.i4059_1_lut_LC_16_21_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__26399),
            .in3(_gnd_net_),
            .lcout(\eeprom.n4903 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2022_2_lut_LC_16_23_0 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2022_2_lut_LC_16_23_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2022_2_lut_LC_16_23_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2022_2_lut_LC_16_23_0  (
            .in0(_gnd_net_),
            .in1(N__26386),
            .in2(_gnd_net_),
            .in3(N__26342),
            .lcout(\eeprom.n3086 ),
            .ltout(),
            .carryin(bfn_16_23_0_),
            .carryout(\eeprom.n3649 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2022_3_lut_LC_16_23_1 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2022_3_lut_LC_16_23_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2022_3_lut_LC_16_23_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2022_3_lut_LC_16_23_1  (
            .in0(_gnd_net_),
            .in1(N__26936),
            .in2(N__26335),
            .in3(N__26300),
            .lcout(\eeprom.n3085 ),
            .ltout(),
            .carryin(\eeprom.n3649 ),
            .carryout(\eeprom.n3650 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2022_4_lut_LC_16_23_2 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2022_4_lut_LC_16_23_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2022_4_lut_LC_16_23_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2022_4_lut_LC_16_23_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__26297),
            .in3(N__26252),
            .lcout(\eeprom.n3084 ),
            .ltout(),
            .carryin(\eeprom.n3650 ),
            .carryout(\eeprom.n3651 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2022_5_lut_LC_16_23_3 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2022_5_lut_LC_16_23_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2022_5_lut_LC_16_23_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2022_5_lut_LC_16_23_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__26249),
            .in3(N__26198),
            .lcout(\eeprom.n3083 ),
            .ltout(),
            .carryin(\eeprom.n3651 ),
            .carryout(\eeprom.n3652 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2022_6_lut_LC_16_23_4 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2022_6_lut_LC_16_23_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2022_6_lut_LC_16_23_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2022_6_lut_LC_16_23_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__26195),
            .in3(N__26153),
            .lcout(\eeprom.n3082 ),
            .ltout(),
            .carryin(\eeprom.n3652 ),
            .carryout(\eeprom.n3653 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2022_7_lut_LC_16_23_5 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2022_7_lut_LC_16_23_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2022_7_lut_LC_16_23_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2022_7_lut_LC_16_23_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__26150),
            .in3(N__26099),
            .lcout(\eeprom.n3081 ),
            .ltout(),
            .carryin(\eeprom.n3653 ),
            .carryout(\eeprom.n3654 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2022_8_lut_LC_16_23_6 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2022_8_lut_LC_16_23_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2022_8_lut_LC_16_23_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2022_8_lut_LC_16_23_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__26096),
            .in3(N__26060),
            .lcout(\eeprom.n3080 ),
            .ltout(),
            .carryin(\eeprom.n3654 ),
            .carryout(\eeprom.n3655 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2022_9_lut_LC_16_23_7 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2022_9_lut_LC_16_23_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2022_9_lut_LC_16_23_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2022_9_lut_LC_16_23_7  (
            .in0(_gnd_net_),
            .in1(N__26937),
            .in2(N__26705),
            .in3(N__26675),
            .lcout(\eeprom.n3079 ),
            .ltout(),
            .carryin(\eeprom.n3655 ),
            .carryout(\eeprom.n3656 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2022_10_lut_LC_16_24_0 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2022_10_lut_LC_16_24_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2022_10_lut_LC_16_24_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2022_10_lut_LC_16_24_0  (
            .in0(_gnd_net_),
            .in1(N__26672),
            .in2(N__27073),
            .in3(N__26642),
            .lcout(\eeprom.n3078 ),
            .ltout(),
            .carryin(bfn_16_24_0_),
            .carryout(\eeprom.n3657 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2022_11_lut_LC_16_24_1 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2022_11_lut_LC_16_24_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2022_11_lut_LC_16_24_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2022_11_lut_LC_16_24_1  (
            .in0(_gnd_net_),
            .in1(N__26885),
            .in2(N__26634),
            .in3(N__26597),
            .lcout(\eeprom.n3077 ),
            .ltout(),
            .carryin(\eeprom.n3657 ),
            .carryout(\eeprom.n3658 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2022_12_lut_LC_16_24_2 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2022_12_lut_LC_16_24_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2022_12_lut_LC_16_24_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2022_12_lut_LC_16_24_2  (
            .in0(_gnd_net_),
            .in1(N__26586),
            .in2(N__27074),
            .in3(N__26546),
            .lcout(\eeprom.n3076 ),
            .ltout(),
            .carryin(\eeprom.n3658 ),
            .carryout(\eeprom.n3659 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2022_13_lut_LC_16_24_3 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2022_13_lut_LC_16_24_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2022_13_lut_LC_16_24_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2022_13_lut_LC_16_24_3  (
            .in0(_gnd_net_),
            .in1(N__26538),
            .in2(N__27077),
            .in3(N__26516),
            .lcout(\eeprom.n3075 ),
            .ltout(),
            .carryin(\eeprom.n3659 ),
            .carryout(\eeprom.n3660 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2022_14_lut_LC_16_24_4 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2022_14_lut_LC_16_24_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2022_14_lut_LC_16_24_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2022_14_lut_LC_16_24_4  (
            .in0(_gnd_net_),
            .in1(N__26511),
            .in2(N__27075),
            .in3(N__26471),
            .lcout(\eeprom.n3074 ),
            .ltout(),
            .carryin(\eeprom.n3660 ),
            .carryout(\eeprom.n3661 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2022_15_lut_LC_16_24_5 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2022_15_lut_LC_16_24_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2022_15_lut_LC_16_24_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2022_15_lut_LC_16_24_5  (
            .in0(_gnd_net_),
            .in1(N__26467),
            .in2(N__27078),
            .in3(N__26429),
            .lcout(\eeprom.n3073 ),
            .ltout(),
            .carryin(\eeprom.n3661 ),
            .carryout(\eeprom.n3662 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2022_16_lut_LC_16_24_6 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2022_16_lut_LC_16_24_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2022_16_lut_LC_16_24_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2022_16_lut_LC_16_24_6  (
            .in0(_gnd_net_),
            .in1(N__26426),
            .in2(N__27076),
            .in3(N__28076),
            .lcout(\eeprom.n3072 ),
            .ltout(),
            .carryin(\eeprom.n3662 ),
            .carryout(\eeprom.n3663 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2022_17_lut_LC_16_24_7 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2022_17_lut_LC_16_24_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2022_17_lut_LC_16_24_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2022_17_lut_LC_16_24_7  (
            .in0(_gnd_net_),
            .in1(N__28073),
            .in2(N__27079),
            .in3(N__28037),
            .lcout(\eeprom.n3071 ),
            .ltout(),
            .carryin(\eeprom.n3663 ),
            .carryout(\eeprom.n3664 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2022_18_lut_LC_16_25_0 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2022_18_lut_LC_16_25_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2022_18_lut_LC_16_25_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2022_18_lut_LC_16_25_0  (
            .in0(_gnd_net_),
            .in1(N__28034),
            .in2(N__26880),
            .in3(N__27998),
            .lcout(\eeprom.n3070 ),
            .ltout(),
            .carryin(bfn_16_25_0_),
            .carryout(\eeprom.n3665 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2022_19_lut_LC_16_25_1 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2022_19_lut_LC_16_25_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2022_19_lut_LC_16_25_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2022_19_lut_LC_16_25_1  (
            .in0(_gnd_net_),
            .in1(N__27995),
            .in2(N__26881),
            .in3(N__27950),
            .lcout(\eeprom.n3069 ),
            .ltout(),
            .carryin(\eeprom.n3665 ),
            .carryout(\eeprom.n3666 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2022_20_lut_LC_16_25_2 .C_ON=1'b0;
    defparam \eeprom.rem_4_add_2022_20_lut_LC_16_25_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2022_20_lut_LC_16_25_2 .LUT_INIT=16'b1001000001100000;
    LogicCell40 \eeprom.rem_4_add_2022_20_lut_LC_16_25_2  (
            .in0(N__26764),
            .in1(N__27947),
            .in2(N__27920),
            .in3(N__27809),
            .lcout(\eeprom.n3100 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam CONSTANT_ONE_LUT4_LC_16_26_0.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_16_26_0.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_16_26_0.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_16_26_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
endmodule // TinyFPGA_B
