// Verilog netlist produced by program LSE :  version Diamond Version 0.0.0
// Netlist written on Fri Feb 28 12:45:14 2020
//
// Verilog Description of module TinyFPGA_B
//

module TinyFPGA_B (CLK, LED, USBPU, ENCODER0_A, ENCODER0_B, ENCODER1_A, 
            ENCODER1_B, HALL1, HALL2, HALL3, FAULT_N, NEOPXL, DE, 
            TX, RX, CS_CLK, CS, CS_MISO, SCL, SDA, INLC, INHC, 
            INLB, INHB, INLA, INHA) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(2[8:18])
    input CLK;   // verilog/TinyFPGA_B.v(3[9:12])
    output LED;   // verilog/TinyFPGA_B.v(4[10:13])
    output USBPU;   // verilog/TinyFPGA_B.v(5[10:15])
    input ENCODER0_A;   // verilog/TinyFPGA_B.v(6[9:19])
    input ENCODER0_B;   // verilog/TinyFPGA_B.v(7[9:19])
    input ENCODER1_A;   // verilog/TinyFPGA_B.v(8[9:19])
    input ENCODER1_B;   // verilog/TinyFPGA_B.v(9[9:19])
    input HALL1 /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(10[9:14])
    input HALL2 /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(11[9:14])
    input HALL3 /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(12[9:14])
    input FAULT_N;   // verilog/TinyFPGA_B.v(13[9:16])
    output NEOPXL;   // verilog/TinyFPGA_B.v(14[10:16])
    output DE;   // verilog/TinyFPGA_B.v(15[10:12])
    output TX /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(16[10:12])
    input RX;   // verilog/TinyFPGA_B.v(17[9:11])
    output CS_CLK;   // verilog/TinyFPGA_B.v(18[10:16])
    output CS;   // verilog/TinyFPGA_B.v(19[10:12])
    input CS_MISO;   // verilog/TinyFPGA_B.v(20[9:16])
    inout SCL /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(21[9:12])
    inout SDA /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(22[9:12])
    output INLC;   // verilog/TinyFPGA_B.v(23[10:14])
    output INHC;   // verilog/TinyFPGA_B.v(24[10:14])
    output INLB;   // verilog/TinyFPGA_B.v(25[10:14])
    output INHB;   // verilog/TinyFPGA_B.v(26[10:14])
    output INLA;   // verilog/TinyFPGA_B.v(27[10:14])
    output INHA;   // verilog/TinyFPGA_B.v(28[10:14])
    
    wire clk16MHz /* synthesis SET_AS_NETWORK=clk16MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[16:24])
    
    wire GND_net, VCC_net, LED_c, ENCODER0_A_N, ENCODER0_B_N, ENCODER1_A_N, 
        ENCODER1_B_N, NEOPXL_c, DE_c, RX_c, CS_CLK_c, CS_c, CS_MISO_c, 
        INLC_c_0, INHC_c_0, INLB_c_0, INHB_c_0, INLA_c_0, INHA_c_0;
    wire [7:0]ID;   // verilog/TinyFPGA_B.v(46[11:13])
    wire [23:0]neopxl_color;   // verilog/TinyFPGA_B.v(48[13:25])
    
    wire hall1, hall2, hall3, pwm_out, dir, GHA, n44069, GHB, 
        GHC;
    wire [23:0]pwm_setpoint;   // verilog/TinyFPGA_B.v(94[20:32])
    wire [23:0]duty;   // verilog/TinyFPGA_B.v(95[21:25])
    wire [7:0]commutation_state;   // verilog/TinyFPGA_B.v(131[12:29])
    wire [7:0]commutation_state_prev;   // verilog/TinyFPGA_B.v(132[12:34])
    
    wire dti;
    wire [7:0]dti_counter;   // verilog/TinyFPGA_B.v(141[12:23])
    
    wire tx_o, tx_enable;
    wire [23:0]encoder0_position_scaled;   // verilog/TinyFPGA_B.v(238[21:45])
    wire [23:0]encoder1_position_scaled;   // verilog/TinyFPGA_B.v(240[21:45])
    wire [23:0]displacement;   // verilog/TinyFPGA_B.v(241[21:33])
    wire [23:0]setpoint;   // verilog/TinyFPGA_B.v(242[22:30])
    wire [23:0]Kp;   // verilog/TinyFPGA_B.v(243[22:24])
    wire [23:0]Ki;   // verilog/TinyFPGA_B.v(244[22:24])
    
    wire n43614, n44068, n44067, n44066, n44065;
    wire [7:0]control_mode;   // verilog/TinyFPGA_B.v(246[14:26])
    wire [23:0]PWMLimit;   // verilog/TinyFPGA_B.v(247[22:30])
    wire [23:0]IntegralLimit;   // verilog/TinyFPGA_B.v(248[22:35])
    wire [23:0]deadband;   // verilog/TinyFPGA_B.v(249[22:30])
    wire [15:0]current;   // verilog/TinyFPGA_B.v(250[22:29])
    
    wire n15;
    wire [15:0]current_limit;   // verilog/TinyFPGA_B.v(251[22:35])
    wire [23:0]motor_state;   // verilog/TinyFPGA_B.v(280[22:33])
    
    wire n44064, n29524, n29523, n6;
    wire [7:0]data;   // verilog/TinyFPGA_B.v(337[14:18])
    
    wire data_ready, sda_out, sda_enable, scl, scl_enable;
    wire [31:0]delay_counter;   // verilog/TinyFPGA_B.v(361[11:24])
    
    wire read;
    wire [2:0]\ID_READOUT_FSM.state ;   // verilog/TinyFPGA_B.v(369[15:20])
    
    wire pwm_setpoint_23__N_263, n209, n211, n249, n250, n251, n252, 
        n253, n254, n255, n256, n257, n258, n259, n260, n261, 
        n262, n263, n264, n265, n266, n267, n268, n269, n270, 
        n55695, n296, n44063, n44062, n55694, n330, n334, n335, 
        n336, n337, n338, n339, n340, n341, n342, n343, n344, 
        n345, n8;
    wire [31:0]encoder0_position;   // verilog/TinyFPGA_B.v(237[11:28])
    
    wire n356, n379, n44061, n44060, n418, n419, n420, n421, 
        n422, n423, n424, n425, n426, n427, n428, n429, n430, 
        n431, n432, n433, n434, n435, n436, n437, n438, n439, 
        n440, n441, n7;
    wire [23:0]pwm_setpoint_23__N_11;
    
    wire n43613;
    wire [7:0]commutation_state_7__N_264;
    
    wire commutation_state_7__N_272, n29522, n29521;
    wire [31:0]encoder1_position;   // verilog/TinyFPGA_B.v(239[11:28])
    
    wire n43612, n4, n50654, GHA_N_478, GLA_N_495, GHB_N_500, GLB_N_509, 
        GHC_N_514, GLC_N_523, dti_N_527, n29520, n29519, n29518, 
        n29516, n29515, RX_N_10;
    wire [31:0]motor_state_23__N_123;
    wire [31:0]encoder0_position_scaled_23__N_327;
    wire [32:0]encoder0_position_scaled_23__N_51;
    
    wire encoder1_position_scaled_23__N_359;
    wire [31:0]encoder1_position_scaled_23__N_75;
    wire [23:0]displacement_23__N_99;
    
    wire n2274, n43610, n43611, n44059, n43558, n44058, n37376, 
        n44057, n1532, n1533, n1534, n1535, n1536, n1537, n1538, 
        n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, 
        n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, 
        n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, 
        n1563, n44056, n55625, n55623, n55622, n8581, n8582, n8583, 
        n8584, n1650, n8585, n8586, n51321, n56688, n56676, n2091, 
        n2233;
    wire [31:0]timer;   // verilog/neopixel.v(9[12:17])
    wire [3:0]state;   // verilog/neopixel.v(16[20:25])
    wire [31:0]\neo_pixel_transmitter.t0 ;   // verilog/neopixel.v(28[14:16])
    
    wire n27100, n5, n50932, n44055;
    wire [3:0]state_3__N_639;
    
    wire n44054, n56814, n56808, n56802, n29514, n21005, n7936, 
        n50148, n4929, n29513, n29512, n29511, n29510, n29509, 
        n29508, n4928, n4927, n44053, n56862, n53125, n4_adj_5443, 
        n4926, n4925, n4924, n4923, n4922, n4921, n4920, n4919, 
        n4918, n4917, n4916, n4915, n4914, n29507, n29506, n44052, 
        n625, n623, n622, n621, n10, n44051, n4913, n29505, 
        n29504, n29503, n29502, n29501, n29500, n4_adj_5444, n415, 
        n414, n413, n412, n411, n407, n29499, n4748, n4_adj_5445, 
        n44050, n44049, n3, n4_adj_5446, n5_adj_5447, n6_adj_5448, 
        n7_adj_5449, n8_adj_5450, n9, n10_adj_5451, n11, n12, n13, 
        n14, n15_adj_5452, n16, n17, n18, n19, n20, n21, n22, 
        n23, n24, n25, n2, n29498, n14_adj_5453, n15_adj_5454, 
        n16_adj_5455, n17_adj_5456, n18_adj_5457, n19_adj_5458, n20_adj_5459, 
        n21_adj_5460, n22_adj_5461, n23_adj_5462, n24_adj_5463, n25_adj_5464, 
        n27093, n29497, n29496, rx_data_ready;
    wire [7:0]rx_data;   // verilog/coms.v(92[13:20])
    wire [7:0]\data_in[3] ;   // verilog/coms.v(96[12:19])
    wire [7:0]\data_in[2] ;   // verilog/coms.v(96[12:19])
    wire [7:0]\data_in[1] ;   // verilog/coms.v(96[12:19])
    wire [7:0]\data_in[0] ;   // verilog/coms.v(96[12:19])
    wire [7:0]\data_in_frame[21] ;   // verilog/coms.v(97[12:25])
    wire [7:0]\data_in_frame[20] ;   // verilog/coms.v(97[12:25])
    wire [7:0]\data_in_frame[16] ;   // verilog/coms.v(97[12:25])
    wire [7:0]\data_in_frame[15] ;   // verilog/coms.v(97[12:25])
    wire [7:0]\data_in_frame[14] ;   // verilog/coms.v(97[12:25])
    wire [7:0]\data_in_frame[13] ;   // verilog/coms.v(97[12:25])
    wire [7:0]\data_in_frame[12] ;   // verilog/coms.v(97[12:25])
    wire [7:0]\data_in_frame[11] ;   // verilog/coms.v(97[12:25])
    wire [7:0]\data_in_frame[10] ;   // verilog/coms.v(97[12:25])
    wire [7:0]\data_in_frame[9] ;   // verilog/coms.v(97[12:25])
    wire [7:0]\data_in_frame[8] ;   // verilog/coms.v(97[12:25])
    wire [7:0]\data_in_frame[5] ;   // verilog/coms.v(97[12:25])
    wire [7:0]\data_in_frame[4] ;   // verilog/coms.v(97[12:25])
    wire [7:0]\data_in_frame[3] ;   // verilog/coms.v(97[12:25])
    wire [7:0]\data_in_frame[2] ;   // verilog/coms.v(97[12:25])
    wire [7:0]\data_in_frame[1] ;   // verilog/coms.v(97[12:25])
    wire [7:0]\data_out_frame[25] ;   // verilog/coms.v(98[12:26])
    wire [7:0]\data_out_frame[24] ;   // verilog/coms.v(98[12:26])
    wire [7:0]\data_out_frame[23] ;   // verilog/coms.v(98[12:26])
    wire [7:0]\data_out_frame[22] ;   // verilog/coms.v(98[12:26])
    wire [7:0]\data_out_frame[21] ;   // verilog/coms.v(98[12:26])
    wire [7:0]\data_out_frame[20] ;   // verilog/coms.v(98[12:26])
    wire [7:0]\data_out_frame[19] ;   // verilog/coms.v(98[12:26])
    wire [7:0]\data_out_frame[18] ;   // verilog/coms.v(98[12:26])
    wire [7:0]\data_out_frame[17] ;   // verilog/coms.v(98[12:26])
    wire [7:0]\data_out_frame[16] ;   // verilog/coms.v(98[12:26])
    wire [7:0]\data_out_frame[15] ;   // verilog/coms.v(98[12:26])
    wire [7:0]\data_out_frame[14] ;   // verilog/coms.v(98[12:26])
    wire [7:0]\data_out_frame[13] ;   // verilog/coms.v(98[12:26])
    wire [7:0]\data_out_frame[12] ;   // verilog/coms.v(98[12:26])
    wire [7:0]\data_out_frame[11] ;   // verilog/coms.v(98[12:26])
    wire [7:0]\data_out_frame[10] ;   // verilog/coms.v(98[12:26])
    wire [7:0]\data_out_frame[9] ;   // verilog/coms.v(98[12:26])
    wire [7:0]\data_out_frame[8] ;   // verilog/coms.v(98[12:26])
    wire [7:0]\data_out_frame[7] ;   // verilog/coms.v(98[12:26])
    wire [7:0]\data_out_frame[6] ;   // verilog/coms.v(98[12:26])
    wire [7:0]\data_out_frame[5] ;   // verilog/coms.v(98[12:26])
    wire [7:0]\data_out_frame[4] ;   // verilog/coms.v(98[12:26])
    
    wire n24210, tx_active;
    wire [31:0]\FRAME_MATCHER.state ;   // verilog/coms.v(113[11:16])
    
    wire n44048, n122, n43542, n19602, n44047, n44046, n44045, 
        n44044, n44043, n43557, n44042, n43556, n44041, n44040, 
        n44039, n44038, n44037, n44036, n44035, n44034, n4912, 
        n4911, n29495, n29494, n44033, n44032, n44031, n44030, 
        n44029, n44028, n44027, n44026, n44025, n44024, n44023, 
        n44022, n44021, n44020, n44019, n44018, n44017, n44016, 
        n44015, n44014, n56784, n56778, n56772, n56766, n56760, 
        n56754, n44013, n44012, n44011, n44010, n44009, n44447, 
        n44446, n44008, n44445, n44444, n44007, n44443, n44442, 
        n44006, n44005, n44004, n44441, n44440, n44439, n44003, 
        n44002, n44438, n44001, n44437, n44000, n44436, n43999, 
        n44435, n44434, n44433, n43998, n43997, n43996, n44432, 
        n44431, n44430, n43995, n43994, n44429, n43993, n44428, 
        n44427, n44426, n43992, n544, n543, n542, n541, n540, 
        n539, n538, n537, n536, n535, n534, n533, n43991, n44425, 
        n43990, n44424, n43989, n43988, n44423, n24_adj_5465, n20_adj_5466, 
        n15_adj_5467, n14_adj_5468, n55624, n55141, n43987, n43986, 
        n44422, n44421, n44420, n44419, n43985, n44418, n43984, 
        n44417, n56086, n44416, n44415, n43983, n43982, n44414, 
        n56233, n32464, n44413, n43981, n43980, n44412, n44411, 
        n44410, n44409, n43979, n44408, n43978, n44407, n44406, 
        n43977, n43541, n37372, n44405, n44404, n43976, n44403, 
        n44402, n44401, n44400, n43975, n44399, n44398, n43974, 
        n44397, n44396, n43973, n43972, n37186, n37346, n44395, 
        n44394, n43971, n43970, n43969, n44393, n44392, n43968, 
        n44391, n43967, n43966, n43965, n44390, n44389, n37342, 
        n43964, n44388, n37340, n37338, n44387, n44386, n43963, 
        n43962, n44385, n44384, n44383, n44382, n44381, n44380, 
        n44379, n44378, n43555, n44377, n44376, n37334, n44375, 
        n44374, n44373, n44372, n43954, n44371, n44370, n43953, 
        n44369, n44368, n43554, n43952, n44367, n37328, n44366, 
        n44365, n44364, n44363, n44362, n43951, n44361, n44360, 
        n43950, n44359, n43949, n4_adj_5469, n532, n29493, n29492, 
        n43948, n44358, n531, n530, n529, n29491, n27198, n29490, 
        n44357, n43947, n3303;
    wire [31:0]\FRAME_MATCHER.state_31__N_3007 ;
    
    wire n44356, n43946, n44355, n43945, n44354, n43944, n44353, 
        n44352, n44351, n37316, n44350, n44349, n43943, n43942, 
        n43941, n43940, n44348, n44347, n43939, n44346, n44345, 
        n43540, n43938, n43553, n37382, n37308, n37306, n44344, 
        n44343, n44342, n43937, n44341, n43936, n44340, n43935, 
        n44339, n44338, n44337, n44336, n43934, n44335, n44334, 
        n44333, n37302, n44332, n37298, n44331, n43539, n43933, 
        n44330, n44329, n44328, n43932, n44327, n44326, n44325, 
        n44324, n44323, n44322, n44321, n44320, n44319, n44318, 
        n44317, n44316, n44315, n44314, n44313, n44312, n44311, 
        n44310, n44309, n37296, n44308, n44307, n44306, n44305, 
        n44304, n27219, n44303, n15_adj_5470, n44302, n29486, n44301, 
        n44300, n44299, n56498, n44298, n44297, n44296, n44295, 
        n44294, n44293, n44292, n44291, n44290, n44289, n44288, 
        n44287, n44286, n44285, n44284, n44283, n44282, n44281, 
        n36544, n36542, n55009, n44280, n44279, n44278, n44277, 
        n43922, n44276, n44275, n44274, n43921, n44273, n43920, 
        n55005, n44272, n44271, n44270, n44269, n44268, n43919, 
        n44267, n43918, n44266, n43917, n43916, n44265, n44264, 
        n43915, n44263, n43914, n43913, n44262, n43912, n44261, 
        n44260, n44259, n43911, n43538, n36528, n55003, n44258, 
        n54995, n37482, n43910, n43909, n44257, n44256, n43908, 
        n44255, n44254, n44253, n43907, n43906, n43905, n44252, 
        n43904, n43552, n44251, n43903, n44250, n44249, n50003, 
        n49995, n43902, n43901, n44248, n43900, n43899, n44247, 
        n43898, n44246, n44245, n44244, n43551, n49998, n43897, 
        n44243, n43896, n44242, n43895, n44241, n43894, n36556, 
        n36554, n54989, n36436, n54987, n54975, n29485, n29484, 
        n43893, n44240, n43892, n44239, n43891, n43890, n43889, 
        n44238, n516, n29483, n29482, n29481, n29480, n29479, 
        n29478, n29477, n29476, n15_adj_5471, n49919, n51223, n49779, 
        n36659, n4_adj_5472, n4_adj_5473, n49757, n49755, n49753, 
        n49751, n49748, n33, n32, n31, n30, n29, n28, n27, 
        n26, n25_adj_5474, n24_adj_5475, n23_adj_5476, n22_adj_5477, 
        n21_adj_5478, n20_adj_5479, n19_adj_5480, n18_adj_5481, n17_adj_5482, 
        n16_adj_5483, n15_adj_5484, n14_adj_5485, n13_adj_5486, n12_adj_5487, 
        n11_adj_5488, n10_adj_5489, n9_adj_5490, n8_adj_5491, n7_adj_5492, 
        n6_adj_5493, n5_adj_5494, n4_adj_5495, n3_adj_5496, n2_adj_5497, 
        n44237, n27232, n25_adj_5498, n24_adj_5499, n23_adj_5500, 
        n22_adj_5501, n21_adj_5502, n20_adj_5503, n19_adj_5504, n18_adj_5505, 
        n17_adj_5506, n16_adj_5507, n15_adj_5508, n14_adj_5509, n13_adj_5510, 
        n12_adj_5511, n11_adj_5512, n10_adj_5513, n9_adj_5514, n8_adj_5515, 
        n7_adj_5516, n6_adj_5517, n5_adj_5518, n4_adj_5519, n3_adj_5520, 
        n2_adj_5521, n14_adj_5522, n43888, n43887, n44236, n2573, 
        n48558, n44235, n43886, n30067, n30066, n44234, n30059, 
        n30058, n30057, n30056, n30055, n30054, n6272, n30053, 
        n30052, n30051, n30050, n30049, n30048, n30047, n6_adj_5523, 
        n30046, n30045, n30044, n44233, n30043, n44232, n30042, 
        n30041, n30040, n30039, n30038, n30037, n5_adj_5524, n30036, 
        n30035, n30034, n30033, n30032, n30031, n30030, n30029, 
        n44231, n49749, n43885, n44230, n43884, n43883, n43882, 
        n44229, n43881, n43880, n43879, n44228, n44227, n30028, 
        control_update;
    wire [23:0]\PID_CONTROLLER.integral ;   // verilog/motorControl.v(35[23:31])
    
    wire n30027, n30026, n30025, n30024, n29472, n29471, n30023, 
        n30022, n29470, n44226, n29469, n29468, n29467, n29466, 
        n29465, n30021, n30020;
    wire [23:0]\PID_CONTROLLER.integral_23__N_3996 ;
    
    wire n363, n40, n32_adj_5525, n44225, n44224;
    wire [1:0]a_new;   // vhdl/quadrature_decoder.vhd(39[9:14])
    
    wire b_prev, n30019, n30018, n30017, n30016, n44223, n30015, 
        position_31__N_4108, n30014, n30013, n30012, n30011, n30010, 
        n30009, n30008, n30007, n30006, n30005, n30004, n30003, 
        n24553, n30002, n30001, n30000, n29999, n29998, n29997, 
        n29996, n29995, n29994, n29993, n29992, n29991, n4910, 
        n4909, n4908, n4907, n4906, n4904, n4903, n4902, n4901, 
        n4900, n4899, n4898, n4897, n4896, n4895, n4894, n4893, 
        n4892, n4891, n4890, n4889, n4888, n4887, n4886, n4885, 
        n4884, n4883, n29990, n29989, n29988, n29464, n29987, 
        n29463, n29986, n29985, n29984, n29983, n29982, n29981, 
        n29980, n29979, n29978;
    wire [1:0]a_new_adj_5692;   // vhdl/quadrature_decoder.vhd(39[9:14])
    
    wire b_prev_adj_5527, n29977, n29976, n29975, n29974, n29973, 
        position_31__N_4108_adj_5528, n29972, n29971, n29970, n29969, 
        n29968, n29967, n14_adj_5529, n50075, n29962, n29961, n29960, 
        n29959, n29958, n29957, n29956, n10_adj_5530, n29955, n29954, 
        n29953, n29952, n29951, n29950, n29949, n29948, n29947, 
        n29946, n29945, n29944, n29462, n29280, n29461, n29460, 
        n29943, n29942, n29941, n44222, n29940, n50770, rw;
    wire [7:0]state_adj_5705;   // verilog/eeprom.v(23[11:16])
    
    wire n43664, n44221, n29939, n29938, n29937, n29936, n29935, 
        n29934, n19_adj_5533, n17_adj_5534, n16_adj_5535, n15_adj_5536, 
        n13_adj_5537, n11_adj_5538, n9_adj_5539, n8_adj_5540, n7_adj_5541, 
        n6_adj_5542, n5_adj_5543, n4_adj_5544, n29933, clk_out;
    wire [15:0]data_adj_5711;   // verilog/tli4970.v(27[14:18])
    
    wire n29932, n29931, n29930;
    wire [7:0]state_adj_5713;   // verilog/tli4970.v(29[13:18])
    
    wire n29929, n29928, n29927, n29456, n29455, n29454, n29453, 
        n29926, n4_adj_5555, n28885, n29925, n29923, n29922, n29921, 
        n43550, n44220, n63, n6_adj_5556, n29920, n29919, n29918, 
        n29916, n29915, n29914, n29913, n29912, n29911, n29910, 
        n29909, n29908, n29907, n29906, n29905, n29904, n29903, 
        n29902, n50822, n44219, n44218, n43663, n29901, n29900, 
        n29899, n50825, n43662, n5_adj_5557, n29898, n29897, n29896, 
        n29895, n29894, n29893, state_7__N_4499, n29892, n29452, 
        n29451, n29450, n29891, n29890, n29889, n29888, n29887, 
        n29886, n29885, n29884, n29883, n29882, n29881, n29880, 
        n29879, n29878, n29877, n24_adj_5558, n55782, n19_adj_5559, 
        n17_adj_5560, n16_adj_5561, n15_adj_5562, n29876, n24_adj_5563, 
        n55778, n19_adj_5564, n17_adj_5565, n16_adj_5566, n15_adj_5567, 
        n13_adj_5568, n50836, r_Rx_Data;
    wire [2:0]r_Bit_Index;   // verilog/uart_rx.v(33[17:28])
    wire [2:0]r_SM_Main;   // verilog/uart_rx.v(36[17:26])
    
    wire n29874, n28852, n29873, n29872, n29871, n29870, n29869, 
        n29868, n29867, n29866, n29865, n43661, n44217, n29864, 
        n29863, n44216, n43660, n43537, n29862, n29449, n29861, 
        n11_adj_5569, n9_adj_5570;
    wire [2:0]r_SM_Main_2__N_3777;
    
    wire n29860, n29448, n29856, n29850, n29849, n29845;
    wire [2:0]r_SM_Main_adj_5723;   // verilog/uart_tx.v(31[16:25])
    wire [2:0]r_Bit_Index_adj_5725;   // verilog/uart_tx.v(33[16:27])
    wire [2:0]r_SM_Main_2__N_3848;
    
    wire n26_adj_5575, n29842, n29447, n28848, n43549, n29839, n29838, 
        n29835, n29834, n29833, n29832, n29831, n29830, n29829, 
        n29827, n29826, n29825, n29824, n29823, n29821, n29820, 
        n29446;
    wire [7:0]state_adj_5736;   // verilog/i2c_controller.v(33[12:17])
    
    wire n29819, n29818;
    wire [7:0]saved_addr;   // verilog/i2c_controller.v(34[12:22])
    
    wire n29445, n29817, n29816, enable_slow_N_4393, n29815, n7_adj_5577, 
        n43659, n43578, n29814, n43658;
    wire [7:0]state_7__N_4290;
    
    wire n8_adj_5578, n7_adj_5579, n6_adj_5580, n5_adj_5581, n29813, 
        n29444, n7354, n29812, n29811, n29443, n43657, n29810, 
        n29809, n29808, n29807, n29806, n29805, n29804;
    wire [7:0]state_7__N_4306;
    
    wire n29442, n29803, n44215, n29802, n29801, n29800, n29799, 
        n29798, n29797, n29796, n29145, n13_adj_5582, n11_adj_5583, 
        n9_adj_5584, n8_adj_5585, n7_adj_5586, n6_adj_5587, n29795, 
        n5_adj_5588, n29794, n29793, n29441, n29440, n29439, n29438, 
        n29437, n29436, n29435, n29434, n4_adj_5589, n29792, n4_adj_5590, 
        n7974, n29791, n29790, n29789, n44214, n29788, n29433, 
        n29432, n29431, n29430, n29429, n29428, n29427, n29426, 
        n29425, n29424, n29423, n29785, n29422, n29784, n29783, 
        n29782, n10_adj_5591, n29352, n29759, n29758, n44213, n7593, 
        n44212, n29421, n51078, n834, n833, n832, n831, n830, 
        n829, n828, n28778, n861, n29420, n896, n897, n898, 
        n899, n900, n901, n927, n928, n929, n930, n931, n932, 
        n933, n934, n935, n29419, n941, n942, n44211, n44210, 
        n960, n51149, n49720, n56736, n995, n996, n997, n998, 
        n999, n1000, n1001, n1026, n1027, n1028, n1029, n1030, 
        n1031, n1032, n1033, n1059, n1093, n1094, n1095, n1096, 
        n1097, n1098, n1099, n1100, n1101, n51076, n1125, n1126, 
        n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1158, 
        n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, 
        n1201, n1224, n1225, n1226, n1227, n1228, n1229, n1230, 
        n1231, n1232, n1233, n1257, n1292, n1293, n1294, n1295, 
        n1296, n1297, n1298, n1299, n1300, n1301, n1323, n1324, 
        n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, 
        n1333, n1356, n50741, n40_adj_5592, n21_adj_5593, n1391, 
        n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, 
        n1400, n1401, n1422, n1423, n1424, n1425, n1426, n1427, 
        n1428, n1429, n1430, n1431, n1432, n1433, n1455, n5_adj_5594, 
        n56730, n1490, n1491, n1492, n1493, n1494, n1495, n1496, 
        n1497, n1498, n1499, n1500, n1501, n1521, n1522, n1523, 
        n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, 
        n1532_adj_5595, n1533_adj_5596, n1554_adj_5597, n1589, n1590, 
        n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, 
        n1599, n1600, n1601, n1620, n1621, n1622, n1623, n1624, 
        n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, 
        n1633, n29418, n1653, n1688, n1689, n1690, n1691, n1692, 
        n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, 
        n1701, n1719, n1720, n1721, n1722, n1723, n1724, n1725, 
        n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, 
        n44209, n43656, n1752, n1787, n1788, n1789, n1790, n1791, 
        n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, 
        n1800, n1801, n1818, n1819, n1820, n1821, n1822, n1823, 
        n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, 
        n1832, n1833, n56328, n1851, n56724, n1886, n1887, n1888, 
        n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, 
        n1897, n1898, n1899, n1900, n1901, n1917, n1918, n1919, 
        n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, 
        n1928, n1929, n1930, n1931, n1932, n1933, n1950, n1985, 
        n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, 
        n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, 
        n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, 
        n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, 
        n2032, n2033, n2049, n48957, n2084, n2085, n2086, n2087, 
        n2088, n2089, n2090, n2091_adj_5598, n2092, n2093, n2094, 
        n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2115, 
        n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, 
        n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, 
        n2132, n2133, n2148, n43655, n44208, n44207, n43654, n2183, 
        n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, 
        n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, 
        n2200, n2201, n43577, n2214, n2215, n2216, n2217, n2218, 
        n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, 
        n2227, n2228, n2229, n2230, n2231, n2232, n2233_adj_5599, 
        n56237, n2247, n56718, n2282, n2283, n2284, n2285, n2286, 
        n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, 
        n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2313, 
        n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, 
        n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, 
        n2330, n2331, n2332, n2333, n2346, n2381, n2382, n2383, 
        n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, 
        n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, 
        n2400, n2401, n2412, n2413, n2414, n2415, n2416, n2417, 
        n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, 
        n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, 
        n56595, n2445, n2480, n2481, n2482, n2483, n2484, n2485, 
        n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, 
        n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, 
        n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, 
        n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526, 
        n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2544, 
        n44206, n2579, n2580, n2581, n2582, n2583, n2584, n2585, 
        n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, 
        n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, 
        n28753, n2610, n2611, n2612, n2613, n2614, n2615, n2616, 
        n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, 
        n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, 
        n2633, n2643, n2678, n2679, n2680, n2681, n2682, n2683, 
        n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, 
        n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699, 
        n2700, n2701, n2709, n2710, n2711, n2712, n2713, n2714, 
        n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, 
        n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, 
        n2731, n2732, n2733, n2742, n2776, n2777, n2778, n2779, 
        n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, 
        n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795, 
        n2796, n2797, n2798, n2799, n2800, n2801, n2808, n2809, 
        n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, 
        n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825, 
        n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, 
        n48068, n27203, n2841, n27261, n2876, n2877, n2878, n2879, 
        n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887, 
        n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895, 
        n2896, n2897, n2898, n2899, n2900, n2901, n2907, n2908, 
        n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916, 
        n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, 
        n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, 
        n2933, n2940, n2975, n2976, n2977, n2978, n2979, n2980, 
        n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, 
        n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, 
        n2997, n2998, n2999, n3000, n3001, n3006, n3007, n3008, 
        n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, 
        n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024, 
        n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, 
        n3033, n3039, n3074, n3075, n3076, n3077, n3078, n3079, 
        n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, 
        n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095, 
        n3096, n3097, n3098, n3099, n3100, n3101, n3105, n3106, 
        n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114, 
        n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, 
        n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, 
        n3131, n3132, n3133, n3138, n56706, n3173, n3174, n3175, 
        n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, 
        n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, 
        n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199, 
        n3200, n3201, n3204, n3205, n3206, n3207, n3208, n3209, 
        n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, 
        n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225, 
        n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, 
        n3237, n3272, n3273, n3274, n3275, n3276, n3277, n3278, 
        n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, 
        n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, 
        n3295, n3296, n3298, n3299, n3300, n3301, n12_adj_5600, 
        n49838, n9_adj_5601, n48522, n56658, n56652, n56628, n48670, 
        n24_adj_5602, n28729, n50886, n50888, n62, n27116, n27119, 
        n47790, n4_adj_5603, n52298, n27243, n29417, n56200, n52278, 
        n29242, n28672, n52270, n56561, n28648, n43576, n52264, 
        n12_adj_5604, n52258, n63_adj_5605, n52252, n52246, n56056, 
        n51396, n52244, n29416, n52242, n27271, n27264, n52232, 
        n54660, n52222, n52220, n22875, n5_adj_5606, n52214, n29282, 
        n52208, n4_adj_5607, n52200, n52196, n27113, n55569, n56171, 
        n52190, n52184, n27258, n52182, n52168, n52162, n52156, 
        n52150, n48947, n54624, n52144, n52142, n29415, n55137, 
        n54622, n52132, n52126, n56025, n52120, n52114, n52112, 
        n7_adj_5608, n8_adj_5609, n27218, n29414, n29413, n29412, 
        n29411, n29410, n29408, n52102, n54609, n52096, n56622, 
        n56616, n48, n49, n50, n51, n52, n53, n54, n55, n29407, 
        n52092, n44205, n56490, n10829, n10_adj_5610, n56458, n52086, 
        n52084, n44204, n43653, n44203, n52070, n52066, n52060, 
        n44202, n52054, n52048, n52046, n52040, n52038, n29406, 
        n29405, n29404, n29403, n29402, n29401, n29400, n48526, 
        n29398, n29397, n29396, n29395, n29394, n29393, n29391, 
        n29390, n29389, n29388, n29387, n29386, n29385, n29384, 
        n29383, n29382, n29381, n29380, n29379, n29378, n29375, 
        n44201, n43575, n43652, n43651, n44200, n43574, n43650, 
        n44199, n43548, n43649, n43573, n43648, n51081, n52026, 
        n44198, n52020, n43647, n43572, n43571, n44197, n43570, 
        n56444, n52012, n52010, n29374, n29371, n29370, n29369, 
        n29368, n52000, n29364, n29363, n29362, n29361, n29360, 
        n29359, n29358, n29571, n51998, n51996, n43646, n43569, 
        n51990, n54594, n51986, n43645, n50021, n29570, n29569, 
        n29568, n29567, n29566, n29565, n29564, n29563, n29562, 
        n29561, n29560, n29559, n29558, n29557, n29556, n29555, 
        n29554, n29553, n29552, n29551, n29550, n29549, n29546, 
        n29545, n29544, n29543, n29542, n29541, n29540, n29539, 
        n43644, n44196, n29538, n29537, n29536, n29534, n29533, 
        n44195, n29356, n29355, n29532, n29531, n29530, n29529, 
        n29528, n29527, n29526, n29525, n43643, n56430, n43642, 
        n51980, n43641, n50013, n43640, n43547, n43568, n2_adj_5611, 
        n3_adj_5612, n4_adj_5613, n5_adj_5614, n6_adj_5615, n7_adj_5616, 
        n8_adj_5617, n9_adj_5618, n10_adj_5619, n11_adj_5620, n12_adj_5621, 
        n13_adj_5622, n14_adj_5623, n15_adj_5624, n16_adj_5625, n17_adj_5626, 
        n18_adj_5627, n19_adj_5628, n20_adj_5629, n21_adj_5630, n22_adj_5631, 
        n23_adj_5632, n24_adj_5633, n25_adj_5634, n26_adj_5635, n27_adj_5636, 
        n28_adj_5637, n29_adj_5638, n30_adj_5639, n31_adj_5640, n32_adj_5641, 
        n33_adj_5642, n54589, n43639, n43567, n43566, n43638, n43565, 
        n29354, n56415, n43564, n44194, n44193, n5_adj_5643, n51960, 
        n4_adj_5644, n44192, n44191, n44190, n44189, n51954, n51952, 
        n44188, n54586, n44187, n44186, n44185, n51946, n44184, 
        n44183, n44182, n44181, n44180, n50829, n44179, n44178, 
        n37418, n44177, n44696, n44695, n44176, n44694, n44693, 
        n44175, n44174, n44173, n44692, n44691, n37416, n44172, 
        n51936, n44171, n44170, n44690, n44689, n44169, n44168, 
        n44167, n44166, n44688, n51930, n44687, n44686, n44165, 
        n44685, n44164, n44684, n44163, n44162, n44683, n44682, 
        n44681, n44161, n44680, n44679, n44160, n44159, n6_adj_5645, 
        n44158, n44157, n51918, n44678, n44677, n44676, n44675, 
        n44674, n44156, n44155, n44154, n51914, n37412, n44673, 
        n44672, n44671, n44670, n44669, n44668, n44153, n44667, 
        n44152, n44151, n44150, n44149, n27208, n44148, n56399, 
        n44147, n44666, n43637, n44146, n44145, n50144, n44144, 
        n44143, n51902, n44142, n44141, n44140, n43563, n51896, 
        n44139, n44138, n44137, n44136, n44135, n44134, n50130, 
        n44133, n44132, n43562, n56142, n44131, n44130, n44129, 
        n44128, n44127, n44126, n44125, n44124, n44123, n53094, 
        n43636, n43536, n44122, n51890, n29353, n44121, n37404, 
        n43546, n44120, n44119, n44118, n44117, n44116, n44115, 
        n43561, n44114, n44113, n44112, n44111, n44110, n44109, 
        n51886, n44108, n43635, n44107, n44106, n44105, n43634, 
        n44104, n43633, n51880, n43632, n44103, n43545, n44102, 
        n51878, n44101, n44100, n43631, n51876, n44099, n44098, 
        n43630, n44097, n50043, n43629, n44096, n44095, n43544, 
        n44094, n44093, n44092, n44091, n27238, n43794, n43793, 
        n43792, n43628, n43627, n43791, n37400, n37398, n43626, 
        n44090, n44089, n37394, n43790, n43625, n44088, n43789, 
        n43624, n44087, n43560, n43788, n43787, n44086, n8_adj_5646, 
        n43786, n44085, n44084, n43623, n44083, n43785, n43784, 
        n43622, n43783, n51860, n43621, n19728, n43782, n43781, 
        n43620, n44082, n44081, n43780, n44080, n43779, n43559, 
        n43778, n43619, n43777, n43535, n44079, n51856, n37392, 
        n43776, n44078, n43543, n37390, n37388, n57033, n43618, 
        n51850, n44077, n43775, n43774, n44076, n44075, n44074, 
        n43773, n44073, n43772, n44072, n53086, n44071, n57032, 
        n37386, n43617, n51842, n44070, n43616, n27094, n7_adj_5647, 
        n15_adj_5648, n17_adj_5649, n19_adj_5650, n21_adj_5651, n51834, 
        n27_adj_5652, n53084, n31_adj_5653, n35, n59, n61, n43615, 
        n51828, n51826, n56382, n51820, n51812, n8_adj_5654, n51806, 
        n51800, n51794, n51792, n56364, n50081, n51780, n51772, 
        n55806, n51766, n51760, n51750, n48878, n51744, n51509, 
        n54553, n51740, n51734, n51732, n51722, n51716, n51714, 
        n51712, n51706, n51702, n51700, n54552, n54551, n54550, 
        n54549, n51694, n53127, n54548, n54547, n53069, n51491, 
        n51690, n51682, n7_adj_5655, n51680, n51678, n51676, n51674, 
        n51672, n56115, n51014, n51670, n51668, n51666, n51664, 
        n51662, n51660, n51658, n51654, n56323, n51646, n51644, 
        n51642, n51640, n51638, n55885, n55884, n54539, n51632, 
        n56874, n55869, n55865, n55863, n51626, n51624, n56302, 
        n55862, n55864, n48778, n55823, n54531, n56614, n51618, 
        n51614, n56280, n55592, n51610, n53036, n53032, n53025, 
        n56868, n6_adj_5656;
    
    VCC i2 (.Y(VCC_net));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1838_23_lut (.I0(GND_net), 
            .I1(n2713), .I2(VCC_net), .I3(n44272), .O(n2780)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1838_23_lut.LUT_INIT = 16'hC33C;
    SB_IO hall2_input (.PACKAGE_PIN(HALL2), .LATCH_INPUT_VALUE(GND_net), 
          .INPUT_CLK(GND_net), .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_1(GND_net), .D_OUT_0(GND_net), .D_IN_0(hall2)) /* synthesis syn_instantiated=1 */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam hall2_input.PIN_TYPE = 6'b000001;
    defparam hall2_input.PULLUP = 1'b1;
    defparam hall2_input.NEG_TRIGGER = 1'b0;
    defparam hall2_input.IO_STANDARD = "SB_LVCMOS";
    SB_IO hall3_input (.PACKAGE_PIN(HALL3), .LATCH_INPUT_VALUE(GND_net), 
          .INPUT_CLK(GND_net), .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_1(GND_net), .D_OUT_0(GND_net), .D_IN_0(hall3)) /* synthesis syn_instantiated=1 */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam hall3_input.PIN_TYPE = 6'b000001;
    defparam hall3_input.PULLUP = 1'b1;
    defparam hall3_input.NEG_TRIGGER = 1'b0;
    defparam hall3_input.IO_STANDARD = "SB_LVCMOS";
    SB_IO tx_output (.PACKAGE_PIN(TX), .LATCH_INPUT_VALUE(GND_net), .INPUT_CLK(GND_net), 
          .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(tx_enable), .D_OUT_1(GND_net), 
          .D_OUT_0(tx_o)) /* synthesis syn_instantiated=1 */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam tx_output.PIN_TYPE = 6'b101001;
    defparam tx_output.PULLUP = 1'b1;
    defparam tx_output.NEG_TRIGGER = 1'b0;
    defparam tx_output.IO_STANDARD = "SB_LVCMOS";
    SB_DFF commutation_state_prev_i0 (.Q(commutation_state_prev[0]), .C(clk16MHz), 
           .D(commutation_state[0]));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i972_3_lut (.I0(n1425), .I1(n1492), 
            .I2(n1455), .I3(GND_net), .O(n1524));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i972_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_175_31 (.CI(n43638), .I0(delay_counter[29]), .I1(GND_net), 
            .CO(n43639));
    SB_LUT4 i15470_3_lut (.I0(IntegralLimit[22]), .I1(\data_in_frame[11] [6]), 
            .I2(n50654), .I3(GND_net), .O(n29550));   // verilog/coms.v(128[12] 303[6])
    defparam i15470_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_1039_17_lut (.I0(GND_net), .I1(n4889), .I2(n4914), .I3(n43786), 
            .O(n426)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1039_17_lut.LUT_INIT = 16'hC33C;
    SB_DFF dir_205 (.Q(dir), .C(clk16MHz), .D(pwm_setpoint_23__N_263));   // verilog/TinyFPGA_B.v(103[9] 129[5])
    SB_LUT4 add_175_30_lut (.I0(GND_net), .I1(delay_counter[28]), .I2(GND_net), 
            .I3(n43637), .O(n1535)) /* synthesis syn_instantiated=1 */ ;
    defparam add_175_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_967_5 (.CI(n44020), 
            .I0(n1431), .I1(VCC_net), .CO(n44021));
    SB_LUT4 i15471_3_lut (.I0(IntegralLimit[21]), .I1(\data_in_frame[11] [5]), 
            .I2(n50654), .I3(GND_net), .O(n29551));   // verilog/coms.v(128[12] 303[6])
    defparam i15471_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_967_4_lut (.I0(GND_net), 
            .I1(n1432), .I2(GND_net), .I3(n44019), .O(n1499)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_967_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15472_3_lut (.I0(IntegralLimit[20]), .I1(\data_in_frame[11] [4]), 
            .I2(n50654), .I3(GND_net), .O(n29552));   // verilog/coms.v(128[12] 303[6])
    defparam i15472_3_lut.LUT_INIT = 16'hacac;
    SB_DFFE dti_207 (.Q(dti), .C(clk16MHz), .E(n28648), .D(dti_N_527));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_967_4 (.CI(n44019), 
            .I0(n1432), .I1(GND_net), .CO(n44020));
    SB_DFF encoder0_position_scaled_i0 (.Q(encoder0_position_scaled[0]), .C(clk16MHz), 
           .D(encoder0_position_scaled_23__N_51[0]));   // verilog/TinyFPGA_B.v(321[10] 334[6])
    SB_LUT4 i14_3_lut (.I0(hall2), .I1(hall3), .I2(hall1), .I3(GND_net), 
            .O(n6_adj_5656));
    defparam i14_3_lut.LUT_INIT = 16'h7e7e;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1838_23 (.CI(n44272), 
            .I0(n2713), .I1(VCC_net), .CO(n44273));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1838_22_lut (.I0(GND_net), 
            .I1(n2714), .I2(VCC_net), .I3(n44271), .O(n2781)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1838_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1039_17 (.CI(n43786), .I0(n4889), .I1(n4914), .CO(n43787));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_967_3_lut (.I0(GND_net), 
            .I1(n1433), .I2(VCC_net), .I3(n44018), .O(n1500)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_967_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_967_3 (.CI(n44018), 
            .I0(n1433), .I1(VCC_net), .CO(n44019));
    SB_LUT4 add_1039_16_lut (.I0(GND_net), .I1(n4890), .I2(n4915), .I3(n43785), 
            .O(n427)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1039_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1039_16 (.CI(n43785), .I0(n4890), .I1(n4915), .CO(n43786));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1838_22 (.CI(n44271), 
            .I0(n2714), .I1(VCC_net), .CO(n44272));
    SB_LUT4 add_1039_15_lut (.I0(GND_net), .I1(n4891), .I2(n4916), .I3(n43784), 
            .O(n428)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1039_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15473_3_lut (.I0(IntegralLimit[19]), .I1(\data_in_frame[11] [3]), 
            .I2(n50654), .I3(GND_net), .O(n29553));   // verilog/coms.v(128[12] 303[6])
    defparam i15473_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_1039_15 (.CI(n43784), .I0(n4891), .I1(n4916), .CO(n43785));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_967_2_lut (.I0(GND_net), 
            .I1(n414), .I2(GND_net), .I3(VCC_net), .O(n1501)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_967_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_1039_14_lut (.I0(GND_net), .I1(n4892), .I2(n4917), .I3(n43783), 
            .O(n429)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1039_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_mux_3_i23_3_lut (.I0(encoder0_position_scaled_23__N_327[22]), 
            .I1(n11_adj_5488), .I2(encoder0_position_scaled_23__N_327[31]), 
            .I3(GND_net), .O(n411));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_mux_3_i23_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut (.I0(hall3), .I1(hall2), .I2(hall1), .I3(GND_net), 
            .O(commutation_state_7__N_264[0]));   // verilog/TinyFPGA_B.v(163[4] 165[7])
    defparam i1_3_lut.LUT_INIT = 16'h1414;
    SB_DFF encoder1_position_scaled_i0 (.Q(encoder1_position_scaled[0]), .C(clk16MHz), 
           .D(encoder1_position_scaled_23__N_75[0]));   // verilog/TinyFPGA_B.v(321[10] 334[6])
    SB_IO sda_output (.PACKAGE_PIN(SDA), .LATCH_INPUT_VALUE(GND_net), .INPUT_CLK(GND_net), 
          .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(sda_enable), .D_OUT_1(GND_net), 
          .D_OUT_0(sda_out), .D_IN_0(state_7__N_4306[3])) /* synthesis syn_instantiated=1 */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam sda_output.PIN_TYPE = 6'b101001;
    defparam sda_output.PULLUP = 1'b1;
    defparam sda_output.NEG_TRIGGER = 1'b0;
    defparam sda_output.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 i15474_3_lut (.I0(IntegralLimit[18]), .I1(\data_in_frame[11] [2]), 
            .I2(n50654), .I3(GND_net), .O(n29554));   // verilog/coms.v(128[12] 303[6])
    defparam i15474_3_lut.LUT_INIT = 16'hacac;
    SB_DFF displacement_i0 (.Q(displacement[0]), .C(clk16MHz), .D(displacement_23__N_99[0]));   // verilog/TinyFPGA_B.v(321[10] 334[6])
    SB_IO CS_pad (.PACKAGE_PIN(CS), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(CS_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam CS_pad.PIN_TYPE = 6'b011001;
    defparam CS_pad.PULLUP = 1'b0;
    defparam CS_pad.NEG_TRIGGER = 1'b0;
    defparam CS_pad.IO_STANDARD = "SB_LVCMOS";
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_967_2 (.CI(VCC_net), 
            .I0(n414), .I1(GND_net), .CO(n44018));
    SB_IO scl_output (.PACKAGE_PIN(SCL), .LATCH_INPUT_VALUE(GND_net), .INPUT_CLK(GND_net), 
          .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(scl_enable), .D_OUT_1(GND_net), 
          .D_OUT_0(scl)) /* synthesis syn_instantiated=1 */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam scl_output.PIN_TYPE = 6'b101001;
    defparam scl_output.PULLUP = 1'b1;
    defparam scl_output.NEG_TRIGGER = 1'b0;
    defparam scl_output.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 i40311_1_lut (.I0(n2544), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n56142));
    defparam i40311_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1838_21_lut (.I0(GND_net), 
            .I1(n2715), .I2(VCC_net), .I3(n44270), .O(n2782)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1838_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_175_30 (.CI(n43637), .I0(delay_counter[28]), .I1(GND_net), 
            .CO(n43638));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1039_3_lut (.I0(n1524), 
            .I1(n1591), .I2(n1554_adj_5597), .I3(GND_net), .O(n1623));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1039_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1838_21 (.CI(n44270), 
            .I0(n2715), .I1(VCC_net), .CO(n44271));
    SB_IO hall1_input (.PACKAGE_PIN(HALL1), .LATCH_INPUT_VALUE(GND_net), 
          .INPUT_CLK(GND_net), .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_1(GND_net), .D_OUT_0(GND_net), .D_IN_0(hall1)) /* synthesis syn_instantiated=1 */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam hall1_input.PIN_TYPE = 6'b000001;
    defparam hall1_input.PULLUP = 1'b1;
    defparam hall1_input.NEG_TRIGGER = 1'b0;
    defparam hall1_input.IO_STANDARD = "SB_LVCMOS";
    \neopixel(CLOCK_SPEED_HZ=16000000)  nx (.clk16MHz(clk16MHz), .\state[0] (state[0]), 
            .\state[1] (state[1]), .GND_net(GND_net), .\neo_pixel_transmitter.t0 ({\neo_pixel_transmitter.t0 }), 
            .n28778(n28778), .\state_3__N_639[1] (state_3__N_639[1]), .neopxl_color({neopxl_color}), 
            .timer({timer}), .VCC_net(VCC_net), .LED_c(LED_c), .n29354(n29354), 
            .n29829(n29829), .n29814(n29814), .n29813(n29813), .n29812(n29812), 
            .n29811(n29811), .n29810(n29810), .n29809(n29809), .n29808(n29808), 
            .n29807(n29807), .n29806(n29806), .n29805(n29805), .n29804(n29804), 
            .n29803(n29803), .n29802(n29802), .n29801(n29801), .n29800(n29800), 
            .n29799(n29799), .n29798(n29798), .n29797(n29797), .n29796(n29796), 
            .n29795(n29795), .n29794(n29794), .n29793(n29793), .n29792(n29792), 
            .n29791(n29791), .n29790(n29790), .n29789(n29789), .n29788(n29788), 
            .n29785(n29785), .n29784(n29784), .n29783(n29783), .n29782(n29782), 
            .NEOPXL_c(NEOPXL_c), .n47790(n47790)) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(50[24] 56[2])
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1838_20_lut (.I0(GND_net), 
            .I1(n2716), .I2(VCC_net), .I3(n44269), .O(n2783)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1838_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1106_3_lut (.I0(n1623), 
            .I1(n1690), .I2(n1653), .I3(GND_net), .O(n1722));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1106_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1838_20 (.CI(n44269), 
            .I0(n2716), .I1(VCC_net), .CO(n44270));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1838_19_lut (.I0(GND_net), 
            .I1(n2717), .I2(VCC_net), .I3(n44268), .O(n2784)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1838_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_175_29_lut (.I0(GND_net), .I1(delay_counter[27]), .I2(GND_net), 
            .I3(n43636), .O(n1536)) /* synthesis syn_instantiated=1 */ ;
    defparam add_175_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1039_14 (.CI(n43783), .I0(n4892), .I1(n4917), .CO(n43784));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1173_3_lut (.I0(n1722), 
            .I1(n1789), .I2(n1752), .I3(GND_net), .O(n1821));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1173_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_1039_13_lut (.I0(GND_net), .I1(n4893), .I2(n4918), .I3(n43782), 
            .O(n430)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1039_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1838_19 (.CI(n44268), 
            .I0(n2717), .I1(VCC_net), .CO(n44269));
    SB_LUT4 i15475_3_lut (.I0(IntegralLimit[17]), .I1(\data_in_frame[11] [1]), 
            .I2(n50654), .I3(GND_net), .O(n29555));   // verilog/coms.v(128[12] 303[6])
    defparam i15475_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_175_29 (.CI(n43636), .I0(delay_counter[27]), .I1(GND_net), 
            .CO(n43637));
    SB_LUT4 i34086_4_lut (.I0(n26_adj_5575), .I1(state_adj_5705[0]), .I2(n6), 
            .I3(state_adj_5736[0]), .O(n49838));
    defparam i34086_4_lut.LUT_INIT = 16'hccc8;
    SB_LUT4 add_175_28_lut (.I0(GND_net), .I1(delay_counter[26]), .I2(GND_net), 
            .I3(n43635), .O(n1537)) /* synthesis syn_instantiated=1 */ ;
    defparam add_175_28_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_900_13_lut (.I0(n56415), 
            .I1(n1323), .I2(VCC_net), .I3(n44017), .O(n1422)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_900_13_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i15476_3_lut (.I0(IntegralLimit[16]), .I1(\data_in_frame[11] [0]), 
            .I2(n50654), .I3(GND_net), .O(n29556));   // verilog/coms.v(128[12] 303[6])
    defparam i15476_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_175_28 (.CI(n43635), .I0(delay_counter[26]), .I1(GND_net), 
            .CO(n43636));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1838_18_lut (.I0(GND_net), 
            .I1(n2718), .I2(VCC_net), .I3(n44267), .O(n2785)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1838_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15477_3_lut (.I0(IntegralLimit[15]), .I1(\data_in_frame[12] [7]), 
            .I2(n50654), .I3(GND_net), .O(n29557));   // verilog/coms.v(128[12] 303[6])
    defparam i15477_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1838_18 (.CI(n44267), 
            .I0(n2718), .I1(VCC_net), .CO(n44268));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1838_17_lut (.I0(GND_net), 
            .I1(n2719), .I2(VCC_net), .I3(n44266), .O(n2786)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1838_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1838_17 (.CI(n44266), 
            .I0(n2719), .I1(VCC_net), .CO(n44267));
    SB_LUT4 i1_3_lut_adj_1712 (.I0(state_adj_5705[1]), .I1(read), .I2(n49919), 
            .I3(GND_net), .O(n12_adj_5600));   // verilog/eeprom.v(26[8] 58[4])
    defparam i1_3_lut_adj_1712.LUT_INIT = 16'ha2a2;
    SB_LUT4 i1_4_lut (.I0(n36659), .I1(n12_adj_5600), .I2(state_adj_5705[0]), 
            .I3(n49919), .O(n48526));   // verilog/eeprom.v(26[8] 58[4])
    defparam i1_4_lut.LUT_INIT = 16'h88a8;
    SB_CARRY add_261_16 (.CI(n43571), .I0(duty[17]), .I1(n56614), .CO(n43572));
    SB_LUT4 i15478_3_lut (.I0(IntegralLimit[14]), .I1(\data_in_frame[12] [6]), 
            .I2(n50654), .I3(GND_net), .O(n29558));   // verilog/coms.v(128[12] 303[6])
    defparam i15478_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_175_27_lut (.I0(GND_net), .I1(delay_counter[25]), .I2(GND_net), 
            .I3(n43634), .O(n1538)) /* synthesis syn_instantiated=1 */ ;
    defparam add_175_27_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15479_3_lut (.I0(IntegralLimit[13]), .I1(\data_in_frame[12] [5]), 
            .I2(n50654), .I3(GND_net), .O(n29559));   // verilog/coms.v(128[12] 303[6])
    defparam i15479_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15396_3_lut (.I0(\data_in[1] [2]), .I1(\data_in[2] [2]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n29476));   // verilog/coms.v(128[12] 303[6])
    defparam i15396_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1838_16_lut (.I0(GND_net), 
            .I1(n2720), .I2(VCC_net), .I3(n44265), .O(n2787)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1838_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1838_16 (.CI(n44265), 
            .I0(n2720), .I1(VCC_net), .CO(n44266));
    SB_LUT4 add_261_15_lut (.I0(current[15]), .I1(duty[16]), .I2(n56614), 
            .I3(n43570), .O(n257)) /* synthesis syn_instantiated=1 */ ;
    defparam add_261_15_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY add_1039_13 (.CI(n43782), .I0(n4893), .I1(n4918), .CO(n43783));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1838_15_lut (.I0(GND_net), 
            .I1(n2721), .I2(VCC_net), .I3(n44264), .O(n2788)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1838_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1838_15 (.CI(n44264), 
            .I0(n2721), .I1(VCC_net), .CO(n44265));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1838_14_lut (.I0(GND_net), 
            .I1(n2722), .I2(VCC_net), .I3(n44263), .O(n2789)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1838_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_900_12_lut (.I0(GND_net), 
            .I1(n1324), .I2(VCC_net), .I3(n44016), .O(n1391)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_900_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_175_27 (.CI(n43634), .I0(delay_counter[25]), .I1(GND_net), 
            .CO(n43635));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_900_12 (.CI(n44016), 
            .I0(n1324), .I1(VCC_net), .CO(n44017));
    SB_LUT4 i15480_3_lut (.I0(IntegralLimit[12]), .I1(\data_in_frame[12] [4]), 
            .I2(n50654), .I3(GND_net), .O(n29560));   // verilog/coms.v(128[12] 303[6])
    defparam i15480_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1838_14 (.CI(n44263), 
            .I0(n2722), .I1(VCC_net), .CO(n44264));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1838_13_lut (.I0(GND_net), 
            .I1(n2723), .I2(VCC_net), .I3(n44262), .O(n2790)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1838_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1240_3_lut (.I0(n1821), 
            .I1(n1888), .I2(n1851), .I3(GND_net), .O(n1920));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1240_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_263_5_lut (.I0(GND_net), .I1(encoder1_position[6]), .I2(GND_net), 
            .I3(n43537), .O(encoder1_position_scaled_23__N_75[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_263_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_1039_12_lut (.I0(GND_net), .I1(n4894), .I2(n4919), .I3(n43781), 
            .O(n431)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1039_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1039_12 (.CI(n43781), .I0(n4894), .I1(n4919), .CO(n43782));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1838_13 (.CI(n44262), 
            .I0(n2723), .I1(VCC_net), .CO(n44263));
    SB_LUT4 add_263_13_lut (.I0(GND_net), .I1(encoder1_position[14]), .I2(GND_net), 
            .I3(n43545), .O(encoder1_position_scaled_23__N_75[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_263_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_900_11_lut (.I0(GND_net), 
            .I1(n1325), .I2(VCC_net), .I3(n44015), .O(n1392)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_900_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1838_12_lut (.I0(GND_net), 
            .I1(n2724), .I2(VCC_net), .I3(n44261), .O(n2791)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1838_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_261_15 (.CI(n43570), .I0(duty[16]), .I1(n56614), .CO(n43571));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_900_11 (.CI(n44015), 
            .I0(n1325), .I1(VCC_net), .CO(n44016));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1307_3_lut (.I0(n1920), 
            .I1(n1987), .I2(n1950), .I3(GND_net), .O(n2019));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1307_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1838_12 (.CI(n44261), 
            .I0(n2724), .I1(VCC_net), .CO(n44262));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1838_11_lut (.I0(GND_net), 
            .I1(n2725), .I2(VCC_net), .I3(n44260), .O(n2792)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1838_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_263_5 (.CI(n43537), .I0(encoder1_position[6]), .I1(GND_net), 
            .CO(n43538));
    SB_LUT4 add_1039_11_lut (.I0(GND_net), .I1(n4895), .I2(n4920), .I3(n43780), 
            .O(n432)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1039_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1838_11 (.CI(n44260), 
            .I0(n2725), .I1(VCC_net), .CO(n44261));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1838_10_lut (.I0(GND_net), 
            .I1(n2726), .I2(VCC_net), .I3(n44259), .O(n2793)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1838_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1838_10 (.CI(n44259), 
            .I0(n2726), .I1(VCC_net), .CO(n44260));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1838_9_lut (.I0(GND_net), 
            .I1(n2727), .I2(VCC_net), .I3(n44258), .O(n2794)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1838_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1039_11 (.CI(n43780), .I0(n4895), .I1(n4920), .CO(n43781));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1838_9 (.CI(n44258), 
            .I0(n2727), .I1(VCC_net), .CO(n44259));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1838_8_lut (.I0(GND_net), 
            .I1(n2728), .I2(VCC_net), .I3(n44257), .O(n2795)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1838_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15481_3_lut (.I0(IntegralLimit[11]), .I1(\data_in_frame[12] [3]), 
            .I2(n50654), .I3(GND_net), .O(n29561));   // verilog/coms.v(128[12] 303[6])
    defparam i15481_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1374_3_lut (.I0(n2019), 
            .I1(n2086), .I2(n2049), .I3(GND_net), .O(n2118));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1374_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1838_8 (.CI(n44257), 
            .I0(n2728), .I1(VCC_net), .CO(n44258));
    SB_LUT4 add_175_26_lut (.I0(GND_net), .I1(delay_counter[24]), .I2(GND_net), 
            .I3(n43633), .O(n1539)) /* synthesis syn_instantiated=1 */ ;
    defparam add_175_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_900_10_lut (.I0(GND_net), 
            .I1(n1326), .I2(VCC_net), .I3(n44014), .O(n1393)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_900_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1838_7_lut (.I0(GND_net), 
            .I1(n2729), .I2(GND_net), .I3(n44256), .O(n2796)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1838_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15482_3_lut (.I0(IntegralLimit[10]), .I1(\data_in_frame[12] [2]), 
            .I2(n50654), .I3(GND_net), .O(n29562));   // verilog/coms.v(128[12] 303[6])
    defparam i15482_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1838_7 (.CI(n44256), 
            .I0(n2729), .I1(GND_net), .CO(n44257));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_900_10 (.CI(n44014), 
            .I0(n1326), .I1(VCC_net), .CO(n44015));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_900_9_lut (.I0(GND_net), 
            .I1(n1327), .I2(VCC_net), .I3(n44013), .O(n1394)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_900_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1838_6_lut (.I0(GND_net), 
            .I1(n2730), .I2(GND_net), .I3(n44255), .O(n2797)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1838_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1838_6 (.CI(n44255), 
            .I0(n2730), .I1(GND_net), .CO(n44256));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_900_9 (.CI(n44013), 
            .I0(n1327), .I1(VCC_net), .CO(n44014));
    SB_LUT4 add_1039_10_lut (.I0(GND_net), .I1(n4896), .I2(n4921), .I3(n43779), 
            .O(n433)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1039_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1838_5_lut (.I0(GND_net), 
            .I1(n2731), .I2(VCC_net), .I3(n44254), .O(n2798)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1838_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_900_8_lut (.I0(GND_net), 
            .I1(n1328), .I2(VCC_net), .I3(n44012), .O(n1395)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_900_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1838_5 (.CI(n44254), 
            .I0(n2731), .I1(VCC_net), .CO(n44255));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1838_4_lut (.I0(GND_net), 
            .I1(n2732), .I2(GND_net), .I3(n44253), .O(n2799)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1838_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1838_4 (.CI(n44253), 
            .I0(n2732), .I1(GND_net), .CO(n44254));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1838_3_lut (.I0(GND_net), 
            .I1(n2733), .I2(VCC_net), .I3(n44252), .O(n2800)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1838_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1838_3 (.CI(n44252), 
            .I0(n2733), .I1(VCC_net), .CO(n44253));
    SB_CARRY add_1039_10 (.CI(n43779), .I0(n4896), .I1(n4921), .CO(n43780));
    SB_LUT4 i15483_3_lut (.I0(IntegralLimit[9]), .I1(\data_in_frame[12] [1]), 
            .I2(n50654), .I3(GND_net), .O(n29563));   // verilog/coms.v(128[12] 303[6])
    defparam i15483_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_900_8 (.CI(n44012), 
            .I0(n1328), .I1(VCC_net), .CO(n44013));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1838_2_lut (.I0(GND_net), 
            .I1(n538), .I2(GND_net), .I3(VCC_net), .O(n2801)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1838_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1838_2 (.CI(VCC_net), 
            .I0(n538), .I1(GND_net), .CO(n44252));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1771_26_lut (.I0(n56115), 
            .I1(n2610), .I2(VCC_net), .I3(n44251), .O(n2709)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1771_26_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1771_25_lut (.I0(GND_net), 
            .I1(n2611), .I2(VCC_net), .I3(n44250), .O(n2678)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1771_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1771_25 (.CI(n44250), 
            .I0(n2611), .I1(VCC_net), .CO(n44251));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_900_7_lut (.I0(GND_net), 
            .I1(n1329), .I2(GND_net), .I3(n44011), .O(n1396)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_900_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_900_7 (.CI(n44011), 
            .I0(n1329), .I1(GND_net), .CO(n44012));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_900_6_lut (.I0(GND_net), 
            .I1(n1330), .I2(GND_net), .I3(n44010), .O(n1397)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_900_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_1039_9_lut (.I0(GND_net), .I1(n4897), .I2(n4922), .I3(n43778), 
            .O(n434)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1039_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1771_24_lut (.I0(GND_net), 
            .I1(n2612), .I2(VCC_net), .I3(n44249), .O(n2679)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1771_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1039_9 (.CI(n43778), .I0(n4897), .I1(n4922), .CO(n43779));
    SB_LUT4 i15397_3_lut (.I0(\data_in[1] [1]), .I1(\data_in[2] [1]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n29477));   // verilog/coms.v(128[12] 303[6])
    defparam i15397_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1771_24 (.CI(n44249), 
            .I0(n2612), .I1(VCC_net), .CO(n44250));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1771_23_lut (.I0(GND_net), 
            .I1(n2613), .I2(VCC_net), .I3(n44248), .O(n2680)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1771_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1771_23 (.CI(n44248), 
            .I0(n2613), .I1(VCC_net), .CO(n44249));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_900_6 (.CI(n44010), 
            .I0(n1330), .I1(GND_net), .CO(n44011));
    SB_CARRY add_175_26 (.CI(n43633), .I0(delay_counter[24]), .I1(GND_net), 
            .CO(n43634));
    SB_LUT4 add_1039_8_lut (.I0(GND_net), .I1(n4898), .I2(n4923), .I3(n43777), 
            .O(n435)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1039_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1771_22_lut (.I0(GND_net), 
            .I1(n2614), .I2(VCC_net), .I3(n44247), .O(n2681)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1771_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1771_22 (.CI(n44247), 
            .I0(n2614), .I1(VCC_net), .CO(n44248));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1771_21_lut (.I0(GND_net), 
            .I1(n2615), .I2(VCC_net), .I3(n44246), .O(n2682)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1771_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_900_5_lut (.I0(GND_net), 
            .I1(n1331), .I2(VCC_net), .I3(n44009), .O(n1398)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_900_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1771_21 (.CI(n44246), 
            .I0(n2615), .I1(VCC_net), .CO(n44247));
    SB_LUT4 add_261_14_lut (.I0(current[15]), .I1(duty[15]), .I2(n56614), 
            .I3(n43569), .O(n258)) /* synthesis syn_instantiated=1 */ ;
    defparam add_261_14_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 i15398_3_lut (.I0(\data_in[1] [0]), .I1(\data_in[2] [0]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n29478));   // verilog/coms.v(128[12] 303[6])
    defparam i15398_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15399_3_lut (.I0(\data_in[0] [7]), .I1(\data_in[1] [7]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n29479));   // verilog/coms.v(128[12] 303[6])
    defparam i15399_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_261_14 (.CI(n43569), .I0(duty[15]), .I1(n56614), .CO(n43570));
    SB_CARRY add_1039_8 (.CI(n43777), .I0(n4898), .I1(n4923), .CO(n43778));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_900_5 (.CI(n44009), 
            .I0(n1331), .I1(VCC_net), .CO(n44010));
    SB_LUT4 i15484_3_lut (.I0(IntegralLimit[8]), .I1(\data_in_frame[12] [0]), 
            .I2(n50654), .I3(GND_net), .O(n29564));   // verilog/coms.v(128[12] 303[6])
    defparam i15484_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15485_3_lut (.I0(IntegralLimit[7]), .I1(\data_in_frame[13] [7]), 
            .I2(n50654), .I3(GND_net), .O(n29565));   // verilog/coms.v(128[12] 303[6])
    defparam i15485_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_1039_7_lut (.I0(GND_net), .I1(n4899), .I2(n4924), .I3(n43776), 
            .O(n436)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1039_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15400_3_lut (.I0(\data_in[0] [6]), .I1(\data_in[1] [6]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n29480));   // verilog/coms.v(128[12] 303[6])
    defparam i15400_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15486_3_lut (.I0(IntegralLimit[6]), .I1(\data_in_frame[13] [6]), 
            .I2(n50654), .I3(GND_net), .O(n29566));   // verilog/coms.v(128[12] 303[6])
    defparam i15486_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15401_3_lut (.I0(\data_in[0] [5]), .I1(\data_in[1] [5]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n29481));   // verilog/coms.v(128[12] 303[6])
    defparam i15401_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15487_3_lut (.I0(IntegralLimit[5]), .I1(\data_in_frame[13] [5]), 
            .I2(n50654), .I3(GND_net), .O(n29567));   // verilog/coms.v(128[12] 303[6])
    defparam i15487_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15402_3_lut (.I0(\data_in[0] [4]), .I1(\data_in[1] [4]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n29482));   // verilog/coms.v(128[12] 303[6])
    defparam i15402_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15403_3_lut (.I0(\data_in[0] [3]), .I1(\data_in[1] [3]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n29483));   // verilog/coms.v(128[12] 303[6])
    defparam i15403_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15404_3_lut (.I0(\data_in[0] [2]), .I1(\data_in[1] [2]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n29484));   // verilog/coms.v(128[12] 303[6])
    defparam i15404_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15488_3_lut (.I0(IntegralLimit[4]), .I1(\data_in_frame[13] [4]), 
            .I2(n50654), .I3(GND_net), .O(n29568));   // verilog/coms.v(128[12] 303[6])
    defparam i15488_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15405_3_lut (.I0(\data_in[0] [1]), .I1(\data_in[1] [1]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n29485));   // verilog/coms.v(128[12] 303[6])
    defparam i15405_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15406_3_lut (.I0(Ki[15]), .I1(\data_in_frame[4] [7]), .I2(n50654), 
            .I3(GND_net), .O(n29486));   // verilog/coms.v(128[12] 303[6])
    defparam i15406_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1375_3_lut (.I0(n2020), 
            .I1(n2087), .I2(n2049), .I3(GND_net), .O(n2119));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1375_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1443_3_lut (.I0(n2120), 
            .I1(n2187), .I2(n2148), .I3(GND_net), .O(n2219));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1443_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1442_3_lut (.I0(n2119), 
            .I1(n2186), .I2(n2148), .I3(GND_net), .O(n2218));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1442_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i3_4_lut (.I0(\ID_READOUT_FSM.state [1]), .I1(n62), .I2(delay_counter[31]), 
            .I3(\ID_READOUT_FSM.state [0]), .O(n51491));
    defparam i3_4_lut.LUT_INIT = 16'h0004;
    SB_LUT4 i15848_3_lut (.I0(PWMLimit[13]), .I1(\data_in_frame[9] [5]), 
            .I2(n50654), .I3(GND_net), .O(n29928));   // verilog/coms.v(128[12] 303[6])
    defparam i15848_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1441_3_lut (.I0(n2118), 
            .I1(n2185), .I2(n2148), .I3(GND_net), .O(n2217));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1441_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15489_3_lut (.I0(IntegralLimit[3]), .I1(\data_in_frame[13] [3]), 
            .I2(n50654), .I3(GND_net), .O(n29569));   // verilog/coms.v(128[12] 303[6])
    defparam i15489_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15849_3_lut (.I0(PWMLimit[12]), .I1(\data_in_frame[9] [4]), 
            .I2(n50654), .I3(GND_net), .O(n29929));   // verilog/coms.v(128[12] 303[6])
    defparam i15849_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15410_3_lut (.I0(Ki[14]), .I1(\data_in_frame[4] [6]), .I2(n50654), 
            .I3(GND_net), .O(n29490));   // verilog/coms.v(128[12] 303[6])
    defparam i15410_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15411_3_lut (.I0(Ki[13]), .I1(\data_in_frame[4] [5]), .I2(n50654), 
            .I3(GND_net), .O(n29491));   // verilog/coms.v(128[12] 303[6])
    defparam i15411_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15490_3_lut (.I0(IntegralLimit[2]), .I1(\data_in_frame[13] [2]), 
            .I2(n50654), .I3(GND_net), .O(n29570));   // verilog/coms.v(128[12] 303[6])
    defparam i15490_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15850_3_lut (.I0(PWMLimit[11]), .I1(\data_in_frame[9] [3]), 
            .I2(n50654), .I3(GND_net), .O(n29930));   // verilog/coms.v(128[12] 303[6])
    defparam i15850_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15412_3_lut (.I0(Ki[12]), .I1(\data_in_frame[4] [4]), .I2(n50654), 
            .I3(GND_net), .O(n29492));   // verilog/coms.v(128[12] 303[6])
    defparam i15412_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15413_3_lut (.I0(Ki[11]), .I1(\data_in_frame[4] [3]), .I2(n50654), 
            .I3(GND_net), .O(n29493));   // verilog/coms.v(128[12] 303[6])
    defparam i15413_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15491_3_lut (.I0(IntegralLimit[1]), .I1(\data_in_frame[13] [1]), 
            .I2(n50654), .I3(GND_net), .O(n29571));   // verilog/coms.v(128[12] 303[6])
    defparam i15491_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i23248_3_lut (.I0(n414), .I1(n1432), .I2(n1433), .I3(GND_net), 
            .O(n37338));
    defparam i23248_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i1_2_lut (.I0(n1427), .I1(n1428), .I2(GND_net), .I3(GND_net), 
            .O(n51930));
    defparam i1_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_1713 (.I0(n1429), .I1(n37338), .I2(n1430), .I3(n1431), 
            .O(n50013));
    defparam i1_4_lut_adj_1713.LUT_INIT = 16'ha080;
    SB_LUT4 i15851_3_lut (.I0(PWMLimit[10]), .I1(\data_in_frame[9] [2]), 
            .I2(n50654), .I3(GND_net), .O(n29931));   // verilog/coms.v(128[12] 303[6])
    defparam i15851_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15852_3_lut (.I0(PWMLimit[9]), .I1(\data_in_frame[9] [1]), 
            .I2(n50654), .I3(GND_net), .O(n29932));   // verilog/coms.v(128[12] 303[6])
    defparam i15852_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15414_3_lut (.I0(Ki[10]), .I1(\data_in_frame[4] [2]), .I2(n50654), 
            .I3(GND_net), .O(n29494));   // verilog/coms.v(128[12] 303[6])
    defparam i15414_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15415_3_lut (.I0(Ki[9]), .I1(\data_in_frame[4] [1]), .I2(n50654), 
            .I3(GND_net), .O(n29495));   // verilog/coms.v(128[12] 303[6])
    defparam i15415_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1714 (.I0(n1424), .I1(n1425), .I2(n1426), .I3(n51930), 
            .O(n51936));
    defparam i1_4_lut_adj_1714.LUT_INIT = 16'hfffe;
    SB_LUT4 i40572_4_lut (.I0(n1423), .I1(n1422), .I2(n51936), .I3(n50013), 
            .O(n1455));
    defparam i40572_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i15059_2_lut (.I0(n28672), .I1(dti), .I2(GND_net), .I3(GND_net), 
            .O(n29145));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    defparam i15059_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i40063_4_lut (.I0(commutation_state[1]), .I1(n24553), .I2(dti), 
            .I3(commutation_state[2]), .O(n28672));
    defparam i40063_4_lut.LUT_INIT = 16'hc5cf;
    SB_LUT4 i15416_3_lut (.I0(Ki[8]), .I1(\data_in_frame[4] [0]), .I2(n50654), 
            .I3(GND_net), .O(n29496));   // verilog/coms.v(128[12] 303[6])
    defparam i15416_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15853_3_lut (.I0(PWMLimit[8]), .I1(\data_in_frame[9] [0]), 
            .I2(n50654), .I3(GND_net), .O(n29933));   // verilog/coms.v(128[12] 303[6])
    defparam i15853_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i903_3_lut (.I0(n1324), .I1(n1391), 
            .I2(n1356), .I3(GND_net), .O(n1423));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i903_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_adj_1715 (.I0(n1528), .I1(n1527), .I2(GND_net), .I3(GND_net), 
            .O(n51820));
    defparam i1_2_lut_adj_1715.LUT_INIT = 16'heeee;
    SB_LUT4 i15417_3_lut (.I0(Ki[7]), .I1(\data_in_frame[5] [7]), .I2(n50654), 
            .I3(GND_net), .O(n29497));   // verilog/coms.v(128[12] 303[6])
    defparam i15417_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15418_3_lut (.I0(Ki[6]), .I1(\data_in_frame[5] [6]), .I2(n50654), 
            .I3(GND_net), .O(n29498));   // verilog/coms.v(128[12] 303[6])
    defparam i15418_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i23314_4_lut (.I0(n415), .I1(n1531), .I2(n1532_adj_5595), 
            .I3(n1533_adj_5596), .O(n37404));
    defparam i23314_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 i1_4_lut_adj_1716 (.I0(n1524), .I1(n1525), .I2(n1526), .I3(n51820), 
            .O(n51826));
    defparam i1_4_lut_adj_1716.LUT_INIT = 16'hfffe;
    SB_LUT4 i15278_4_lut (.I0(state_7__N_4306[3]), .I1(data[1]), .I2(n10_adj_5610), 
            .I3(n27243), .O(n29358));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i15278_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i15279_4_lut (.I0(state_7__N_4306[3]), .I1(data[2]), .I2(n4_adj_5555), 
            .I3(n27238), .O(n29359));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i15279_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i15419_3_lut (.I0(Ki[5]), .I1(\data_in_frame[5] [5]), .I2(n50654), 
            .I3(GND_net), .O(n29499));   // verilog/coms.v(128[12] 303[6])
    defparam i15419_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15280_4_lut (.I0(state_7__N_4306[3]), .I1(data[3]), .I2(n4_adj_5555), 
            .I3(n27243), .O(n29360));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i15280_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i1_4_lut_adj_1717 (.I0(n1529), .I1(n51826), .I2(n37404), .I3(n1530), 
            .O(n51828));
    defparam i1_4_lut_adj_1717.LUT_INIT = 16'heccc;
    SB_LUT4 i40555_4_lut (.I0(n1522), .I1(n1521), .I2(n51828), .I3(n1523), 
            .O(n1554_adj_5597));
    defparam i40555_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i40568_1_lut (.I0(n1455), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n56399));
    defparam i40568_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i970_3_lut (.I0(n1423), .I1(n1490), 
            .I2(n1455), .I3(GND_net), .O(n1522));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i970_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15281_4_lut (.I0(state_7__N_4306[3]), .I1(data[4]), .I2(n4), 
            .I3(n27238), .O(n29361));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i15281_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i15282_4_lut (.I0(state_7__N_4306[3]), .I1(data[5]), .I2(n4), 
            .I3(n27243), .O(n29362));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i15282_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i23244_3_lut (.I0(n941), .I1(n1632), .I2(n1633), .I3(GND_net), 
            .O(n37334));
    defparam i23244_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i15283_4_lut (.I0(state_7__N_4306[3]), .I1(data[6]), .I2(n36542), 
            .I3(n27238), .O(n29363));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i15283_4_lut.LUT_INIT = 16'hccac;
    SB_LUT4 i15284_4_lut (.I0(state_7__N_4306[3]), .I1(data[7]), .I2(n36542), 
            .I3(n27243), .O(n29364));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i15284_4_lut.LUT_INIT = 16'hccac;
    SB_LUT4 i15422_3_lut (.I0(Ki[4]), .I1(\data_in_frame[5] [4]), .I2(n50654), 
            .I3(GND_net), .O(n29502));   // verilog/coms.v(128[12] 303[6])
    defparam i15422_3_lut.LUT_INIT = 16'hacac;
    SB_DFFESR delay_counter_i0_i1 (.Q(delay_counter[1]), .C(clk16MHz), .E(n7593), 
            .D(n1562), .R(n29242));   // verilog/TinyFPGA_B.v(368[10] 396[6])
    SB_LUT4 i15423_3_lut (.I0(Ki[3]), .I1(\data_in_frame[5] [3]), .I2(n50654), 
            .I3(GND_net), .O(n29503));   // verilog/coms.v(128[12] 303[6])
    defparam i15423_3_lut.LUT_INIT = 16'hacac;
    SB_DFFESR delay_counter_i0_i2 (.Q(delay_counter[2]), .C(clk16MHz), .E(n7593), 
            .D(n1561), .R(n29242));   // verilog/TinyFPGA_B.v(368[10] 396[6])
    SB_DFFESR delay_counter_i0_i3 (.Q(delay_counter[3]), .C(clk16MHz), .E(n7593), 
            .D(n1560), .R(n29242));   // verilog/TinyFPGA_B.v(368[10] 396[6])
    SB_DFFESR delay_counter_i0_i4 (.Q(delay_counter[4]), .C(clk16MHz), .E(n7593), 
            .D(n1559), .R(n29242));   // verilog/TinyFPGA_B.v(368[10] 396[6])
    SB_DFFESR delay_counter_i0_i5 (.Q(delay_counter[5]), .C(clk16MHz), .E(n7593), 
            .D(n1558), .R(n29242));   // verilog/TinyFPGA_B.v(368[10] 396[6])
    SB_DFFESR delay_counter_i0_i6 (.Q(delay_counter[6]), .C(clk16MHz), .E(n7593), 
            .D(n1557), .R(n29242));   // verilog/TinyFPGA_B.v(368[10] 396[6])
    SB_DFFESR delay_counter_i0_i7 (.Q(delay_counter[7]), .C(clk16MHz), .E(n7593), 
            .D(n1556), .R(n29242));   // verilog/TinyFPGA_B.v(368[10] 396[6])
    SB_DFFESR delay_counter_i0_i8 (.Q(delay_counter[8]), .C(clk16MHz), .E(n7593), 
            .D(n1555), .R(n29242));   // verilog/TinyFPGA_B.v(368[10] 396[6])
    SB_DFFESR delay_counter_i0_i9 (.Q(delay_counter[9]), .C(clk16MHz), .E(n7593), 
            .D(n1554), .R(n29242));   // verilog/TinyFPGA_B.v(368[10] 396[6])
    SB_DFFESR delay_counter_i0_i10 (.Q(delay_counter[10]), .C(clk16MHz), 
            .E(n7593), .D(n1553), .R(n29242));   // verilog/TinyFPGA_B.v(368[10] 396[6])
    SB_DFFESR delay_counter_i0_i11 (.Q(delay_counter[11]), .C(clk16MHz), 
            .E(n7593), .D(n1552), .R(n29242));   // verilog/TinyFPGA_B.v(368[10] 396[6])
    SB_LUT4 i15288_3_lut (.I0(IntegralLimit[0]), .I1(\data_in_frame[13] [0]), 
            .I2(n50654), .I3(GND_net), .O(n29368));   // verilog/coms.v(128[12] 303[6])
    defparam i15288_3_lut.LUT_INIT = 16'hacac;
    SB_DFFESR delay_counter_i0_i12 (.Q(delay_counter[12]), .C(clk16MHz), 
            .E(n7593), .D(n1551), .R(n29242));   // verilog/TinyFPGA_B.v(368[10] 396[6])
    SB_DFFESR delay_counter_i0_i13 (.Q(delay_counter[13]), .C(clk16MHz), 
            .E(n7593), .D(n1550), .R(n29242));   // verilog/TinyFPGA_B.v(368[10] 396[6])
    SB_LUT4 i15424_3_lut (.I0(Ki[2]), .I1(\data_in_frame[5] [2]), .I2(n50654), 
            .I3(GND_net), .O(n29504));   // verilog/coms.v(128[12] 303[6])
    defparam i15424_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1718 (.I0(n1629), .I1(n37334), .I2(n1630), .I3(n1631), 
            .O(n50021));
    defparam i1_4_lut_adj_1718.LUT_INIT = 16'ha080;
    SB_DFFESR delay_counter_i0_i14 (.Q(delay_counter[14]), .C(clk16MHz), 
            .E(n7593), .D(n1549), .R(n29242));   // verilog/TinyFPGA_B.v(368[10] 396[6])
    SB_LUT4 i15289_3_lut (.I0(Kp[0]), .I1(\data_in_frame[3] [0]), .I2(n50654), 
            .I3(GND_net), .O(n29369));   // verilog/coms.v(128[12] 303[6])
    defparam i15289_3_lut.LUT_INIT = 16'hacac;
    SB_DFFESR delay_counter_i0_i15 (.Q(delay_counter[15]), .C(clk16MHz), 
            .E(n7593), .D(n1548), .R(n29242));   // verilog/TinyFPGA_B.v(368[10] 396[6])
    SB_DFFESR delay_counter_i0_i16 (.Q(delay_counter[16]), .C(clk16MHz), 
            .E(n7593), .D(n1547), .R(n29242));   // verilog/TinyFPGA_B.v(368[10] 396[6])
    SB_LUT4 i15290_3_lut (.I0(Ki[0]), .I1(\data_in_frame[5] [0]), .I2(n50654), 
            .I3(GND_net), .O(n29370));   // verilog/coms.v(128[12] 303[6])
    defparam i15290_3_lut.LUT_INIT = 16'hacac;
    SB_DFFESR delay_counter_i0_i17 (.Q(delay_counter[17]), .C(clk16MHz), 
            .E(n7593), .D(n1546), .R(n29242));   // verilog/TinyFPGA_B.v(368[10] 396[6])
    SB_DFFESR delay_counter_i0_i18 (.Q(delay_counter[18]), .C(clk16MHz), 
            .E(n7593), .D(n1545), .R(n29242));   // verilog/TinyFPGA_B.v(368[10] 396[6])
    SB_DFFESR delay_counter_i0_i19 (.Q(delay_counter[19]), .C(clk16MHz), 
            .E(n7593), .D(n1544), .R(n29242));   // verilog/TinyFPGA_B.v(368[10] 396[6])
    SB_LUT4 i1_4_lut_adj_1719 (.I0(n1623), .I1(n50021), .I2(n1625), .I3(n1628), 
            .O(n51960));
    defparam i1_4_lut_adj_1719.LUT_INIT = 16'hfffe;
    SB_DFFESR delay_counter_i0_i20 (.Q(delay_counter[20]), .C(clk16MHz), 
            .E(n7593), .D(n1543), .R(n29242));   // verilog/TinyFPGA_B.v(368[10] 396[6])
    SB_DFFESR delay_counter_i0_i21 (.Q(delay_counter[21]), .C(clk16MHz), 
            .E(n7593), .D(n1542), .R(n29242));   // verilog/TinyFPGA_B.v(368[10] 396[6])
    SB_DFFESR delay_counter_i0_i22 (.Q(delay_counter[22]), .C(clk16MHz), 
            .E(n7593), .D(n1541), .R(n29242));   // verilog/TinyFPGA_B.v(368[10] 396[6])
    SB_DFFESR delay_counter_i0_i23 (.Q(delay_counter[23]), .C(clk16MHz), 
            .E(n7593), .D(n1540), .R(n29242));   // verilog/TinyFPGA_B.v(368[10] 396[6])
    SB_LUT4 i15291_3_lut (.I0(\data_in[0] [0]), .I1(\data_in[1] [0]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n29371));   // verilog/coms.v(128[12] 303[6])
    defparam i15291_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFESR delay_counter_i0_i24 (.Q(delay_counter[24]), .C(clk16MHz), 
            .E(n7593), .D(n1539), .R(n29242));   // verilog/TinyFPGA_B.v(368[10] 396[6])
    SB_DFFESR delay_counter_i0_i25 (.Q(delay_counter[25]), .C(clk16MHz), 
            .E(n7593), .D(n1538), .R(n29242));   // verilog/TinyFPGA_B.v(368[10] 396[6])
    SB_DFFESR delay_counter_i0_i26 (.Q(delay_counter[26]), .C(clk16MHz), 
            .E(n7593), .D(n1537), .R(n29242));   // verilog/TinyFPGA_B.v(368[10] 396[6])
    SB_DFFESR delay_counter_i0_i27 (.Q(delay_counter[27]), .C(clk16MHz), 
            .E(n7593), .D(n1536), .R(n29242));   // verilog/TinyFPGA_B.v(368[10] 396[6])
    SB_DFFESR delay_counter_i0_i28 (.Q(delay_counter[28]), .C(clk16MHz), 
            .E(n7593), .D(n1535), .R(n29242));   // verilog/TinyFPGA_B.v(368[10] 396[6])
    SB_DFFESR delay_counter_i0_i29 (.Q(delay_counter[29]), .C(clk16MHz), 
            .E(n7593), .D(n1534), .R(n29242));   // verilog/TinyFPGA_B.v(368[10] 396[6])
    SB_DFFESR delay_counter_i0_i30 (.Q(delay_counter[30]), .C(clk16MHz), 
            .E(n7593), .D(n1533), .R(n29242));   // verilog/TinyFPGA_B.v(368[10] 396[6])
    SB_DFFESR delay_counter_i0_i31 (.Q(delay_counter[31]), .C(clk16MHz), 
            .E(n7593), .D(n1532), .R(n29242));   // verilog/TinyFPGA_B.v(368[10] 396[6])
    SB_LUT4 i15425_3_lut (.I0(Ki[1]), .I1(\data_in_frame[5] [1]), .I2(n50654), 
            .I3(GND_net), .O(n29505));   // verilog/coms.v(128[12] 303[6])
    defparam i15425_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15294_3_lut (.I0(control_mode[0]), .I1(\data_in_frame[1] [0]), 
            .I2(n50654), .I3(GND_net), .O(n29374));   // verilog/coms.v(128[12] 303[6])
    defparam i15294_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1720 (.I0(n1624), .I1(n1622), .I2(n1626), .I3(n1627), 
            .O(n51149));
    defparam i1_4_lut_adj_1720.LUT_INIT = 16'hfffe;
    SB_LUT4 i40537_4_lut (.I0(n51149), .I1(n1620), .I2(n1621), .I3(n51960), 
            .O(n1653));
    defparam i40537_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1037_3_lut (.I0(n1522), 
            .I1(n1589), .I2(n1554_adj_5597), .I3(GND_net), .O(n1621));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1037_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15295_3_lut (.I0(current_limit[0]), .I1(\data_in_frame[21] [0]), 
            .I2(n50654), .I3(GND_net), .O(n29375));   // verilog/coms.v(128[12] 303[6])
    defparam i15295_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15426_3_lut (.I0(Kp[15]), .I1(\data_in_frame[2] [7]), .I2(n50654), 
            .I3(GND_net), .O(n29506));   // verilog/coms.v(128[12] 303[6])
    defparam i15426_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_3_lut_adj_1721 (.I0(n1726), .I1(n1728), .I2(n1727), .I3(GND_net), 
            .O(n51850));
    defparam i1_3_lut_adj_1721.LUT_INIT = 16'hfefe;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_mux_3_i25_3_lut (.I0(encoder0_position_scaled_23__N_327[24]), 
            .I1(n9_adj_5490), .I2(encoder0_position_scaled_23__N_327[31]), 
            .I3(GND_net), .O(n934));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_mux_3_i25_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i641_3_lut (.I0(n934), .I1(n1001), 
            .I2(n960), .I3(GND_net), .O(n1033));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i641_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i708_3_lut (.I0(n1033), .I1(n1100), 
            .I2(n1059), .I3(GND_net), .O(n1132));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i708_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i23310_4_lut (.I0(n942), .I1(n1731), .I2(n1732), .I3(n1733), 
            .O(n37400));
    defparam i23310_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 i1_4_lut_adj_1722 (.I0(n1723), .I1(n1724), .I2(n51850), .I3(n1725), 
            .O(n51856));
    defparam i1_4_lut_adj_1722.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_adj_1723 (.I0(n1729), .I1(n1730), .I2(GND_net), .I3(GND_net), 
            .O(n51954));
    defparam i1_2_lut_adj_1723.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut_adj_1724 (.I0(n51954), .I1(n1722), .I2(n51856), .I3(n37400), 
            .O(n51860));
    defparam i1_4_lut_adj_1724.LUT_INIT = 16'hfefc;
    SB_LUT4 i40518_4_lut (.I0(n1720), .I1(n1719), .I2(n1721), .I3(n51860), 
            .O(n1752));
    defparam i40518_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1104_3_lut (.I0(n1621), 
            .I1(n1688), .I2(n1653), .I3(GND_net), .O(n1720));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1104_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1725 (.I0(n1827), .I1(n1826), .I2(n1825), .I3(n1828), 
            .O(n51980));
    defparam i1_4_lut_adj_1725.LUT_INIT = 16'hfffe;
    SB_LUT4 i23308_4_lut (.I0(n529), .I1(n1831), .I2(n1832), .I3(n1833), 
            .O(n37398));
    defparam i23308_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 i1_4_lut_adj_1726 (.I0(n1822), .I1(n1823), .I2(n1824), .I3(n51980), 
            .O(n51986));
    defparam i1_4_lut_adj_1726.LUT_INIT = 16'hfffe;
    SB_LUT4 i15427_3_lut (.I0(Kp[14]), .I1(\data_in_frame[2] [6]), .I2(n50654), 
            .I3(GND_net), .O(n29507));   // verilog/coms.v(128[12] 303[6])
    defparam i15427_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_adj_1727 (.I0(n1829), .I1(n1830), .I2(GND_net), .I3(GND_net), 
            .O(n52132));
    defparam i1_2_lut_adj_1727.LUT_INIT = 16'h8888;
    SB_LUT4 mux_1037_i1_4_lut (.I0(n54531), .I1(duty[0]), .I2(n296), .I3(n356), 
            .O(n4929));   // verilog/TinyFPGA_B.v(123[17] 125[11])
    defparam mux_1037_i1_4_lut.LUT_INIT = 16'h3a30;
    SB_LUT4 i1_4_lut_adj_1728 (.I0(n1821), .I1(n52132), .I2(n51986), .I3(n37398), 
            .O(n51990));
    defparam i1_4_lut_adj_1728.LUT_INIT = 16'hfefa;
    SB_LUT4 i15428_3_lut (.I0(Kp[13]), .I1(\data_in_frame[2] [5]), .I2(n50654), 
            .I3(GND_net), .O(n29508));   // verilog/coms.v(128[12] 303[6])
    defparam i15428_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15429_3_lut (.I0(Kp[12]), .I1(\data_in_frame[2] [4]), .I2(n50654), 
            .I3(GND_net), .O(n29509));   // verilog/coms.v(128[12] 303[6])
    defparam i15429_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i34007_3_lut (.I0(n6_adj_5493), .I1(n8585), .I2(n49748), .I3(GND_net), 
            .O(n49755));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam i34007_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34008_3_lut (.I0(encoder0_position_scaled_23__N_327[27]), .I1(n49755), 
            .I2(encoder0_position_scaled_23__N_327[31]), .I3(GND_net), .O(n832));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam i34008_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i571_3_lut (.I0(n832), .I1(n899), 
            .I2(n861), .I3(GND_net), .O(n931));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i571_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i638_3_lut (.I0(n931), .I1(n998), 
            .I2(n960), .I3(GND_net), .O(n1030));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i638_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i40496_4_lut (.I0(n1819), .I1(n1818), .I2(n1820), .I3(n51990), 
            .O(n1851));
    defparam i40496_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i705_3_lut (.I0(n1030), .I1(n1097), 
            .I2(n1059), .I3(GND_net), .O(n1129));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i705_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1171_3_lut (.I0(n1720), 
            .I1(n1787), .I2(n1752), .I3(GND_net), .O(n1819));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1171_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1729 (.I0(n1928), .I1(n1925), .I2(n1927), .I3(n1926), 
            .O(n51760));
    defparam i1_4_lut_adj_1729.LUT_INIT = 16'hfffe;
    SB_LUT4 i15430_3_lut (.I0(Kp[11]), .I1(\data_in_frame[2] [3]), .I2(n50654), 
            .I3(GND_net), .O(n29510));   // verilog/coms.v(128[12] 303[6])
    defparam i15430_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15431_3_lut (.I0(Kp[10]), .I1(\data_in_frame[2] [2]), .I2(n50654), 
            .I3(GND_net), .O(n29511));   // verilog/coms.v(128[12] 303[6])
    defparam i15431_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i34005_3_lut (.I0(n5_adj_5494), .I1(n8584), .I2(n49748), .I3(GND_net), 
            .O(n49753));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam i34005_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34006_3_lut (.I0(encoder0_position_scaled_23__N_327[28]), .I1(n49753), 
            .I2(encoder0_position_scaled_23__N_327[31]), .I3(GND_net), .O(n831));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam i34006_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i570_3_lut (.I0(n831), .I1(n898), 
            .I2(n861), .I3(GND_net), .O(n930));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i570_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i637_3_lut (.I0(n930), .I1(n997), 
            .I2(n960), .I3(GND_net), .O(n1029));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i637_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i704_3_lut (.I0(n1029), .I1(n1096), 
            .I2(n1059), .I3(GND_net), .O(n1128));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i704_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i23238_3_lut (.I0(n530), .I1(n1932), .I2(n1933), .I3(GND_net), 
            .O(n37328));
    defparam i23238_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i1_4_lut_adj_1730 (.I0(n1922), .I1(n1923), .I2(n51760), .I3(n1924), 
            .O(n51766));
    defparam i1_4_lut_adj_1730.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1731 (.I0(n1929), .I1(n37328), .I2(n1930), .I3(n1931), 
            .O(n50043));
    defparam i1_4_lut_adj_1731.LUT_INIT = 16'ha080;
    SB_LUT4 i1_4_lut_adj_1732 (.I0(n1920), .I1(n50043), .I2(n1921), .I3(n51766), 
            .O(n51772));
    defparam i1_4_lut_adj_1732.LUT_INIT = 16'hfffe;
    SB_LUT4 i40475_4_lut (.I0(n1918), .I1(n1917), .I2(n1919), .I3(n51772), 
            .O(n1950));
    defparam i40475_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1238_3_lut (.I0(n1819), 
            .I1(n1886), .I2(n1851), .I3(GND_net), .O(n1918));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1238_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 RX_I_0_1_lut (.I0(RX_c), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(RX_N_10));   // verilog/TinyFPGA_B.v(260[10:13])
    defparam RX_I_0_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i23304_4_lut (.I0(n531), .I1(n2031), .I2(n2032), .I3(n2033), 
            .O(n37394));
    defparam i23304_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 i1_3_lut_adj_1733 (.I0(n2025), .I1(n2027), .I2(n2024), .I3(GND_net), 
            .O(n52010));
    defparam i1_3_lut_adj_1733.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_2_lut_adj_1734 (.I0(n2028), .I1(n2026), .I2(GND_net), .I3(GND_net), 
            .O(n52020));
    defparam i1_2_lut_adj_1734.LUT_INIT = 16'heeee;
    SB_LUT4 i22679_2_lut (.I0(duty[1]), .I1(n296), .I2(GND_net), .I3(GND_net), 
            .O(n4928));   // verilog/TinyFPGA_B.v(123[17] 125[11])
    defparam i22679_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i1_4_lut_adj_1735 (.I0(n2021), .I1(n2022), .I2(n2023), .I3(n52020), 
            .O(n52026));
    defparam i1_4_lut_adj_1735.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1736 (.I0(n2029), .I1(n52010), .I2(n37394), .I3(n2030), 
            .O(n52012));
    defparam i1_4_lut_adj_1736.LUT_INIT = 16'heccc;
    SB_LUT4 i1_4_lut_adj_1737 (.I0(n48957), .I1(\FRAME_MATCHER.state [0]), 
            .I2(n4_adj_5472), .I3(n22875), .O(n40_adj_5592));   // verilog/coms.v(128[12] 303[6])
    defparam i1_4_lut_adj_1737.LUT_INIT = 16'hc8fa;
    SB_LUT4 i1_4_lut_adj_1738 (.I0(n2019), .I1(n2018), .I2(n2020), .I3(n52026), 
            .O(n50932));
    defparam i1_4_lut_adj_1738.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_3_lut_adj_1739 (.I0(n27219), .I1(n48947), .I2(n3303), .I3(GND_net), 
            .O(n21_adj_5593));   // verilog/coms.v(128[12] 303[6])
    defparam i1_3_lut_adj_1739.LUT_INIT = 16'hcdcd;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i973_3_lut (.I0(n1426), .I1(n1493), 
            .I2(n1455), .I3(GND_net), .O(n1525));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i973_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i40453_4_lut (.I0(n2017), .I1(n2016), .I2(n50932), .I3(n52012), 
            .O(n2049));
    defparam i40453_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1305_3_lut (.I0(n1918), 
            .I1(n1985), .I2(n1950), .I3(GND_net), .O(n2017));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1305_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1740 (.I0(n40_adj_5592), .I1(\FRAME_MATCHER.state [3]), 
            .I2(n6_adj_5645), .I3(\FRAME_MATCHER.state [0]), .O(n4_adj_5473));   // verilog/coms.v(128[12] 303[6])
    defparam i1_4_lut_adj_1740.LUT_INIT = 16'haaae;
    SB_LUT4 i15835_3_lut (.I0(\PID_CONTROLLER.integral [1]), .I1(\PID_CONTROLLER.integral_23__N_3996 [1]), 
            .I2(control_update), .I3(GND_net), .O(n29915));   // verilog/motorControl.v(41[14] 61[8])
    defparam i15835_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2_4_lut (.I0(\FRAME_MATCHER.state [0]), .I1(n4_adj_5473), .I2(n21_adj_5593), 
            .I3(n22875), .O(n50741));   // verilog/coms.v(128[12] 303[6])
    defparam i2_4_lut.LUT_INIT = 16'hecfc;
    SB_LUT4 unary_minus_18_inv_0_i2_1_lut (.I0(duty[1]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n24));   // verilog/TinyFPGA_B.v(119[24:29])
    defparam unary_minus_18_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_2_lut_adj_1741 (.I0(n2126), .I1(n2127), .I2(GND_net), .I3(GND_net), 
            .O(n51614));
    defparam i1_2_lut_adj_1741.LUT_INIT = 16'heeee;
    SB_LUT4 i40613_1_lut (.I0(n1158), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n56444));
    defparam i40613_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i701_3_lut (.I0(n1026), .I1(n1093), 
            .I2(n1059), .I3(GND_net), .O(n1125));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i701_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_unary_minus_2_inv_0_i1_1_lut (.I0(encoder0_position[0]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n33_adj_5642));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_unary_minus_2_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_4_lut_adj_1742 (.I0(n2125), .I1(n51614), .I2(n2124), .I3(n2128), 
            .O(n51618));
    defparam i1_4_lut_adj_1742.LUT_INIT = 16'hfffe;
    SB_LUT4 i23302_4_lut (.I0(n532), .I1(n2131), .I2(n2132), .I3(n2133), 
            .O(n37392));
    defparam i23302_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 i15836_4_lut (.I0(CS_MISO_c), .I1(data_adj_5711[9]), .I2(n5_adj_5557), 
            .I3(n27198), .O(n29916));   // verilog/tli4970.v(35[10] 68[6])
    defparam i15836_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i15298_3_lut (.I0(\data_out_frame[11] [4]), .I1(encoder1_position_scaled[4]), 
            .I2(n24210), .I3(GND_net), .O(n29378));   // verilog/coms.v(128[12] 303[6])
    defparam i15298_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_281_i23_4_lut (.I0(encoder1_position_scaled[22]), .I1(displacement[22]), 
            .I2(n15), .I3(n15_adj_5471), .O(motor_state_23__N_123[22]));   // verilog/TinyFPGA_B.v(284[5] 286[10])
    defparam mux_281_i23_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i15299_3_lut (.I0(\data_out_frame[11] [3]), .I1(encoder1_position_scaled[3]), 
            .I2(n24210), .I3(GND_net), .O(n29379));   // verilog/coms.v(128[12] 303[6])
    defparam i15299_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15300_3_lut (.I0(\data_out_frame[11] [2]), .I1(encoder1_position_scaled[2]), 
            .I2(n24210), .I3(GND_net), .O(n29380));   // verilog/coms.v(128[12] 303[6])
    defparam i15300_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15301_3_lut (.I0(\PID_CONTROLLER.integral [0]), .I1(\PID_CONTROLLER.integral_23__N_3996 [0]), 
            .I2(control_update), .I3(GND_net), .O(n29381));   // verilog/motorControl.v(41[14] 61[8])
    defparam i15301_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15302_3_lut (.I0(\data_out_frame[11] [1]), .I1(encoder1_position_scaled[1]), 
            .I2(n24210), .I3(GND_net), .O(n29382));   // verilog/coms.v(128[12] 303[6])
    defparam i15302_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15303_3_lut (.I0(\data_out_frame[11] [0]), .I1(encoder1_position_scaled[0]), 
            .I2(n24210), .I3(GND_net), .O(n29383));   // verilog/coms.v(128[12] 303[6])
    defparam i15303_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15304_3_lut (.I0(\data_out_frame[10] [7]), .I1(encoder1_position_scaled[15]), 
            .I2(n24210), .I3(GND_net), .O(n29384));   // verilog/coms.v(128[12] 303[6])
    defparam i15304_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1743 (.I0(n2121), .I1(n2122), .I2(n51618), .I3(n2123), 
            .O(n51624));
    defparam i1_4_lut_adj_1743.LUT_INIT = 16'hfffe;
    SB_LUT4 i15305_3_lut (.I0(\data_out_frame[10] [6]), .I1(encoder1_position_scaled[14]), 
            .I2(n24210), .I3(GND_net), .O(n29385));   // verilog/coms.v(128[12] 303[6])
    defparam i15305_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15306_3_lut (.I0(\data_out_frame[10] [5]), .I1(encoder1_position_scaled[13]), 
            .I2(n24210), .I3(GND_net), .O(n29386));   // verilog/coms.v(128[12] 303[6])
    defparam i15306_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15307_3_lut (.I0(\data_out_frame[10] [4]), .I1(encoder1_position_scaled[12]), 
            .I2(n24210), .I3(GND_net), .O(n29387));   // verilog/coms.v(128[12] 303[6])
    defparam i15307_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15308_3_lut (.I0(\data_out_frame[10] [3]), .I1(encoder1_position_scaled[11]), 
            .I2(n24210), .I3(GND_net), .O(n29388));   // verilog/coms.v(128[12] 303[6])
    defparam i15308_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1744 (.I0(n2129), .I1(n51624), .I2(n37392), .I3(n2130), 
            .O(n51626));
    defparam i1_4_lut_adj_1744.LUT_INIT = 16'heccc;
    SB_LUT4 i15854_3_lut (.I0(PWMLimit[7]), .I1(\data_in_frame[10] [7]), 
            .I2(n50654), .I3(GND_net), .O(n29934));   // verilog/coms.v(128[12] 303[6])
    defparam i15854_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1745 (.I0(n27218), .I1(n63_adj_5605), .I2(n19602), 
            .I3(n48957), .O(n5_adj_5594));   // verilog/coms.v(128[12] 303[6])
    defparam i1_4_lut_adj_1745.LUT_INIT = 16'hdc50;
    SB_LUT4 i3_4_lut_adj_1746 (.I0(n7_adj_5608), .I1(\FRAME_MATCHER.state_31__N_3007 [2]), 
            .I2(n8_adj_5609), .I3(n27219), .O(n8_adj_5646));   // verilog/coms.v(128[12] 303[6])
    defparam i3_4_lut_adj_1746.LUT_INIT = 16'hfafe;
    SB_LUT4 i22678_2_lut (.I0(duty[2]), .I1(n296), .I2(GND_net), .I3(GND_net), 
            .O(n4927));   // verilog/TinyFPGA_B.v(123[17] 125[11])
    defparam i22678_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i1_4_lut_adj_1747 (.I0(n2118), .I1(n2119), .I2(n2120), .I3(n51626), 
            .O(n51632));
    defparam i1_4_lut_adj_1747.LUT_INIT = 16'hfffe;
    SB_LUT4 i15855_3_lut (.I0(PWMLimit[6]), .I1(\data_in_frame[10] [6]), 
            .I2(n50654), .I3(GND_net), .O(n29935));   // verilog/coms.v(128[12] 303[6])
    defparam i15855_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i4_4_lut (.I0(n122), .I1(n8_adj_5646), .I2(n63), .I3(n5_adj_5594), 
            .O(n57033));   // verilog/coms.v(128[12] 303[6])
    defparam i4_4_lut.LUT_INIT = 16'hefcf;
    SB_LUT4 i40430_4_lut (.I0(n2116), .I1(n2115), .I2(n2117), .I3(n51632), 
            .O(n2148));
    defparam i40430_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1771_20_lut (.I0(GND_net), 
            .I1(n2616), .I2(VCC_net), .I3(n44245), .O(n2683)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1771_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1771_20 (.CI(n44245), 
            .I0(n2616), .I1(VCC_net), .CO(n44246));
    SB_LUT4 i15856_3_lut (.I0(PWMLimit[5]), .I1(\data_in_frame[10] [5]), 
            .I2(n50654), .I3(GND_net), .O(n29936));   // verilog/coms.v(128[12] 303[6])
    defparam i15856_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15857_3_lut (.I0(PWMLimit[4]), .I1(\data_in_frame[10] [4]), 
            .I2(n50654), .I3(GND_net), .O(n29937));   // verilog/coms.v(128[12] 303[6])
    defparam i15857_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1372_3_lut (.I0(n2017), 
            .I1(n2084), .I2(n2049), .I3(GND_net), .O(n2116));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1372_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15309_3_lut (.I0(\data_out_frame[10] [2]), .I1(encoder1_position_scaled[10]), 
            .I2(n24210), .I3(GND_net), .O(n29389));   // verilog/coms.v(128[12] 303[6])
    defparam i15309_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15858_3_lut (.I0(PWMLimit[3]), .I1(\data_in_frame[10] [3]), 
            .I2(n50654), .I3(GND_net), .O(n29938));   // verilog/coms.v(128[12] 303[6])
    defparam i15858_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1440_3_lut (.I0(n2117), 
            .I1(n2184), .I2(n2148), .I3(GND_net), .O(n2216));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1440_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1439_3_lut (.I0(n2116), 
            .I1(n2183), .I2(n2148), .I3(GND_net), .O(n2215));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1439_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15310_3_lut (.I0(\data_out_frame[10] [1]), .I1(encoder1_position_scaled[9]), 
            .I2(n24210), .I3(GND_net), .O(n29390));   // verilog/coms.v(128[12] 303[6])
    defparam i15310_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15859_3_lut (.I0(PWMLimit[2]), .I1(\data_in_frame[10] [2]), 
            .I2(n50654), .I3(GND_net), .O(n29939));   // verilog/coms.v(128[12] 303[6])
    defparam i15859_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15860_3_lut (.I0(PWMLimit[1]), .I1(\data_in_frame[10] [1]), 
            .I2(n50654), .I3(GND_net), .O(n29940));   // verilog/coms.v(128[12] 303[6])
    defparam i15860_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15838_3_lut (.I0(PWMLimit[23]), .I1(\data_in_frame[8] [7]), 
            .I2(n50654), .I3(GND_net), .O(n29918));   // verilog/coms.v(128[12] 303[6])
    defparam i15838_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15861_3_lut (.I0(current_limit[15]), .I1(\data_in_frame[20] [7]), 
            .I2(n50654), .I3(GND_net), .O(n29941));   // verilog/coms.v(128[12] 303[6])
    defparam i15861_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15862_3_lut (.I0(current_limit[14]), .I1(\data_in_frame[20] [6]), 
            .I2(n50654), .I3(GND_net), .O(n29942));   // verilog/coms.v(128[12] 303[6])
    defparam i15862_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15839_3_lut (.I0(PWMLimit[22]), .I1(\data_in_frame[8] [6]), 
            .I2(n50654), .I3(GND_net), .O(n29919));   // verilog/coms.v(128[12] 303[6])
    defparam i15839_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15863_3_lut (.I0(current_limit[13]), .I1(\data_in_frame[20] [5]), 
            .I2(n50654), .I3(GND_net), .O(n29943));   // verilog/coms.v(128[12] 303[6])
    defparam i15863_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15864_3_lut (.I0(current_limit[12]), .I1(\data_in_frame[20] [4]), 
            .I2(n50654), .I3(GND_net), .O(n29944));   // verilog/coms.v(128[12] 303[6])
    defparam i15864_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15432_3_lut (.I0(Kp[9]), .I1(\data_in_frame[2] [1]), .I2(n50654), 
            .I3(GND_net), .O(n29512));   // verilog/coms.v(128[12] 303[6])
    defparam i15432_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i22677_2_lut (.I0(duty[3]), .I1(n296), .I2(GND_net), .I3(GND_net), 
            .O(n4926));   // verilog/TinyFPGA_B.v(123[17] 125[11])
    defparam i22677_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i15311_3_lut (.I0(current[0]), .I1(data_adj_5711[0]), .I2(n28729), 
            .I3(GND_net), .O(n29391));   // verilog/tli4970.v(35[10] 68[6])
    defparam i15311_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15865_3_lut (.I0(current_limit[11]), .I1(\data_in_frame[20] [3]), 
            .I2(n50654), .I3(GND_net), .O(n29945));   // verilog/coms.v(128[12] 303[6])
    defparam i15865_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15866_3_lut (.I0(current_limit[10]), .I1(\data_in_frame[20] [2]), 
            .I2(n50654), .I3(GND_net), .O(n29946));   // verilog/coms.v(128[12] 303[6])
    defparam i15866_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1748 (.I0(control_mode[3]), .I1(control_mode[4]), 
            .I2(control_mode[2]), .I3(control_mode[6]), .O(n52298));   // verilog/TinyFPGA_B.v(284[5:22])
    defparam i1_4_lut_adj_1748.LUT_INIT = 16'hfffe;
    SB_LUT4 i15867_3_lut (.I0(current_limit[9]), .I1(\data_in_frame[20] [1]), 
            .I2(n50654), .I3(GND_net), .O(n29947));   // verilog/coms.v(128[12] 303[6])
    defparam i15867_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_3_lut_adj_1749 (.I0(n52298), .I1(control_mode[7]), .I2(control_mode[5]), 
            .I3(GND_net), .O(n27261));   // verilog/TinyFPGA_B.v(284[5:22])
    defparam i1_3_lut_adj_1749.LUT_INIT = 16'hfefe;
    SB_LUT4 i15868_3_lut (.I0(current_limit[8]), .I1(\data_in_frame[20] [0]), 
            .I2(n50654), .I3(GND_net), .O(n29948));   // verilog/coms.v(128[12] 303[6])
    defparam i15868_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15869_3_lut (.I0(current_limit[7]), .I1(\data_in_frame[21] [7]), 
            .I2(n50654), .I3(GND_net), .O(n29949));   // verilog/coms.v(128[12] 303[6])
    defparam i15869_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1750 (.I0(n2224), .I1(n2228), .I2(n2223), .I3(n2226), 
            .O(n52038));
    defparam i1_4_lut_adj_1750.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_3_lut_adj_1751 (.I0(n52038), .I1(n2227), .I2(n2225), .I3(GND_net), 
            .O(n52040));
    defparam i1_3_lut_adj_1751.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_2_lut_adj_1752 (.I0(n27100), .I1(control_mode[1]), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_5471));   // verilog/TinyFPGA_B.v(285[5:22])
    defparam i1_2_lut_adj_1752.LUT_INIT = 16'hbbbb;
    SB_LUT4 i15870_3_lut (.I0(current_limit[6]), .I1(\data_in_frame[21] [6]), 
            .I2(n50654), .I3(GND_net), .O(n29950));   // verilog/coms.v(128[12] 303[6])
    defparam i15870_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_3_lut_adj_1753 (.I0(control_mode[0]), .I1(n27261), .I2(control_mode[1]), 
            .I3(GND_net), .O(n15));   // verilog/TinyFPGA_B.v(284[5:22])
    defparam i1_3_lut_adj_1753.LUT_INIT = 16'hfdfd;
    SB_LUT4 i23300_4_lut (.I0(n533), .I1(n2231), .I2(n2232), .I3(n2233_adj_5599), 
            .O(n37390));
    defparam i23300_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 i1_4_lut_adj_1754 (.I0(n2220), .I1(n2221), .I2(n52040), .I3(n2222), 
            .O(n52046));
    defparam i1_4_lut_adj_1754.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1755 (.I0(n2229), .I1(n52046), .I2(n37390), .I3(n2230), 
            .O(n52048));
    defparam i1_4_lut_adj_1755.LUT_INIT = 16'heccc;
    SB_LUT4 i1_4_lut_adj_1756 (.I0(n2217), .I1(n2218), .I2(n2219), .I3(n52048), 
            .O(n52054));
    defparam i1_4_lut_adj_1756.LUT_INIT = 16'hfffe;
    SB_LUT4 i15871_3_lut (.I0(current_limit[5]), .I1(\data_in_frame[21] [5]), 
            .I2(n50654), .I3(GND_net), .O(n29951));   // verilog/coms.v(128[12] 303[6])
    defparam i15871_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_281_i24_4_lut (.I0(encoder1_position_scaled[23]), .I1(displacement[23]), 
            .I2(n15), .I3(n15_adj_5471), .O(motor_state_23__N_123[23]));   // verilog/TinyFPGA_B.v(284[5] 286[10])
    defparam mux_281_i24_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i15872_3_lut (.I0(current_limit[4]), .I1(\data_in_frame[21] [4]), 
            .I2(n50654), .I3(GND_net), .O(n29952));   // verilog/coms.v(128[12] 303[6])
    defparam i15872_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i40405_4_lut (.I0(n2215), .I1(n2214), .I2(n2216), .I3(n52054), 
            .O(n2247));
    defparam i40405_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1450_rep_28_3_lut (.I0(n2127), 
            .I1(n2194), .I2(n2148), .I3(GND_net), .O(n2226));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1450_rep_28_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15433_3_lut (.I0(Kp[8]), .I1(\data_in_frame[2] [0]), .I2(n50654), 
            .I3(GND_net), .O(n29513));   // verilog/coms.v(128[12] 303[6])
    defparam i15433_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1518_3_lut (.I0(n2227), 
            .I1(n2294), .I2(n2247), .I3(GND_net), .O(n2326));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1518_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15873_3_lut (.I0(current_limit[3]), .I1(\data_in_frame[21] [3]), 
            .I2(n50654), .I3(GND_net), .O(n29953));   // verilog/coms.v(128[12] 303[6])
    defparam i15873_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15840_3_lut (.I0(PWMLimit[21]), .I1(\data_in_frame[8] [5]), 
            .I2(n50654), .I3(GND_net), .O(n29920));   // verilog/coms.v(128[12] 303[6])
    defparam i15840_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15874_3_lut (.I0(current_limit[2]), .I1(\data_in_frame[21] [2]), 
            .I2(n50654), .I3(GND_net), .O(n29954));   // verilog/coms.v(128[12] 303[6])
    defparam i15874_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15841_3_lut (.I0(PWMLimit[20]), .I1(\data_in_frame[8] [4]), 
            .I2(n50654), .I3(GND_net), .O(n29921));   // verilog/coms.v(128[12] 303[6])
    defparam i15841_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15275_3_lut (.I0(deadband[0]), .I1(\data_in_frame[16] [0]), 
            .I2(n50654), .I3(GND_net), .O(n29355));   // verilog/coms.v(128[12] 303[6])
    defparam i15275_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15875_3_lut (.I0(current_limit[1]), .I1(\data_in_frame[21] [1]), 
            .I2(n50654), .I3(GND_net), .O(n29955));   // verilog/coms.v(128[12] 303[6])
    defparam i15875_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15876_3_lut (.I0(control_mode[7]), .I1(\data_in_frame[1] [7]), 
            .I2(n50654), .I3(GND_net), .O(n29956));   // verilog/coms.v(128[12] 303[6])
    defparam i15876_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i22676_2_lut (.I0(duty[4]), .I1(n296), .I2(GND_net), .I3(GND_net), 
            .O(n4925));   // verilog/TinyFPGA_B.v(123[17] 125[11])
    defparam i22676_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i15276_3_lut (.I0(\data_out_frame[11] [5]), .I1(encoder1_position_scaled[5]), 
            .I2(n24210), .I3(GND_net), .O(n29356));   // verilog/coms.v(128[12] 303[6])
    defparam i15276_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15877_3_lut (.I0(control_mode[6]), .I1(\data_in_frame[1] [6]), 
            .I2(n50654), .I3(GND_net), .O(n29957));   // verilog/coms.v(128[12] 303[6])
    defparam i15877_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i40599_1_lut (.I0(n1257), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n56430));
    defparam i40599_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i15878_3_lut (.I0(control_mode[5]), .I1(\data_in_frame[1] [5]), 
            .I2(n50654), .I3(GND_net), .O(n29958));   // verilog/coms.v(128[12] 303[6])
    defparam i15878_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15879_3_lut (.I0(control_mode[4]), .I1(\data_in_frame[1] [4]), 
            .I2(n50654), .I3(GND_net), .O(n29959));   // verilog/coms.v(128[12] 303[6])
    defparam i15879_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15880_3_lut (.I0(control_mode[3]), .I1(\data_in_frame[1] [3]), 
            .I2(n50654), .I3(GND_net), .O(n29960));   // verilog/coms.v(128[12] 303[6])
    defparam i15880_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1757 (.I0(n2323), .I1(n2327), .I2(n2326), .I3(n2325), 
            .O(n51732));
    defparam i1_4_lut_adj_1757.LUT_INIT = 16'hfffe;
    SB_LUT4 i15881_3_lut (.I0(control_mode[2]), .I1(\data_in_frame[1] [2]), 
            .I2(n50654), .I3(GND_net), .O(n29961));   // verilog/coms.v(128[12] 303[6])
    defparam i15881_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_3_lut_adj_1758 (.I0(n51732), .I1(n2328), .I2(n2324), .I3(GND_net), 
            .O(n51734));
    defparam i1_3_lut_adj_1758.LUT_INIT = 16'hfefe;
    SB_LUT4 i23298_4_lut (.I0(n534), .I1(n2331), .I2(n2332), .I3(n2333), 
            .O(n37388));
    defparam i23298_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 i15882_3_lut (.I0(control_mode[1]), .I1(\data_in_frame[1] [1]), 
            .I2(n50654), .I3(GND_net), .O(n29962));   // verilog/coms.v(128[12] 303[6])
    defparam i15882_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1759 (.I0(n2320), .I1(n2321), .I2(n51734), .I3(n2322), 
            .O(n51740));
    defparam i1_4_lut_adj_1759.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_unary_minus_2_inv_0_i2_1_lut (.I0(encoder0_position_scaled_23__N_327[1]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n32_adj_5641));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_unary_minus_2_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i40449_1_lut (.I0(n2049), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n56280));
    defparam i40449_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i15887_3_lut (.I0(\data_out_frame[23] [2]), .I1(neopxl_color[18]), 
            .I2(n24210), .I3(GND_net), .O(n29967));   // verilog/coms.v(128[12] 303[6])
    defparam i15887_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15888_3_lut (.I0(\data_out_frame[23] [1]), .I1(neopxl_color[17]), 
            .I2(n24210), .I3(GND_net), .O(n29968));   // verilog/coms.v(128[12] 303[6])
    defparam i15888_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_1760 (.I0(n2329), .I1(n2330), .I2(GND_net), .I3(GND_net), 
            .O(n52060));
    defparam i1_2_lut_adj_1760.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut_adj_1761 (.I0(n2319), .I1(n52060), .I2(n51740), .I3(n37388), 
            .O(n51744));
    defparam i1_4_lut_adj_1761.LUT_INIT = 16'hfefa;
    SB_LUT4 i1_4_lut_adj_1762 (.I0(n2316), .I1(n2317), .I2(n2318), .I3(n51744), 
            .O(n51750));
    defparam i1_4_lut_adj_1762.LUT_INIT = 16'hfffe;
    SB_LUT4 i40374_4_lut (.I0(n2314), .I1(n2313), .I2(n2315), .I3(n51750), 
            .O(n2346));
    defparam i40374_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1517_rep_19_3_lut (.I0(n2293), 
            .I1(n2392), .I2(n2346), .I3(GND_net), .O(n53086));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1517_rep_19_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i39145_2_lut (.I0(n2346), .I1(n2247), .I2(GND_net), .I3(GND_net), 
            .O(n54975));
    defparam i39145_2_lut.LUT_INIT = 16'h7777;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1584_rep_17_3_lut (.I0(n53086), 
            .I1(n2491), .I2(n2445), .I3(GND_net), .O(n53084));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1584_rep_17_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i39761_4_lut (.I0(n53084), .I1(n2226), .I2(n2445), .I3(n54975), 
            .O(n55592));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam i39761_4_lut.LUT_INIT = 16'haaca;
    SB_LUT4 i15889_3_lut (.I0(\data_out_frame[23] [0]), .I1(neopxl_color[16]), 
            .I2(n24210), .I3(GND_net), .O(n29969));   // verilog/coms.v(128[12] 303[6])
    defparam i15889_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15890_3_lut (.I0(\data_out_frame[22] [7]), .I1(current[7]), 
            .I2(n24210), .I3(GND_net), .O(n29970));   // verilog/coms.v(128[12] 303[6])
    defparam i15890_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i39762_3_lut (.I0(n55592), .I1(n2590), .I2(n2544), .I3(GND_net), 
            .O(n2622));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam i39762_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15891_3_lut (.I0(\data_out_frame[22] [6]), .I1(current[6]), 
            .I2(n24210), .I3(GND_net), .O(n29971));   // verilog/coms.v(128[12] 303[6])
    defparam i15891_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15892_3_lut (.I0(\data_out_frame[22] [5]), .I1(current[5]), 
            .I2(n24210), .I3(GND_net), .O(n29972));   // verilog/coms.v(128[12] 303[6])
    defparam i15892_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15893_3_lut (.I0(\data_out_frame[22] [4]), .I1(current[4]), 
            .I2(n24210), .I3(GND_net), .O(n29973));   // verilog/coms.v(128[12] 303[6])
    defparam i15893_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15894_3_lut (.I0(\data_out_frame[22] [3]), .I1(current[3]), 
            .I2(n24210), .I3(GND_net), .O(n29974));   // verilog/coms.v(128[12] 303[6])
    defparam i15894_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1717_3_lut (.I0(n2522), 
            .I1(n2589), .I2(n2544), .I3(GND_net), .O(n2621));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1717_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_adj_1763 (.I0(n2621), .I1(n2622), .I2(GND_net), .I3(GND_net), 
            .O(n52112));
    defparam i1_2_lut_adj_1763.LUT_INIT = 16'heeee;
    SB_LUT4 i1_3_lut_adj_1764 (.I0(n2624), .I1(n2628), .I2(n2626), .I3(GND_net), 
            .O(n52114));
    defparam i1_3_lut_adj_1764.LUT_INIT = 16'hfefe;
    SB_LUT4 i23292_4_lut (.I0(n537), .I1(n2631), .I2(n2632), .I3(n2633), 
            .O(n37382));
    defparam i23292_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 i1_4_lut_adj_1765 (.I0(n2619), .I1(n2625), .I2(n2627), .I3(n2623), 
            .O(n52220));
    defparam i1_4_lut_adj_1765.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1766 (.I0(n2629), .I1(n52220), .I2(n37382), .I3(n2630), 
            .O(n52222));
    defparam i1_4_lut_adj_1766.LUT_INIT = 16'heccc;
    SB_LUT4 unary_minus_18_inv_0_i1_1_lut (.I0(duty[0]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n25));   // verilog/TinyFPGA_B.v(119[24:29])
    defparam unary_minus_18_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i15434_3_lut (.I0(Kp[7]), .I1(\data_in_frame[3] [7]), .I2(n50654), 
            .I3(GND_net), .O(n29514));   // verilog/coms.v(128[12] 303[6])
    defparam i15434_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1767 (.I0(n2618), .I1(n2620), .I2(n52114), .I3(n52112), 
            .O(n52120));
    defparam i1_4_lut_adj_1767.LUT_INIT = 16'hfffe;
    SB_LUT4 i15435_3_lut (.I0(Kp[6]), .I1(\data_in_frame[3] [6]), .I2(n50654), 
            .I3(GND_net), .O(n29515));   // verilog/coms.v(128[12] 303[6])
    defparam i15435_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 unary_minus_19_inv_0_i1_1_lut (.I0(current[0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_5464));   // verilog/TinyFPGA_B.v(121[16:24])
    defparam unary_minus_19_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i15895_3_lut (.I0(\data_out_frame[22] [2]), .I1(current[2]), 
            .I2(n24210), .I3(GND_net), .O(n29975));   // verilog/coms.v(128[12] 303[6])
    defparam i15895_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1768 (.I0(n2616), .I1(n2615), .I2(n2617), .I3(n52222), 
            .O(n51396));
    defparam i1_4_lut_adj_1768.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1769 (.I0(n2613), .I1(n2614), .I2(n51396), .I3(n52120), 
            .O(n52126));
    defparam i1_4_lut_adj_1769.LUT_INIT = 16'hfffe;
    SB_LUT4 i40287_4_lut (.I0(n2611), .I1(n2610), .I2(n2612), .I3(n52126), 
            .O(n2643));
    defparam i40287_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1711_3_lut (.I0(n2516), 
            .I1(n2583), .I2(n2544), .I3(GND_net), .O(n2615));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1711_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1778_3_lut (.I0(n2615), 
            .I1(n2682), .I2(n2643), .I3(GND_net), .O(n2714));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1778_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15439_3_lut (.I0(Kp[3]), .I1(\data_in_frame[3] [3]), .I2(n50654), 
            .I3(GND_net), .O(n29519));   // verilog/coms.v(128[12] 303[6])
    defparam i15439_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15440_3_lut (.I0(Kp[2]), .I1(\data_in_frame[3] [2]), .I2(n50654), 
            .I3(GND_net), .O(n29520));   // verilog/coms.v(128[12] 303[6])
    defparam i15440_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15441_3_lut (.I0(Kp[1]), .I1(\data_in_frame[3] [1]), .I2(n50654), 
            .I3(GND_net), .O(n29521));   // verilog/coms.v(128[12] 303[6])
    defparam i15441_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i40667_1_lut (.I0(n3237), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n56498));
    defparam i40667_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_4_lut_adj_1770 (.I0(commutation_state[2]), .I1(commutation_state[1]), 
            .I2(commutation_state_prev[2]), .I3(commutation_state_prev[1]), 
            .O(n4_adj_5607));   // verilog/TinyFPGA_B.v(146[7:48])
    defparam i1_4_lut_adj_1770.LUT_INIT = 16'h7bde;
    SB_LUT4 i1_4_lut_adj_1771 (.I0(enable_slow_N_4393), .I1(data_ready), 
            .I2(state_adj_5705[1]), .I3(state_adj_5705[0]), .O(n48670));   // verilog/eeprom.v(26[8] 58[4])
    defparam i1_4_lut_adj_1771.LUT_INIT = 16'hccd0;
    SB_LUT4 i15313_4_lut (.I0(rw), .I1(state_adj_5705[0]), .I2(state_adj_5705[1]), 
            .I3(n6272), .O(n29393));   // verilog/eeprom.v(26[8] 58[4])
    defparam i15313_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i2_2_lut (.I0(dti_counter[1]), .I1(dti_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n10_adj_5591));   // verilog/TinyFPGA_B.v(171[9:23])
    defparam i2_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i6_4_lut (.I0(dti_counter[7]), .I1(dti_counter[4]), .I2(dti_counter[5]), 
            .I3(dti_counter[6]), .O(n14_adj_5522));   // verilog/TinyFPGA_B.v(171[9:23])
    defparam i6_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_4_lut (.I0(dti_counter[0]), .I1(n14_adj_5522), .I2(n10_adj_5591), 
            .I3(dti_counter[3]), .O(n24553));   // verilog/TinyFPGA_B.v(171[9:23])
    defparam i7_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i40655_2_lut (.I0(n24553), .I1(dti), .I2(GND_net), .I3(GND_net), 
            .O(dti_N_527));
    defparam i40655_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i912_3_lut (.I0(n1333), .I1(n1400), 
            .I2(n1356), .I3(GND_net), .O(n1432));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i912_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15442_3_lut (.I0(deadband[23]), .I1(\data_in_frame[14] [7]), 
            .I2(n50654), .I3(GND_net), .O(n29522));   // verilog/coms.v(128[12] 303[6])
    defparam i15442_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_263_13 (.CI(n43545), .I0(encoder1_position[14]), .I1(GND_net), 
            .CO(n43546));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1771_19_lut (.I0(GND_net), 
            .I1(n2617), .I2(VCC_net), .I3(n44244), .O(n2684)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1771_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1771_19 (.CI(n44244), 
            .I0(n2617), .I1(VCC_net), .CO(n44245));
    SB_LUT4 add_261_13_lut (.I0(current[11]), .I1(duty[14]), .I2(n56614), 
            .I3(n43568), .O(n259)) /* synthesis syn_instantiated=1 */ ;
    defparam add_261_13_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1771_18_lut (.I0(GND_net), 
            .I1(n2618), .I2(VCC_net), .I3(n44243), .O(n2685)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1771_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_900_4_lut (.I0(GND_net), 
            .I1(n1332), .I2(GND_net), .I3(n44008), .O(n1399)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_900_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1771_18 (.CI(n44243), 
            .I0(n2618), .I1(VCC_net), .CO(n44244));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1771_17_lut (.I0(GND_net), 
            .I1(n2619), .I2(VCC_net), .I3(n44242), .O(n2686)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1771_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_900_4 (.CI(n44008), 
            .I0(n1332), .I1(GND_net), .CO(n44009));
    SB_LUT4 add_175_25_lut (.I0(GND_net), .I1(delay_counter[23]), .I2(GND_net), 
            .I3(n43632), .O(n1540)) /* synthesis syn_instantiated=1 */ ;
    defparam add_175_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1771_17 (.CI(n44242), 
            .I0(n2619), .I1(VCC_net), .CO(n44243));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_900_3_lut (.I0(GND_net), 
            .I1(n1333), .I2(VCC_net), .I3(n44007), .O(n1400)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_900_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_900_3 (.CI(n44007), 
            .I0(n1333), .I1(VCC_net), .CO(n44008));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_900_2_lut (.I0(GND_net), 
            .I1(n413), .I2(GND_net), .I3(VCC_net), .O(n1401)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_900_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_900_2 (.CI(VCC_net), 
            .I0(n413), .I1(GND_net), .CO(n44007));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_833_12_lut (.I0(n56430), 
            .I1(n1224), .I2(VCC_net), .I3(n44006), .O(n1323)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_833_12_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_833_11_lut (.I0(GND_net), 
            .I1(n1225), .I2(VCC_net), .I3(n44005), .O(n1292)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_833_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_833_11 (.CI(n44005), 
            .I0(n1225), .I1(VCC_net), .CO(n44006));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_833_10_lut (.I0(GND_net), 
            .I1(n1226), .I2(VCC_net), .I3(n44004), .O(n1293)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_833_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_833_10 (.CI(n44004), 
            .I0(n1226), .I1(VCC_net), .CO(n44005));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_833_9_lut (.I0(GND_net), 
            .I1(n1227), .I2(VCC_net), .I3(n44003), .O(n1294)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_833_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1039_7 (.CI(n43776), .I0(n4899), .I1(n4924), .CO(n43777));
    SB_LUT4 add_1039_6_lut (.I0(GND_net), .I1(n4900), .I2(n4925), .I3(n43775), 
            .O(n437)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1039_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1771_16_lut (.I0(GND_net), 
            .I1(n2620), .I2(VCC_net), .I3(n44241), .O(n2687)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1771_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_833_9 (.CI(n44003), 
            .I0(n1227), .I1(VCC_net), .CO(n44004));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1040_3_lut (.I0(n1525), 
            .I1(n1592), .I2(n1554_adj_5597), .I3(GND_net), .O(n1624));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1040_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_mux_3_i1_3_lut (.I0(encoder0_position[0]), 
            .I1(n33), .I2(encoder0_position_scaled_23__N_327[31]), .I3(GND_net), 
            .O(n544));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_mux_3_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_833_8_lut (.I0(GND_net), 
            .I1(n1228), .I2(VCC_net), .I3(n44002), .O(n1295)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_833_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1039_6 (.CI(n43775), .I0(n4900), .I1(n4925), .CO(n43776));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1771_16 (.CI(n44241), 
            .I0(n2620), .I1(VCC_net), .CO(n44242));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_833_8 (.CI(n44002), 
            .I0(n1228), .I1(VCC_net), .CO(n44003));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_833_7_lut (.I0(GND_net), 
            .I1(n1229), .I2(GND_net), .I3(n44001), .O(n1296)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_833_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1771_15_lut (.I0(GND_net), 
            .I1(n2621), .I2(VCC_net), .I3(n44240), .O(n2688)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1771_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_833_7 (.CI(n44001), 
            .I0(n1229), .I1(GND_net), .CO(n44002));
    SB_CARRY add_175_25 (.CI(n43632), .I0(delay_counter[23]), .I1(GND_net), 
            .CO(n43633));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_833_6_lut (.I0(GND_net), 
            .I1(n1230), .I2(GND_net), .I3(n44000), .O(n1297)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_833_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_833_6 (.CI(n44000), 
            .I0(n1230), .I1(GND_net), .CO(n44001));
    SB_LUT4 add_175_24_lut (.I0(GND_net), .I1(delay_counter[22]), .I2(GND_net), 
            .I3(n43631), .O(n1541)) /* synthesis syn_instantiated=1 */ ;
    defparam add_175_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1771_15 (.CI(n44240), 
            .I0(n2621), .I1(VCC_net), .CO(n44241));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1771_14_lut (.I0(GND_net), 
            .I1(n2622), .I2(VCC_net), .I3(n44239), .O(n2689)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1771_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i40659_1_lut (.I0(n37482), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n56490));
    defparam i40659_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_1039_5_lut (.I0(GND_net), .I1(n4901), .I2(n4926), .I3(n43774), 
            .O(n438)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1039_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_833_5_lut (.I0(GND_net), 
            .I1(n1231), .I2(VCC_net), .I3(n43999), .O(n1298)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_833_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_833_5 (.CI(n43999), 
            .I0(n1231), .I1(VCC_net), .CO(n44000));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i2193_3_lut (.I0(n3222), 
            .I1(n3289), .I2(n3237), .I3(GND_net), .O(n27_adj_5652));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i2193_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_261_13 (.CI(n43568), .I0(duty[14]), .I1(n56614), .CO(n43569));
    SB_LUT4 i15314_3_lut (.I0(\data_out_frame[10] [0]), .I1(encoder1_position_scaled[8]), 
            .I2(n24210), .I3(GND_net), .O(n29394));   // verilog/coms.v(128[12] 303[6])
    defparam i15314_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_833_4_lut (.I0(GND_net), 
            .I1(n1232), .I2(GND_net), .I3(n43998), .O(n1299)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_833_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1771_14 (.CI(n44239), 
            .I0(n2622), .I1(VCC_net), .CO(n44240));
    SB_LUT4 i15315_3_lut (.I0(\data_out_frame[9] [7]), .I1(encoder1_position_scaled[23]), 
            .I2(n24210), .I3(GND_net), .O(n29395));   // verilog/coms.v(128[12] 303[6])
    defparam i15315_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_833_4 (.CI(n43998), 
            .I0(n1232), .I1(GND_net), .CO(n43999));
    SB_CARRY add_1039_5 (.CI(n43774), .I0(n4901), .I1(n4926), .CO(n43775));
    SB_CARRY add_175_24 (.CI(n43631), .I0(delay_counter[22]), .I1(GND_net), 
            .CO(n43632));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1771_13_lut (.I0(GND_net), 
            .I1(n2623), .I2(VCC_net), .I3(n44238), .O(n2690)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1771_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15316_3_lut (.I0(\data_out_frame[9] [6]), .I1(encoder1_position_scaled[22]), 
            .I2(n24210), .I3(GND_net), .O(n29396));   // verilog/coms.v(128[12] 303[6])
    defparam i15316_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_175_23_lut (.I0(GND_net), .I1(delay_counter[21]), .I2(GND_net), 
            .I3(n43630), .O(n1542)) /* synthesis syn_instantiated=1 */ ;
    defparam add_175_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_833_3_lut (.I0(GND_net), 
            .I1(n1233), .I2(VCC_net), .I3(n43997), .O(n1300)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_833_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1771_13 (.CI(n44238), 
            .I0(n2623), .I1(VCC_net), .CO(n44239));
    SB_LUT4 add_1039_4_lut (.I0(GND_net), .I1(n4902), .I2(n4927), .I3(n43773), 
            .O(n439)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1039_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_833_3 (.CI(n43997), 
            .I0(n1233), .I1(VCC_net), .CO(n43998));
    SB_CARRY add_175_23 (.CI(n43630), .I0(delay_counter[21]), .I1(GND_net), 
            .CO(n43631));
    SB_LUT4 add_175_22_lut (.I0(GND_net), .I1(delay_counter[20]), .I2(GND_net), 
            .I3(n43629), .O(n1543)) /* synthesis syn_instantiated=1 */ ;
    defparam add_175_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_261_12_lut (.I0(current[10]), .I1(duty[13]), .I2(n56614), 
            .I3(n43567), .O(n260)) /* synthesis syn_instantiated=1 */ ;
    defparam add_261_12_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY add_1039_4 (.CI(n43773), .I0(n4902), .I1(n4927), .CO(n43774));
    SB_LUT4 i15317_3_lut (.I0(\data_out_frame[9] [5]), .I1(encoder1_position_scaled[21]), 
            .I2(n24210), .I3(GND_net), .O(n29397));   // verilog/coms.v(128[12] 303[6])
    defparam i15317_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_833_2_lut (.I0(GND_net), 
            .I1(n412), .I2(GND_net), .I3(VCC_net), .O(n1301)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_833_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_833_2 (.CI(VCC_net), 
            .I0(n412), .I1(GND_net), .CO(n43997));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i2198_3_lut (.I0(n3227), 
            .I1(n3294), .I2(n3237), .I3(GND_net), .O(n17_adj_5649));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i2198_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_766_11_lut (.I0(n56444), 
            .I1(n1125), .I2(VCC_net), .I3(n43996), .O(n1224)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_766_11_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i15318_3_lut (.I0(CS_c), .I1(state_adj_5713[0]), .I2(state_adj_5713[1]), 
            .I3(GND_net), .O(n29398));   // verilog/tli4970.v(35[10] 68[6])
    defparam i15318_3_lut.LUT_INIT = 16'ha3a3;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_766_10_lut (.I0(GND_net), 
            .I1(n1126), .I2(VCC_net), .I3(n43995), .O(n1193)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_766_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_261_12 (.CI(n43567), .I0(duty[13]), .I1(n56614), .CO(n43568));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1771_12_lut (.I0(GND_net), 
            .I1(n2624), .I2(VCC_net), .I3(n44237), .O(n2691)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1771_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_766_10 (.CI(n43995), 
            .I0(n1126), .I1(VCC_net), .CO(n43996));
    SB_LUT4 add_1039_3_lut (.I0(GND_net), .I1(n4903), .I2(n4928), .I3(n43772), 
            .O(n440)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1039_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1771_12 (.CI(n44237), 
            .I0(n2624), .I1(VCC_net), .CO(n44238));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1771_11_lut (.I0(GND_net), 
            .I1(n2625), .I2(VCC_net), .I3(n44236), .O(n2692)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1771_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_766_9_lut (.I0(GND_net), 
            .I1(n1127), .I2(VCC_net), .I3(n43994), .O(n1194)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_766_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_261_11_lut (.I0(current[9]), .I1(duty[12]), .I2(n56614), 
            .I3(n43566), .O(n261)) /* synthesis syn_instantiated=1 */ ;
    defparam add_261_11_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_unary_minus_2_inv_0_i3_1_lut (.I0(encoder0_position_scaled_23__N_327[2]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n31_adj_5640));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_unary_minus_2_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_175_22 (.CI(n43629), .I0(delay_counter[20]), .I1(GND_net), 
            .CO(n43630));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i2196_3_lut (.I0(n3225), 
            .I1(n3292), .I2(n3237), .I3(GND_net), .O(n21_adj_5651));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i2196_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_261_16_lut (.I0(current[15]), .I1(duty[17]), .I2(n56614), 
            .I3(n43571), .O(n256)) /* synthesis syn_instantiated=1 */ ;
    defparam add_261_16_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 unary_minus_19_inv_0_i2_1_lut (.I0(current[1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n24_adj_5463));   // verilog/TinyFPGA_B.v(121[16:24])
    defparam unary_minus_19_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i23102_4_lut (.I0(n544), .I1(n543), .I2(n3301), .I3(n3237), 
            .O(n37186));
    defparam i23102_4_lut.LUT_INIT = 16'heefa;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i2191_3_lut (.I0(n3220), 
            .I1(n3287), .I2(n3237), .I3(GND_net), .O(n31_adj_5653));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i2191_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i40776_4_lut (.I0(n15_adj_5470), .I1(clk_out), .I2(state_adj_5713[0]), 
            .I3(state_adj_5713[1]), .O(n9_adj_5601));   // verilog/tli4970.v(35[10] 68[6])
    defparam i40776_4_lut.LUT_INIT = 16'hc8fc;
    SB_LUT4 i15320_3_lut (.I0(\data_out_frame[9] [4]), .I1(encoder1_position_scaled[20]), 
            .I2(n24210), .I3(GND_net), .O(n29400));   // verilog/coms.v(128[12] 303[6])
    defparam i15320_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15321_3_lut (.I0(\data_out_frame[9] [3]), .I1(encoder1_position_scaled[19]), 
            .I2(n24210), .I3(GND_net), .O(n29401));   // verilog/coms.v(128[12] 303[6])
    defparam i15321_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1771_11 (.CI(n44236), 
            .I0(n2625), .I1(VCC_net), .CO(n44237));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_unary_minus_2_inv_0_i4_1_lut (.I0(encoder0_position_scaled_23__N_327[3]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n30_adj_5639));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_unary_minus_2_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1771_10_lut (.I0(GND_net), 
            .I1(n2626), .I2(VCC_net), .I3(n44235), .O(n2693)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1771_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i2197_3_lut (.I0(n3226), 
            .I1(n3293), .I2(n3237), .I3(GND_net), .O(n19_adj_5650));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i2197_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_766_9 (.CI(n43994), 
            .I0(n1127), .I1(VCC_net), .CO(n43995));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_766_8_lut (.I0(GND_net), 
            .I1(n1128), .I2(VCC_net), .I3(n43993), .O(n1195)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_766_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1771_10 (.CI(n44235), 
            .I0(n2626), .I1(VCC_net), .CO(n44236));
    SB_LUT4 i15322_3_lut (.I0(\data_out_frame[9] [2]), .I1(encoder1_position_scaled[18]), 
            .I2(n24210), .I3(GND_net), .O(n29402));   // verilog/coms.v(128[12] 303[6])
    defparam i15322_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1771_9_lut (.I0(GND_net), 
            .I1(n2627), .I2(VCC_net), .I3(n44234), .O(n2694)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1771_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15323_3_lut (.I0(\data_out_frame[9] [1]), .I1(encoder1_position_scaled[17]), 
            .I2(n24210), .I3(GND_net), .O(n29403));   // verilog/coms.v(128[12] 303[6])
    defparam i15323_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_766_8 (.CI(n43993), 
            .I0(n1128), .I1(VCC_net), .CO(n43994));
    SB_CARRY add_1039_3 (.CI(n43772), .I0(n4903), .I1(n4928), .CO(n43773));
    SB_LUT4 i1_4_lut_adj_1772 (.I0(n3219), .I1(n27_adj_5652), .I2(n3286), 
            .I3(n3237), .O(n51638));
    defparam i1_4_lut_adj_1772.LUT_INIT = 16'heefc;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1771_9 (.CI(n44234), 
            .I0(n2627), .I1(VCC_net), .CO(n44235));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_766_7_lut (.I0(GND_net), 
            .I1(n1129), .I2(GND_net), .I3(n43992), .O(n1196)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_766_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15324_3_lut (.I0(\data_out_frame[9] [0]), .I1(encoder1_position_scaled[16]), 
            .I2(n24210), .I3(GND_net), .O(n29404));   // verilog/coms.v(128[12] 303[6])
    defparam i15324_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_1039_2_lut (.I0(GND_net), .I1(n4904), .I2(n4929), .I3(GND_net), 
            .O(n441)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1039_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1771_8_lut (.I0(GND_net), 
            .I1(n2628), .I2(VCC_net), .I3(n44233), .O(n2695)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1771_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i2199_3_lut (.I0(n3228), 
            .I1(n3295), .I2(n3237), .I3(GND_net), .O(n15_adj_5648));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i2199_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15325_3_lut (.I0(\data_out_frame[8] [7]), .I1(encoder0_position_scaled[7]), 
            .I2(n24210), .I3(GND_net), .O(n29405));   // verilog/coms.v(128[12] 303[6])
    defparam i15325_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_766_7 (.CI(n43992), 
            .I0(n1129), .I1(GND_net), .CO(n43993));
    SB_LUT4 add_175_21_lut (.I0(GND_net), .I1(delay_counter[19]), .I2(GND_net), 
            .I3(n43628), .O(n1544)) /* synthesis syn_instantiated=1 */ ;
    defparam add_175_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1773 (.I0(n3223), .I1(n31_adj_5653), .I2(n3290), 
            .I3(n3237), .O(n51646));
    defparam i1_4_lut_adj_1773.LUT_INIT = 16'heefc;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1771_8 (.CI(n44233), 
            .I0(n2628), .I1(VCC_net), .CO(n44234));
    SB_LUT4 i15326_3_lut (.I0(\data_out_frame[8] [6]), .I1(encoder0_position_scaled[6]), 
            .I2(n24210), .I3(GND_net), .O(n29406));   // verilog/coms.v(128[12] 303[6])
    defparam i15326_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12_4_lut (.I0(\ID_READOUT_FSM.state [1]), .I1(n7974), .I2(n28885), 
            .I3(\ID_READOUT_FSM.state [0]), .O(n48068));   // verilog/TinyFPGA_B.v(368[10] 396[6])
    defparam i12_4_lut.LUT_INIT = 16'h3a0a;
    SB_LUT4 i15327_4_lut (.I0(CS_MISO_c), .I1(data_adj_5711[15]), .I2(n36528), 
            .I3(n27264), .O(n29407));   // verilog/tli4970.v(35[10] 68[6])
    defparam i15327_4_lut.LUT_INIT = 16'hccac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1771_7_lut (.I0(GND_net), 
            .I1(n2629), .I2(GND_net), .I3(n44232), .O(n2696)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1771_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_766_6_lut (.I0(GND_net), 
            .I1(n1130), .I2(GND_net), .I3(n43991), .O(n1197)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_766_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_766_6 (.CI(n43991), 
            .I0(n1130), .I1(GND_net), .CO(n43992));
    SB_LUT4 i15328_3_lut (.I0(\data_out_frame[8] [5]), .I1(encoder0_position_scaled[5]), 
            .I2(n24210), .I3(GND_net), .O(n29408));   // verilog/coms.v(128[12] 303[6])
    defparam i15328_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_1039_2 (.CI(GND_net), .I0(n4904), .I1(n4929), .CO(n43772));
    SB_LUT4 i1_4_lut_adj_1774 (.I0(n3224), .I1(n19_adj_5650), .I2(n3291), 
            .I3(n3237), .O(n51642));
    defparam i1_4_lut_adj_1774.LUT_INIT = 16'heefc;
    SB_LUT4 i15330_3_lut (.I0(\data_out_frame[8] [4]), .I1(encoder0_position_scaled[4]), 
            .I2(n24210), .I3(GND_net), .O(n29410));   // verilog/coms.v(128[12] 303[6])
    defparam i15330_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_18_inv_0_i3_1_lut (.I0(duty[2]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n23));   // verilog/TinyFPGA_B.v(119[24:29])
    defparam unary_minus_18_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_766_5_lut (.I0(GND_net), 
            .I1(n1131), .I2(VCC_net), .I3(n43990), .O(n1198)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_766_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_766_5 (.CI(n43990), 
            .I0(n1131), .I1(VCC_net), .CO(n43991));
    SB_LUT4 i15443_3_lut (.I0(deadband[22]), .I1(\data_in_frame[14] [6]), 
            .I2(n50654), .I3(GND_net), .O(n29523));   // verilog/coms.v(128[12] 303[6])
    defparam i15443_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1775 (.I0(n3221), .I1(n17_adj_5649), .I2(n3288), 
            .I3(n3237), .O(n51644));
    defparam i1_4_lut_adj_1775.LUT_INIT = 16'heefc;
    SB_LUT4 i15331_3_lut (.I0(\data_out_frame[8] [3]), .I1(encoder0_position_scaled[3]), 
            .I2(n24210), .I3(GND_net), .O(n29411));   // verilog/coms.v(128[12] 303[6])
    defparam i15331_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1771_7 (.CI(n44232), 
            .I0(n2629), .I1(GND_net), .CO(n44233));
    SB_LUT4 i15332_3_lut (.I0(\data_out_frame[8] [2]), .I1(encoder0_position_scaled[2]), 
            .I2(n24210), .I3(GND_net), .O(n29412));   // verilog/coms.v(128[12] 303[6])
    defparam i15332_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1771_6_lut (.I0(GND_net), 
            .I1(n2630), .I2(GND_net), .I3(n44231), .O(n2697)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1771_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1776 (.I0(n3229), .I1(n21_adj_5651), .I2(n3296), 
            .I3(n3237), .O(n51640));
    defparam i1_4_lut_adj_1776.LUT_INIT = 16'heefc;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1771_6 (.CI(n44231), 
            .I0(n2630), .I1(GND_net), .CO(n44232));
    SB_LUT4 i1_4_lut_adj_1777 (.I0(n51642), .I1(n51646), .I2(n15_adj_5648), 
            .I3(n51638), .O(n51654));
    defparam i1_4_lut_adj_1777.LUT_INIT = 16'hfffe;
    SB_LUT4 i15333_4_lut (.I0(tx_active), .I1(r_SM_Main_adj_5723[1]), .I2(n19728), 
            .I3(n4_adj_5644), .O(n29413));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i15333_4_lut.LUT_INIT = 16'h32aa;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_766_4_lut (.I0(GND_net), 
            .I1(n1132), .I2(GND_net), .I3(n43989), .O(n1199)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_766_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_unary_minus_2_inv_0_i5_1_lut (.I0(encoder0_position_scaled_23__N_327[4]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n29_adj_5638));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_unary_minus_2_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1771_5_lut (.I0(GND_net), 
            .I1(n2631), .I2(VCC_net), .I3(n44230), .O(n2698)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1771_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1771_5 (.CI(n44230), 
            .I0(n2631), .I1(VCC_net), .CO(n44231));
    SB_CARRY add_175_21 (.CI(n43628), .I0(delay_counter[19]), .I1(GND_net), 
            .CO(n43629));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i843_3_lut (.I0(n1232), .I1(n1299), 
            .I2(n1257), .I3(GND_net), .O(n1331));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i843_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i2189_3_lut (.I0(n3218), 
            .I1(n3285), .I2(n3237), .I3(GND_net), .O(n35));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i2189_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1778 (.I0(n35), .I1(n51654), .I2(n51640), .I3(n51644), 
            .O(n51658));
    defparam i1_4_lut_adj_1778.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i842_3_lut (.I0(n1231), .I1(n1298), 
            .I2(n1257), .I3(GND_net), .O(n1330));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i842_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_766_4 (.CI(n43989), 
            .I0(n1132), .I1(GND_net), .CO(n43990));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i841_3_lut (.I0(n1230), .I1(n1297), 
            .I2(n1257), .I3(GND_net), .O(n1329));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i841_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15334_3_lut (.I0(\data_out_frame[8] [1]), .I1(encoder0_position_scaled[1]), 
            .I2(n24210), .I3(GND_net), .O(n29414));   // verilog/coms.v(128[12] 303[6])
    defparam i15334_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1779 (.I0(n3217), .I1(n51658), .I2(n3284), .I3(n3237), 
            .O(n51660));
    defparam i1_4_lut_adj_1779.LUT_INIT = 16'heefc;
    SB_LUT4 i15335_3_lut (.I0(\data_out_frame[8] [0]), .I1(encoder0_position_scaled[0]), 
            .I2(n24210), .I3(GND_net), .O(n29415));   // verilog/coms.v(128[12] 303[6])
    defparam i15335_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15336_3_lut (.I0(\data_out_frame[7] [7]), .I1(encoder0_position_scaled[15]), 
            .I2(n24210), .I3(GND_net), .O(n29416));   // verilog/coms.v(128[12] 303[6])
    defparam i15336_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1771_4_lut (.I0(GND_net), 
            .I1(n2632), .I2(GND_net), .I3(n44229), .O(n2699)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1771_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i2203_3_lut (.I0(n3232), 
            .I1(n3299), .I2(n3237), .I3(GND_net), .O(n7_adj_5647));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i2203_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16_4_lut (.I0(n3231), .I1(n54589), .I2(n3237), .I3(n3230), 
            .O(n5_adj_5606));
    defparam i16_4_lut.LUT_INIT = 16'hac0c;
    SB_GB_IO CLK_pad (.PACKAGE_PIN(CLK), .OUTPUT_ENABLE(VCC_net), .GLOBAL_BUFFER_OUTPUT(clk16MHz));   // verilog/TinyFPGA_B.v(3[9:12])
    defparam CLK_pad.PIN_TYPE = 6'b000001;
    defparam CLK_pad.PULLUP = 1'b0;
    defparam CLK_pad.NEG_TRIGGER = 1'b0;
    defparam CLK_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 i1_4_lut_adj_1780 (.I0(n3216), .I1(n51660), .I2(n3283), .I3(n3237), 
            .O(n51662));
    defparam i1_4_lut_adj_1780.LUT_INIT = 16'heefc;
    SB_LUT4 i23207_4_lut (.I0(n37186), .I1(n3233), .I2(n3300), .I3(n3237), 
            .O(n37296));
    defparam i23207_4_lut.LUT_INIT = 16'h88a0;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_766_3_lut (.I0(GND_net), 
            .I1(n1133), .I2(VCC_net), .I3(n43988), .O(n1200)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_766_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1771_4 (.CI(n44229), 
            .I0(n2632), .I1(GND_net), .CO(n44230));
    SB_LUT4 i1_4_lut_adj_1781 (.I0(n37296), .I1(n51662), .I2(n5_adj_5606), 
            .I3(n7_adj_5647), .O(n51664));
    defparam i1_4_lut_adj_1781.LUT_INIT = 16'hfcec;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1771_3_lut (.I0(GND_net), 
            .I1(n2633), .I2(VCC_net), .I3(n44228), .O(n2700)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1771_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i836_3_lut (.I0(n1225), .I1(n1292), 
            .I2(n1257), .I3(GND_net), .O(n1324));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i836_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i840_3_lut (.I0(n1229), .I1(n1296), 
            .I2(n1257), .I3(GND_net), .O(n1328));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i840_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1771_3 (.CI(n44228), 
            .I0(n2633), .I1(VCC_net), .CO(n44229));
    SB_LUT4 i1_4_lut_adj_1782 (.I0(n3215), .I1(n51664), .I2(n3282), .I3(n3237), 
            .O(n51666));
    defparam i1_4_lut_adj_1782.LUT_INIT = 16'heefc;
    SB_LUT4 i1_4_lut_adj_1783 (.I0(n3214), .I1(n51666), .I2(n3281), .I3(n3237), 
            .O(n51668));
    defparam i1_4_lut_adj_1783.LUT_INIT = 16'heefc;
    SB_LUT4 unary_minus_19_inv_0_i3_1_lut (.I0(current[2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_5462));   // verilog/TinyFPGA_B.v(121[16:24])
    defparam unary_minus_19_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_4_lut_adj_1784 (.I0(n3213), .I1(n51668), .I2(n3280), .I3(n3237), 
            .O(n51670));
    defparam i1_4_lut_adj_1784.LUT_INIT = 16'heefc;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1771_2_lut (.I0(GND_net), 
            .I1(n537), .I2(GND_net), .I3(VCC_net), .O(n2701)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1771_2_lut.LUT_INIT = 16'hC33C;
    SB_DFF read_221 (.Q(read), .C(clk16MHz), .D(n51491));   // verilog/TinyFPGA_B.v(368[10] 396[6])
    SB_LUT4 i1_4_lut_adj_1785 (.I0(n3212), .I1(n51670), .I2(n3279), .I3(n3237), 
            .O(n51672));
    defparam i1_4_lut_adj_1785.LUT_INIT = 16'heefc;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_unary_minus_2_inv_0_i6_1_lut (.I0(encoder0_position_scaled_23__N_327[5]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n28_adj_5637));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_unary_minus_2_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1771_2 (.CI(VCC_net), 
            .I0(n537), .I1(GND_net), .CO(n44228));
    SB_LUT4 i1_4_lut_adj_1786 (.I0(n3211), .I1(n51672), .I2(n3278), .I3(n3237), 
            .O(n51674));
    defparam i1_4_lut_adj_1786.LUT_INIT = 16'heefc;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_766_3 (.CI(n43988), 
            .I0(n1133), .I1(VCC_net), .CO(n43989));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_unary_minus_2_inv_0_i7_1_lut (.I0(encoder0_position_scaled_23__N_327[6]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n27_adj_5636));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_unary_minus_2_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_4_lut_adj_1787 (.I0(n3210), .I1(n51674), .I2(n3277), .I3(n3237), 
            .O(n51676));
    defparam i1_4_lut_adj_1787.LUT_INIT = 16'heefc;
    SB_LUT4 i1_4_lut_adj_1788 (.I0(n3209), .I1(n51676), .I2(n3276), .I3(n3237), 
            .O(n51678));
    defparam i1_4_lut_adj_1788.LUT_INIT = 16'heefc;
    SB_LUT4 unary_minus_18_inv_0_i4_1_lut (.I0(duty[3]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n22));   // verilog/TinyFPGA_B.v(119[24:29])
    defparam unary_minus_18_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_19_inv_0_i4_1_lut (.I0(current[3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n22_adj_5461));   // verilog/TinyFPGA_B.v(121[16:24])
    defparam unary_minus_19_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_19_inv_0_i5_1_lut (.I0(current[4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_5460));   // verilog/TinyFPGA_B.v(121[16:24])
    defparam unary_minus_19_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_unary_minus_2_inv_0_i8_1_lut (.I0(encoder0_position_scaled_23__N_327[7]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n26_adj_5635));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_unary_minus_2_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i15337_3_lut (.I0(\data_out_frame[7] [6]), .I1(encoder0_position_scaled[14]), 
            .I2(n24210), .I3(GND_net), .O(n29417));   // verilog/coms.v(128[12] 303[6])
    defparam i15337_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1789 (.I0(n3208), .I1(n51678), .I2(n3275), .I3(n3237), 
            .O(n51680));
    defparam i1_4_lut_adj_1789.LUT_INIT = 16'heefc;
    SB_LUT4 unary_minus_19_inv_0_i6_1_lut (.I0(current[5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n20_adj_5459));   // verilog/TinyFPGA_B.v(121[16:24])
    defparam unary_minus_19_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_19_inv_0_i7_1_lut (.I0(current[6]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_5458));   // verilog/TinyFPGA_B.v(121[16:24])
    defparam unary_minus_19_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_4_lut_adj_1790 (.I0(n3207), .I1(n51680), .I2(n3274), .I3(n3237), 
            .O(n51682));
    defparam i1_4_lut_adj_1790.LUT_INIT = 16'heefc;
    SB_LUT4 unary_minus_19_inv_0_i8_1_lut (.I0(current[7]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n18_adj_5457));   // verilog/TinyFPGA_B.v(121[16:24])
    defparam unary_minus_19_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i2177_3_lut (.I0(n3206), 
            .I1(n3273), .I2(n3237), .I3(GND_net), .O(n59));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i2177_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i2176_3_lut (.I0(n3205), 
            .I1(n3272), .I2(n3237), .I3(GND_net), .O(n61));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i2176_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15896_3_lut (.I0(\data_out_frame[22] [1]), .I1(current[1]), 
            .I2(n24210), .I3(GND_net), .O(n29976));   // verilog/coms.v(128[12] 303[6])
    defparam i15896_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15897_3_lut (.I0(\data_out_frame[22] [0]), .I1(current[0]), 
            .I2(n24210), .I3(GND_net), .O(n29977));   // verilog/coms.v(128[12] 303[6])
    defparam i15897_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i40662_4_lut (.I0(n61), .I1(n53025), .I2(n59), .I3(n51682), 
            .O(n37482));
    defparam i40662_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i15898_3_lut (.I0(\data_out_frame[21] [7]), .I1(current[15]), 
            .I2(n24210), .I3(GND_net), .O(n29978));   // verilog/coms.v(128[12] 303[6])
    defparam i15898_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i2110_3_lut (.I0(n3107), 
            .I1(n3174), .I2(n3138), .I3(GND_net), .O(n3206));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i2110_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 unary_minus_18_inv_0_i5_1_lut (.I0(duty[4]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n21));   // verilog/TinyFPGA_B.v(119[24:29])
    defparam unary_minus_18_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i2109_3_lut (.I0(n3106), 
            .I1(n3173), .I2(n3138), .I3(GND_net), .O(n3205));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i2109_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15899_3_lut (.I0(\data_out_frame[21] [6]), .I1(current[15]), 
            .I2(n24210), .I3(GND_net), .O(n29979));   // verilog/coms.v(128[12] 303[6])
    defparam i15899_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i2113_3_lut (.I0(n3110), 
            .I1(n3177), .I2(n3138), .I3(GND_net), .O(n3209));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i2113_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15900_3_lut (.I0(\data_out_frame[21] [5]), .I1(current[15]), 
            .I2(n24210), .I3(GND_net), .O(n29980));   // verilog/coms.v(128[12] 303[6])
    defparam i15900_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15901_3_lut (.I0(\data_out_frame[21] [4]), .I1(current[15]), 
            .I2(n24210), .I3(GND_net), .O(n29981));   // verilog/coms.v(128[12] 303[6])
    defparam i15901_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15902_3_lut (.I0(\data_out_frame[21] [3]), .I1(current[11]), 
            .I2(n24210), .I3(GND_net), .O(n29982));   // verilog/coms.v(128[12] 303[6])
    defparam i15902_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i2112_3_lut (.I0(n3109), 
            .I1(n3176), .I2(n3138), .I3(GND_net), .O(n3208));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i2112_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i2111_3_lut (.I0(n3108), 
            .I1(n3175), .I2(n3138), .I3(GND_net), .O(n3207));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i2111_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i2135_3_lut (.I0(n3132), 
            .I1(n3199), .I2(n3138), .I3(GND_net), .O(n3231));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i2135_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15903_3_lut (.I0(\data_out_frame[21] [2]), .I1(current[10]), 
            .I2(n24210), .I3(GND_net), .O(n29983));   // verilog/coms.v(128[12] 303[6])
    defparam i15903_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15904_3_lut (.I0(\data_out_frame[21] [1]), .I1(current[9]), 
            .I2(n24210), .I3(GND_net), .O(n29984));   // verilog/coms.v(128[12] 303[6])
    defparam i15904_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i2134_3_lut (.I0(n3131), 
            .I1(n3198), .I2(n3138), .I3(GND_net), .O(n3230));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i2134_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i2133_3_lut (.I0(n3130), 
            .I1(n3197), .I2(n3138), .I3(GND_net), .O(n3229));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i2133_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i2116_3_lut (.I0(n3113), 
            .I1(n3180), .I2(n3138), .I3(GND_net), .O(n3212));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i2116_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i2115_3_lut (.I0(n3112), 
            .I1(n3179), .I2(n3138), .I3(GND_net), .O(n3211));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i2115_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i2114_3_lut (.I0(n3111), 
            .I1(n3178), .I2(n3138), .I3(GND_net), .O(n3210));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i2114_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i2118_3_lut (.I0(n3115), 
            .I1(n3182), .I2(n3138), .I3(GND_net), .O(n3214));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i2118_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i2117_3_lut (.I0(n3114), 
            .I1(n3181), .I2(n3138), .I3(GND_net), .O(n3213));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i2117_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i2120_3_lut (.I0(n3117), 
            .I1(n3184), .I2(n3138), .I3(GND_net), .O(n3216));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i2120_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i2119_3_lut (.I0(n3116), 
            .I1(n3183), .I2(n3138), .I3(GND_net), .O(n3215));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i2119_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i2137_3_lut (.I0(n542), .I1(n3201), 
            .I2(n3138), .I3(GND_net), .O(n3233));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i2137_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i2136_3_lut (.I0(n3133), 
            .I1(n3200), .I2(n3138), .I3(GND_net), .O(n3232));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i2136_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_mux_3_i2_3_lut (.I0(encoder0_position_scaled_23__N_327[1]), 
            .I1(n32), .I2(encoder0_position_scaled_23__N_327[31]), .I3(GND_net), 
            .O(n543));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_mux_3_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i2131_3_lut (.I0(n3128), 
            .I1(n3195), .I2(n3138), .I3(GND_net), .O(n3227));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i2131_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15905_3_lut (.I0(\data_out_frame[21] [0]), .I1(current[8]), 
            .I2(n24210), .I3(GND_net), .O(n29985));   // verilog/coms.v(128[12] 303[6])
    defparam i15905_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15906_3_lut (.I0(\data_out_frame[20] [7]), .I1(displacement[7]), 
            .I2(n24210), .I3(GND_net), .O(n29986));   // verilog/coms.v(128[12] 303[6])
    defparam i15906_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1107_3_lut (.I0(n1624), 
            .I1(n1691), .I2(n1653), .I3(GND_net), .O(n1723));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1107_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i2124_3_lut (.I0(n3121), 
            .I1(n3188), .I2(n3138), .I3(GND_net), .O(n3220));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i2124_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i2123_3_lut (.I0(n3120), 
            .I1(n3187), .I2(n3138), .I3(GND_net), .O(n3219));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i2123_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15907_3_lut (.I0(\data_out_frame[20] [6]), .I1(displacement[6]), 
            .I2(n24210), .I3(GND_net), .O(n29987));   // verilog/coms.v(128[12] 303[6])
    defparam i15907_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1704_25_lut (.I0(n56142), 
            .I1(n2511), .I2(VCC_net), .I3(n44227), .O(n2610)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1704_25_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1704_24_lut (.I0(GND_net), 
            .I1(n2512), .I2(VCC_net), .I3(n44226), .O(n2579)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1704_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1704_24 (.CI(n44226), 
            .I0(n2512), .I1(VCC_net), .CO(n44227));
    SB_LUT4 add_175_20_lut (.I0(GND_net), .I1(delay_counter[18]), .I2(GND_net), 
            .I3(n43627), .O(n1545)) /* synthesis syn_instantiated=1 */ ;
    defparam add_175_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1704_23_lut (.I0(GND_net), 
            .I1(n2513), .I2(VCC_net), .I3(n44225), .O(n2580)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1704_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i2125_3_lut (.I0(n3122), 
            .I1(n3189), .I2(n3138), .I3(GND_net), .O(n3221));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i2125_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15908_3_lut (.I0(\data_out_frame[20] [5]), .I1(displacement[5]), 
            .I2(n24210), .I3(GND_net), .O(n29988));   // verilog/coms.v(128[12] 303[6])
    defparam i15908_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1704_23 (.CI(n44225), 
            .I0(n2513), .I1(VCC_net), .CO(n44226));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i839_3_lut (.I0(n1228), .I1(n1295), 
            .I2(n1257), .I3(GND_net), .O(n1327));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i839_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1704_22_lut (.I0(GND_net), 
            .I1(n2514), .I2(VCC_net), .I3(n44224), .O(n2581)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1704_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15909_3_lut (.I0(\data_out_frame[20] [4]), .I1(displacement[4]), 
            .I2(n24210), .I3(GND_net), .O(n29989));   // verilog/coms.v(128[12] 303[6])
    defparam i15909_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15910_3_lut (.I0(\data_out_frame[20] [3]), .I1(displacement[3]), 
            .I2(n24210), .I3(GND_net), .O(n29990));   // verilog/coms.v(128[12] 303[6])
    defparam i15910_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i2122_3_lut (.I0(n3119), 
            .I1(n3186), .I2(n3138), .I3(GND_net), .O(n3218));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i2122_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i838_3_lut (.I0(n1227), .I1(n1294), 
            .I2(n1257), .I3(GND_net), .O(n1326));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i838_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i2129_3_lut (.I0(n3126), 
            .I1(n3193), .I2(n3138), .I3(GND_net), .O(n3225));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i2129_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15911_3_lut (.I0(\data_out_frame[20] [2]), .I1(displacement[2]), 
            .I2(n24210), .I3(GND_net), .O(n29991));   // verilog/coms.v(128[12] 303[6])
    defparam i15911_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i2130_3_lut (.I0(n3127), 
            .I1(n3194), .I2(n3138), .I3(GND_net), .O(n3226));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i2130_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i2132_3_lut (.I0(n3129), 
            .I1(n3196), .I2(n3138), .I3(GND_net), .O(n3228));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i2132_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15912_3_lut (.I0(\data_out_frame[20] [1]), .I1(displacement[1]), 
            .I2(n24210), .I3(GND_net), .O(n29992));   // verilog/coms.v(128[12] 303[6])
    defparam i15912_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15913_3_lut (.I0(\data_out_frame[20] [0]), .I1(displacement[0]), 
            .I2(n24210), .I3(GND_net), .O(n29993));   // verilog/coms.v(128[12] 303[6])
    defparam i15913_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i837_3_lut (.I0(n1226), .I1(n1293), 
            .I2(n1257), .I3(GND_net), .O(n1325));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i837_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1704_22 (.CI(n44224), 
            .I0(n2514), .I1(VCC_net), .CO(n44225));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1704_21_lut (.I0(GND_net), 
            .I1(n2515), .I2(VCC_net), .I3(n44223), .O(n2582)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1704_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1704_21 (.CI(n44223), 
            .I0(n2515), .I1(VCC_net), .CO(n44224));
    SB_LUT4 i34003_3_lut (.I0(n4_adj_5495), .I1(n8583), .I2(n49748), .I3(GND_net), 
            .O(n49751));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam i34003_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i2128_3_lut (.I0(n3125), 
            .I1(n3192), .I2(n3138), .I3(GND_net), .O(n3224));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i2128_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i2127_3_lut (.I0(n3124), 
            .I1(n3191), .I2(n3138), .I3(GND_net), .O(n3223));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i2127_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15914_3_lut (.I0(\data_out_frame[19] [7]), .I1(displacement[15]), 
            .I2(n24210), .I3(GND_net), .O(n29994));   // verilog/coms.v(128[12] 303[6])
    defparam i15914_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i2121_3_lut (.I0(n3118), 
            .I1(n3185), .I2(n3138), .I3(GND_net), .O(n3217));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i2121_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i2126_3_lut (.I0(n3123), 
            .I1(n3190), .I2(n3138), .I3(GND_net), .O(n3222));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i2126_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1704_20_lut (.I0(GND_net), 
            .I1(n2516), .I2(VCC_net), .I3(n44222), .O(n2583)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1704_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1791 (.I0(n3225), .I1(n3218), .I2(n3221), .I3(n3219), 
            .O(n52242));
    defparam i1_4_lut_adj_1791.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_adj_1792 (.I0(n3220), .I1(n3227), .I2(GND_net), .I3(GND_net), 
            .O(n52232));
    defparam i1_2_lut_adj_1792.LUT_INIT = 16'heeee;
    SB_LUT4 i15915_3_lut (.I0(\data_out_frame[19] [6]), .I1(displacement[14]), 
            .I2(n24210), .I3(GND_net), .O(n29995));   // verilog/coms.v(128[12] 303[6])
    defparam i15915_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15916_3_lut (.I0(\data_out_frame[19] [5]), .I1(displacement[13]), 
            .I2(n24210), .I3(GND_net), .O(n29996));   // verilog/coms.v(128[12] 303[6])
    defparam i15916_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15917_3_lut (.I0(\data_out_frame[19] [4]), .I1(displacement[12]), 
            .I2(n24210), .I3(GND_net), .O(n29997));   // verilog/coms.v(128[12] 303[6])
    defparam i15917_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_175_20 (.CI(n43627), .I0(delay_counter[18]), .I1(GND_net), 
            .CO(n43628));
    SB_LUT4 i1_4_lut_adj_1793 (.I0(n3222), .I1(n3217), .I2(n52232), .I3(n3223), 
            .O(n52244));
    defparam i1_4_lut_adj_1793.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_766_2_lut (.I0(GND_net), 
            .I1(n411), .I2(GND_net), .I3(VCC_net), .O(n1201)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_766_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_766_2 (.CI(VCC_net), 
            .I0(n411), .I1(GND_net), .CO(n43988));
    SB_LUT4 i1_4_lut_adj_1794 (.I0(n52242), .I1(n3224), .I2(n3228), .I3(n3226), 
            .O(n52246));
    defparam i1_4_lut_adj_1794.LUT_INIT = 16'hfffe;
    SB_LUT4 i23209_3_lut (.I0(n543), .I1(n3232), .I2(n3233), .I3(GND_net), 
            .O(n37298));
    defparam i23209_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i1_4_lut_adj_1795 (.I0(n3215), .I1(n3216), .I2(n52246), .I3(n52244), 
            .O(n52252));
    defparam i1_4_lut_adj_1795.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1796 (.I0(n3229), .I1(n37298), .I2(n3230), .I3(n3231), 
            .O(n50148));
    defparam i1_4_lut_adj_1796.LUT_INIT = 16'ha080;
    SB_LUT4 unary_minus_19_inv_0_i9_1_lut (.I0(current[8]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_5456));   // verilog/TinyFPGA_B.v(121[16:24])
    defparam unary_minus_19_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_4_lut_adj_1797 (.I0(n3213), .I1(n3214), .I2(n50148), .I3(n52252), 
            .O(n52258));
    defparam i1_4_lut_adj_1797.LUT_INIT = 16'hfffe;
    SB_LUT4 unary_minus_19_inv_0_i10_1_lut (.I0(current[9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n16_adj_5455));   // verilog/TinyFPGA_B.v(121[16:24])
    defparam unary_minus_19_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i15918_3_lut (.I0(\data_out_frame[19] [3]), .I1(displacement[11]), 
            .I2(n24210), .I3(GND_net), .O(n29998));   // verilog/coms.v(128[12] 303[6])
    defparam i15918_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15919_3_lut (.I0(\data_out_frame[19] [2]), .I1(displacement[10]), 
            .I2(n24210), .I3(GND_net), .O(n29999));   // verilog/coms.v(128[12] 303[6])
    defparam i15919_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1798 (.I0(n3210), .I1(n3211), .I2(n3212), .I3(n52258), 
            .O(n52264));
    defparam i1_4_lut_adj_1798.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1799 (.I0(n3207), .I1(n3208), .I2(n3209), .I3(n52264), 
            .O(n52270));
    defparam i1_4_lut_adj_1799.LUT_INIT = 16'hfffe;
    SB_LUT4 i15920_3_lut (.I0(\data_out_frame[19] [1]), .I1(displacement[9]), 
            .I2(n24210), .I3(GND_net), .O(n30000));   // verilog/coms.v(128[12] 303[6])
    defparam i15920_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15921_3_lut (.I0(\data_out_frame[19] [0]), .I1(displacement[8]), 
            .I2(n24210), .I3(GND_net), .O(n30001));   // verilog/coms.v(128[12] 303[6])
    defparam i15921_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15922_3_lut (.I0(\data_out_frame[18] [7]), .I1(displacement[23]), 
            .I2(n24210), .I3(GND_net), .O(n30002));   // verilog/coms.v(128[12] 303[6])
    defparam i15922_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i40700_4_lut (.I0(n3205), .I1(n3204), .I2(n3206), .I3(n52270), 
            .O(n3237));
    defparam i40700_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i2043_3_lut (.I0(n3008), 
            .I1(n3075), .I2(n3039), .I3(GND_net), .O(n3107));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i2043_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15923_3_lut (.I0(\data_out_frame[18] [6]), .I1(displacement[22]), 
            .I2(n24210), .I3(GND_net), .O(n30003));   // verilog/coms.v(128[12] 303[6])
    defparam i15923_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15924_3_lut (.I0(\data_out_frame[18] [5]), .I1(displacement[21]), 
            .I2(n24210), .I3(GND_net), .O(n30004));   // verilog/coms.v(128[12] 303[6])
    defparam i15924_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15925_3_lut (.I0(\data_out_frame[18] [4]), .I1(displacement[20]), 
            .I2(n24210), .I3(GND_net), .O(n30005));   // verilog/coms.v(128[12] 303[6])
    defparam i15925_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1704_20 (.CI(n44222), 
            .I0(n2516), .I1(VCC_net), .CO(n44223));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i2042_3_lut (.I0(n3007), 
            .I1(n3074), .I2(n3039), .I3(GND_net), .O(n3106));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i2042_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15926_3_lut (.I0(\data_out_frame[18] [3]), .I1(displacement[19]), 
            .I2(n24210), .I3(GND_net), .O(n30006));   // verilog/coms.v(128[12] 303[6])
    defparam i15926_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1704_19_lut (.I0(GND_net), 
            .I1(n2517), .I2(VCC_net), .I3(n44221), .O(n2584)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1704_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15927_3_lut (.I0(\data_out_frame[18] [2]), .I1(displacement[18]), 
            .I2(n24210), .I3(GND_net), .O(n30007));   // verilog/coms.v(128[12] 303[6])
    defparam i15927_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15928_3_lut (.I0(\data_out_frame[18] [1]), .I1(displacement[17]), 
            .I2(n24210), .I3(GND_net), .O(n30008));   // verilog/coms.v(128[12] 303[6])
    defparam i15928_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_699_10_lut (.I0(GND_net), 
            .I1(n1026), .I2(VCC_net), .I3(n43987), .O(n1093)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_699_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i2045_3_lut (.I0(n3010), 
            .I1(n3077), .I2(n3039), .I3(GND_net), .O(n3109));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i2045_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i2044_3_lut (.I0(n3009), 
            .I1(n3076), .I2(n3039), .I3(GND_net), .O(n3108));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i2044_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15929_3_lut (.I0(\data_out_frame[18] [0]), .I1(displacement[16]), 
            .I2(n24210), .I3(GND_net), .O(n30009));   // verilog/coms.v(128[12] 303[6])
    defparam i15929_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_699_9_lut (.I0(GND_net), 
            .I1(n1027), .I2(VCC_net), .I3(n43986), .O(n1094)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_699_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15930_3_lut (.I0(\data_out_frame[17] [7]), .I1(pwm_setpoint[7]), 
            .I2(n24210), .I3(GND_net), .O(n30010));   // verilog/coms.v(128[12] 303[6])
    defparam i15930_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i2050_3_lut (.I0(n3015), 
            .I1(n3082), .I2(n3039), .I3(GND_net), .O(n3114));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i2050_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1704_19 (.CI(n44221), 
            .I0(n2517), .I1(VCC_net), .CO(n44222));
    SB_LUT4 i15931_3_lut (.I0(\data_out_frame[17] [6]), .I1(pwm_setpoint[6]), 
            .I2(n24210), .I3(GND_net), .O(n30011));   // verilog/coms.v(128[12] 303[6])
    defparam i15931_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1704_18_lut (.I0(GND_net), 
            .I1(n2518), .I2(VCC_net), .I3(n44220), .O(n2585)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1704_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1704_18 (.CI(n44220), 
            .I0(n2518), .I1(VCC_net), .CO(n44221));
    SB_LUT4 unary_minus_19_inv_0_i11_1_lut (.I0(current[10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_5454));   // verilog/TinyFPGA_B.v(121[16:24])
    defparam unary_minus_19_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i2049_3_lut (.I0(n3014), 
            .I1(n3081), .I2(n3039), .I3(GND_net), .O(n3113));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i2049_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i2046_3_lut (.I0(n3011), 
            .I1(n3078), .I2(n3039), .I3(GND_net), .O(n3110));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i2046_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i2054_3_lut (.I0(n3019), 
            .I1(n3086), .I2(n3039), .I3(GND_net), .O(n3118));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i2054_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1704_17_lut (.I0(GND_net), 
            .I1(n2519), .I2(VCC_net), .I3(n44219), .O(n2586)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1704_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i2053_3_lut (.I0(n3018), 
            .I1(n3085), .I2(n3039), .I3(GND_net), .O(n3117));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i2053_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15932_3_lut (.I0(\data_out_frame[17] [5]), .I1(pwm_setpoint[5]), 
            .I2(n24210), .I3(GND_net), .O(n30012));   // verilog/coms.v(128[12] 303[6])
    defparam i15932_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i2048_3_lut (.I0(n3013), 
            .I1(n3080), .I2(n3039), .I3(GND_net), .O(n3112));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i2048_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15933_3_lut (.I0(\data_out_frame[17] [4]), .I1(pwm_setpoint[4]), 
            .I2(n24210), .I3(GND_net), .O(n30013));   // verilog/coms.v(128[12] 303[6])
    defparam i15933_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15934_3_lut (.I0(\data_out_frame[17] [3]), .I1(pwm_setpoint[3]), 
            .I2(n24210), .I3(GND_net), .O(n30014));   // verilog/coms.v(128[12] 303[6])
    defparam i15934_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i2055_3_lut (.I0(n3020), 
            .I1(n3087), .I2(n3039), .I3(GND_net), .O(n3119));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i2055_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_699_9 (.CI(n43986), 
            .I0(n1027), .I1(VCC_net), .CO(n43987));
    SB_LUT4 i15935_3_lut (.I0(\data_out_frame[17] [2]), .I1(pwm_setpoint[2]), 
            .I2(n24210), .I3(GND_net), .O(n30015));   // verilog/coms.v(128[12] 303[6])
    defparam i15935_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15936_3_lut (.I0(\data_out_frame[17] [1]), .I1(pwm_setpoint[1]), 
            .I2(n24210), .I3(GND_net), .O(n30016));   // verilog/coms.v(128[12] 303[6])
    defparam i15936_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_699_8_lut (.I0(GND_net), 
            .I1(n1028), .I2(VCC_net), .I3(n43985), .O(n1095)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_699_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15937_3_lut (.I0(\data_out_frame[17] [0]), .I1(pwm_setpoint[0]), 
            .I2(n24210), .I3(GND_net), .O(n30017));   // verilog/coms.v(128[12] 303[6])
    defparam i15937_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i2056_3_lut (.I0(n3021), 
            .I1(n3088), .I2(n3039), .I3(GND_net), .O(n3120));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i2056_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i2069_3_lut (.I0(n541), .I1(n3101), 
            .I2(n3039), .I3(GND_net), .O(n3133));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i2069_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15938_3_lut (.I0(\data_out_frame[16] [7]), .I1(pwm_setpoint[15]), 
            .I2(n24210), .I3(GND_net), .O(n30018));   // verilog/coms.v(128[12] 303[6])
    defparam i15938_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15939_3_lut (.I0(\data_out_frame[16] [6]), .I1(pwm_setpoint[14]), 
            .I2(n24210), .I3(GND_net), .O(n30019));   // verilog/coms.v(128[12] 303[6])
    defparam i15939_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i2068_3_lut (.I0(n3033), 
            .I1(n3100), .I2(n3039), .I3(GND_net), .O(n3132));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i2068_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15940_3_lut (.I0(\data_out_frame[16] [5]), .I1(pwm_setpoint[13]), 
            .I2(n24210), .I3(GND_net), .O(n30020));   // verilog/coms.v(128[12] 303[6])
    defparam i15940_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1704_17 (.CI(n44219), 
            .I0(n2519), .I1(VCC_net), .CO(n44220));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_699_8 (.CI(n43985), 
            .I0(n1028), .I1(VCC_net), .CO(n43986));
    SB_LUT4 i15941_3_lut (.I0(\data_out_frame[16] [4]), .I1(pwm_setpoint[12]), 
            .I2(n24210), .I3(GND_net), .O(n30021));   // verilog/coms.v(128[12] 303[6])
    defparam i15941_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i2067_3_lut (.I0(n3032), 
            .I1(n3099), .I2(n3039), .I3(GND_net), .O(n3131));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i2067_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1704_16_lut (.I0(GND_net), 
            .I1(n2520), .I2(VCC_net), .I3(n44218), .O(n2587)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1704_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_mux_3_i3_3_lut (.I0(encoder0_position_scaled_23__N_327[2]), 
            .I1(n31), .I2(encoder0_position_scaled_23__N_327[31]), .I3(GND_net), 
            .O(n542));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_mux_3_i3_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15942_3_lut (.I0(\data_out_frame[16] [3]), .I1(pwm_setpoint[11]), 
            .I2(n24210), .I3(GND_net), .O(n30022));   // verilog/coms.v(128[12] 303[6])
    defparam i15942_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15943_3_lut (.I0(\data_out_frame[16] [2]), .I1(pwm_setpoint[10]), 
            .I2(n24210), .I3(GND_net), .O(n30023));   // verilog/coms.v(128[12] 303[6])
    defparam i15943_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1704_16 (.CI(n44218), 
            .I0(n2520), .I1(VCC_net), .CO(n44219));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_699_7_lut (.I0(GND_net), 
            .I1(n1029), .I2(GND_net), .I3(n43984), .O(n1096)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_699_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i2063_3_lut (.I0(n3028), 
            .I1(n3095), .I2(n3039), .I3(GND_net), .O(n3127));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i2063_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15944_3_lut (.I0(\data_out_frame[16] [1]), .I1(pwm_setpoint[9]), 
            .I2(n24210), .I3(GND_net), .O(n30024));   // verilog/coms.v(128[12] 303[6])
    defparam i15944_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1704_15_lut (.I0(GND_net), 
            .I1(n2521), .I2(VCC_net), .I3(n44217), .O(n2588)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1704_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1704_15 (.CI(n44217), 
            .I0(n2521), .I1(VCC_net), .CO(n44218));
    SB_LUT4 unary_minus_19_inv_0_i12_1_lut (.I0(current[11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n14_adj_5453));   // verilog/TinyFPGA_B.v(121[16:24])
    defparam unary_minus_19_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_699_7 (.CI(n43984), 
            .I0(n1029), .I1(GND_net), .CO(n43985));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i2058_3_lut (.I0(n3023), 
            .I1(n3090), .I2(n3039), .I3(GND_net), .O(n3122));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i2058_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15945_3_lut (.I0(\data_out_frame[16] [0]), .I1(pwm_setpoint[8]), 
            .I2(n24210), .I3(GND_net), .O(n30025));   // verilog/coms.v(128[12] 303[6])
    defparam i15945_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15946_3_lut (.I0(\data_out_frame[15] [7]), .I1(pwm_setpoint[23]), 
            .I2(n24210), .I3(GND_net), .O(n30026));   // verilog/coms.v(128[12] 303[6])
    defparam i15946_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i2057_3_lut (.I0(n3022), 
            .I1(n3089), .I2(n3039), .I3(GND_net), .O(n3121));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i2057_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_699_6_lut (.I0(GND_net), 
            .I1(n1030), .I2(GND_net), .I3(n43983), .O(n1097)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_699_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15947_3_lut (.I0(\data_out_frame[15] [6]), .I1(pwm_setpoint[22]), 
            .I2(n24210), .I3(GND_net), .O(n30027));   // verilog/coms.v(128[12] 303[6])
    defparam i15947_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15948_3_lut (.I0(\data_out_frame[15] [5]), .I1(pwm_setpoint[21]), 
            .I2(n24210), .I3(GND_net), .O(n30028));   // verilog/coms.v(128[12] 303[6])
    defparam i15948_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15678_4_lut (.I0(CS_MISO_c), .I1(data_adj_5711[1]), .I2(n6_adj_5556), 
            .I3(n27271), .O(n29758));   // verilog/tli4970.v(35[10] 68[6])
    defparam i15678_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i2047_3_lut (.I0(n3012), 
            .I1(n3079), .I2(n3039), .I3(GND_net), .O(n3111));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i2047_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15949_3_lut (.I0(\data_out_frame[15] [4]), .I1(pwm_setpoint[20]), 
            .I2(n24210), .I3(GND_net), .O(n30029));   // verilog/coms.v(128[12] 303[6])
    defparam i15949_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15679_4_lut (.I0(r_Rx_Data), .I1(rx_data[1]), .I2(n4_adj_5443), 
            .I3(n27203), .O(n29759));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i15679_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i15950_3_lut (.I0(\data_out_frame[15] [3]), .I1(pwm_setpoint[19]), 
            .I2(n24210), .I3(GND_net), .O(n30030));   // verilog/coms.v(128[12] 303[6])
    defparam i15950_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1704_14_lut (.I0(GND_net), 
            .I1(n2522), .I2(VCC_net), .I3(n44216), .O(n2589)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1704_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_699_6 (.CI(n43983), 
            .I0(n1030), .I1(GND_net), .CO(n43984));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_unary_minus_2_inv_0_i9_1_lut (.I0(encoder0_position_scaled_23__N_327[8]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n25_adj_5634));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_unary_minus_2_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i2051_3_lut (.I0(n3016), 
            .I1(n3083), .I2(n3039), .I3(GND_net), .O(n3115));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i2051_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15951_3_lut (.I0(\data_out_frame[15] [2]), .I1(pwm_setpoint[18]), 
            .I2(n24210), .I3(GND_net), .O(n30031));   // verilog/coms.v(128[12] 303[6])
    defparam i15951_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15952_3_lut (.I0(\data_out_frame[15] [1]), .I1(pwm_setpoint[17]), 
            .I2(n24210), .I3(GND_net), .O(n30032));   // verilog/coms.v(128[12] 303[6])
    defparam i15952_3_lut.LUT_INIT = 16'hcaca;
    SB_IO CS_MISO_pad (.PACKAGE_PIN(CS_MISO), .OUTPUT_ENABLE(VCC_net), .D_IN_0(CS_MISO_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam CS_MISO_pad.PIN_TYPE = 6'b000001;
    defparam CS_MISO_pad.PULLUP = 1'b0;
    defparam CS_MISO_pad.NEG_TRIGGER = 1'b0;
    defparam CS_MISO_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_699_5_lut (.I0(GND_net), 
            .I1(n1031), .I2(VCC_net), .I3(n43982), .O(n1098)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_699_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_699_5 (.CI(n43982), 
            .I0(n1031), .I1(VCC_net), .CO(n43983));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i2062_3_lut (.I0(n3027), 
            .I1(n3094), .I2(n3039), .I3(GND_net), .O(n3126));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i2062_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15953_3_lut (.I0(\data_out_frame[15] [0]), .I1(pwm_setpoint[16]), 
            .I2(n24210), .I3(GND_net), .O(n30033));   // verilog/coms.v(128[12] 303[6])
    defparam i15953_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15954_3_lut (.I0(\data_out_frame[14] [7]), .I1(setpoint[7]), 
            .I2(n24210), .I3(GND_net), .O(n30034));   // verilog/coms.v(128[12] 303[6])
    defparam i15954_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_699_4_lut (.I0(GND_net), 
            .I1(n1032), .I2(GND_net), .I3(n43981), .O(n1099)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_699_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1704_14 (.CI(n44216), 
            .I0(n2522), .I1(VCC_net), .CO(n44217));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_699_4 (.CI(n43981), 
            .I0(n1032), .I1(GND_net), .CO(n43982));
    SB_LUT4 add_175_19_lut (.I0(GND_net), .I1(delay_counter[17]), .I2(GND_net), 
            .I3(n43626), .O(n1546)) /* synthesis syn_instantiated=1 */ ;
    defparam add_175_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1704_13_lut (.I0(GND_net), 
            .I1(n2523), .I2(VCC_net), .I3(n44215), .O(n2590)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1704_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_699_3_lut (.I0(GND_net), 
            .I1(n1033), .I2(VCC_net), .I3(n43980), .O(n1100)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_699_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_699_3 (.CI(n43980), 
            .I0(n1033), .I1(VCC_net), .CO(n43981));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i2059_3_lut (.I0(n3024), 
            .I1(n3091), .I2(n3039), .I3(GND_net), .O(n3123));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i2059_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15955_3_lut (.I0(\data_out_frame[14] [6]), .I1(setpoint[6]), 
            .I2(n24210), .I3(GND_net), .O(n30035));   // verilog/coms.v(128[12] 303[6])
    defparam i15955_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i2061_3_lut (.I0(n3026), 
            .I1(n3093), .I2(n3039), .I3(GND_net), .O(n3125));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i2061_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i2052_3_lut (.I0(n3017), 
            .I1(n3084), .I2(n3039), .I3(GND_net), .O(n3116));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i2052_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1704_13 (.CI(n44215), 
            .I0(n2523), .I1(VCC_net), .CO(n44216));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1704_12_lut (.I0(GND_net), 
            .I1(n2524), .I2(VCC_net), .I3(n44214), .O(n2591)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1704_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_699_2_lut (.I0(GND_net), 
            .I1(n935), .I2(GND_net), .I3(VCC_net), .O(n1101)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_699_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15956_3_lut (.I0(\data_out_frame[14] [5]), .I1(setpoint[5]), 
            .I2(n24210), .I3(GND_net), .O(n30036));   // verilog/coms.v(128[12] 303[6])
    defparam i15956_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i2066_3_lut (.I0(n3031), 
            .I1(n3098), .I2(n3039), .I3(GND_net), .O(n3130));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i2066_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i34004_3_lut (.I0(encoder0_position_scaled_23__N_327[29]), .I1(n49751), 
            .I2(encoder0_position_scaled_23__N_327[31]), .I3(GND_net), .O(n830));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam i34004_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_699_2 (.CI(VCC_net), 
            .I0(n935), .I1(GND_net), .CO(n43980));
    SB_LUT4 i15957_3_lut (.I0(\data_out_frame[14] [4]), .I1(setpoint[4]), 
            .I2(n24210), .I3(GND_net), .O(n30037));   // verilog/coms.v(128[12] 303[6])
    defparam i15957_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1704_12 (.CI(n44214), 
            .I0(n2524), .I1(VCC_net), .CO(n44215));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1704_11_lut (.I0(GND_net), 
            .I1(n2525), .I2(VCC_net), .I3(n44213), .O(n2592)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1704_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_632_9_lut (.I0(n960), 
            .I1(n927), .I2(VCC_net), .I3(n43979), .O(n1026)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_632_9_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_632_8_lut (.I0(GND_net), 
            .I1(n928), .I2(VCC_net), .I3(n43978), .O(n995)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_632_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15958_3_lut (.I0(\data_out_frame[14] [3]), .I1(setpoint[3]), 
            .I2(n24210), .I3(GND_net), .O(n30038));   // verilog/coms.v(128[12] 303[6])
    defparam i15958_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i569_3_lut (.I0(n830), .I1(n897), 
            .I2(n861), .I3(GND_net), .O(n929));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i569_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_632_8 (.CI(n43978), 
            .I0(n928), .I1(VCC_net), .CO(n43979));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1704_11 (.CI(n44213), 
            .I0(n2525), .I1(VCC_net), .CO(n44214));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i2065_3_lut (.I0(n3030), 
            .I1(n3097), .I2(n3039), .I3(GND_net), .O(n3129));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i2065_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10_1_lut (.I0(current[15]), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n2));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_632_7_lut (.I0(GND_net), 
            .I1(n929), .I2(GND_net), .I3(n43977), .O(n996)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_632_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1704_10_lut (.I0(GND_net), 
            .I1(n2526), .I2(VCC_net), .I3(n44212), .O(n2593)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1704_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i2064_3_lut (.I0(n3029), 
            .I1(n3096), .I2(n3039), .I3(GND_net), .O(n3128));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i2064_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15959_3_lut (.I0(\data_out_frame[14] [2]), .I1(setpoint[2]), 
            .I2(n24210), .I3(GND_net), .O(n30039));   // verilog/coms.v(128[12] 303[6])
    defparam i15959_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15960_3_lut (.I0(\data_out_frame[14] [1]), .I1(setpoint[1]), 
            .I2(n24210), .I3(GND_net), .O(n30040));   // verilog/coms.v(128[12] 303[6])
    defparam i15960_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i636_3_lut (.I0(n929), .I1(n996), 
            .I2(n960), .I3(GND_net), .O(n1028));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i636_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15961_3_lut (.I0(\data_out_frame[14] [0]), .I1(setpoint[0]), 
            .I2(n24210), .I3(GND_net), .O(n30041));   // verilog/coms.v(128[12] 303[6])
    defparam i15961_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i2060_3_lut (.I0(n3025), 
            .I1(n3092), .I2(n3039), .I3(GND_net), .O(n3124));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i2060_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15962_3_lut (.I0(\data_out_frame[13] [7]), .I1(setpoint[15]), 
            .I2(n24210), .I3(GND_net), .O(n30042));   // verilog/coms.v(128[12] 303[6])
    defparam i15962_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i703_3_lut (.I0(n1028), .I1(n1095), 
            .I2(n1059), .I3(GND_net), .O(n1127));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i703_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i40730_1_lut (.I0(n3138), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n56561));
    defparam i40730_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_2_lut_adj_1800 (.I0(n3124), .I1(n3128), .I2(GND_net), .I3(GND_net), 
            .O(n51690));
    defparam i1_2_lut_adj_1800.LUT_INIT = 16'heeee;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1704_10 (.CI(n44212), 
            .I0(n2526), .I1(VCC_net), .CO(n44213));
    SB_LUT4 i1_4_lut_adj_1801 (.I0(n3121), .I1(n51690), .I2(n3122), .I3(n3127), 
            .O(n51694));
    defparam i1_4_lut_adj_1801.LUT_INIT = 16'hfffe;
    SB_LUT4 i23282_4_lut (.I0(n542), .I1(n3131), .I2(n3132), .I3(n3133), 
            .O(n37372));
    defparam i23282_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1704_9_lut (.I0(GND_net), 
            .I1(n2527), .I2(VCC_net), .I3(n44211), .O(n2594)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1704_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1704_9 (.CI(n44211), 
            .I0(n2527), .I1(VCC_net), .CO(n44212));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_632_7 (.CI(n43977), 
            .I0(n929), .I1(GND_net), .CO(n43978));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1704_8_lut (.I0(GND_net), 
            .I1(n2528), .I2(VCC_net), .I3(n44210), .O(n2595)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1704_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_adj_1802 (.I0(n3120), .I1(n3119), .I2(GND_net), .I3(GND_net), 
            .O(n51998));
    defparam i1_2_lut_adj_1802.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_1803 (.I0(n3129), .I1(n51998), .I2(n37372), .I3(n3130), 
            .O(n52000));
    defparam i1_4_lut_adj_1803.LUT_INIT = 16'heccc;
    SB_LUT4 i15963_3_lut (.I0(\data_out_frame[13] [6]), .I1(setpoint[14]), 
            .I2(n24210), .I3(GND_net), .O(n30043));   // verilog/coms.v(128[12] 303[6])
    defparam i15963_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1804 (.I0(n3112), .I1(n3117), .I2(n51694), .I3(n3118), 
            .O(n51700));
    defparam i1_4_lut_adj_1804.LUT_INIT = 16'hfffe;
    SB_LUT4 i15964_3_lut (.I0(\data_out_frame[13] [5]), .I1(setpoint[13]), 
            .I2(n24210), .I3(GND_net), .O(n30044));   // verilog/coms.v(128[12] 303[6])
    defparam i15964_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15965_3_lut (.I0(\data_out_frame[13] [4]), .I1(setpoint[12]), 
            .I2(n24210), .I3(GND_net), .O(n30045));   // verilog/coms.v(128[12] 303[6])
    defparam i15965_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1704_8 (.CI(n44210), 
            .I0(n2528), .I1(VCC_net), .CO(n44211));
    SB_LUT4 i15966_3_lut (.I0(\data_out_frame[13] [3]), .I1(setpoint[11]), 
            .I2(n24210), .I3(GND_net), .O(n30046));   // verilog/coms.v(128[12] 303[6])
    defparam i15966_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1805 (.I0(n3116), .I1(n3125), .I2(n3123), .I3(n3126), 
            .O(n51946));
    defparam i1_4_lut_adj_1805.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1806 (.I0(n3115), .I1(n51700), .I2(n3111), .I3(n52000), 
            .O(n51702));
    defparam i1_4_lut_adj_1806.LUT_INIT = 16'hfffe;
    SB_LUT4 i15967_3_lut (.I0(\data_out_frame[13] [2]), .I1(setpoint[10]), 
            .I2(n24210), .I3(GND_net), .O(n30047));   // verilog/coms.v(128[12] 303[6])
    defparam i15967_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1807 (.I0(n3110), .I1(n3113), .I2(n3114), .I3(n51946), 
            .O(n51952));
    defparam i1_4_lut_adj_1807.LUT_INIT = 16'hfffe;
    SB_LUT4 i15968_3_lut (.I0(\data_out_frame[13] [1]), .I1(setpoint[9]), 
            .I2(n24210), .I3(GND_net), .O(n30048));   // verilog/coms.v(128[12] 303[6])
    defparam i15968_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1704_7_lut (.I0(GND_net), 
            .I1(n2529), .I2(GND_net), .I3(n44209), .O(n2596)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1704_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15969_3_lut (.I0(\data_out_frame[13] [0]), .I1(setpoint[8]), 
            .I2(n24210), .I3(GND_net), .O(n30049));   // verilog/coms.v(128[12] 303[6])
    defparam i15969_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_175_19 (.CI(n43626), .I0(delay_counter[17]), .I1(GND_net), 
            .CO(n43627));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1704_7 (.CI(n44209), 
            .I0(n2529), .I1(GND_net), .CO(n44210));
    SB_LUT4 i15970_3_lut (.I0(\data_out_frame[12] [7]), .I1(setpoint[23]), 
            .I2(n24210), .I3(GND_net), .O(n30050));   // verilog/coms.v(128[12] 303[6])
    defparam i15970_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15971_3_lut (.I0(\data_out_frame[12] [6]), .I1(setpoint[22]), 
            .I2(n24210), .I3(GND_net), .O(n30051));   // verilog/coms.v(128[12] 303[6])
    defparam i15971_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1704_6_lut (.I0(GND_net), 
            .I1(n2530), .I2(GND_net), .I3(n44208), .O(n2597)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1704_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_632_6_lut (.I0(GND_net), 
            .I1(n930), .I2(GND_net), .I3(n43976), .O(n997)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_632_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1704_6 (.CI(n44208), 
            .I0(n2530), .I1(GND_net), .CO(n44209));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1704_5_lut (.I0(GND_net), 
            .I1(n2531), .I2(VCC_net), .I3(n44207), .O(n2598)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1704_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_632_6 (.CI(n43976), 
            .I0(n930), .I1(GND_net), .CO(n43977));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1704_5 (.CI(n44207), 
            .I0(n2531), .I1(VCC_net), .CO(n44208));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1704_4_lut (.I0(GND_net), 
            .I1(n2532), .I2(GND_net), .I3(n44206), .O(n2599)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1704_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_632_5_lut (.I0(GND_net), 
            .I1(n931), .I2(VCC_net), .I3(n43975), .O(n998)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_632_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1704_4 (.CI(n44206), 
            .I0(n2532), .I1(GND_net), .CO(n44207));
    SB_LUT4 i15702_3_lut (.I0(\neo_pixel_transmitter.t0 [31]), .I1(timer[31]), 
            .I2(n47790), .I3(GND_net), .O(n29782));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15702_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15703_3_lut (.I0(\neo_pixel_transmitter.t0 [30]), .I1(timer[30]), 
            .I2(n47790), .I3(GND_net), .O(n29783));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15703_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_175_18_lut (.I0(GND_net), .I1(delay_counter[16]), .I2(GND_net), 
            .I3(n43625), .O(n1547)) /* synthesis syn_instantiated=1 */ ;
    defparam add_175_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15704_3_lut (.I0(\neo_pixel_transmitter.t0 [29]), .I1(timer[29]), 
            .I2(n47790), .I3(GND_net), .O(n29784));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15704_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15972_3_lut (.I0(\data_out_frame[12] [5]), .I1(setpoint[21]), 
            .I2(n24210), .I3(GND_net), .O(n30052));   // verilog/coms.v(128[12] 303[6])
    defparam i15972_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1808 (.I0(n3108), .I1(n51952), .I2(n51702), .I3(n3109), 
            .O(n51706));
    defparam i1_4_lut_adj_1808.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1704_3_lut (.I0(GND_net), 
            .I1(n2533), .I2(VCC_net), .I3(n44205), .O(n2600)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1704_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i40734_4_lut (.I0(n3106), .I1(n3105), .I2(n3107), .I3(n51706), 
            .O(n3138));
    defparam i40734_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i15973_3_lut (.I0(\data_out_frame[12] [4]), .I1(setpoint[20]), 
            .I2(n24210), .I3(GND_net), .O(n30053));   // verilog/coms.v(128[12] 303[6])
    defparam i15973_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15705_3_lut (.I0(\neo_pixel_transmitter.t0 [28]), .I1(timer[28]), 
            .I2(n47790), .I3(GND_net), .O(n29785));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15705_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15974_3_lut (.I0(\data_out_frame[12] [3]), .I1(setpoint[19]), 
            .I2(n24210), .I3(GND_net), .O(n30054));   // verilog/coms.v(128[12] 303[6])
    defparam i15974_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1976_3_lut (.I0(n2909), 
            .I1(n2976), .I2(n2940), .I3(GND_net), .O(n3008));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1976_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15975_3_lut (.I0(\data_out_frame[12] [2]), .I1(setpoint[18]), 
            .I2(n24210), .I3(GND_net), .O(n30055));   // verilog/coms.v(128[12] 303[6])
    defparam i15975_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_632_5 (.CI(n43975), 
            .I0(n931), .I1(VCC_net), .CO(n43976));
    SB_LUT4 i15976_3_lut (.I0(\data_out_frame[12] [1]), .I1(setpoint[17]), 
            .I2(n24210), .I3(GND_net), .O(n30056));   // verilog/coms.v(128[12] 303[6])
    defparam i15976_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1704_3 (.CI(n44205), 
            .I0(n2533), .I1(VCC_net), .CO(n44206));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1704_2_lut (.I0(GND_net), 
            .I1(n536), .I2(GND_net), .I3(VCC_net), .O(n2601)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1704_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15977_3_lut (.I0(\data_out_frame[12] [0]), .I1(setpoint[16]), 
            .I2(n24210), .I3(GND_net), .O(n30057));   // verilog/coms.v(128[12] 303[6])
    defparam i15977_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_175_18 (.CI(n43625), .I0(delay_counter[16]), .I1(GND_net), 
            .CO(n43626));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1704_2 (.CI(VCC_net), 
            .I0(n536), .I1(GND_net), .CO(n44205));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1637_24_lut (.I0(n56171), 
            .I1(n2412), .I2(VCC_net), .I3(n44204), .O(n2511)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1637_24_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i15708_3_lut (.I0(\neo_pixel_transmitter.t0 [27]), .I1(timer[27]), 
            .I2(n47790), .I3(GND_net), .O(n29788));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15708_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15709_3_lut (.I0(\neo_pixel_transmitter.t0 [26]), .I1(timer[26]), 
            .I2(n47790), .I3(GND_net), .O(n29789));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15709_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1975_3_lut (.I0(n2908), 
            .I1(n2975), .I2(n2940), .I3(GND_net), .O(n3007));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1975_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1979_3_lut (.I0(n2912), 
            .I1(n2979), .I2(n2940), .I3(GND_net), .O(n3011));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1979_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1637_23_lut (.I0(GND_net), 
            .I1(n2413), .I2(VCC_net), .I3(n44203), .O(n2480)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1637_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15710_3_lut (.I0(\neo_pixel_transmitter.t0 [25]), .I1(timer[25]), 
            .I2(n47790), .I3(GND_net), .O(n29790));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15710_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15711_3_lut (.I0(\neo_pixel_transmitter.t0 [24]), .I1(timer[24]), 
            .I2(n47790), .I3(GND_net), .O(n29791));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15711_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15978_3_lut (.I0(\data_out_frame[11] [7]), .I1(encoder1_position_scaled[7]), 
            .I2(n24210), .I3(GND_net), .O(n30058));   // verilog/coms.v(128[12] 303[6])
    defparam i15978_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15712_3_lut (.I0(\neo_pixel_transmitter.t0 [23]), .I1(timer[23]), 
            .I2(n47790), .I3(GND_net), .O(n29792));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15712_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1978_3_lut (.I0(n2911), 
            .I1(n2978), .I2(n2940), .I3(GND_net), .O(n3010));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1978_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15979_4_lut (.I0(CS_MISO_c), .I1(data_adj_5711[10]), .I2(n5), 
            .I3(n27198), .O(n30059));   // verilog/tli4970.v(35[10] 68[6])
    defparam i15979_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_632_4_lut (.I0(GND_net), 
            .I1(n932), .I2(GND_net), .I3(n43974), .O(n999)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_632_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1977_3_lut (.I0(n2910), 
            .I1(n2977), .I2(n2940), .I3(GND_net), .O(n3009));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1977_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1982_3_lut (.I0(n2915), 
            .I1(n2982), .I2(n2940), .I3(GND_net), .O(n3014));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1982_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1981_3_lut (.I0(n2914), 
            .I1(n2981), .I2(n2940), .I3(GND_net), .O(n3013));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1981_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15713_3_lut (.I0(\neo_pixel_transmitter.t0 [22]), .I1(timer[22]), 
            .I2(n47790), .I3(GND_net), .O(n29793));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15713_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_175_17_lut (.I0(GND_net), .I1(delay_counter[15]), .I2(GND_net), 
            .I3(n43624), .O(n1548)) /* synthesis syn_instantiated=1 */ ;
    defparam add_175_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_632_4 (.CI(n43974), 
            .I0(n932), .I1(GND_net), .CO(n43975));
    SB_CARRY add_175_17 (.CI(n43624), .I0(delay_counter[15]), .I1(GND_net), 
            .CO(n43625));
    SB_LUT4 i15714_3_lut (.I0(\neo_pixel_transmitter.t0 [21]), .I1(timer[21]), 
            .I2(n47790), .I3(GND_net), .O(n29794));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15714_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1980_3_lut (.I0(n2913), 
            .I1(n2980), .I2(n2940), .I3(GND_net), .O(n3012));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1980_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1995_3_lut (.I0(n2928), 
            .I1(n2995), .I2(n2940), .I3(GND_net), .O(n3027));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1995_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15715_3_lut (.I0(\neo_pixel_transmitter.t0 [20]), .I1(timer[20]), 
            .I2(n47790), .I3(GND_net), .O(n29795));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15715_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1991_3_lut (.I0(n2924), 
            .I1(n2991), .I2(n2940), .I3(GND_net), .O(n3023));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1991_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15716_3_lut (.I0(\neo_pixel_transmitter.t0 [19]), .I1(timer[19]), 
            .I2(n47790), .I3(GND_net), .O(n29796));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15716_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15717_3_lut (.I0(\neo_pixel_transmitter.t0 [18]), .I1(timer[18]), 
            .I2(n47790), .I3(GND_net), .O(n29797));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15717_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1987_3_lut (.I0(n2920), 
            .I1(n2987), .I2(n2940), .I3(GND_net), .O(n3019));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1987_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1809 (.I0(n7974), .I1(n21005), .I2(data_ready), 
            .I3(\ID_READOUT_FSM.state [0]), .O(n49720));
    defparam i1_4_lut_adj_1809.LUT_INIT = 16'heaee;
    SB_LUT4 i15718_3_lut (.I0(\neo_pixel_transmitter.t0 [17]), .I1(timer[17]), 
            .I2(n47790), .I3(GND_net), .O(n29798));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15718_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1984_3_lut (.I0(n2917), 
            .I1(n2984), .I2(n2940), .I3(GND_net), .O(n3016));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1984_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i2_4_lut_adj_1810 (.I0(\ID_READOUT_FSM.state [0]), .I1(n36436), 
            .I2(\ID_READOUT_FSM.state [1]), .I3(n49720), .O(n28885));
    defparam i2_4_lut_adj_1810.LUT_INIT = 16'h4c00;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1983_3_lut (.I0(n2916), 
            .I1(n2983), .I2(n2940), .I3(GND_net), .O(n3015));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1983_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15776_3_lut (.I0(n28885), .I1(\ID_READOUT_FSM.state [0]), .I2(n7974), 
            .I3(GND_net), .O(n29856));   // verilog/TinyFPGA_B.v(368[10] 396[6])
    defparam i15776_3_lut.LUT_INIT = 16'h4646;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1999_3_lut (.I0(n2932), 
            .I1(n2999), .I2(n2940), .I3(GND_net), .O(n3031));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1999_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15719_3_lut (.I0(\neo_pixel_transmitter.t0 [16]), .I1(timer[16]), 
            .I2(n47790), .I3(GND_net), .O(n29799));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15719_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1811 (.I0(n36659), .I1(n49919), .I2(state_adj_5705[0]), 
            .I3(read), .O(n48558));   // verilog/eeprom.v(26[8] 58[4])
    defparam i1_4_lut_adj_1811.LUT_INIT = 16'h8280;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_632_3_lut (.I0(GND_net), 
            .I1(n933), .I2(VCC_net), .I3(n43973), .O(n1000)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_632_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1637_23 (.CI(n44203), 
            .I0(n2413), .I1(VCC_net), .CO(n44204));
    SB_LUT4 i15720_3_lut (.I0(\neo_pixel_transmitter.t0 [15]), .I1(timer[15]), 
            .I2(n47790), .I3(GND_net), .O(n29800));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15720_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1998_3_lut (.I0(n2931), 
            .I1(n2998), .I2(n2940), .I3(GND_net), .O(n3030));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1998_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15721_3_lut (.I0(\neo_pixel_transmitter.t0 [14]), .I1(timer[14]), 
            .I2(n47790), .I3(GND_net), .O(n29801));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15721_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1997_3_lut (.I0(n2930), 
            .I1(n2997), .I2(n2940), .I3(GND_net), .O(n3029));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1997_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1986_3_lut (.I0(n2919), 
            .I1(n2986), .I2(n2940), .I3(GND_net), .O(n3018));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1986_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1985_3_lut (.I0(n2918), 
            .I1(n2985), .I2(n2940), .I3(GND_net), .O(n3017));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1985_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15722_3_lut (.I0(\neo_pixel_transmitter.t0 [13]), .I1(timer[13]), 
            .I2(n47790), .I3(GND_net), .O(n29802));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15722_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15765_3_lut (.I0(n29282), .I1(r_Bit_Index[0]), .I2(n28852), 
            .I3(GND_net), .O(n29845));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i15765_3_lut.LUT_INIT = 16'h1414;
    SB_LUT4 i15762_3_lut (.I0(n29280), .I1(r_Bit_Index_adj_5725[0]), .I2(n28848), 
            .I3(GND_net), .O(n29842));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i15762_3_lut.LUT_INIT = 16'h1414;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1989_3_lut (.I0(n2922), 
            .I1(n2989), .I2(n2940), .I3(GND_net), .O(n3021));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1989_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15723_3_lut (.I0(\neo_pixel_transmitter.t0 [12]), .I1(timer[12]), 
            .I2(n47790), .I3(GND_net), .O(n29803));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15723_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15986_4_lut (.I0(CS_MISO_c), .I1(data_adj_5711[11]), .I2(n36554), 
            .I3(n27198), .O(n30066));   // verilog/tli4970.v(35[10] 68[6])
    defparam i15986_4_lut.LUT_INIT = 16'hccac;
    SB_LUT4 i15724_3_lut (.I0(\neo_pixel_transmitter.t0 [11]), .I1(timer[11]), 
            .I2(n47790), .I3(GND_net), .O(n29804));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15724_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1990_3_lut (.I0(n2923), 
            .I1(n2990), .I2(n2940), .I3(GND_net), .O(n3022));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1990_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1988_3_lut (.I0(n2921), 
            .I1(n2988), .I2(n2940), .I3(GND_net), .O(n3020));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1988_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15725_3_lut (.I0(\neo_pixel_transmitter.t0 [10]), .I1(timer[10]), 
            .I2(n47790), .I3(GND_net), .O(n29805));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15725_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i2001_3_lut (.I0(n540), .I1(n3001), 
            .I2(n2940), .I3(GND_net), .O(n3033));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i2001_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i2000_3_lut (.I0(n2933), 
            .I1(n3000), .I2(n2940), .I3(GND_net), .O(n3032));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i2000_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_mux_3_i4_3_lut (.I0(encoder0_position_scaled_23__N_327[3]), 
            .I1(n30), .I2(encoder0_position_scaled_23__N_327[31]), .I3(GND_net), 
            .O(n541));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_mux_3_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1996_3_lut (.I0(n2929), 
            .I1(n2996), .I2(n2940), .I3(GND_net), .O(n3028));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1996_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15726_3_lut (.I0(\neo_pixel_transmitter.t0 [9]), .I1(timer[9]), 
            .I2(n47790), .I3(GND_net), .O(n29806));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15726_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1993_3_lut (.I0(n2926), 
            .I1(n2993), .I2(n2940), .I3(GND_net), .O(n3025));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1993_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1637_22_lut (.I0(GND_net), 
            .I1(n2414), .I2(VCC_net), .I3(n44202), .O(n2481)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1637_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15727_3_lut (.I0(\neo_pixel_transmitter.t0 [8]), .I1(timer[8]), 
            .I2(n47790), .I3(GND_net), .O(n29807));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15727_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15728_3_lut (.I0(\neo_pixel_transmitter.t0 [7]), .I1(timer[7]), 
            .I2(n47790), .I3(GND_net), .O(n29808));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15728_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15729_3_lut (.I0(\neo_pixel_transmitter.t0 [6]), .I1(timer[6]), 
            .I2(n47790), .I3(GND_net), .O(n29809));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15729_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1637_22 (.CI(n44202), 
            .I0(n2414), .I1(VCC_net), .CO(n44203));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1637_21_lut (.I0(GND_net), 
            .I1(n2415), .I2(VCC_net), .I3(n44201), .O(n2482)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1637_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1637_21 (.CI(n44201), 
            .I0(n2415), .I1(VCC_net), .CO(n44202));
    SB_LUT4 i15730_3_lut (.I0(\neo_pixel_transmitter.t0 [5]), .I1(timer[5]), 
            .I2(n47790), .I3(GND_net), .O(n29810));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15730_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_632_3 (.CI(n43973), 
            .I0(n933), .I1(VCC_net), .CO(n43974));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1994_3_lut (.I0(n2927), 
            .I1(n2994), .I2(n2940), .I3(GND_net), .O(n3026));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1994_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_632_2_lut (.I0(GND_net), 
            .I1(n934), .I2(GND_net), .I3(VCC_net), .O(n1001)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_632_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15731_3_lut (.I0(\neo_pixel_transmitter.t0 [4]), .I1(timer[4]), 
            .I2(n47790), .I3(GND_net), .O(n29811));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15731_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1992_3_lut (.I0(n2925), 
            .I1(n2992), .I2(n2940), .I3(GND_net), .O(n3024));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1992_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_632_2 (.CI(VCC_net), 
            .I0(n934), .I1(GND_net), .CO(n43973));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_565_8_lut (.I0(n861), 
            .I1(n828), .I2(VCC_net), .I3(n43972), .O(n927)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_565_8_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i15732_3_lut (.I0(\neo_pixel_transmitter.t0 [3]), .I1(timer[3]), 
            .I2(n47790), .I3(GND_net), .O(n29812));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15732_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1637_20_lut (.I0(GND_net), 
            .I1(n2416), .I2(VCC_net), .I3(n44200), .O(n2483)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1637_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_565_7_lut (.I0(GND_net), 
            .I1(n829), .I2(GND_net), .I3(n43971), .O(n896)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_565_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_565_7 (.CI(n43971), 
            .I0(n829), .I1(GND_net), .CO(n43972));
    SB_LUT4 i40764_1_lut (.I0(n3039), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n56595));
    defparam i40764_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_565_6_lut (.I0(GND_net), 
            .I1(n830), .I2(GND_net), .I3(n43970), .O(n897)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_565_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1637_20 (.CI(n44200), 
            .I0(n2416), .I1(VCC_net), .CO(n44201));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_565_6 (.CI(n43970), 
            .I0(n830), .I1(GND_net), .CO(n43971));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1637_19_lut (.I0(GND_net), 
            .I1(n2417), .I2(VCC_net), .I3(n44199), .O(n2484)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1637_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15733_3_lut (.I0(\neo_pixel_transmitter.t0 [2]), .I1(timer[2]), 
            .I2(n47790), .I3(GND_net), .O(n29813));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15733_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_565_5_lut (.I0(GND_net), 
            .I1(n831), .I2(VCC_net), .I3(n43969), .O(n898)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_565_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_3_lut_adj_1812 (.I0(n3020), .I1(n3022), .I2(n3021), .I3(GND_net), 
            .O(n52142));
    defparam i1_3_lut_adj_1812.LUT_INIT = 16'hfefe;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_565_5 (.CI(n43969), 
            .I0(n831), .I1(VCC_net), .CO(n43970));
    SB_LUT4 i1_4_lut_adj_1813 (.I0(n3024), .I1(n3026), .I2(n3025), .I3(n3028), 
            .O(n52144));
    defparam i1_4_lut_adj_1813.LUT_INIT = 16'hfffe;
    SB_LUT4 i15734_3_lut (.I0(\neo_pixel_transmitter.t0 [1]), .I1(timer[1]), 
            .I2(n47790), .I3(GND_net), .O(n29814));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15734_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1637_19 (.CI(n44199), 
            .I0(n2417), .I1(VCC_net), .CO(n44200));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1637_18_lut (.I0(GND_net), 
            .I1(n2418), .I2(VCC_net), .I3(n44198), .O(n2485)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1637_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15987_4_lut (.I0(CS_MISO_c), .I1(data_adj_5711[12]), .I2(n36528), 
            .I3(n27232), .O(n30067));   // verilog/tli4970.v(35[10] 68[6])
    defparam i15987_4_lut.LUT_INIT = 16'hccac;
    SB_LUT4 add_175_16_lut (.I0(GND_net), .I1(delay_counter[14]), .I2(GND_net), 
            .I3(n43623), .O(n1549)) /* synthesis syn_instantiated=1 */ ;
    defparam add_175_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1637_18 (.CI(n44198), 
            .I0(n2418), .I1(VCC_net), .CO(n44199));
    SB_LUT4 i15735_3_lut (.I0(ID[7]), .I1(data[7]), .I2(n51509), .I3(GND_net), 
            .O(n29815));   // verilog/TinyFPGA_B.v(368[10] 396[6])
    defparam i15735_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1637_17_lut (.I0(GND_net), 
            .I1(n2419), .I2(VCC_net), .I3(n44197), .O(n2486)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1637_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1637_17 (.CI(n44197), 
            .I0(n2419), .I1(VCC_net), .CO(n44198));
    SB_LUT4 i23213_3_lut (.I0(n541), .I1(n3032), .I2(n3033), .I3(GND_net), 
            .O(n37302));
    defparam i23213_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i1_4_lut_adj_1814 (.I0(n3029), .I1(n37302), .I2(n3030), .I3(n3031), 
            .O(n50144));
    defparam i1_4_lut_adj_1814.LUT_INIT = 16'ha080;
    SB_LUT4 i1_4_lut_adj_1815 (.I0(n3017), .I1(n52144), .I2(n52142), .I3(n3018), 
            .O(n52150));
    defparam i1_4_lut_adj_1815.LUT_INIT = 16'hfffe;
    SB_LUT4 i15736_3_lut (.I0(ID[6]), .I1(data[6]), .I2(n51509), .I3(GND_net), 
            .O(n29816));   // verilog/TinyFPGA_B.v(368[10] 396[6])
    defparam i15736_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15737_3_lut (.I0(ID[5]), .I1(data[5]), .I2(n51509), .I3(GND_net), 
            .O(n29817));   // verilog/TinyFPGA_B.v(368[10] 396[6])
    defparam i15737_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1816 (.I0(n3019), .I1(n50144), .I2(n3023), .I3(n3027), 
            .O(n51223));
    defparam i1_4_lut_adj_1816.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1817 (.I0(n51223), .I1(n3015), .I2(n3016), .I3(n52150), 
            .O(n52156));
    defparam i1_4_lut_adj_1817.LUT_INIT = 16'hfffe;
    SB_LUT4 i15738_3_lut (.I0(ID[4]), .I1(data[4]), .I2(n51509), .I3(GND_net), 
            .O(n29818));   // verilog/TinyFPGA_B.v(368[10] 396[6])
    defparam i15738_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15739_3_lut (.I0(ID[3]), .I1(data[3]), .I2(n51509), .I3(GND_net), 
            .O(n29819));   // verilog/TinyFPGA_B.v(368[10] 396[6])
    defparam i15739_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1818 (.I0(n3012), .I1(n3013), .I2(n52156), .I3(n3014), 
            .O(n52162));
    defparam i1_4_lut_adj_1818.LUT_INIT = 16'hfffe;
    SB_LUT4 i15740_3_lut (.I0(ID[2]), .I1(data[2]), .I2(n51509), .I3(GND_net), 
            .O(n29820));   // verilog/TinyFPGA_B.v(368[10] 396[6])
    defparam i15740_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1819 (.I0(n3009), .I1(n3010), .I2(n3011), .I3(n52162), 
            .O(n52168));
    defparam i1_4_lut_adj_1819.LUT_INIT = 16'hfffe;
    SB_LUT4 i40767_4_lut (.I0(n3007), .I1(n3006), .I2(n3008), .I3(n52168), 
            .O(n3039));
    defparam i40767_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i2_3_lut (.I0(data_ready), .I1(\ID_READOUT_FSM.state [1]), .I2(\ID_READOUT_FSM.state [0]), 
            .I3(GND_net), .O(n51509));
    defparam i2_3_lut.LUT_INIT = 16'hdfdf;
    SB_LUT4 i15741_3_lut (.I0(ID[1]), .I1(data[1]), .I2(n51509), .I3(GND_net), 
            .O(n29821));   // verilog/TinyFPGA_B.v(368[10] 396[6])
    defparam i15741_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15743_4_lut (.I0(CS_MISO_c), .I1(data_adj_5711[2]), .I2(n6_adj_5556), 
            .I3(n27258), .O(n29823));   // verilog/tli4970.v(35[10] 68[6])
    defparam i15743_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1909_3_lut (.I0(n2810), 
            .I1(n2877), .I2(n2841), .I3(GND_net), .O(n2909));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1909_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1908_3_lut (.I0(n2809), 
            .I1(n2876), .I2(n2841), .I3(GND_net), .O(n2908));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1908_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15744_3_lut (.I0(\data_out_frame[25] [7]), .I1(neopxl_color[7]), 
            .I2(n24210), .I3(GND_net), .O(n29824));   // verilog/coms.v(128[12] 303[6])
    defparam i15744_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1912_3_lut (.I0(n2813), 
            .I1(n2880), .I2(n2841), .I3(GND_net), .O(n2912));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1912_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1911_3_lut (.I0(n2812), 
            .I1(n2879), .I2(n2841), .I3(GND_net), .O(n2911));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1911_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1910_3_lut (.I0(n2811), 
            .I1(n2878), .I2(n2841), .I3(GND_net), .O(n2910));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1910_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15745_3_lut (.I0(\data_out_frame[25] [6]), .I1(neopxl_color[6]), 
            .I2(n24210), .I3(GND_net), .O(n29825));   // verilog/coms.v(128[12] 303[6])
    defparam i15745_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15746_3_lut (.I0(\data_out_frame[25] [5]), .I1(neopxl_color[5]), 
            .I2(n24210), .I3(GND_net), .O(n29826));   // verilog/coms.v(128[12] 303[6])
    defparam i15746_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1915_3_lut (.I0(n2816), 
            .I1(n2883), .I2(n2841), .I3(GND_net), .O(n2915));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1915_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15747_3_lut (.I0(\data_out_frame[25] [4]), .I1(neopxl_color[4]), 
            .I2(n24210), .I3(GND_net), .O(n29827));   // verilog/coms.v(128[12] 303[6])
    defparam i15747_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15750_3_lut (.I0(\data_out_frame[25] [3]), .I1(neopxl_color[3]), 
            .I2(n24210), .I3(GND_net), .O(n29830));   // verilog/coms.v(128[12] 303[6])
    defparam i15750_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15338_3_lut (.I0(\data_out_frame[7] [5]), .I1(encoder0_position_scaled[13]), 
            .I2(n24210), .I3(GND_net), .O(n29418));   // verilog/coms.v(128[12] 303[6])
    defparam i15338_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34001_3_lut (.I0(n3_adj_5496), .I1(n8582), .I2(n49748), .I3(GND_net), 
            .O(n49749));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam i34001_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34002_rep_60_3_lut (.I0(encoder0_position_scaled_23__N_327[30]), 
            .I1(n896), .I2(n861), .I3(GND_net), .O(n53127));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam i34002_rep_60_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1914_3_lut (.I0(n2815), 
            .I1(n2882), .I2(n2841), .I3(GND_net), .O(n2914));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1914_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15751_3_lut (.I0(\data_out_frame[25] [2]), .I1(neopxl_color[2]), 
            .I2(n24210), .I3(GND_net), .O(n29831));   // verilog/coms.v(128[12] 303[6])
    defparam i15751_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15752_3_lut (.I0(\data_out_frame[25] [1]), .I1(neopxl_color[1]), 
            .I2(n24210), .I3(GND_net), .O(n29832));   // verilog/coms.v(128[12] 303[6])
    defparam i15752_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15753_3_lut (.I0(\data_out_frame[25] [0]), .I1(neopxl_color[0]), 
            .I2(n24210), .I3(GND_net), .O(n29833));   // verilog/coms.v(128[12] 303[6])
    defparam i15753_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15754_3_lut (.I0(\data_out_frame[24] [7]), .I1(neopxl_color[15]), 
            .I2(n24210), .I3(GND_net), .O(n29834));   // verilog/coms.v(128[12] 303[6])
    defparam i15754_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15755_4_lut (.I0(state_7__N_4306[3]), .I1(data[0]), .I2(n10_adj_5610), 
            .I3(n27238), .O(n29835));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i15755_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1913_3_lut (.I0(n2814), 
            .I1(n2881), .I2(n2841), .I3(GND_net), .O(n2913));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1913_3_lut.LUT_INIT = 16'hacac;
    SB_DFF dti_counter_2279__i7 (.Q(dti_counter[7]), .C(clk16MHz), .D(n48));   // verilog/TinyFPGA_B.v(174[23:37])
    SB_DFF dti_counter_2279__i6 (.Q(dti_counter[6]), .C(clk16MHz), .D(n49));   // verilog/TinyFPGA_B.v(174[23:37])
    SB_DFF dti_counter_2279__i5 (.Q(dti_counter[5]), .C(clk16MHz), .D(n50));   // verilog/TinyFPGA_B.v(174[23:37])
    SB_DFF dti_counter_2279__i4 (.Q(dti_counter[4]), .C(clk16MHz), .D(n51));   // verilog/TinyFPGA_B.v(174[23:37])
    SB_DFF dti_counter_2279__i3 (.Q(dti_counter[3]), .C(clk16MHz), .D(n52));   // verilog/TinyFPGA_B.v(174[23:37])
    SB_DFF dti_counter_2279__i2 (.Q(dti_counter[2]), .C(clk16MHz), .D(n53));   // verilog/TinyFPGA_B.v(174[23:37])
    SB_DFF dti_counter_2279__i1 (.Q(dti_counter[1]), .C(clk16MHz), .D(n54));   // verilog/TinyFPGA_B.v(174[23:37])
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_565_4_lut (.I0(GND_net), 
            .I1(n832), .I2(GND_net), .I3(n43968), .O(n899)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_565_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1918_3_lut (.I0(n2819), 
            .I1(n2886), .I2(n2841), .I3(GND_net), .O(n2918));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1918_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15758_4_lut (.I0(CS_MISO_c), .I1(data_adj_5711[3]), .I2(n6_adj_5556), 
            .I3(n27264), .O(n29838));   // verilog/tli4970.v(35[10] 68[6])
    defparam i15758_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1917_3_lut (.I0(n2818), 
            .I1(n2885), .I2(n2841), .I3(GND_net), .O(n2917));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1917_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1933_3_lut (.I0(n539), .I1(n2901), 
            .I2(n2841), .I3(GND_net), .O(n2933));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1933_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15759_4_lut (.I0(CS_MISO_c), .I1(data_adj_5711[4]), .I2(n6_adj_5523), 
            .I3(n27232), .O(n29839));   // verilog/tli4970.v(35[10] 68[6])
    defparam i15759_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1637_16_lut (.I0(GND_net), 
            .I1(n2420), .I2(VCC_net), .I3(n44196), .O(n2487)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1637_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_175_16 (.CI(n43623), .I0(delay_counter[14]), .I1(GND_net), 
            .CO(n43624));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1932_3_lut (.I0(n2833), 
            .I1(n2900), .I2(n2841), .I3(GND_net), .O(n2932));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1932_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_565_4 (.CI(n43968), 
            .I0(n832), .I1(GND_net), .CO(n43969));
    SB_LUT4 i15769_4_lut (.I0(r_Rx_Data), .I1(rx_data[0]), .I2(n4_adj_5443), 
            .I3(n27208), .O(n29849));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i15769_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_unary_minus_2_inv_0_i10_1_lut (.I0(encoder0_position_scaled_23__N_327[9]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n24_adj_5633));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_unary_minus_2_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1637_16 (.CI(n44196), 
            .I0(n2420), .I1(VCC_net), .CO(n44197));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1637_15_lut (.I0(GND_net), 
            .I1(n2421), .I2(VCC_net), .I3(n44195), .O(n2488)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1637_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15770_4_lut (.I0(CS_MISO_c), .I1(data_adj_5711[0]), .I2(n7_adj_5577), 
            .I3(state_7__N_4499), .O(n29850));   // verilog/tli4970.v(35[10] 68[6])
    defparam i15770_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 add_263_12_lut (.I0(GND_net), .I1(encoder1_position[13]), .I2(GND_net), 
            .I3(n43544), .O(encoder1_position_scaled_23__N_75[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_263_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_565_3_lut (.I0(GND_net), 
            .I1(n833), .I2(VCC_net), .I3(n43967), .O(n900)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_565_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_175_15_lut (.I0(GND_net), .I1(delay_counter[13]), .I2(GND_net), 
            .I3(n43622), .O(n1550)) /* synthesis syn_instantiated=1 */ ;
    defparam add_175_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_565_3 (.CI(n43967), 
            .I0(n833), .I1(VCC_net), .CO(n43968));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1637_15 (.CI(n44195), 
            .I0(n2421), .I1(VCC_net), .CO(n44196));
    SB_LUT4 i15780_4_lut (.I0(r_Rx_Data), .I1(rx_data[7]), .I2(n36556), 
            .I3(n27203), .O(n29860));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i15780_4_lut.LUT_INIT = 16'hccac;
    SB_CARRY add_261_11 (.CI(n43566), .I0(duty[12]), .I1(n56614), .CO(n43567));
    SB_LUT4 i15781_3_lut (.I0(\data_out_frame[24] [6]), .I1(neopxl_color[14]), 
            .I2(n24210), .I3(GND_net), .O(n29861));   // verilog/coms.v(128[12] 303[6])
    defparam i15781_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1931_3_lut (.I0(n2832), 
            .I1(n2899), .I2(n2841), .I3(GND_net), .O(n2931));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1931_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15782_3_lut (.I0(\data_out_frame[24] [5]), .I1(neopxl_color[13]), 
            .I2(n24210), .I3(GND_net), .O(n29862));   // verilog/coms.v(128[12] 303[6])
    defparam i15782_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1637_14_lut (.I0(GND_net), 
            .I1(n2422), .I2(VCC_net), .I3(n44194), .O(n2489)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1637_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_mux_3_i5_3_lut (.I0(encoder0_position_scaled_23__N_327[4]), 
            .I1(n29), .I2(encoder0_position_scaled_23__N_327[31]), .I3(GND_net), 
            .O(n540));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_mux_3_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15783_3_lut (.I0(\data_out_frame[24] [4]), .I1(neopxl_color[12]), 
            .I2(n24210), .I3(GND_net), .O(n29863));   // verilog/coms.v(128[12] 303[6])
    defparam i15783_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1924_3_lut (.I0(n2825), 
            .I1(n2892), .I2(n2841), .I3(GND_net), .O(n2924));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1924_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i1_1_lut (.I0(encoder1_position_scaled[0]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n25_adj_5498));   // verilog/TinyFPGA_B.v(324[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_565_2_lut (.I0(GND_net), 
            .I1(n834), .I2(GND_net), .I3(VCC_net), .O(n901)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_565_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i635_3_lut (.I0(n928), .I1(n995), 
            .I2(n960), .I3(GND_net), .O(n1027));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i635_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15784_3_lut (.I0(\data_out_frame[24] [3]), .I1(neopxl_color[11]), 
            .I2(n24210), .I3(GND_net), .O(n29864));   // verilog/coms.v(128[12] 303[6])
    defparam i15784_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15785_3_lut (.I0(\data_out_frame[24] [2]), .I1(neopxl_color[10]), 
            .I2(n24210), .I3(GND_net), .O(n29865));   // verilog/coms.v(128[12] 303[6])
    defparam i15785_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1921_3_lut (.I0(n2822), 
            .I1(n2889), .I2(n2841), .I3(GND_net), .O(n2921));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1921_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15786_3_lut (.I0(\data_out_frame[24] [1]), .I1(neopxl_color[9]), 
            .I2(n24210), .I3(GND_net), .O(n29866));   // verilog/coms.v(128[12] 303[6])
    defparam i15786_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_565_2 (.CI(VCC_net), 
            .I0(n834), .I1(GND_net), .CO(n43967));
    SB_LUT4 i15787_3_lut (.I0(\data_out_frame[24] [0]), .I1(neopxl_color[8]), 
            .I2(n24210), .I3(GND_net), .O(n29867));   // verilog/coms.v(128[12] 303[6])
    defparam i15787_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_175_15 (.CI(n43622), .I0(delay_counter[13]), .I1(GND_net), 
            .CO(n43623));
    SB_LUT4 i15788_3_lut (.I0(\data_out_frame[23] [7]), .I1(neopxl_color[23]), 
            .I2(n24210), .I3(GND_net), .O(n29868));   // verilog/coms.v(128[12] 303[6])
    defparam i15788_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1920_3_lut (.I0(n2821), 
            .I1(n2888), .I2(n2841), .I3(GND_net), .O(n2920));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1920_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1926_3_lut (.I0(n2827), 
            .I1(n2894), .I2(n2841), .I3(GND_net), .O(n2926));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1926_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i702_3_lut (.I0(n1027), .I1(n1094), 
            .I2(n1059), .I3(GND_net), .O(n1126));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i702_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i2_1_lut (.I0(encoder1_position_scaled[1]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n24_adj_5499));   // verilog/TinyFPGA_B.v(324[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i40369_1_lut (.I0(n2346), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n56200));
    defparam i40369_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i769_rep_54_3_lut (.I0(n1126), 
            .I1(n1193), .I2(n1158), .I3(GND_net), .O(n1225));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i769_rep_54_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_mux_3_i27_3_lut (.I0(encoder0_position_scaled_23__N_327[26]), 
            .I1(n7_adj_5492), .I2(encoder0_position_scaled_23__N_327[31]), 
            .I3(GND_net), .O(n407));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_mux_3_i27_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15789_4_lut (.I0(CS_MISO_c), .I1(data_adj_5711[5]), .I2(n6_adj_5523), 
            .I3(n27271), .O(n29869));   // verilog/tli4970.v(35[10] 68[6])
    defparam i15789_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 add_2747_7_lut (.I0(GND_net), .I1(n621), .I2(GND_net), .I3(n43966), 
            .O(n8581)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2747_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2747_6_lut (.I0(GND_net), .I1(n622), .I2(GND_net), .I3(n43965), 
            .O(n8582)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2747_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1637_14 (.CI(n44194), 
            .I0(n2422), .I1(VCC_net), .CO(n44195));
    SB_CARRY add_2747_6 (.CI(n43965), .I0(n622), .I1(GND_net), .CO(n43966));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1637_13_lut (.I0(GND_net), 
            .I1(n2423), .I2(VCC_net), .I3(n44193), .O(n2490)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1637_13_lut.LUT_INIT = 16'hC33C;
    SB_IO RX_pad (.PACKAGE_PIN(RX), .OUTPUT_ENABLE(VCC_net), .D_IN_0(RX_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam RX_pad.PIN_TYPE = 6'b000001;
    defparam RX_pad.PULLUP = 1'b0;
    defparam RX_pad.NEG_TRIGGER = 1'b0;
    defparam RX_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO ENCODER1_B_pad (.PACKAGE_PIN(ENCODER1_B), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(ENCODER1_B_N));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ENCODER1_B_pad.PIN_TYPE = 6'b000001;
    defparam ENCODER1_B_pad.PULLUP = 1'b0;
    defparam ENCODER1_B_pad.NEG_TRIGGER = 1'b0;
    defparam ENCODER1_B_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO ENCODER1_A_pad (.PACKAGE_PIN(ENCODER1_A), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(ENCODER1_A_N));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ENCODER1_A_pad.PIN_TYPE = 6'b000001;
    defparam ENCODER1_A_pad.PULLUP = 1'b0;
    defparam ENCODER1_A_pad.NEG_TRIGGER = 1'b0;
    defparam ENCODER1_A_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO ENCODER0_B_pad (.PACKAGE_PIN(ENCODER0_B), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(ENCODER0_B_N));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ENCODER0_B_pad.PIN_TYPE = 6'b000001;
    defparam ENCODER0_B_pad.PULLUP = 1'b0;
    defparam ENCODER0_B_pad.NEG_TRIGGER = 1'b0;
    defparam ENCODER0_B_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO ENCODER0_A_pad (.PACKAGE_PIN(ENCODER0_A), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(ENCODER0_A_N));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ENCODER0_A_pad.PIN_TYPE = 6'b000001;
    defparam ENCODER0_A_pad.PULLUP = 1'b0;
    defparam ENCODER0_A_pad.NEG_TRIGGER = 1'b0;
    defparam ENCODER0_A_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO INHA_pad (.PACKAGE_PIN(INHA), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INHA_c_0));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INHA_pad.PIN_TYPE = 6'b011001;
    defparam INHA_pad.PULLUP = 1'b0;
    defparam INHA_pad.NEG_TRIGGER = 1'b0;
    defparam INHA_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO INLC_pad (.PACKAGE_PIN(INLC), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INLC_c_0));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INLC_pad.PIN_TYPE = 6'b011001;
    defparam INLC_pad.PULLUP = 1'b0;
    defparam INLC_pad.NEG_TRIGGER = 1'b0;
    defparam INLC_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO INLA_pad (.PACKAGE_PIN(INLA), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INLA_c_0));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INLA_pad.PIN_TYPE = 6'b011001;
    defparam INLA_pad.PULLUP = 1'b0;
    defparam INLA_pad.NEG_TRIGGER = 1'b0;
    defparam INLA_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO INHB_pad (.PACKAGE_PIN(INHB), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INHB_c_0));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INHB_pad.PIN_TYPE = 6'b011001;
    defparam INHB_pad.PULLUP = 1'b0;
    defparam INHB_pad.NEG_TRIGGER = 1'b0;
    defparam INHB_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO INLB_pad (.PACKAGE_PIN(INLB), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INLB_c_0));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INLB_pad.PIN_TYPE = 6'b011001;
    defparam INLB_pad.PULLUP = 1'b0;
    defparam INLB_pad.NEG_TRIGGER = 1'b0;
    defparam INLB_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO INHC_pad (.PACKAGE_PIN(INHC), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INHC_c_0));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INHC_pad.PIN_TYPE = 6'b011001;
    defparam INHC_pad.PULLUP = 1'b0;
    defparam INHC_pad.NEG_TRIGGER = 1'b0;
    defparam INHC_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO CS_CLK_pad (.PACKAGE_PIN(CS_CLK), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(CS_CLK_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam CS_CLK_pad.PIN_TYPE = 6'b011001;
    defparam CS_CLK_pad.PULLUP = 1'b0;
    defparam CS_CLK_pad.NEG_TRIGGER = 1'b0;
    defparam CS_CLK_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 add_175_14_lut (.I0(GND_net), .I1(delay_counter[12]), .I2(GND_net), 
            .I3(n43621), .O(n1551)) /* synthesis syn_instantiated=1 */ ;
    defparam add_175_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1637_13 (.CI(n44193), 
            .I0(n2423), .I1(VCC_net), .CO(n44194));
    SB_LUT4 add_2747_5_lut (.I0(GND_net), .I1(n623), .I2(VCC_net), .I3(n43964), 
            .O(n8583)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2747_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1637_12_lut (.I0(GND_net), 
            .I1(n2424), .I2(VCC_net), .I3(n44192), .O(n2491)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1637_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_261_10_lut (.I0(current[8]), .I1(duty[11]), .I2(n56614), 
            .I3(n43565), .O(n262)) /* synthesis syn_instantiated=1 */ ;
    defparam add_261_10_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1637_12 (.CI(n44192), 
            .I0(n2424), .I1(VCC_net), .CO(n44193));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1637_11_lut (.I0(GND_net), 
            .I1(n2425), .I2(VCC_net), .I3(n44191), .O(n2492)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1637_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1637_11 (.CI(n44191), 
            .I0(n2425), .I1(VCC_net), .CO(n44192));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1637_10_lut (.I0(GND_net), 
            .I1(n2426), .I2(VCC_net), .I3(n44190), .O(n2493)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1637_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1637_10 (.CI(n44190), 
            .I0(n2426), .I1(VCC_net), .CO(n44191));
    SB_CARRY add_175_14 (.CI(n43621), .I0(delay_counter[12]), .I1(GND_net), 
            .CO(n43622));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1637_9_lut (.I0(GND_net), 
            .I1(n2427), .I2(VCC_net), .I3(n44189), .O(n2494)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1637_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_175_13_lut (.I0(GND_net), .I1(delay_counter[11]), .I2(GND_net), 
            .I3(n43620), .O(n1552)) /* synthesis syn_instantiated=1 */ ;
    defparam add_175_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2747_5 (.CI(n43964), .I0(n623), .I1(VCC_net), .CO(n43965));
    SB_LUT4 add_2747_4_lut (.I0(GND_net), .I1(n516), .I2(GND_net), .I3(n43963), 
            .O(n8584)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2747_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1820 (.I0(n4_adj_5495), .I1(n5_adj_5494), .I2(n407), 
            .I3(n6_adj_5493), .O(n5_adj_5643));
    defparam i1_4_lut_adj_1820.LUT_INIT = 16'heeea;
    SB_LUT4 i15790_3_lut (.I0(\data_out_frame[23] [6]), .I1(neopxl_color[22]), 
            .I2(n24210), .I3(GND_net), .O(n29870));   // verilog/coms.v(128[12] 303[6])
    defparam i15790_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1923_3_lut (.I0(n2824), 
            .I1(n2891), .I2(n2841), .I3(GND_net), .O(n2923));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1923_3_lut.LUT_INIT = 16'hacac;
    SB_IO DE_pad (.PACKAGE_PIN(DE), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DE_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DE_pad.PIN_TYPE = 6'b011001;
    defparam DE_pad.PULLUP = 1'b0;
    defparam DE_pad.NEG_TRIGGER = 1'b0;
    defparam DE_pad.IO_STANDARD = "SB_LVCMOS";
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1637_9 (.CI(n44189), 
            .I0(n2427), .I1(VCC_net), .CO(n44190));
    SB_CARRY add_2747_4 (.CI(n43963), .I0(n516), .I1(GND_net), .CO(n43964));
    SB_LUT4 add_2747_3_lut (.I0(GND_net), .I1(n625), .I2(VCC_net), .I3(n43962), 
            .O(n8585)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2747_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 n10829_bdd_4_lut (.I0(n10829), .I1(n418), .I2(current[15]), 
            .I3(duty[23]), .O(n56874));
    defparam n10829_bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n56874_bdd_3_lut (.I0(n56874), .I1(duty[23]), .I2(n249), .I3(GND_net), 
            .O(pwm_setpoint_23__N_11[23]));
    defparam n56874_bdd_3_lut.LUT_INIT = 16'h9898;
    SB_LUT4 n10829_bdd_4_lut_40999 (.I0(n10829), .I1(n419), .I2(current[15]), 
            .I3(duty[23]), .O(n56868));
    defparam n10829_bdd_4_lut_40999.LUT_INIT = 16'he4aa;
    SB_LUT4 n56868_bdd_4_lut (.I0(n56868), .I1(duty[22]), .I2(n249), .I3(duty[23]), 
            .O(pwm_setpoint_23__N_11[22]));
    defparam n56868_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n10829_bdd_4_lut_40994 (.I0(n10829), .I1(n420), .I2(current[15]), 
            .I3(duty[23]), .O(n56862));
    defparam n10829_bdd_4_lut_40994.LUT_INIT = 16'he4aa;
    SB_LUT4 n56862_bdd_4_lut (.I0(n56862), .I1(duty[21]), .I2(n249), .I3(duty[23]), 
            .O(pwm_setpoint_23__N_11[21]));
    defparam n56862_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1637_8_lut (.I0(GND_net), 
            .I1(n2428), .I2(VCC_net), .I3(n44188), .O(n2495)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1637_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15791_4_lut (.I0(r_Rx_Data), .I1(rx_data[2]), .I2(n4_adj_5469), 
            .I3(n27208), .O(n29871));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i15791_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 unary_minus_18_inv_0_i6_1_lut (.I0(duty[5]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n20));   // verilog/TinyFPGA_B.v(119[24:29])
    defparam unary_minus_18_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_2747_3 (.CI(n43962), .I0(n625), .I1(VCC_net), .CO(n43963));
    SB_LUT4 add_2747_2_lut (.I0(GND_net), .I1(n407), .I2(GND_net), .I3(VCC_net), 
            .O(n8586)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2747_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1928_3_lut (.I0(n2829), 
            .I1(n2896), .I2(n2841), .I3(GND_net), .O(n2928));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1928_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_2747_2 (.CI(VCC_net), .I0(n407), .I1(GND_net), .CO(n43962));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1637_8 (.CI(n44188), 
            .I0(n2428), .I1(VCC_net), .CO(n44189));
    SB_LUT4 i15792_3_lut (.I0(\data_out_frame[23] [5]), .I1(neopxl_color[21]), 
            .I2(n24210), .I3(GND_net), .O(n29872));   // verilog/coms.v(128[12] 303[6])
    defparam i15792_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34009_3_lut (.I0(n7_adj_5492), .I1(n8586), .I2(n49748), .I3(GND_net), 
            .O(n49757));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam i34009_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15793_3_lut (.I0(\data_out_frame[23] [4]), .I1(neopxl_color[20]), 
            .I2(n24210), .I3(GND_net), .O(n29873));   // verilog/coms.v(128[12] 303[6])
    defparam i15793_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15794_3_lut (.I0(\data_out_frame[23] [3]), .I1(neopxl_color[19]), 
            .I2(n24210), .I3(GND_net), .O(n29874));   // verilog/coms.v(128[12] 303[6])
    defparam i15794_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34010_rep_58_3_lut (.I0(encoder0_position_scaled_23__N_327[26]), 
            .I1(n900), .I2(n861), .I3(GND_net), .O(n53125));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam i34010_rep_58_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1821 (.I0(hall3), .I1(commutation_state[1]), .I2(hall2), 
            .I3(hall1), .O(n48778));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    defparam i1_4_lut_adj_1821.LUT_INIT = 16'hd054;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1916_3_lut (.I0(n2817), 
            .I1(n2884), .I2(n2841), .I3(GND_net), .O(n2916));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1916_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_175_13 (.CI(n43620), .I0(delay_counter[11]), .I1(GND_net), 
            .CO(n43621));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1930_3_lut (.I0(n2831), 
            .I1(n2898), .I2(n2841), .I3(GND_net), .O(n2930));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1930_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_175_12_lut (.I0(GND_net), .I1(delay_counter[10]), .I2(GND_net), 
            .I3(n43619), .O(n1553)) /* synthesis syn_instantiated=1 */ ;
    defparam add_175_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1637_7_lut (.I0(GND_net), 
            .I1(n2429), .I2(GND_net), .I3(n44187), .O(n2496)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1637_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1637_7 (.CI(n44187), 
            .I0(n2429), .I1(GND_net), .CO(n44188));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i639_3_lut (.I0(n932), .I1(n999), 
            .I2(n960), .I3(GND_net), .O(n1031));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i639_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1637_6_lut (.I0(GND_net), 
            .I1(n2430), .I2(GND_net), .I3(n44186), .O(n2497)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1637_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1637_6 (.CI(n44186), 
            .I0(n2430), .I1(GND_net), .CO(n44187));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1929_3_lut (.I0(n2830), 
            .I1(n2897), .I2(n2841), .I3(GND_net), .O(n2929));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1929_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i23328_4_lut (.I0(n834), .I1(n831), .I2(n832), .I3(n833), 
            .O(n37418));
    defparam i23328_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 i23400_4_lut (.I0(n829), .I1(n828), .I2(n37418), .I3(n830), 
            .O(n861));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam i23400_4_lut.LUT_INIT = 16'heccc;
    SB_LUT4 i15796_4_lut (.I0(CS_MISO_c), .I1(data_adj_5711[6]), .I2(n6_adj_5523), 
            .I3(n27258), .O(n29876));   // verilog/tli4970.v(35[10] 68[6])
    defparam i15796_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1927_3_lut (.I0(n2828), 
            .I1(n2895), .I2(n2841), .I3(GND_net), .O(n2927));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1927_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15797_4_lut (.I0(r_Rx_Data), .I1(rx_data[3]), .I2(n4_adj_5469), 
            .I3(n27203), .O(n29877));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i15797_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1925_3_lut (.I0(n2826), 
            .I1(n2893), .I2(n2841), .I3(GND_net), .O(n2925));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1925_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1922_3_lut (.I0(n2823), 
            .I1(n2890), .I2(n2841), .I3(GND_net), .O(n2922));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1922_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1919_3_lut (.I0(n2820), 
            .I1(n2887), .I2(n2841), .I3(GND_net), .O(n2919));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1919_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15798_4_lut (.I0(r_Rx_Data), .I1(rx_data[4]), .I2(n4_adj_5445), 
            .I3(n27208), .O(n29878));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i15798_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_mux_3_i26_3_lut (.I0(encoder0_position_scaled_23__N_327[25]), 
            .I1(n8_adj_5491), .I2(encoder0_position_scaled_23__N_327[31]), 
            .I3(GND_net), .O(n834));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_mux_3_i26_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_18_inv_0_i7_1_lut (.I0(duty[6]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n19));   // verilog/TinyFPGA_B.v(119[24:29])
    defparam unary_minus_18_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1637_5_lut (.I0(GND_net), 
            .I1(n2431), .I2(VCC_net), .I3(n44185), .O(n2498)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1637_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_175_12 (.CI(n43619), .I0(delay_counter[10]), .I1(GND_net), 
            .CO(n43620));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1637_5 (.CI(n44185), 
            .I0(n2431), .I1(VCC_net), .CO(n44186));
    SB_CARRY add_261_10 (.CI(n43565), .I0(duty[11]), .I1(n56614), .CO(n43566));
    SB_LUT4 add_175_11_lut (.I0(GND_net), .I1(delay_counter[9]), .I2(GND_net), 
            .I3(n43618), .O(n1554)) /* synthesis syn_instantiated=1 */ ;
    defparam add_175_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_261_9_lut (.I0(current[7]), .I1(duty[10]), .I2(n56614), 
            .I3(n43564), .O(n263)) /* synthesis syn_instantiated=1 */ ;
    defparam add_261_9_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY add_263_12 (.CI(n43544), .I0(encoder1_position[13]), .I1(GND_net), 
            .CO(n43545));
    SB_CARRY add_175_11 (.CI(n43618), .I0(delay_counter[9]), .I1(GND_net), 
            .CO(n43619));
    SB_LUT4 i23326_4_lut (.I0(n934), .I1(n931), .I2(n932), .I3(n933), 
            .O(n37416));
    defparam i23326_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 i1_2_lut_adj_1822 (.I0(n929), .I1(n930), .I2(GND_net), .I3(GND_net), 
            .O(n51834));
    defparam i1_2_lut_adj_1822.LUT_INIT = 16'h8888;
    SB_LUT4 i15799_4_lut (.I0(CS_MISO_c), .I1(data_adj_5711[7]), .I2(n6_adj_5523), 
            .I3(n27264), .O(n29879));   // verilog/tli4970.v(35[10] 68[6])
    defparam i15799_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i1_4_lut_adj_1823 (.I0(n927), .I1(n51834), .I2(n928), .I3(n37416), 
            .O(n960));
    defparam i1_4_lut_adj_1823.LUT_INIT = 16'hfefa;
    SB_LUT4 i40194_1_lut (.I0(n2940), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n56025));
    defparam i40194_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i573_3_lut (.I0(n834), .I1(n901), 
            .I2(n861), .I3(GND_net), .O(n933));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i573_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1824 (.I0(n2928), .I1(n2923), .I2(n2926), .I3(n2920), 
            .O(n51876));
    defparam i1_4_lut_adj_1824.LUT_INIT = 16'hfffe;
    SB_LUT4 add_175_10_lut (.I0(GND_net), .I1(delay_counter[8]), .I2(GND_net), 
            .I3(n43617), .O(n1555)) /* synthesis syn_instantiated=1 */ ;
    defparam add_175_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_175_10 (.CI(n43617), .I0(delay_counter[8]), .I1(GND_net), 
            .CO(n43618));
    SB_LUT4 add_175_9_lut (.I0(GND_net), .I1(delay_counter[7]), .I2(GND_net), 
            .I3(n43616), .O(n1556)) /* synthesis syn_instantiated=1 */ ;
    defparam add_175_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_175_9 (.CI(n43616), .I0(delay_counter[7]), .I1(GND_net), 
            .CO(n43617));
    SB_LUT4 add_263_4_lut (.I0(GND_net), .I1(encoder1_position[5]), .I2(GND_net), 
            .I3(n43536), .O(encoder1_position_scaled_23__N_75[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_263_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15800_4_lut (.I0(r_Rx_Data), .I1(rx_data[5]), .I2(n4_adj_5445), 
            .I3(n27203), .O(n29880));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i15800_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_25_lut (.I0(GND_net), .I1(encoder0_position_scaled[23]), 
            .I2(n2_adj_5521), .I3(n43954), .O(displacement_23__N_99[23])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_3_lut_adj_1825 (.I0(n51876), .I1(n2921), .I2(n2924), .I3(GND_net), 
            .O(n51878));
    defparam i1_3_lut_adj_1825.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_4_lut_adj_1826 (.I0(n2919), .I1(n2922), .I2(n2925), .I3(n2927), 
            .O(n51880));
    defparam i1_4_lut_adj_1826.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i640_3_lut (.I0(n933), .I1(n1000), 
            .I2(n960), .I3(GND_net), .O(n1032));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i640_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i707_3_lut (.I0(n1032), .I1(n1099), 
            .I2(n1059), .I3(GND_net), .O(n1131));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i707_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15801_3_lut (.I0(current[11]), .I1(data_adj_5711[11]), .I2(n28729), 
            .I3(GND_net), .O(n29881));   // verilog/tli4970.v(35[10] 68[6])
    defparam i15801_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i23286_4_lut (.I0(n540), .I1(n2931), .I2(n2932), .I3(n2933), 
            .O(n37376));
    defparam i23286_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 i15802_3_lut (.I0(current[10]), .I1(data_adj_5711[10]), .I2(n28729), 
            .I3(GND_net), .O(n29882));   // verilog/tli4970.v(35[10] 68[6])
    defparam i15802_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15803_3_lut (.I0(current[9]), .I1(data_adj_5711[9]), .I2(n28729), 
            .I3(GND_net), .O(n29883));   // verilog/tli4970.v(35[10] 68[6])
    defparam i15803_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15804_3_lut (.I0(current[8]), .I1(data_adj_5711[8]), .I2(n28729), 
            .I3(GND_net), .O(n29884));   // verilog/tli4970.v(35[10] 68[6])
    defparam i15804_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i706_3_lut (.I0(n1031), .I1(n1098), 
            .I2(n1059), .I3(GND_net), .O(n1130));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i706_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1827 (.I0(n2917), .I1(n2918), .I2(n51880), .I3(n51878), 
            .O(n51886));
    defparam i1_4_lut_adj_1827.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_24_lut (.I0(GND_net), .I1(encoder0_position_scaled[22]), 
            .I2(n3_adj_5520), .I3(n43953), .O(displacement_23__N_99[22])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_175_8_lut (.I0(GND_net), .I1(delay_counter[6]), .I2(GND_net), 
            .I3(n43615), .O(n1557)) /* synthesis syn_instantiated=1 */ ;
    defparam add_175_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_24 (.CI(n43953), .I0(encoder0_position_scaled[22]), 
            .I1(n3_adj_5520), .CO(n43954));
    SB_LUT4 i15805_3_lut (.I0(current[7]), .I1(data_adj_5711[7]), .I2(n28729), 
            .I3(GND_net), .O(n29885));   // verilog/tli4970.v(35[10] 68[6])
    defparam i15805_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_23_lut (.I0(GND_net), .I1(encoder0_position_scaled[21]), 
            .I2(n4_adj_5519), .I3(n43952), .O(displacement_23__N_99[21])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_23 (.CI(n43952), .I0(encoder0_position_scaled[21]), 
            .I1(n4_adj_5519), .CO(n43953));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1637_4_lut (.I0(GND_net), 
            .I1(n2432), .I2(GND_net), .I3(n44184), .O(n2499)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1637_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15806_3_lut (.I0(current[6]), .I1(data_adj_5711[6]), .I2(n28729), 
            .I3(GND_net), .O(n29886));   // verilog/tli4970.v(35[10] 68[6])
    defparam i15806_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_22_lut (.I0(GND_net), .I1(encoder0_position_scaled[20]), 
            .I2(n5_adj_5518), .I3(n43951), .O(displacement_23__N_99[20])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i775_3_lut (.I0(n1132), .I1(n1199), 
            .I2(n1158), .I3(GND_net), .O(n1231));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i775_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 unary_minus_18_inv_0_i8_1_lut (.I0(duty[7]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n18));   // verilog/TinyFPGA_B.v(119[24:29])
    defparam unary_minus_18_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_2_lut_adj_1828 (.I0(n2929), .I1(n2930), .I2(GND_net), .I3(GND_net), 
            .O(n52200));
    defparam i1_2_lut_adj_1828.LUT_INIT = 16'h8888;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_22 (.CI(n43951), .I0(encoder0_position_scaled[20]), 
            .I1(n5_adj_5518), .CO(n43952));
    SB_LUT4 i15807_3_lut (.I0(current[5]), .I1(data_adj_5711[5]), .I2(n28729), 
            .I3(GND_net), .O(n29887));   // verilog/tli4970.v(35[10] 68[6])
    defparam i15807_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_21_lut (.I0(GND_net), .I1(encoder0_position_scaled[19]), 
            .I2(n6_adj_5517), .I3(n43950), .O(displacement_23__N_99[19])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i774_3_lut (.I0(n1131), .I1(n1198), 
            .I2(n1158), .I3(GND_net), .O(n1230));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i774_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_21 (.CI(n43950), .I0(encoder0_position_scaled[19]), 
            .I1(n6_adj_5517), .CO(n43951));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_20_lut (.I0(GND_net), .I1(encoder0_position_scaled[18]), 
            .I2(n7_adj_5516), .I3(n43949), .O(displacement_23__N_99[18])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i773_3_lut (.I0(n1130), .I1(n1197), 
            .I2(n1158), .I3(GND_net), .O(n1229));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i773_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_20 (.CI(n43949), .I0(encoder0_position_scaled[18]), 
            .I1(n7_adj_5516), .CO(n43950));
    SB_LUT4 i1_4_lut_adj_1829 (.I0(n2916), .I1(n52200), .I2(n51886), .I3(n37376), 
            .O(n51890));
    defparam i1_4_lut_adj_1829.LUT_INIT = 16'hfefa;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i3_1_lut (.I0(encoder1_position_scaled[2]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n23_adj_5500));   // verilog/TinyFPGA_B.v(324[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_175_8 (.CI(n43615), .I0(delay_counter[6]), .I1(GND_net), 
            .CO(n43616));
    SB_LUT4 i15808_3_lut (.I0(current[4]), .I1(data_adj_5711[4]), .I2(n28729), 
            .I3(GND_net), .O(n29888));   // verilog/tli4970.v(35[10] 68[6])
    defparam i15808_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_175_7_lut (.I0(GND_net), .I1(delay_counter[5]), .I2(GND_net), 
            .I3(n43614), .O(n1558)) /* synthesis syn_instantiated=1 */ ;
    defparam add_175_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15809_3_lut (.I0(current[3]), .I1(data_adj_5711[3]), .I2(n28729), 
            .I3(GND_net), .O(n29889));   // verilog/tli4970.v(35[10] 68[6])
    defparam i15809_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_19_lut (.I0(GND_net), .I1(encoder0_position_scaled[17]), 
            .I2(n8_adj_5515), .I3(n43948), .O(displacement_23__N_99[17])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_19 (.CI(n43948), .I0(encoder0_position_scaled[17]), 
            .I1(n8_adj_5515), .CO(n43949));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_18_lut (.I0(GND_net), .I1(encoder0_position_scaled[16]), 
            .I2(n9_adj_5514), .I3(n43947), .O(displacement_23__N_99[16])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_18 (.CI(n43947), .I0(encoder0_position_scaled[16]), 
            .I1(n9_adj_5514), .CO(n43948));
    SB_LUT4 unary_minus_18_inv_0_i9_1_lut (.I0(duty[8]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n17));   // verilog/TinyFPGA_B.v(119[24:29])
    defparam unary_minus_18_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_17_lut (.I0(GND_net), .I1(encoder0_position_scaled[15]), 
            .I2(n10_adj_5513), .I3(n43946), .O(displacement_23__N_99[15])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_175_7 (.CI(n43614), .I0(delay_counter[5]), .I1(GND_net), 
            .CO(n43615));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_unary_minus_2_inv_0_i11_1_lut (.I0(encoder0_position_scaled_23__N_327[10]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n23_adj_5632));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_unary_minus_2_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_175_6_lut (.I0(GND_net), .I1(delay_counter[4]), .I2(GND_net), 
            .I3(n43613), .O(n1559)) /* synthesis syn_instantiated=1 */ ;
    defparam add_175_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_17 (.CI(n43946), .I0(encoder0_position_scaled[15]), 
            .I1(n10_adj_5513), .CO(n43947));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_16_lut (.I0(GND_net), .I1(encoder0_position_scaled[14]), 
            .I2(n11_adj_5512), .I3(n43945), .O(displacement_23__N_99[14])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1637_4 (.CI(n44184), 
            .I0(n2432), .I1(GND_net), .CO(n44185));
    SB_LUT4 i1_4_lut_adj_1830 (.I0(n2913), .I1(n2914), .I2(n2915), .I3(n51890), 
            .O(n51896));
    defparam i1_4_lut_adj_1830.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1831 (.I0(n2910), .I1(n2911), .I2(n2912), .I3(n51896), 
            .O(n51902));
    defparam i1_4_lut_adj_1831.LUT_INIT = 16'hfffe;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_16 (.CI(n43945), .I0(encoder0_position_scaled[14]), 
            .I1(n11_adj_5512), .CO(n43946));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_15_lut (.I0(GND_net), .I1(encoder0_position_scaled[13]), 
            .I2(n12_adj_5511), .I3(n43944), .O(displacement_23__N_99[13])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_15 (.CI(n43944), .I0(encoder0_position_scaled[13]), 
            .I1(n12_adj_5511), .CO(n43945));
    SB_LUT4 i40197_4_lut (.I0(n2908), .I1(n2907), .I2(n2909), .I3(n51902), 
            .O(n2940));
    defparam i40197_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_14_lut (.I0(GND_net), .I1(encoder0_position_scaled[12]), 
            .I2(n13_adj_5510), .I3(n43943), .O(displacement_23__N_99[12])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_14 (.CI(n43943), .I0(encoder0_position_scaled[12]), 
            .I1(n13_adj_5510), .CO(n43944));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_13_lut (.I0(GND_net), .I1(encoder0_position_scaled[11]), 
            .I2(n14_adj_5509), .I3(n43942), .O(displacement_23__N_99[11])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_175_6 (.CI(n43613), .I0(delay_counter[4]), .I1(GND_net), 
            .CO(n43614));
    SB_LUT4 add_175_5_lut (.I0(GND_net), .I1(delay_counter[3]), .I2(GND_net), 
            .I3(n43612), .O(n1560)) /* synthesis syn_instantiated=1 */ ;
    defparam add_175_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_13 (.CI(n43942), .I0(encoder0_position_scaled[11]), 
            .I1(n14_adj_5509), .CO(n43943));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_12_lut (.I0(GND_net), .I1(encoder0_position_scaled[10]), 
            .I2(n15_adj_5508), .I3(n43941), .O(displacement_23__N_99[10])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_12 (.CI(n43941), .I0(encoder0_position_scaled[10]), 
            .I1(n15_adj_5508), .CO(n43942));
    SB_LUT4 unary_minus_18_inv_0_i10_1_lut (.I0(duty[9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n16));   // verilog/TinyFPGA_B.v(119[24:29])
    defparam unary_minus_18_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_11_lut (.I0(GND_net), .I1(encoder0_position_scaled[9]), 
            .I2(n16_adj_5507), .I3(n43940), .O(displacement_23__N_99[9])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_175_5 (.CI(n43612), .I0(delay_counter[3]), .I1(GND_net), 
            .CO(n43613));
    SB_LUT4 add_175_4_lut (.I0(GND_net), .I1(delay_counter[2]), .I2(GND_net), 
            .I3(n43611), .O(n1561)) /* synthesis syn_instantiated=1 */ ;
    defparam add_175_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_175_4 (.CI(n43611), .I0(delay_counter[2]), .I1(GND_net), 
            .CO(n43612));
    SB_LUT4 i40551_1_lut (.I0(n1554_adj_5597), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n56382));
    defparam i40551_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1842_3_lut (.I0(n2711), 
            .I1(n2778), .I2(n2742), .I3(GND_net), .O(n2810));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1842_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_unary_minus_2_inv_0_i12_1_lut (.I0(encoder0_position_scaled_23__N_327[11]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n22_adj_5631));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_unary_minus_2_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_unary_minus_2_inv_0_i13_1_lut (.I0(encoder0_position_scaled_23__N_327[12]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n21_adj_5630));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_unary_minus_2_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_unary_minus_2_inv_0_i14_1_lut (.I0(encoder0_position_scaled_23__N_327[13]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n20_adj_5629));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_unary_minus_2_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_11 (.CI(n43940), .I0(encoder0_position_scaled[9]), 
            .I1(n16_adj_5507), .CO(n43941));
    SB_LUT4 add_175_3_lut (.I0(GND_net), .I1(delay_counter[1]), .I2(GND_net), 
            .I3(n43610), .O(n1562)) /* synthesis syn_instantiated=1 */ ;
    defparam add_175_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_263_11_lut (.I0(GND_net), .I1(encoder1_position[12]), .I2(GND_net), 
            .I3(n43543), .O(encoder1_position_scaled_23__N_75[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_263_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1637_3_lut (.I0(GND_net), 
            .I1(n2433), .I2(VCC_net), .I3(n44183), .O(n2500)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1637_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_10_lut (.I0(GND_net), .I1(encoder0_position_scaled[8]), 
            .I2(n17_adj_5506), .I3(n43939), .O(displacement_23__N_99[8])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_10 (.CI(n43939), .I0(encoder0_position_scaled[8]), 
            .I1(n17_adj_5506), .CO(n43940));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1637_3 (.CI(n44183), 
            .I0(n2433), .I1(VCC_net), .CO(n44184));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1840_3_lut (.I0(n2709), 
            .I1(n2776), .I2(n2742), .I3(GND_net), .O(n2808));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1840_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_unary_minus_2_inv_0_i15_1_lut (.I0(encoder0_position_scaled_23__N_327[14]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n19_adj_5628));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_unary_minus_2_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1848_3_lut (.I0(n2717), 
            .I1(n2784), .I2(n2742), .I3(GND_net), .O(n2816));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1848_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i40225_1_lut (.I0(n2841), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n56056));
    defparam i40225_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_175_3 (.CI(n43610), .I0(delay_counter[1]), .I1(GND_net), 
            .CO(n43611));
    SB_LUT4 add_175_2_lut (.I0(GND_net), .I1(delay_counter[0]), .I2(GND_net), 
            .I3(VCC_net), .O(n1563)) /* synthesis syn_instantiated=1 */ ;
    defparam add_175_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_261_9 (.CI(n43564), .I0(duty[10]), .I1(n56614), .CO(n43565));
    SB_CARRY add_263_4 (.CI(n43536), .I0(encoder1_position[5]), .I1(GND_net), 
            .CO(n43537));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_9_lut (.I0(GND_net), .I1(encoder0_position_scaled[7]), 
            .I2(n18_adj_5505), .I3(n43938), .O(displacement_23__N_99[7])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_9 (.CI(n43938), .I0(encoder0_position_scaled[7]), 
            .I1(n18_adj_5505), .CO(n43939));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_8_lut (.I0(GND_net), .I1(encoder0_position_scaled[6]), 
            .I2(n19_adj_5504), .I3(n43937), .O(displacement_23__N_99[6])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_8 (.CI(n43937), .I0(encoder0_position_scaled[6]), 
            .I1(n19_adj_5504), .CO(n43938));
    SB_CARRY add_175_2 (.CI(VCC_net), .I0(delay_counter[0]), .I1(GND_net), 
            .CO(n43610));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_7_lut (.I0(GND_net), .I1(encoder0_position_scaled[5]), 
            .I2(n20_adj_5503), .I3(n43936), .O(displacement_23__N_99[5])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_7 (.CI(n43936), .I0(encoder0_position_scaled[5]), 
            .I1(n20_adj_5503), .CO(n43937));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_6_lut (.I0(GND_net), .I1(encoder0_position_scaled[4]), 
            .I2(n21_adj_5502), .I3(n43935), .O(displacement_23__N_99[4])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_6 (.CI(n43935), .I0(encoder0_position_scaled[4]), 
            .I1(n21_adj_5502), .CO(n43936));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1174_3_lut (.I0(n1723), 
            .I1(n1790), .I2(n1752), .I3(GND_net), .O(n1822));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1174_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_5_lut (.I0(GND_net), .I1(encoder0_position_scaled[3]), 
            .I2(n22_adj_5501), .I3(n43934), .O(displacement_23__N_99[3])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_unary_minus_2_inv_0_i16_1_lut (.I0(encoder0_position_scaled_23__N_327[15]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n18_adj_5627));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_unary_minus_2_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1637_2_lut (.I0(GND_net), 
            .I1(n535), .I2(GND_net), .I3(VCC_net), .O(n2501)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1637_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_5 (.CI(n43934), .I0(encoder0_position_scaled[3]), 
            .I1(n22_adj_5501), .CO(n43935));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_4_lut (.I0(GND_net), .I1(encoder0_position_scaled[2]), 
            .I2(n23_adj_5500), .I3(n43933), .O(displacement_23__N_99[2])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_4 (.CI(n43933), .I0(encoder0_position_scaled[2]), 
            .I1(n23_adj_5500), .CO(n43934));
    SB_CARRY add_263_11 (.CI(n43543), .I0(encoder1_position[12]), .I1(GND_net), 
            .CO(n43544));
    SB_LUT4 add_261_8_lut (.I0(current[6]), .I1(duty[9]), .I2(n56614), 
            .I3(n43563), .O(n264)) /* synthesis syn_instantiated=1 */ ;
    defparam add_261_8_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1841_3_lut (.I0(n2710), 
            .I1(n2777), .I2(n2742), .I3(GND_net), .O(n2809));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1841_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1845_3_lut (.I0(n2714), 
            .I1(n2781), .I2(n2742), .I3(GND_net), .O(n2813));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1845_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1844_3_lut (.I0(n2713), 
            .I1(n2780), .I2(n2742), .I3(GND_net), .O(n2812));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1844_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i4_1_lut (.I0(encoder1_position_scaled[3]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n22_adj_5501));   // verilog/TinyFPGA_B.v(324[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1843_3_lut (.I0(n2712), 
            .I1(n2779), .I2(n2742), .I3(GND_net), .O(n2811));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1843_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15810_3_lut (.I0(current[2]), .I1(data_adj_5711[2]), .I2(n28729), 
            .I3(GND_net), .O(n29890));   // verilog/tli4970.v(35[10] 68[6])
    defparam i15810_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_unary_minus_2_inv_0_i17_1_lut (.I0(encoder0_position_scaled_23__N_327[16]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n17_adj_5626));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_unary_minus_2_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1863_3_lut (.I0(n2732), 
            .I1(n2799), .I2(n2742), .I3(GND_net), .O(n2831));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1863_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1862_3_lut (.I0(n2731), 
            .I1(n2798), .I2(n2742), .I3(GND_net), .O(n2830));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1862_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i23256_3_lut (.I0(n935), .I1(n1032), .I2(n1033), .I3(GND_net), 
            .O(n37346));
    defparam i23256_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_unary_minus_2_inv_0_i18_1_lut (.I0(encoder0_position_scaled_23__N_327[17]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n16_adj_5625));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_unary_minus_2_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_18_inv_0_i11_1_lut (.I0(duty[10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_5452));   // verilog/TinyFPGA_B.v(119[24:29])
    defparam unary_minus_18_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i5_1_lut (.I0(encoder1_position_scaled[4]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n21_adj_5502));   // verilog/TinyFPGA_B.v(324[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1861_3_lut (.I0(n2730), 
            .I1(n2797), .I2(n2742), .I3(GND_net), .O(n2829));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1861_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1637_2 (.CI(VCC_net), 
            .I0(n535), .I1(GND_net), .CO(n44183));
    SB_DFF displacement_i23 (.Q(displacement[23]), .C(clk16MHz), .D(displacement_23__N_99[23]));   // verilog/TinyFPGA_B.v(321[10] 334[6])
    SB_DFF displacement_i22 (.Q(displacement[22]), .C(clk16MHz), .D(displacement_23__N_99[22]));   // verilog/TinyFPGA_B.v(321[10] 334[6])
    SB_LUT4 encoder0_position_scaled_23__I_0_227_unary_minus_2_inv_0_i19_1_lut (.I0(encoder0_position_scaled_23__N_327[18]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n15_adj_5624));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_unary_minus_2_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_18_inv_0_i12_1_lut (.I0(duty[11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n14));   // verilog/TinyFPGA_B.v(119[24:29])
    defparam unary_minus_18_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1865_3_lut (.I0(n538), .I1(n2801), 
            .I2(n2742), .I3(GND_net), .O(n2833));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1865_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1864_3_lut (.I0(n2733), 
            .I1(n2800), .I2(n2742), .I3(GND_net), .O(n2832));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1864_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i6_1_lut (.I0(encoder1_position_scaled[5]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n20_adj_5503));   // verilog/TinyFPGA_B.v(324[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1570_23_lut (.I0(n56200), 
            .I1(n2313), .I2(VCC_net), .I3(n44182), .O(n2412)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1570_23_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_3_lut (.I0(GND_net), .I1(encoder0_position_scaled[1]), 
            .I2(n24_adj_5499), .I3(n43932), .O(displacement_23__N_99[1])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_261_8 (.CI(n43563), .I0(duty[9]), .I1(n56614), .CO(n43564));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_mux_3_i6_3_lut (.I0(encoder0_position_scaled_23__N_327[5]), 
            .I1(n28), .I2(encoder0_position_scaled_23__N_327[31]), .I3(GND_net), 
            .O(n539));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_mux_3_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_3 (.CI(n43932), .I0(encoder0_position_scaled[1]), 
            .I1(n24_adj_5499), .CO(n43933));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_2_lut (.I0(GND_net), .I1(encoder0_position_scaled[0]), 
            .I2(n25_adj_5498), .I3(VCC_net), .O(displacement_23__N_99[0])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1570_22_lut (.I0(GND_net), 
            .I1(n2314), .I2(VCC_net), .I3(n44181), .O(n2381)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1570_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1570_22 (.CI(n44181), 
            .I0(n2314), .I1(VCC_net), .CO(n44182));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1570_21_lut (.I0(GND_net), 
            .I1(n2315), .I2(VCC_net), .I3(n44180), .O(n2382)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1570_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_2 (.CI(VCC_net), .I0(encoder0_position_scaled[0]), 
            .I1(n25_adj_5498), .CO(n43932));
    SB_LUT4 add_261_7_lut (.I0(current[5]), .I1(duty[8]), .I2(n56614), 
            .I3(n43562), .O(n265)) /* synthesis syn_instantiated=1 */ ;
    defparam add_261_7_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1570_21 (.CI(n44180), 
            .I0(n2315), .I1(VCC_net), .CO(n44181));
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i7_1_lut (.I0(encoder1_position_scaled[6]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n19_adj_5504));   // verilog/TinyFPGA_B.v(324[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1570_20_lut (.I0(GND_net), 
            .I1(n2316), .I2(VCC_net), .I3(n44179), .O(n2383)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1570_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1860_3_lut (.I0(n2729), 
            .I1(n2796), .I2(n2742), .I3(GND_net), .O(n2828));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1860_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i8_1_lut (.I0(encoder1_position_scaled[7]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n18_adj_5505));   // verilog/TinyFPGA_B.v(324[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1570_20 (.CI(n44179), 
            .I0(n2316), .I1(VCC_net), .CO(n44180));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1570_19_lut (.I0(GND_net), 
            .I1(n2317), .I2(VCC_net), .I3(n44178), .O(n2384)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1570_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15811_3_lut (.I0(current[1]), .I1(data_adj_5711[1]), .I2(n28729), 
            .I3(GND_net), .O(n29891));   // verilog/tli4970.v(35[10] 68[6])
    defparam i15811_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF displacement_i21 (.Q(displacement[21]), .C(clk16MHz), .D(displacement_23__N_99[21]));   // verilog/TinyFPGA_B.v(321[10] 334[6])
    SB_DFF displacement_i20 (.Q(displacement[20]), .C(clk16MHz), .D(displacement_23__N_99[20]));   // verilog/TinyFPGA_B.v(321[10] 334[6])
    SB_DFF displacement_i19 (.Q(displacement[19]), .C(clk16MHz), .D(displacement_23__N_99[19]));   // verilog/TinyFPGA_B.v(321[10] 334[6])
    SB_DFF displacement_i18 (.Q(displacement[18]), .C(clk16MHz), .D(displacement_23__N_99[18]));   // verilog/TinyFPGA_B.v(321[10] 334[6])
    SB_DFF displacement_i17 (.Q(displacement[17]), .C(clk16MHz), .D(displacement_23__N_99[17]));   // verilog/TinyFPGA_B.v(321[10] 334[6])
    SB_DFF displacement_i16 (.Q(displacement[16]), .C(clk16MHz), .D(displacement_23__N_99[16]));   // verilog/TinyFPGA_B.v(321[10] 334[6])
    SB_DFF displacement_i15 (.Q(displacement[15]), .C(clk16MHz), .D(displacement_23__N_99[15]));   // verilog/TinyFPGA_B.v(321[10] 334[6])
    SB_DFF displacement_i14 (.Q(displacement[14]), .C(clk16MHz), .D(displacement_23__N_99[14]));   // verilog/TinyFPGA_B.v(321[10] 334[6])
    SB_DFF displacement_i13 (.Q(displacement[13]), .C(clk16MHz), .D(displacement_23__N_99[13]));   // verilog/TinyFPGA_B.v(321[10] 334[6])
    SB_DFF displacement_i12 (.Q(displacement[12]), .C(clk16MHz), .D(displacement_23__N_99[12]));   // verilog/TinyFPGA_B.v(321[10] 334[6])
    SB_DFF displacement_i11 (.Q(displacement[11]), .C(clk16MHz), .D(displacement_23__N_99[11]));   // verilog/TinyFPGA_B.v(321[10] 334[6])
    SB_DFF displacement_i10 (.Q(displacement[10]), .C(clk16MHz), .D(displacement_23__N_99[10]));   // verilog/TinyFPGA_B.v(321[10] 334[6])
    SB_DFF displacement_i9 (.Q(displacement[9]), .C(clk16MHz), .D(displacement_23__N_99[9]));   // verilog/TinyFPGA_B.v(321[10] 334[6])
    SB_DFF displacement_i8 (.Q(displacement[8]), .C(clk16MHz), .D(displacement_23__N_99[8]));   // verilog/TinyFPGA_B.v(321[10] 334[6])
    SB_DFF displacement_i7 (.Q(displacement[7]), .C(clk16MHz), .D(displacement_23__N_99[7]));   // verilog/TinyFPGA_B.v(321[10] 334[6])
    SB_DFF displacement_i6 (.Q(displacement[6]), .C(clk16MHz), .D(displacement_23__N_99[6]));   // verilog/TinyFPGA_B.v(321[10] 334[6])
    SB_DFF displacement_i5 (.Q(displacement[5]), .C(clk16MHz), .D(displacement_23__N_99[5]));   // verilog/TinyFPGA_B.v(321[10] 334[6])
    SB_DFF displacement_i4 (.Q(displacement[4]), .C(clk16MHz), .D(displacement_23__N_99[4]));   // verilog/TinyFPGA_B.v(321[10] 334[6])
    SB_DFF displacement_i3 (.Q(displacement[3]), .C(clk16MHz), .D(displacement_23__N_99[3]));   // verilog/TinyFPGA_B.v(321[10] 334[6])
    SB_DFF displacement_i2 (.Q(displacement[2]), .C(clk16MHz), .D(displacement_23__N_99[2]));   // verilog/TinyFPGA_B.v(321[10] 334[6])
    SB_DFF displacement_i1 (.Q(displacement[1]), .C(clk16MHz), .D(displacement_23__N_99[1]));   // verilog/TinyFPGA_B.v(321[10] 334[6])
    SB_DFF encoder1_position_scaled_i23 (.Q(encoder1_position_scaled[23]), 
           .C(clk16MHz), .D(encoder1_position_scaled_23__N_75[23]));   // verilog/TinyFPGA_B.v(321[10] 334[6])
    SB_DFF encoder1_position_scaled_i22 (.Q(encoder1_position_scaled[22]), 
           .C(clk16MHz), .D(encoder1_position_scaled_23__N_75[22]));   // verilog/TinyFPGA_B.v(321[10] 334[6])
    SB_DFF encoder1_position_scaled_i21 (.Q(encoder1_position_scaled[21]), 
           .C(clk16MHz), .D(encoder1_position_scaled_23__N_75[21]));   // verilog/TinyFPGA_B.v(321[10] 334[6])
    SB_DFF encoder1_position_scaled_i20 (.Q(encoder1_position_scaled[20]), 
           .C(clk16MHz), .D(encoder1_position_scaled_23__N_75[20]));   // verilog/TinyFPGA_B.v(321[10] 334[6])
    SB_DFF encoder1_position_scaled_i19 (.Q(encoder1_position_scaled[19]), 
           .C(clk16MHz), .D(encoder1_position_scaled_23__N_75[19]));   // verilog/TinyFPGA_B.v(321[10] 334[6])
    SB_DFF encoder1_position_scaled_i18 (.Q(encoder1_position_scaled[18]), 
           .C(clk16MHz), .D(encoder1_position_scaled_23__N_75[18]));   // verilog/TinyFPGA_B.v(321[10] 334[6])
    SB_DFF encoder1_position_scaled_i17 (.Q(encoder1_position_scaled[17]), 
           .C(clk16MHz), .D(encoder1_position_scaled_23__N_75[17]));   // verilog/TinyFPGA_B.v(321[10] 334[6])
    SB_DFF encoder1_position_scaled_i16 (.Q(encoder1_position_scaled[16]), 
           .C(clk16MHz), .D(encoder1_position_scaled_23__N_75[16]));   // verilog/TinyFPGA_B.v(321[10] 334[6])
    SB_DFF encoder1_position_scaled_i15 (.Q(encoder1_position_scaled[15]), 
           .C(clk16MHz), .D(encoder1_position_scaled_23__N_75[15]));   // verilog/TinyFPGA_B.v(321[10] 334[6])
    SB_DFF encoder1_position_scaled_i14 (.Q(encoder1_position_scaled[14]), 
           .C(clk16MHz), .D(encoder1_position_scaled_23__N_75[14]));   // verilog/TinyFPGA_B.v(321[10] 334[6])
    SB_DFF encoder1_position_scaled_i13 (.Q(encoder1_position_scaled[13]), 
           .C(clk16MHz), .D(encoder1_position_scaled_23__N_75[13]));   // verilog/TinyFPGA_B.v(321[10] 334[6])
    SB_DFF encoder1_position_scaled_i12 (.Q(encoder1_position_scaled[12]), 
           .C(clk16MHz), .D(encoder1_position_scaled_23__N_75[12]));   // verilog/TinyFPGA_B.v(321[10] 334[6])
    SB_DFF encoder1_position_scaled_i11 (.Q(encoder1_position_scaled[11]), 
           .C(clk16MHz), .D(encoder1_position_scaled_23__N_75[11]));   // verilog/TinyFPGA_B.v(321[10] 334[6])
    SB_DFF encoder1_position_scaled_i10 (.Q(encoder1_position_scaled[10]), 
           .C(clk16MHz), .D(encoder1_position_scaled_23__N_75[10]));   // verilog/TinyFPGA_B.v(321[10] 334[6])
    SB_DFF encoder1_position_scaled_i9 (.Q(encoder1_position_scaled[9]), .C(clk16MHz), 
           .D(encoder1_position_scaled_23__N_75[9]));   // verilog/TinyFPGA_B.v(321[10] 334[6])
    SB_DFF encoder1_position_scaled_i8 (.Q(encoder1_position_scaled[8]), .C(clk16MHz), 
           .D(encoder1_position_scaled_23__N_75[8]));   // verilog/TinyFPGA_B.v(321[10] 334[6])
    SB_DFF encoder1_position_scaled_i7 (.Q(encoder1_position_scaled[7]), .C(clk16MHz), 
           .D(encoder1_position_scaled_23__N_75[7]));   // verilog/TinyFPGA_B.v(321[10] 334[6])
    SB_DFF encoder1_position_scaled_i6 (.Q(encoder1_position_scaled[6]), .C(clk16MHz), 
           .D(encoder1_position_scaled_23__N_75[6]));   // verilog/TinyFPGA_B.v(321[10] 334[6])
    SB_DFF encoder1_position_scaled_i5 (.Q(encoder1_position_scaled[5]), .C(clk16MHz), 
           .D(encoder1_position_scaled_23__N_75[5]));   // verilog/TinyFPGA_B.v(321[10] 334[6])
    SB_DFF encoder1_position_scaled_i4 (.Q(encoder1_position_scaled[4]), .C(clk16MHz), 
           .D(encoder1_position_scaled_23__N_75[4]));   // verilog/TinyFPGA_B.v(321[10] 334[6])
    SB_DFF encoder1_position_scaled_i3 (.Q(encoder1_position_scaled[3]), .C(clk16MHz), 
           .D(encoder1_position_scaled_23__N_75[3]));   // verilog/TinyFPGA_B.v(321[10] 334[6])
    SB_DFF encoder1_position_scaled_i2 (.Q(encoder1_position_scaled[2]), .C(clk16MHz), 
           .D(encoder1_position_scaled_23__N_75[2]));   // verilog/TinyFPGA_B.v(321[10] 334[6])
    SB_DFF encoder1_position_scaled_i1 (.Q(encoder1_position_scaled[1]), .C(clk16MHz), 
           .D(encoder1_position_scaled_23__N_75[1]));   // verilog/TinyFPGA_B.v(321[10] 334[6])
    SB_DFF encoder0_position_scaled_i23 (.Q(encoder0_position_scaled[23]), 
           .C(clk16MHz), .D(encoder0_position_scaled_23__N_51[23]));   // verilog/TinyFPGA_B.v(321[10] 334[6])
    SB_LUT4 i15812_4_lut (.I0(CS_MISO_c), .I1(data_adj_5711[8]), .I2(n5_adj_5524), 
            .I3(n27198), .O(n29892));   // verilog/tli4970.v(35[10] 68[6])
    defparam i15812_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_unary_minus_2_inv_0_i20_1_lut (.I0(encoder0_position_scaled_23__N_327[19]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n14_adj_5623));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_unary_minus_2_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1856_3_lut (.I0(n2725), 
            .I1(n2792), .I2(n2742), .I3(GND_net), .O(n2824));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1856_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1847_3_lut (.I0(n2716), 
            .I1(n2783), .I2(n2742), .I3(GND_net), .O(n2815));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1847_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1846_3_lut (.I0(n2715), 
            .I1(n2782), .I2(n2742), .I3(GND_net), .O(n2814));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1846_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1858_3_lut (.I0(n2727), 
            .I1(n2794), .I2(n2742), .I3(GND_net), .O(n2826));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1858_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_unary_minus_2_inv_0_i21_1_lut (.I0(encoder0_position_scaled_23__N_327[20]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n13_adj_5622));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_unary_minus_2_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_18_inv_0_i13_1_lut (.I0(duty[12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n13));   // verilog/TinyFPGA_B.v(119[24:29])
    defparam unary_minus_18_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i9_1_lut (.I0(encoder1_position_scaled[8]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n17_adj_5506));   // verilog/TinyFPGA_B.v(324[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_DFF encoder0_position_scaled_i22 (.Q(encoder0_position_scaled[22]), 
           .C(clk16MHz), .D(encoder0_position_scaled_23__N_51[22]));   // verilog/TinyFPGA_B.v(321[10] 334[6])
    SB_LUT4 encoder0_position_scaled_23__I_0_227_unary_minus_2_inv_0_i22_1_lut (.I0(encoder0_position_scaled_23__N_327[21]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n12_adj_5621));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_unary_minus_2_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_unary_minus_2_inv_0_i23_1_lut (.I0(encoder0_position_scaled_23__N_327[22]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n11_adj_5620));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_unary_minus_2_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_DFF encoder0_position_scaled_i21 (.Q(encoder0_position_scaled[21]), 
           .C(clk16MHz), .D(encoder0_position_scaled_23__N_51[21]));   // verilog/TinyFPGA_B.v(321[10] 334[6])
    SB_DFF encoder0_position_scaled_i20 (.Q(encoder0_position_scaled[20]), 
           .C(clk16MHz), .D(encoder0_position_scaled_23__N_51[20]));   // verilog/TinyFPGA_B.v(321[10] 334[6])
    SB_DFF encoder0_position_scaled_i19 (.Q(encoder0_position_scaled[19]), 
           .C(clk16MHz), .D(encoder0_position_scaled_23__N_51[19]));   // verilog/TinyFPGA_B.v(321[10] 334[6])
    SB_DFF encoder0_position_scaled_i18 (.Q(encoder0_position_scaled[18]), 
           .C(clk16MHz), .D(encoder0_position_scaled_23__N_51[18]));   // verilog/TinyFPGA_B.v(321[10] 334[6])
    SB_DFF encoder0_position_scaled_i17 (.Q(encoder0_position_scaled[17]), 
           .C(clk16MHz), .D(encoder0_position_scaled_23__N_51[17]));   // verilog/TinyFPGA_B.v(321[10] 334[6])
    SB_DFF encoder0_position_scaled_i16 (.Q(encoder0_position_scaled[16]), 
           .C(clk16MHz), .D(encoder0_position_scaled_23__N_51[16]));   // verilog/TinyFPGA_B.v(321[10] 334[6])
    SB_DFF encoder0_position_scaled_i15 (.Q(encoder0_position_scaled[15]), 
           .C(clk16MHz), .D(encoder0_position_scaled_23__N_51[15]));   // verilog/TinyFPGA_B.v(321[10] 334[6])
    SB_DFF encoder0_position_scaled_i14 (.Q(encoder0_position_scaled[14]), 
           .C(clk16MHz), .D(encoder0_position_scaled_23__N_51[14]));   // verilog/TinyFPGA_B.v(321[10] 334[6])
    SB_DFF encoder0_position_scaled_i13 (.Q(encoder0_position_scaled[13]), 
           .C(clk16MHz), .D(encoder0_position_scaled_23__N_51[13]));   // verilog/TinyFPGA_B.v(321[10] 334[6])
    SB_DFF encoder0_position_scaled_i12 (.Q(encoder0_position_scaled[12]), 
           .C(clk16MHz), .D(encoder0_position_scaled_23__N_51[12]));   // verilog/TinyFPGA_B.v(321[10] 334[6])
    SB_DFF encoder0_position_scaled_i11 (.Q(encoder0_position_scaled[11]), 
           .C(clk16MHz), .D(encoder0_position_scaled_23__N_51[11]));   // verilog/TinyFPGA_B.v(321[10] 334[6])
    SB_DFF encoder0_position_scaled_i10 (.Q(encoder0_position_scaled[10]), 
           .C(clk16MHz), .D(encoder0_position_scaled_23__N_51[10]));   // verilog/TinyFPGA_B.v(321[10] 334[6])
    SB_DFF encoder0_position_scaled_i9 (.Q(encoder0_position_scaled[9]), .C(clk16MHz), 
           .D(encoder0_position_scaled_23__N_51[9]));   // verilog/TinyFPGA_B.v(321[10] 334[6])
    SB_DFF encoder0_position_scaled_i8 (.Q(encoder0_position_scaled[8]), .C(clk16MHz), 
           .D(encoder0_position_scaled_23__N_51[8]));   // verilog/TinyFPGA_B.v(321[10] 334[6])
    SB_DFF encoder0_position_scaled_i7 (.Q(encoder0_position_scaled[7]), .C(clk16MHz), 
           .D(encoder0_position_scaled_23__N_51[7]));   // verilog/TinyFPGA_B.v(321[10] 334[6])
    SB_DFF encoder0_position_scaled_i6 (.Q(encoder0_position_scaled[6]), .C(clk16MHz), 
           .D(encoder0_position_scaled_23__N_51[6]));   // verilog/TinyFPGA_B.v(321[10] 334[6])
    SB_DFF encoder0_position_scaled_i5 (.Q(encoder0_position_scaled[5]), .C(clk16MHz), 
           .D(encoder0_position_scaled_23__N_51[5]));   // verilog/TinyFPGA_B.v(321[10] 334[6])
    SB_DFF encoder0_position_scaled_i4 (.Q(encoder0_position_scaled[4]), .C(clk16MHz), 
           .D(encoder0_position_scaled_23__N_51[4]));   // verilog/TinyFPGA_B.v(321[10] 334[6])
    SB_DFF encoder0_position_scaled_i3 (.Q(encoder0_position_scaled[3]), .C(clk16MHz), 
           .D(encoder0_position_scaled_23__N_51[3]));   // verilog/TinyFPGA_B.v(321[10] 334[6])
    SB_DFF encoder0_position_scaled_i2 (.Q(encoder0_position_scaled[2]), .C(clk16MHz), 
           .D(encoder0_position_scaled_23__N_51[2]));   // verilog/TinyFPGA_B.v(321[10] 334[6])
    SB_DFF encoder0_position_scaled_i1 (.Q(encoder0_position_scaled[1]), .C(clk16MHz), 
           .D(encoder0_position_scaled_23__N_51[1]));   // verilog/TinyFPGA_B.v(321[10] 334[6])
    SB_LUT4 unary_minus_18_inv_0_i14_1_lut (.I0(duty[13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n12));   // verilog/TinyFPGA_B.v(119[24:29])
    defparam unary_minus_18_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1570_19 (.CI(n44178), 
            .I0(n2317), .I1(VCC_net), .CO(n44179));
    SB_LUT4 unary_minus_18_inv_0_i15_1_lut (.I0(duty[14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n11));   // verilog/TinyFPGA_B.v(119[24:29])
    defparam unary_minus_18_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1570_18_lut (.I0(GND_net), 
            .I1(n2318), .I2(VCC_net), .I3(n44177), .O(n2385)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1570_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1859_3_lut (.I0(n2728), 
            .I1(n2795), .I2(n2742), .I3(GND_net), .O(n2827));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1859_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 unary_minus_18_inv_0_i16_1_lut (.I0(duty[15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n10_adj_5451));   // verilog/TinyFPGA_B.v(119[24:29])
    defparam unary_minus_18_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1851_3_lut (.I0(n2720), 
            .I1(n2787), .I2(n2742), .I3(GND_net), .O(n2819));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1851_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 unary_minus_18_inv_0_i17_1_lut (.I0(duty[16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n9));   // verilog/TinyFPGA_B.v(119[24:29])
    defparam unary_minus_18_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1853_3_lut (.I0(n2722), 
            .I1(n2789), .I2(n2742), .I3(GND_net), .O(n2821));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1853_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15813_3_lut (.I0(\PID_CONTROLLER.integral [23]), .I1(\PID_CONTROLLER.integral_23__N_3996 [23]), 
            .I2(control_update), .I3(GND_net), .O(n29893));   // verilog/motorControl.v(41[14] 61[8])
    defparam i15813_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1570_18 (.CI(n44177), 
            .I0(n2318), .I1(VCC_net), .CO(n44178));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_unary_minus_2_inv_0_i24_1_lut (.I0(encoder0_position_scaled_23__N_327[23]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n10_adj_5619));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_unary_minus_2_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1852_3_lut (.I0(n2721), 
            .I1(n2788), .I2(n2742), .I3(GND_net), .O(n2820));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1852_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_unary_minus_2_inv_0_i25_1_lut (.I0(encoder0_position_scaled_23__N_327[24]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n9_adj_5618));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_unary_minus_2_inv_0_i25_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1570_17_lut (.I0(GND_net), 
            .I1(n2319), .I2(VCC_net), .I3(n44176), .O(n2386)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1570_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_18_inv_0_i18_1_lut (.I0(duty[17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n8_adj_5450));   // verilog/TinyFPGA_B.v(119[24:29])
    defparam unary_minus_18_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_DFF commutation_state_prev_i2 (.Q(commutation_state_prev[2]), .C(clk16MHz), 
           .D(commutation_state[2]));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i10_1_lut (.I0(encoder1_position_scaled[9]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n16_adj_5507));   // verilog/TinyFPGA_B.v(324[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i11_1_lut (.I0(encoder1_position_scaled[10]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n15_adj_5508));   // verilog/TinyFPGA_B.v(324[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_261_7 (.CI(n43562), .I0(duty[8]), .I1(n56614), .CO(n43563));
    SB_LUT4 add_263_10_lut (.I0(GND_net), .I1(encoder1_position[11]), .I2(GND_net), 
            .I3(n43542), .O(encoder1_position_scaled_23__N_75[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_263_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1857_3_lut (.I0(n2726), 
            .I1(n2793), .I2(n2742), .I3(GND_net), .O(n2825));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1857_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15814_3_lut (.I0(\PID_CONTROLLER.integral [22]), .I1(\PID_CONTROLLER.integral_23__N_3996 [22]), 
            .I2(control_update), .I3(GND_net), .O(n29894));   // verilog/motorControl.v(41[14] 61[8])
    defparam i15814_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15815_3_lut (.I0(\PID_CONTROLLER.integral [21]), .I1(\PID_CONTROLLER.integral_23__N_3996 [21]), 
            .I2(control_update), .I3(GND_net), .O(n29895));   // verilog/motorControl.v(41[14] 61[8])
    defparam i15815_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i12_1_lut (.I0(encoder1_position_scaled[11]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n14_adj_5509));   // verilog/TinyFPGA_B.v(324[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i15816_3_lut (.I0(\PID_CONTROLLER.integral [20]), .I1(\PID_CONTROLLER.integral_23__N_3996 [20]), 
            .I2(control_update), .I3(GND_net), .O(n29896));   // verilog/motorControl.v(41[14] 61[8])
    defparam i15816_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1855_3_lut (.I0(n2724), 
            .I1(n2791), .I2(n2742), .I3(GND_net), .O(n2823));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1855_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i13_1_lut (.I0(encoder1_position_scaled[12]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n13_adj_5510));   // verilog/TinyFPGA_B.v(324[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_18_inv_0_i19_1_lut (.I0(duty[18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n7_adj_5449));   // verilog/TinyFPGA_B.v(119[24:29])
    defparam unary_minus_18_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i15817_3_lut (.I0(\PID_CONTROLLER.integral [19]), .I1(\PID_CONTROLLER.integral_23__N_3996 [19]), 
            .I2(control_update), .I3(GND_net), .O(n29897));   // verilog/motorControl.v(41[14] 61[8])
    defparam i15817_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1854_3_lut (.I0(n2723), 
            .I1(n2790), .I2(n2742), .I3(GND_net), .O(n2822));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1854_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1850_3_lut (.I0(n2719), 
            .I1(n2786), .I2(n2742), .I3(GND_net), .O(n2818));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1850_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15818_3_lut (.I0(\PID_CONTROLLER.integral [18]), .I1(\PID_CONTROLLER.integral_23__N_3996 [18]), 
            .I2(control_update), .I3(GND_net), .O(n29898));   // verilog/motorControl.v(41[14] 61[8])
    defparam i15818_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15819_3_lut (.I0(\PID_CONTROLLER.integral [17]), .I1(\PID_CONTROLLER.integral_23__N_3996 [17]), 
            .I2(control_update), .I3(GND_net), .O(n29899));   // verilog/motorControl.v(41[14] 61[8])
    defparam i15819_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5_4_lut (.I0(delay_counter[27]), .I1(delay_counter[29]), .I2(delay_counter[24]), 
            .I3(delay_counter[26]), .O(n12_adj_5604));
    defparam i5_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i6_4_lut_adj_1832 (.I0(delay_counter[28]), .I1(n12_adj_5604), 
            .I2(delay_counter[25]), .I3(delay_counter[30]), .O(n27116));
    defparam i6_4_lut_adj_1832.LUT_INIT = 16'hfffe;
    SB_LUT4 i5_3_lut (.I0(delay_counter[3]), .I1(delay_counter[5]), .I2(delay_counter[4]), 
            .I3(GND_net), .O(n14_adj_5468));
    defparam i5_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 unary_minus_18_inv_0_i20_1_lut (.I0(duty[19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_5448));   // verilog/TinyFPGA_B.v(119[24:29])
    defparam unary_minus_18_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_unary_minus_2_inv_0_i26_1_lut (.I0(encoder0_position_scaled_23__N_327[25]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n8_adj_5617));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_unary_minus_2_inv_0_i26_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1849_3_lut (.I0(n2718), 
            .I1(n2785), .I2(n2742), .I3(GND_net), .O(n2817));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1849_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1833 (.I0(n2822), .I1(n2823), .I2(n2825), .I3(n2820), 
            .O(n52182));
    defparam i1_4_lut_adj_1833.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_unary_minus_2_inv_0_i27_1_lut (.I0(encoder0_position_scaled_23__N_327[26]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n7_adj_5616));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_unary_minus_2_inv_0_i27_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i6_4_lut_adj_1834 (.I0(delay_counter[8]), .I1(delay_counter[7]), 
            .I2(delay_counter[1]), .I3(delay_counter[0]), .O(n15_adj_5467));
    defparam i6_4_lut_adj_1834.LUT_INIT = 16'hfffe;
    SB_LUT4 i8_4_lut (.I0(n15_adj_5467), .I1(delay_counter[2]), .I2(n14_adj_5468), 
            .I3(delay_counter[6]), .O(n27119));
    defparam i8_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 unary_minus_18_inv_0_i21_1_lut (.I0(duty[20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n5_adj_5447));   // verilog/TinyFPGA_B.v(119[24:29])
    defparam unary_minus_18_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i15820_3_lut (.I0(\PID_CONTROLLER.integral [16]), .I1(\PID_CONTROLLER.integral_23__N_3996 [16]), 
            .I2(control_update), .I3(GND_net), .O(n29900));   // verilog/motorControl.v(41[14] 61[8])
    defparam i15820_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15821_3_lut (.I0(\PID_CONTROLLER.integral [15]), .I1(\PID_CONTROLLER.integral_23__N_3996 [15]), 
            .I2(control_update), .I3(GND_net), .O(n29901));   // verilog/motorControl.v(41[14] 61[8])
    defparam i15821_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15822_3_lut (.I0(\PID_CONTROLLER.integral [14]), .I1(\PID_CONTROLLER.integral_23__N_3996 [14]), 
            .I2(control_update), .I3(GND_net), .O(n29902));   // verilog/motorControl.v(41[14] 61[8])
    defparam i15822_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1835 (.I0(n2821), .I1(n2819), .I2(n2827), .I3(n2826), 
            .O(n52184));
    defparam i1_4_lut_adj_1835.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1836 (.I0(n2814), .I1(n2815), .I2(n2824), .I3(n2828), 
            .O(n52208));
    defparam i1_4_lut_adj_1836.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i14_1_lut (.I0(encoder1_position_scaled[13]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n12_adj_5511));   // verilog/TinyFPGA_B.v(324[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i2_3_lut_adj_1837 (.I0(delay_counter[17]), .I1(delay_counter[16]), 
            .I2(delay_counter[15]), .I3(GND_net), .O(n27113));
    defparam i2_3_lut_adj_1837.LUT_INIT = 16'hfefe;
    SB_LUT4 i4655_4_lut (.I0(n27119), .I1(delay_counter[11]), .I2(delay_counter[10]), 
            .I3(delay_counter[9]), .O(n24_adj_5602));
    defparam i4655_4_lut.LUT_INIT = 16'hc8c0;
    SB_LUT4 i2_4_lut_adj_1838 (.I0(n24_adj_5602), .I1(delay_counter[14]), 
            .I2(delay_counter[12]), .I3(delay_counter[13]), .O(n51076));
    defparam i2_4_lut_adj_1838.LUT_INIT = 16'hc800;
    SB_LUT4 i2_3_lut_adj_1839 (.I0(n51076), .I1(delay_counter[18]), .I2(n27113), 
            .I3(GND_net), .O(n51321));
    defparam i2_3_lut_adj_1839.LUT_INIT = 16'hfefe;
    SB_DFF \ID_READOUT_FSM.state__i0  (.Q(\ID_READOUT_FSM.state [0]), .C(clk16MHz), 
           .D(n29856));   // verilog/TinyFPGA_B.v(368[10] 396[6])
    SB_LUT4 i23217_3_lut (.I0(n539), .I1(n2832), .I2(n2833), .I3(GND_net), 
            .O(n37306));
    defparam i23217_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 unary_minus_19_add_3_15_lut (.I0(GND_net), .I1(GND_net), .I2(n2), 
            .I3(n43922), .O(n330)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_19_add_3_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1840 (.I0(n2817), .I1(n2818), .I2(n52184), .I3(n52182), 
            .O(n52190));
    defparam i1_4_lut_adj_1840.LUT_INIT = 16'hfffe;
    SB_LUT4 unary_minus_18_inv_0_i22_1_lut (.I0(duty[21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_5446));   // verilog/TinyFPGA_B.v(119[24:29])
    defparam unary_minus_18_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_19_add_3_14_lut (.I0(GND_net), .I1(GND_net), .I2(n2), 
            .I3(n43921), .O(n334)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_19_add_3_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_unary_minus_2_inv_0_i28_1_lut (.I0(encoder0_position_scaled_23__N_327[27]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n6_adj_5615));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_unary_minus_2_inv_0_i28_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY unary_minus_19_add_3_14 (.CI(n43921), .I0(GND_net), .I1(n2), 
            .CO(n43922));
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i15_1_lut (.I0(encoder1_position_scaled[14]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n11_adj_5512));   // verilog/TinyFPGA_B.v(324[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_19_add_3_13_lut (.I0(GND_net), .I1(GND_net), .I2(n14_adj_5453), 
            .I3(n43920), .O(n335)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_19_add_3_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_19_add_3_13 (.CI(n43920), .I0(GND_net), .I1(n14_adj_5453), 
            .CO(n43921));
    SB_LUT4 i2_4_lut_adj_1841 (.I0(delay_counter[23]), .I1(n51321), .I2(delay_counter[20]), 
            .I3(delay_counter[19]), .O(n7_adj_5655));
    defparam i2_4_lut_adj_1841.LUT_INIT = 16'heaaa;
    SB_LUT4 i1_4_lut_adj_1842 (.I0(n2829), .I1(n37306), .I2(n2830), .I3(n2831), 
            .O(n50130));
    defparam i1_4_lut_adj_1842.LUT_INIT = 16'ha080;
    SB_LUT4 unary_minus_19_add_3_12_lut (.I0(GND_net), .I1(GND_net), .I2(n15_adj_5454), 
            .I3(n43919), .O(n336)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_19_add_3_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_19_add_3_12 (.CI(n43919), .I0(GND_net), .I1(n15_adj_5454), 
            .CO(n43920));
    SB_LUT4 i1_4_lut_adj_1843 (.I0(n2811), .I1(n2812), .I2(n2813), .I3(n52208), 
            .O(n52214));
    defparam i1_4_lut_adj_1843.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i16_1_lut (.I0(encoder1_position_scaled[15]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n10_adj_5513));   // verilog/TinyFPGA_B.v(324[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_19_add_3_11_lut (.I0(GND_net), .I1(GND_net), .I2(n16_adj_5455), 
            .I3(n43918), .O(n337)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_19_add_3_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_19_add_3_11 (.CI(n43918), .I0(GND_net), .I1(n16_adj_5455), 
            .CO(n43919));
    SB_LUT4 unary_minus_19_add_3_10_lut (.I0(GND_net), .I1(GND_net), .I2(n17_adj_5456), 
            .I3(n43917), .O(n338)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_19_add_3_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_unary_minus_2_inv_0_i29_1_lut (.I0(encoder0_position_scaled_23__N_327[28]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n5_adj_5614));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_unary_minus_2_inv_0_i29_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i17_1_lut (.I0(encoder1_position_scaled[16]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n9_adj_5514));   // verilog/TinyFPGA_B.v(324[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i4_4_lut_adj_1844 (.I0(n7_adj_5655), .I1(delay_counter[21]), 
            .I2(delay_counter[22]), .I3(n27116), .O(n62));
    defparam i4_4_lut_adj_1844.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_unary_minus_2_inv_0_i30_1_lut (.I0(encoder0_position_scaled_23__N_327[29]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n4_adj_5613));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_unary_minus_2_inv_0_i30_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1570_17 (.CI(n44176), 
            .I0(n2319), .I1(VCC_net), .CO(n44177));
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i18_1_lut (.I0(encoder1_position_scaled[17]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n8_adj_5515));   // verilog/TinyFPGA_B.v(324[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i5782_3_lut (.I0(n62), .I1(\ID_READOUT_FSM.state [0]), .I2(delay_counter[31]), 
            .I3(GND_net), .O(n21005));
    defparam i5782_3_lut.LUT_INIT = 16'hcece;
    SB_LUT4 i1_2_lut_adj_1845 (.I0(delay_counter[12]), .I1(delay_counter[11]), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_5603));
    defparam i1_2_lut_adj_1845.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_1846 (.I0(n2809), .I1(n50130), .I2(n2816), .I3(n52190), 
            .O(n52196));
    defparam i1_4_lut_adj_1846.LUT_INIT = 16'hfffe;
    SB_CARRY unary_minus_19_add_3_10 (.CI(n43917), .I0(GND_net), .I1(n17_adj_5456), 
            .CO(n43918));
    SB_LUT4 i15823_3_lut (.I0(\PID_CONTROLLER.integral [13]), .I1(\PID_CONTROLLER.integral_23__N_3996 [13]), 
            .I2(control_update), .I3(GND_net), .O(n29903));   // verilog/motorControl.v(41[14] 61[8])
    defparam i15823_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_261_6_lut (.I0(current[4]), .I1(duty[7]), .I2(n56614), 
            .I3(n43561), .O(n266)) /* synthesis syn_instantiated=1 */ ;
    defparam add_261_6_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1570_16_lut (.I0(GND_net), 
            .I1(n2320), .I2(VCC_net), .I3(n44175), .O(n2387)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1570_16_lut.LUT_INIT = 16'hC33C;
    SB_DFF commutation_state_prev_i1 (.Q(commutation_state_prev[1]), .C(clk16MHz), 
           .D(commutation_state[1]));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    SB_DFF pwm_setpoint_i23 (.Q(pwm_setpoint[23]), .C(clk16MHz), .D(pwm_setpoint_23__N_11[23]));   // verilog/TinyFPGA_B.v(103[9] 129[5])
    SB_DFFESR delay_counter_i0_i0 (.Q(delay_counter[0]), .C(clk16MHz), .E(n7593), 
            .D(n1563), .R(n29242));   // verilog/TinyFPGA_B.v(368[10] 396[6])
    SB_DFF pwm_setpoint_i22 (.Q(pwm_setpoint[22]), .C(clk16MHz), .D(pwm_setpoint_23__N_11[22]));   // verilog/TinyFPGA_B.v(103[9] 129[5])
    SB_DFF dti_counter_2279__i0 (.Q(dti_counter[0]), .C(clk16MHz), .D(n55));   // verilog/TinyFPGA_B.v(174[23:37])
    SB_LUT4 i15824_3_lut (.I0(\PID_CONTROLLER.integral [12]), .I1(\PID_CONTROLLER.integral_23__N_3996 [12]), 
            .I2(control_update), .I3(GND_net), .O(n29904));   // verilog/motorControl.v(41[14] 61[8])
    defparam i15824_3_lut.LUT_INIT = 16'hcaca;
    GND i1 (.Y(GND_net));
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i19_1_lut (.I0(encoder1_position_scaled[18]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n7_adj_5516));   // verilog/TinyFPGA_B.v(324[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i15825_3_lut (.I0(\PID_CONTROLLER.integral [11]), .I1(\PID_CONTROLLER.integral_23__N_3996 [11]), 
            .I2(control_update), .I3(GND_net), .O(n29905));   // verilog/motorControl.v(41[14] 61[8])
    defparam i15825_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i20_1_lut (.I0(encoder1_position_scaled[19]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n6_adj_5517));   // verilog/TinyFPGA_B.v(324[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i40228_4_lut (.I0(n52196), .I1(n2808), .I2(n52214), .I3(n2810), 
            .O(n2841));
    defparam i40228_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 unary_minus_19_add_3_9_lut (.I0(GND_net), .I1(GND_net), .I2(n18_adj_5457), 
            .I3(n43916), .O(n339)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_19_add_3_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1570_16 (.CI(n44175), 
            .I0(n2320), .I1(VCC_net), .CO(n44176));
    SB_CARRY unary_minus_19_add_3_9 (.CI(n43916), .I0(GND_net), .I1(n18_adj_5457), 
            .CO(n43917));
    SB_LUT4 unary_minus_19_add_3_8_lut (.I0(GND_net), .I1(GND_net), .I2(n19_adj_5458), 
            .I3(n43915), .O(n340)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_19_add_3_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_261_6 (.CI(n43561), .I0(duty[7]), .I1(n56614), .CO(n43562));
    SB_CARRY unary_minus_19_add_3_8 (.CI(n43915), .I0(GND_net), .I1(n19_adj_5458), 
            .CO(n43916));
    SB_LUT4 unary_minus_19_add_3_7_lut (.I0(GND_net), .I1(GND_net), .I2(n20_adj_5459), 
            .I3(n43914), .O(n341)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_19_add_3_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_19_add_3_7 (.CI(n43914), .I0(GND_net), .I1(n20_adj_5459), 
            .CO(n43915));
    SB_DFF pwm_setpoint_i21 (.Q(pwm_setpoint[21]), .C(clk16MHz), .D(pwm_setpoint_23__N_11[21]));   // verilog/TinyFPGA_B.v(103[9] 129[5])
    SB_DFF pwm_setpoint_i20 (.Q(pwm_setpoint[20]), .C(clk16MHz), .D(pwm_setpoint_23__N_11[20]));   // verilog/TinyFPGA_B.v(103[9] 129[5])
    SB_LUT4 unary_minus_19_add_3_6_lut (.I0(GND_net), .I1(GND_net), .I2(n21_adj_5460), 
            .I3(n43913), .O(n342)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_19_add_3_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_19_add_3_6 (.CI(n43913), .I0(GND_net), .I1(n21_adj_5460), 
            .CO(n43914));
    SB_LUT4 unary_minus_19_add_3_5_lut (.I0(GND_net), .I1(GND_net), .I2(n22_adj_5461), 
            .I3(n43912), .O(n343)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_19_add_3_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_19_add_3_5 (.CI(n43912), .I0(GND_net), .I1(n22_adj_5461), 
            .CO(n43913));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1570_15_lut (.I0(GND_net), 
            .I1(n2321), .I2(VCC_net), .I3(n44174), .O(n2388)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1570_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1570_15 (.CI(n44174), 
            .I0(n2321), .I1(VCC_net), .CO(n44175));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1570_14_lut (.I0(GND_net), 
            .I1(n2322), .I2(VCC_net), .I3(n44173), .O(n2389)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1570_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_19_add_3_4_lut (.I0(GND_net), .I1(GND_net), .I2(n23_adj_5462), 
            .I3(n43911), .O(n344)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_19_add_3_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_19_add_3_4 (.CI(n43911), .I0(GND_net), .I1(n23_adj_5462), 
            .CO(n43912));
    SB_DFF pwm_setpoint_i19 (.Q(pwm_setpoint[19]), .C(clk16MHz), .D(pwm_setpoint_23__N_11[19]));   // verilog/TinyFPGA_B.v(103[9] 129[5])
    SB_DFF pwm_setpoint_i18 (.Q(pwm_setpoint[18]), .C(clk16MHz), .D(pwm_setpoint_23__N_11[18]));   // verilog/TinyFPGA_B.v(103[9] 129[5])
    SB_DFF pwm_setpoint_i17 (.Q(pwm_setpoint[17]), .C(clk16MHz), .D(pwm_setpoint_23__N_11[17]));   // verilog/TinyFPGA_B.v(103[9] 129[5])
    SB_DFF pwm_setpoint_i16 (.Q(pwm_setpoint[16]), .C(clk16MHz), .D(pwm_setpoint_23__N_11[16]));   // verilog/TinyFPGA_B.v(103[9] 129[5])
    SB_DFF pwm_setpoint_i15 (.Q(pwm_setpoint[15]), .C(clk16MHz), .D(pwm_setpoint_23__N_11[15]));   // verilog/TinyFPGA_B.v(103[9] 129[5])
    SB_DFF pwm_setpoint_i14 (.Q(pwm_setpoint[14]), .C(clk16MHz), .D(pwm_setpoint_23__N_11[14]));   // verilog/TinyFPGA_B.v(103[9] 129[5])
    SB_DFF pwm_setpoint_i13 (.Q(pwm_setpoint[13]), .C(clk16MHz), .D(pwm_setpoint_23__N_11[13]));   // verilog/TinyFPGA_B.v(103[9] 129[5])
    SB_DFF pwm_setpoint_i12 (.Q(pwm_setpoint[12]), .C(clk16MHz), .D(pwm_setpoint_23__N_11[12]));   // verilog/TinyFPGA_B.v(103[9] 129[5])
    SB_DFF pwm_setpoint_i11 (.Q(pwm_setpoint[11]), .C(clk16MHz), .D(pwm_setpoint_23__N_11[11]));   // verilog/TinyFPGA_B.v(103[9] 129[5])
    SB_DFF pwm_setpoint_i10 (.Q(pwm_setpoint[10]), .C(clk16MHz), .D(pwm_setpoint_23__N_11[10]));   // verilog/TinyFPGA_B.v(103[9] 129[5])
    SB_DFF pwm_setpoint_i9 (.Q(pwm_setpoint[9]), .C(clk16MHz), .D(pwm_setpoint_23__N_11[9]));   // verilog/TinyFPGA_B.v(103[9] 129[5])
    SB_DFF pwm_setpoint_i8 (.Q(pwm_setpoint[8]), .C(clk16MHz), .D(pwm_setpoint_23__N_11[8]));   // verilog/TinyFPGA_B.v(103[9] 129[5])
    SB_DFF pwm_setpoint_i7 (.Q(pwm_setpoint[7]), .C(clk16MHz), .D(pwm_setpoint_23__N_11[7]));   // verilog/TinyFPGA_B.v(103[9] 129[5])
    SB_DFF pwm_setpoint_i6 (.Q(pwm_setpoint[6]), .C(clk16MHz), .D(pwm_setpoint_23__N_11[6]));   // verilog/TinyFPGA_B.v(103[9] 129[5])
    SB_DFF pwm_setpoint_i5 (.Q(pwm_setpoint[5]), .C(clk16MHz), .D(pwm_setpoint_23__N_11[5]));   // verilog/TinyFPGA_B.v(103[9] 129[5])
    SB_DFF pwm_setpoint_i4 (.Q(pwm_setpoint[4]), .C(clk16MHz), .D(pwm_setpoint_23__N_11[4]));   // verilog/TinyFPGA_B.v(103[9] 129[5])
    SB_LUT4 i1_4_lut_adj_1847 (.I0(n1029), .I1(n37346), .I2(n1030), .I3(n1031), 
            .O(n50003));
    defparam i1_4_lut_adj_1847.LUT_INIT = 16'ha080;
    SB_DFF pwm_setpoint_i3 (.Q(pwm_setpoint[3]), .C(clk16MHz), .D(pwm_setpoint_23__N_11[3]));   // verilog/TinyFPGA_B.v(103[9] 129[5])
    SB_LUT4 i40630_4_lut (.I0(n1026), .I1(n50003), .I2(n1027), .I3(n1028), 
            .O(n1059));
    defparam i40630_4_lut.LUT_INIT = 16'h0001;
    SB_DFF pwm_setpoint_i2 (.Q(pwm_setpoint[2]), .C(clk16MHz), .D(pwm_setpoint_23__N_11[2]));   // verilog/TinyFPGA_B.v(103[9] 129[5])
    SB_LUT4 encoder0_position_scaled_23__I_0_227_mux_3_i24_3_lut (.I0(encoder0_position_scaled_23__N_327[23]), 
            .I1(n10_adj_5489), .I2(encoder0_position_scaled_23__N_327[31]), 
            .I3(GND_net), .O(n935));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_mux_3_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF pwm_setpoint_i1 (.Q(pwm_setpoint[1]), .C(clk16MHz), .D(pwm_setpoint_23__N_11[1]));   // verilog/TinyFPGA_B.v(103[9] 129[5])
    SB_LUT4 i23322_4_lut (.I0(n411), .I1(n1131), .I2(n1132), .I3(n1133), 
            .O(n37412));
    defparam i23322_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 i1_3_lut_adj_1848 (.I0(n1126), .I1(n1127), .I2(n1128), .I3(GND_net), 
            .O(n51780));
    defparam i1_3_lut_adj_1848.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_2_lut_adj_1849 (.I0(n1129), .I1(n1130), .I2(GND_net), .I3(GND_net), 
            .O(n51914));
    defparam i1_2_lut_adj_1849.LUT_INIT = 16'h8888;
    SB_LUT4 i40617_4_lut (.I0(n51914), .I1(n1125), .I2(n51780), .I3(n37412), 
            .O(n1158));
    defparam i40617_4_lut.LUT_INIT = 16'h0103;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_unary_minus_2_inv_0_i31_1_lut (.I0(encoder0_position_scaled_23__N_327[30]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n3_adj_5612));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_unary_minus_2_inv_0_i31_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i709_rep_55_3_lut (.I0(n935), 
            .I1(n1101), .I2(n1059), .I3(GND_net), .O(n1133));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i709_rep_55_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i777_3_lut (.I0(n411), .I1(n1201), 
            .I2(n1158), .I3(GND_net), .O(n1233));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i777_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i776_3_lut (.I0(n1133), .I1(n1200), 
            .I2(n1158), .I3(GND_net), .O(n1232));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i776_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 n10829_bdd_4_lut_40989 (.I0(n10829), .I1(n421), .I2(current[15]), 
            .I3(duty[23]), .O(n56814));
    defparam n10829_bdd_4_lut_40989.LUT_INIT = 16'he4aa;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i772_3_lut (.I0(n1129), .I1(n1196), 
            .I2(n1158), .I3(GND_net), .O(n1228));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i772_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 n56814_bdd_4_lut (.I0(n56814), .I1(duty[20]), .I2(n250), .I3(duty[23]), 
            .O(pwm_setpoint_23__N_11[20]));
    defparam n56814_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i771_3_lut (.I0(n1128), .I1(n1195), 
            .I2(n1158), .I3(GND_net), .O(n1227));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i771_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i770_3_lut (.I0(n1127), .I1(n1194), 
            .I2(n1158), .I3(GND_net), .O(n1226));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i770_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 n10829_bdd_4_lut_40949 (.I0(n10829), .I1(n422), .I2(current[15]), 
            .I3(duty[23]), .O(n56808));
    defparam n10829_bdd_4_lut_40949.LUT_INIT = 16'he4aa;
    SB_LUT4 i23252_3_lut (.I0(n412), .I1(n1232), .I2(n1233), .I3(GND_net), 
            .O(n37342));
    defparam i23252_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 n56808_bdd_4_lut (.I0(n56808), .I1(duty[19]), .I2(n251), .I3(duty[23]), 
            .O(pwm_setpoint_23__N_11[19]));
    defparam n56808_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_3_lut_adj_1850 (.I0(n1226), .I1(n1227), .I2(n1228), .I3(GND_net), 
            .O(n51918));
    defparam i1_3_lut_adj_1850.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_4_lut_adj_1851 (.I0(n1229), .I1(n37342), .I2(n1230), .I3(n1231), 
            .O(n49998));
    defparam i1_4_lut_adj_1851.LUT_INIT = 16'ha080;
    SB_LUT4 n10829_bdd_4_lut_40944 (.I0(n10829), .I1(n423), .I2(current[15]), 
            .I3(duty[23]), .O(n56802));
    defparam n10829_bdd_4_lut_40944.LUT_INIT = 16'he4aa;
    SB_LUT4 i40603_4_lut (.I0(n1225), .I1(n1224), .I2(n49998), .I3(n51918), 
            .O(n1257));
    defparam i40603_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 n56802_bdd_4_lut (.I0(n56802), .I1(duty[18]), .I2(n252), .I3(duty[23]), 
            .O(pwm_setpoint_23__N_11[18]));
    defparam n56802_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_mux_3_i22_3_lut (.I0(encoder0_position_scaled_23__N_327[21]), 
            .I1(n12_adj_5487), .I2(encoder0_position_scaled_23__N_327[31]), 
            .I3(GND_net), .O(n412));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_mux_3_i22_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i845_rep_53_3_lut (.I0(n412), 
            .I1(n1301), .I2(n1257), .I3(GND_net), .O(n1333));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i845_rep_53_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_mux_3_i21_3_lut (.I0(encoder0_position_scaled_23__N_327[20]), 
            .I1(n13_adj_5486), .I2(encoder0_position_scaled_23__N_327[31]), 
            .I3(GND_net), .O(n413));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_mux_3_i21_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i23250_3_lut (.I0(n413), .I1(n1332), .I2(n1333), .I3(GND_net), 
            .O(n37340));
    defparam i23250_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i1_4_lut_adj_1852 (.I0(n1325), .I1(n1326), .I2(n1327), .I3(n1328), 
            .O(n51842));
    defparam i1_4_lut_adj_1852.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1853 (.I0(n1329), .I1(n37340), .I2(n1330), .I3(n1331), 
            .O(n49995));
    defparam i1_4_lut_adj_1853.LUT_INIT = 16'ha080;
    SB_LUT4 n10829_bdd_4_lut_40939 (.I0(n10829), .I1(n424), .I2(current[15]), 
            .I3(duty[23]), .O(n56784));
    defparam n10829_bdd_4_lut_40939.LUT_INIT = 16'he4aa;
    SB_LUT4 unary_minus_19_add_3_3_lut (.I0(GND_net), .I1(GND_net), .I2(n24_adj_5463), 
            .I3(n43910), .O(n345)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_19_add_3_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i2_4_lut_adj_1854 (.I0(delay_counter[9]), .I1(n4_adj_5603), 
            .I2(delay_counter[10]), .I3(n27119), .O(n50770));
    defparam i2_4_lut_adj_1854.LUT_INIT = 16'hfcec;
    SB_CARRY unary_minus_19_add_3_3 (.CI(n43910), .I0(GND_net), .I1(n24_adj_5463), 
            .CO(n43911));
    SB_LUT4 unary_minus_18_inv_0_i23_1_lut (.I0(duty[22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n3));   // verilog/TinyFPGA_B.v(119[24:29])
    defparam unary_minus_18_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i21_1_lut (.I0(encoder1_position_scaled[20]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n5_adj_5518));   // verilog/TinyFPGA_B.v(324[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i15826_3_lut (.I0(\PID_CONTROLLER.integral [10]), .I1(\PID_CONTROLLER.integral_23__N_3996 [10]), 
            .I2(control_update), .I3(GND_net), .O(n29906));   // verilog/motorControl.v(41[14] 61[8])
    defparam i15826_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_19_add_3_2_lut (.I0(n25), .I1(GND_net), .I2(n25_adj_5464), 
            .I3(VCC_net), .O(n54539)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_19_add_3_2_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i15827_3_lut (.I0(\PID_CONTROLLER.integral [9]), .I1(\PID_CONTROLLER.integral_23__N_3996 [9]), 
            .I2(control_update), .I3(GND_net), .O(n29907));   // verilog/motorControl.v(41[14] 61[8])
    defparam i15827_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY unary_minus_19_add_3_2 (.CI(VCC_net), .I0(GND_net), .I1(n25_adj_5464), 
            .CO(n43910));
    SB_LUT4 add_5094_32_lut (.I0(GND_net), .I1(encoder0_position[31]), .I2(VCC_net), 
            .I3(n43909), .O(encoder0_position_scaled_23__N_327[31])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5094_32_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i22_1_lut (.I0(encoder1_position_scaled[21]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n4_adj_5519));   // verilog/TinyFPGA_B.v(324[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 n56784_bdd_4_lut (.I0(n56784), .I1(duty[17]), .I2(n253), .I3(duty[23]), 
            .O(pwm_setpoint_23__N_11[17]));
    defparam n56784_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n10829_bdd_4_lut_40925 (.I0(n10829), .I1(n425), .I2(current[15]), 
            .I3(duty[23]), .O(n56778));
    defparam n10829_bdd_4_lut_40925.LUT_INIT = 16'he4aa;
    SB_LUT4 n56778_bdd_4_lut (.I0(n56778), .I1(duty[16]), .I2(n254), .I3(duty[23]), 
            .O(pwm_setpoint_23__N_11[16]));
    defparam n56778_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i2_4_lut_adj_1855 (.I0(n50770), .I1(n27113), .I2(delay_counter[13]), 
            .I3(delay_counter[14]), .O(n51014));
    defparam i2_4_lut_adj_1855.LUT_INIT = 16'hffec;
    SB_LUT4 n10829_bdd_4_lut_40920 (.I0(n10829), .I1(n426), .I2(current[15]), 
            .I3(duty[23]), .O(n56772));
    defparam n10829_bdd_4_lut_40920.LUT_INIT = 16'he4aa;
    SB_LUT4 n56772_bdd_4_lut (.I0(n56772), .I1(duty[15]), .I2(n255), .I3(duty[23]), 
            .O(pwm_setpoint_23__N_11[15]));
    defparam n56772_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i15828_3_lut (.I0(\PID_CONTROLLER.integral [8]), .I1(\PID_CONTROLLER.integral_23__N_3996 [8]), 
            .I2(control_update), .I3(GND_net), .O(n29908));   // verilog/motorControl.v(41[14] 61[8])
    defparam i15828_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n10829_bdd_4_lut_40915 (.I0(n10829), .I1(n427), .I2(current[15]), 
            .I3(duty[23]), .O(n56766));
    defparam n10829_bdd_4_lut_40915.LUT_INIT = 16'he4aa;
    SB_LUT4 n56766_bdd_4_lut (.I0(n56766), .I1(duty[14]), .I2(n256), .I3(duty[23]), 
            .O(pwm_setpoint_23__N_11[14]));
    defparam n56766_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n10829_bdd_4_lut_40910 (.I0(n10829), .I1(n428), .I2(current[15]), 
            .I3(duty[23]), .O(n56760));
    defparam n10829_bdd_4_lut_40910.LUT_INIT = 16'he4aa;
    SB_LUT4 i3_3_lut (.I0(delay_counter[20]), .I1(delay_counter[21]), .I2(delay_counter[23]), 
            .I3(GND_net), .O(n8));
    defparam i3_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 n56760_bdd_4_lut (.I0(n56760), .I1(duty[13]), .I2(n257), .I3(duty[23]), 
            .O(pwm_setpoint_23__N_11[13]));
    defparam n56760_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n10829_bdd_4_lut_40905 (.I0(n10829), .I1(n429), .I2(current[15]), 
            .I3(duty[23]), .O(n56754));
    defparam n10829_bdd_4_lut_40905.LUT_INIT = 16'he4aa;
    SB_LUT4 n56754_bdd_4_lut (.I0(n56754), .I1(duty[12]), .I2(n258), .I3(duty[23]), 
            .O(pwm_setpoint_23__N_11[12]));
    defparam n56754_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i2_4_lut_adj_1856 (.I0(delay_counter[22]), .I1(n51014), .I2(delay_counter[19]), 
            .I3(delay_counter[18]), .O(n7));
    defparam i2_4_lut_adj_1856.LUT_INIT = 16'ha8a0;
    SB_LUT4 i22581_4_lut (.I0(n7), .I1(delay_counter[31]), .I2(n27116), 
            .I3(n8), .O(n1650));   // verilog/TinyFPGA_B.v(389[14:38])
    defparam i22581_4_lut.LUT_INIT = 16'h3230;
    SB_LUT4 i40533_1_lut (.I0(n1653), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n56364));
    defparam i40533_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 n10829_bdd_4_lut_40900 (.I0(n10829), .I1(n430), .I2(current[11]), 
            .I3(duty[23]), .O(n56736));
    defparam n10829_bdd_4_lut_40900.LUT_INIT = 16'he4aa;
    SB_LUT4 n56736_bdd_4_lut (.I0(n56736), .I1(duty[11]), .I2(n259), .I3(duty[23]), 
            .O(pwm_setpoint_23__N_11[11]));
    defparam n56736_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n10829_bdd_4_lut_40886 (.I0(n10829), .I1(n431), .I2(current[10]), 
            .I3(duty[23]), .O(n56730));
    defparam n10829_bdd_4_lut_40886.LUT_INIT = 16'he4aa;
    SB_LUT4 n56730_bdd_4_lut (.I0(n56730), .I1(duty[10]), .I2(n260), .I3(duty[23]), 
            .O(pwm_setpoint_23__N_11[10]));
    defparam n56730_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n10829_bdd_4_lut_40881 (.I0(n10829), .I1(n432), .I2(current[9]), 
            .I3(duty[23]), .O(n56724));
    defparam n10829_bdd_4_lut_40881.LUT_INIT = 16'he4aa;
    SB_LUT4 n56724_bdd_4_lut (.I0(n56724), .I1(duty[9]), .I2(n261), .I3(duty[23]), 
            .O(pwm_setpoint_23__N_11[9]));
    defparam n56724_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1774_3_lut (.I0(n2611), 
            .I1(n2678), .I2(n2643), .I3(GND_net), .O(n2710));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1774_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1776_3_lut (.I0(n2613), 
            .I1(n2680), .I2(n2643), .I3(GND_net), .O(n2712));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1776_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1775_3_lut (.I0(n2612), 
            .I1(n2679), .I2(n2643), .I3(GND_net), .O(n2711));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1775_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i40255_1_lut (.I0(n2742), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n56086));
    defparam i40255_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_3_lut_adj_1857 (.I0(n2722), .I1(n2726), .I2(n2724), .I3(GND_net), 
            .O(n52066));
    defparam i1_3_lut_adj_1857.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_4_lut_adj_1858 (.I0(n52066), .I1(n2720), .I2(n2728), .I3(n2725), 
            .O(n52070));
    defparam i1_4_lut_adj_1858.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_2_lut_adj_1859 (.I0(ID[2]), .I1(ID[4]), .I2(GND_net), .I3(GND_net), 
            .O(n10_adj_5530));   // verilog/TinyFPGA_B.v(387[12:17])
    defparam i2_2_lut_adj_1859.LUT_INIT = 16'heeee;
    SB_LUT4 i6_4_lut_adj_1860 (.I0(ID[7]), .I1(ID[5]), .I2(ID[1]), .I3(ID[0]), 
            .O(n14_adj_5529));   // verilog/TinyFPGA_B.v(387[12:17])
    defparam i6_4_lut_adj_1860.LUT_INIT = 16'hfffe;
    SB_LUT4 i1021_1_lut (.I0(n296), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n4748));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam i1021_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1570_14 (.CI(n44173), 
            .I0(n2322), .I1(VCC_net), .CO(n44174));
    SB_LUT4 i1_2_lut_adj_1861 (.I0(n2723), .I1(n2727), .I2(GND_net), .I3(GND_net), 
            .O(n51712));
    defparam i1_2_lut_adj_1861.LUT_INIT = 16'heeee;
    SB_LUT4 i7_4_lut_adj_1862 (.I0(ID[3]), .I1(n14_adj_5529), .I2(n10_adj_5530), 
            .I3(ID[6]), .O(n27093));   // verilog/TinyFPGA_B.v(387[12:17])
    defparam i7_4_lut_adj_1862.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1570_13_lut (.I0(GND_net), 
            .I1(n2323), .I2(VCC_net), .I3(n44172), .O(n2390)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1570_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i23219_3_lut (.I0(n538), .I1(n2732), .I2(n2733), .I3(GND_net), 
            .O(n37308));
    defparam i23219_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i1_4_lut_adj_1863 (.I0(n2729), .I1(n37308), .I2(n2730), .I3(n2731), 
            .O(n50081));
    defparam i1_4_lut_adj_1863.LUT_INIT = 16'ha080;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i23_1_lut (.I0(encoder1_position_scaled[22]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n3_adj_5520));   // verilog/TinyFPGA_B.v(324[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_4_lut_adj_1864 (.I0(n2718), .I1(n51712), .I2(n2717), .I3(n52070), 
            .O(n51714));
    defparam i1_4_lut_adj_1864.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1865 (.I0(n2716), .I1(n51714), .I2(n2715), .I3(n50081), 
            .O(n51716));
    defparam i1_4_lut_adj_1865.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i24_1_lut (.I0(encoder1_position_scaled[23]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n2_adj_5521));   // verilog/TinyFPGA_B.v(324[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i15191_4_lut (.I0(n7593), .I1(n1650), .I2(n21005), .I3(n27094), 
            .O(n29242));   // verilog/TinyFPGA_B.v(368[10] 396[6])
    defparam i15191_4_lut.LUT_INIT = 16'ha088;
    SB_LUT4 i1_4_lut_adj_1866 (.I0(n2711), .I1(n2713), .I2(n51716), .I3(n2714), 
            .O(n51722));
    defparam i1_4_lut_adj_1866.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_3_lut_adj_1867 (.I0(n2712), .I1(n2719), .I2(n2721), .I3(GND_net), 
            .O(n51610));
    defparam i1_3_lut_adj_1867.LUT_INIT = 16'hfefe;
    SB_LUT4 i40258_4_lut (.I0(n2709), .I1(n51610), .I2(n51722), .I3(n2710), 
            .O(n2742));
    defparam i40258_4_lut.LUT_INIT = 16'h0001;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1570_13 (.CI(n44172), 
            .I0(n2323), .I1(VCC_net), .CO(n44173));
    SB_LUT4 add_5094_31_lut (.I0(GND_net), .I1(encoder0_position[30]), .I2(VCC_net), 
            .I3(n43908), .O(encoder0_position_scaled_23__N_327[30])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5094_31_lut.LUT_INIT = 16'hC33C;
    SB_IO NEOPXL_pad (.PACKAGE_PIN(NEOPXL), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(NEOPXL_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam NEOPXL_pad.PIN_TYPE = 6'b011001;
    defparam NEOPXL_pad.PULLUP = 1'b0;
    defparam NEOPXL_pad.NEG_TRIGGER = 1'b0;
    defparam NEOPXL_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO USBPU_pad (.PACKAGE_PIN(USBPU), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(GND_net));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam USBPU_pad.PIN_TYPE = 6'b011001;
    defparam USBPU_pad.PULLUP = 1'b0;
    defparam USBPU_pad.NEG_TRIGGER = 1'b0;
    defparam USBPU_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO LED_pad (.PACKAGE_PIN(LED), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(LED_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam LED_pad.PIN_TYPE = 6'b011001;
    defparam LED_pad.PULLUP = 1'b0;
    defparam LED_pad.NEG_TRIGGER = 1'b0;
    defparam LED_pad.IO_STANDARD = "SB_LVCMOS";
    SB_CARRY add_5094_31 (.CI(n43908), .I0(encoder0_position[30]), .I1(VCC_net), 
            .CO(n43909));
    SB_DFFESR GHC_214 (.Q(GHC), .C(clk16MHz), .E(n28672), .D(GHC_N_514), 
            .R(n29145));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1570_12_lut (.I0(GND_net), 
            .I1(n2324), .I2(VCC_net), .I3(n44171), .O(n2391)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1570_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1570_12 (.CI(n44171), 
            .I0(n2324), .I1(VCC_net), .CO(n44172));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1570_11_lut (.I0(GND_net), 
            .I1(n2325), .I2(VCC_net), .I3(n44170), .O(n2392)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1570_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5094_30_lut (.I0(GND_net), .I1(encoder0_position[29]), .I2(VCC_net), 
            .I3(n43907), .O(encoder0_position_scaled_23__N_327[29])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5094_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1570_11 (.CI(n44170), 
            .I0(n2325), .I1(VCC_net), .CO(n44171));
    SB_LUT4 mux_281_i1_4_lut (.I0(encoder1_position_scaled[0]), .I1(displacement[0]), 
            .I2(n15), .I3(n15_adj_5471), .O(motor_state_23__N_123[0]));   // verilog/TinyFPGA_B.v(284[5] 286[10])
    defparam mux_281_i1_4_lut.LUT_INIT = 16'h0aca;
    SB_CARRY add_5094_30 (.CI(n43907), .I0(encoder0_position[29]), .I1(VCC_net), 
            .CO(n43908));
    SB_LUT4 add_5094_29_lut (.I0(GND_net), .I1(encoder0_position[28]), .I2(VCC_net), 
            .I3(n43906), .O(encoder0_position_scaled_23__N_327[28])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5094_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5094_29 (.CI(n43906), .I0(encoder0_position[28]), .I1(VCC_net), 
            .CO(n43907));
    SB_LUT4 add_5094_28_lut (.I0(GND_net), .I1(encoder0_position[27]), .I2(VCC_net), 
            .I3(n43905), .O(encoder0_position_scaled_23__N_327[27])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5094_28_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1570_10_lut (.I0(GND_net), 
            .I1(n2326), .I2(VCC_net), .I3(n44169), .O(n2393)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1570_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1570_10 (.CI(n44169), 
            .I0(n2326), .I1(VCC_net), .CO(n44170));
    SB_CARRY add_5094_28 (.CI(n43905), .I0(encoder0_position[27]), .I1(VCC_net), 
            .CO(n43906));
    SB_LUT4 add_5094_27_lut (.I0(GND_net), .I1(encoder0_position[26]), .I2(VCC_net), 
            .I3(n43904), .O(encoder0_position_scaled_23__N_327[26])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5094_27_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i907_3_lut (.I0(n1328), .I1(n1395), 
            .I2(n1356), .I3(GND_net), .O(n1427));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i907_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i974_3_lut (.I0(n1427), .I1(n1494), 
            .I2(n1455), .I3(GND_net), .O(n1526));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i974_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1041_3_lut (.I0(n1526), 
            .I1(n1593), .I2(n1554_adj_5597), .I3(GND_net), .O(n1625));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1041_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1570_9_lut (.I0(GND_net), 
            .I1(n2327), .I2(VCC_net), .I3(n44168), .O(n2394)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1570_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5094_27 (.CI(n43904), .I0(encoder0_position[26]), .I1(VCC_net), 
            .CO(n43905));
    SB_LUT4 n10829_bdd_4_lut_40876 (.I0(n10829), .I1(n433), .I2(current[8]), 
            .I3(duty[23]), .O(n56718));
    defparam n10829_bdd_4_lut_40876.LUT_INIT = 16'he4aa;
    SB_LUT4 n56718_bdd_4_lut (.I0(n56718), .I1(duty[8]), .I2(n262), .I3(duty[23]), 
            .O(pwm_setpoint_23__N_11[8]));
    defparam n56718_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n10829_bdd_4_lut_40871 (.I0(n10829), .I1(n434), .I2(current[7]), 
            .I3(duty[23]), .O(n56706));
    defparam n10829_bdd_4_lut_40871.LUT_INIT = 16'he4aa;
    SB_LUT4 n56706_bdd_4_lut (.I0(n56706), .I1(duty[7]), .I2(n263), .I3(duty[23]), 
            .O(pwm_setpoint_23__N_11[7]));
    defparam n56706_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n10829_bdd_4_lut_40861 (.I0(n10829), .I1(n435), .I2(current[6]), 
            .I3(duty[23]), .O(n56688));
    defparam n10829_bdd_4_lut_40861.LUT_INIT = 16'he4aa;
    SB_LUT4 n56688_bdd_4_lut (.I0(n56688), .I1(duty[6]), .I2(n264), .I3(duty[23]), 
            .O(pwm_setpoint_23__N_11[6]));
    defparam n56688_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 add_5094_26_lut (.I0(GND_net), .I1(encoder0_position[25]), .I2(VCC_net), 
            .I3(n43903), .O(encoder0_position_scaled_23__N_327[25])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5094_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1108_3_lut (.I0(n1625), 
            .I1(n1692), .I2(n1653), .I3(GND_net), .O(n1724));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1108_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i40588_4_lut (.I0(n49995), .I1(n1323), .I2(n1324), .I3(n51842), 
            .O(n1356));
    defparam i40588_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1175_3_lut (.I0(n1724), 
            .I1(n1791), .I2(n1752), .I3(GND_net), .O(n1823));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1175_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1242_3_lut (.I0(n1823), 
            .I1(n1890), .I2(n1851), .I3(GND_net), .O(n1922));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1242_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_5094_26 (.CI(n43903), .I0(encoder0_position[25]), .I1(VCC_net), 
            .CO(n43904));
    SB_LUT4 mux_281_i2_4_lut (.I0(encoder1_position_scaled[1]), .I1(displacement[1]), 
            .I2(n15), .I3(n15_adj_5471), .O(motor_state_23__N_123[1]));   // verilog/TinyFPGA_B.v(284[5] 286[10])
    defparam mux_281_i2_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1309_3_lut (.I0(n1922), 
            .I1(n1989), .I2(n1950), .I3(GND_net), .O(n2021));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1309_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_5094_25_lut (.I0(GND_net), .I1(encoder0_position[24]), .I2(VCC_net), 
            .I3(n43902), .O(encoder0_position_scaled_23__N_327[24])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5094_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5094_25 (.CI(n43902), .I0(encoder0_position[24]), .I1(VCC_net), 
            .CO(n43903));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1376_3_lut (.I0(n2021), 
            .I1(n2088), .I2(n2049), .I3(GND_net), .O(n2120));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1376_3_lut.LUT_INIT = 16'hacac;
    SB_DFFESR GHB_212 (.Q(GHB), .C(clk16MHz), .E(n28672), .D(GHB_N_500), 
            .R(n29145));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1570_9 (.CI(n44168), 
            .I0(n2327), .I1(VCC_net), .CO(n44169));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1570_8_lut (.I0(GND_net), 
            .I1(n2328), .I2(VCC_net), .I3(n44167), .O(n2395)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1570_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1570_8 (.CI(n44167), 
            .I0(n2328), .I1(VCC_net), .CO(n44168));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1570_7_lut (.I0(GND_net), 
            .I1(n2329), .I2(GND_net), .I3(n44166), .O(n2396)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1570_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5094_24_lut (.I0(GND_net), .I1(encoder0_position[23]), .I2(VCC_net), 
            .I3(n43901), .O(encoder0_position_scaled_23__N_327[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5094_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5094_24 (.CI(n43901), .I0(encoder0_position[23]), .I1(VCC_net), 
            .CO(n43902));
    SB_LUT4 add_5094_23_lut (.I0(GND_net), .I1(encoder0_position[22]), .I2(VCC_net), 
            .I3(n43900), .O(encoder0_position_scaled_23__N_327[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5094_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5094_23 (.CI(n43900), .I0(encoder0_position[22]), .I1(VCC_net), 
            .CO(n43901));
    SB_LUT4 i15829_3_lut (.I0(\PID_CONTROLLER.integral [7]), .I1(\PID_CONTROLLER.integral_23__N_3996 [7]), 
            .I2(control_update), .I3(GND_net), .O(n29909));   // verilog/motorControl.v(41[14] 61[8])
    defparam i15829_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_5094_22_lut (.I0(GND_net), .I1(encoder0_position[21]), .I2(VCC_net), 
            .I3(n43899), .O(encoder0_position_scaled_23__N_327[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5094_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5094_22 (.CI(n43899), .I0(encoder0_position[21]), .I1(VCC_net), 
            .CO(n43900));
    SB_LUT4 add_5094_21_lut (.I0(GND_net), .I1(encoder0_position[20]), .I2(VCC_net), 
            .I3(n43898), .O(encoder0_position_scaled_23__N_327[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5094_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5094_21 (.CI(n43898), .I0(encoder0_position[20]), .I1(VCC_net), 
            .CO(n43899));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1570_7 (.CI(n44166), 
            .I0(n2329), .I1(GND_net), .CO(n44167));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1570_6_lut (.I0(GND_net), 
            .I1(n2330), .I2(GND_net), .I3(n44165), .O(n2397)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1570_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5094_20_lut (.I0(GND_net), .I1(encoder0_position[19]), .I2(VCC_net), 
            .I3(n43897), .O(encoder0_position_scaled_23__N_327[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5094_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5094_20 (.CI(n43897), .I0(encoder0_position[19]), .I1(VCC_net), 
            .CO(n43898));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1570_6 (.CI(n44165), 
            .I0(n2330), .I1(GND_net), .CO(n44166));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1570_5_lut (.I0(GND_net), 
            .I1(n2331), .I2(VCC_net), .I3(n44164), .O(n2398)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1570_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5094_19_lut (.I0(GND_net), .I1(encoder0_position[18]), .I2(VCC_net), 
            .I3(n43896), .O(encoder0_position_scaled_23__N_327[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5094_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5094_19 (.CI(n43896), .I0(encoder0_position[18]), .I1(VCC_net), 
            .CO(n43897));
    SB_LUT4 add_5094_18_lut (.I0(GND_net), .I1(encoder0_position[17]), .I2(VCC_net), 
            .I3(n43895), .O(encoder0_position_scaled_23__N_327[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5094_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1570_5 (.CI(n44164), 
            .I0(n2331), .I1(VCC_net), .CO(n44165));
    SB_CARRY add_5094_18 (.CI(n43895), .I0(encoder0_position[17]), .I1(VCC_net), 
            .CO(n43896));
    SB_LUT4 add_5094_17_lut (.I0(GND_net), .I1(encoder0_position[16]), .I2(VCC_net), 
            .I3(n43894), .O(encoder0_position_scaled_23__N_327[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5094_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1570_4_lut (.I0(GND_net), 
            .I1(n2332), .I2(GND_net), .I3(n44163), .O(n2399)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1570_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1570_4 (.CI(n44163), 
            .I0(n2332), .I1(GND_net), .CO(n44164));
    SB_CARRY add_5094_17 (.CI(n43894), .I0(encoder0_position[16]), .I1(VCC_net), 
            .CO(n43895));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1570_3_lut (.I0(GND_net), 
            .I1(n2333), .I2(VCC_net), .I3(n44162), .O(n2400)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1570_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1570_3 (.CI(n44162), 
            .I0(n2333), .I1(VCC_net), .CO(n44163));
    SB_LUT4 add_5094_16_lut (.I0(GND_net), .I1(encoder0_position[15]), .I2(VCC_net), 
            .I3(n43893), .O(encoder0_position_scaled_23__N_327[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5094_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_281_i3_4_lut (.I0(encoder1_position_scaled[2]), .I1(displacement[2]), 
            .I2(n15), .I3(n15_adj_5471), .O(motor_state_23__N_123[2]));   // verilog/TinyFPGA_B.v(284[5] 286[10])
    defparam mux_281_i3_4_lut.LUT_INIT = 16'h0aca;
    SB_CARRY add_5094_16 (.CI(n43893), .I0(encoder0_position[15]), .I1(VCC_net), 
            .CO(n43894));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1570_2_lut (.I0(GND_net), 
            .I1(n534), .I2(GND_net), .I3(VCC_net), .O(n2401)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1570_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5094_15_lut (.I0(GND_net), .I1(encoder0_position[14]), .I2(VCC_net), 
            .I3(n43892), .O(encoder0_position_scaled_23__N_327[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5094_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1570_2 (.CI(VCC_net), 
            .I0(n534), .I1(GND_net), .CO(n44162));
    SB_LUT4 i40284_1_lut (.I0(n2643), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n56115));
    defparam i40284_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_5094_15 (.CI(n43892), .I0(encoder0_position[14]), .I1(VCC_net), 
            .CO(n43893));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1503_22_lut (.I0(n56233), 
            .I1(n2214), .I2(VCC_net), .I3(n44161), .O(n2313)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1503_22_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mux_281_i4_4_lut (.I0(encoder1_position_scaled[3]), .I1(displacement[3]), 
            .I2(n15), .I3(n15_adj_5471), .O(motor_state_23__N_123[3]));   // verilog/TinyFPGA_B.v(284[5] 286[10])
    defparam mux_281_i4_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1503_21_lut (.I0(GND_net), 
            .I1(n2215), .I2(VCC_net), .I3(n44160), .O(n2282)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1503_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5094_14_lut (.I0(GND_net), .I1(encoder0_position[13]), .I2(VCC_net), 
            .I3(n43891), .O(encoder0_position_scaled_23__N_327[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5094_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5094_14 (.CI(n43891), .I0(encoder0_position[13]), .I1(VCC_net), 
            .CO(n43892));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1503_21 (.CI(n44160), 
            .I0(n2215), .I1(VCC_net), .CO(n44161));
    SB_LUT4 add_5094_13_lut (.I0(GND_net), .I1(encoder0_position[12]), .I2(VCC_net), 
            .I3(n43890), .O(encoder0_position_scaled_23__N_327[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5094_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5094_13 (.CI(n43890), .I0(encoder0_position[12]), .I1(VCC_net), 
            .CO(n43891));
    SB_LUT4 add_5094_12_lut (.I0(GND_net), .I1(encoder0_position[11]), .I2(VCC_net), 
            .I3(n43889), .O(encoder0_position_scaled_23__N_327[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5094_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1503_20_lut (.I0(GND_net), 
            .I1(n2216), .I2(VCC_net), .I3(n44159), .O(n2283)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1503_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1503_20 (.CI(n44159), 
            .I0(n2216), .I1(VCC_net), .CO(n44160));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i904_rep_52_3_lut (.I0(n1325), 
            .I1(n1392), .I2(n1356), .I3(GND_net), .O(n1424));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i904_rep_52_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1503_19_lut (.I0(GND_net), 
            .I1(n2217), .I2(VCC_net), .I3(n44158), .O(n2284)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1503_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1503_19 (.CI(n44158), 
            .I0(n2217), .I1(VCC_net), .CO(n44159));
    SB_LUT4 i15436_3_lut (.I0(Kp[5]), .I1(\data_in_frame[3] [5]), .I2(n50654), 
            .I3(GND_net), .O(n29516));   // verilog/coms.v(128[12] 303[6])
    defparam i15436_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_5094_12 (.CI(n43889), .I0(encoder0_position[11]), .I1(VCC_net), 
            .CO(n43890));
    SB_LUT4 add_5094_11_lut (.I0(GND_net), .I1(encoder0_position[10]), .I2(VCC_net), 
            .I3(n43888), .O(encoder0_position_scaled_23__N_327[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5094_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1503_18_lut (.I0(GND_net), 
            .I1(n2218), .I2(VCC_net), .I3(n44157), .O(n2285)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1503_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1503_18 (.CI(n44157), 
            .I0(n2218), .I1(VCC_net), .CO(n44158));
    SB_CARRY add_5094_11 (.CI(n43888), .I0(encoder0_position[10]), .I1(VCC_net), 
            .CO(n43889));
    SB_DFFESR GHA_210 (.Q(GHA), .C(clk16MHz), .E(n28672), .D(GHA_N_478), 
            .R(n29145));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1503_17_lut (.I0(GND_net), 
            .I1(n2219), .I2(VCC_net), .I3(n44156), .O(n2286)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1503_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1503_17 (.CI(n44156), 
            .I0(n2219), .I1(VCC_net), .CO(n44157));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1503_16_lut (.I0(GND_net), 
            .I1(n2220), .I2(VCC_net), .I3(n44155), .O(n2287)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1503_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5094_10_lut (.I0(GND_net), .I1(encoder0_position[9]), .I2(VCC_net), 
            .I3(n43887), .O(encoder0_position_scaled_23__N_327[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5094_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1503_16 (.CI(n44155), 
            .I0(n2220), .I1(VCC_net), .CO(n44156));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1503_15_lut (.I0(GND_net), 
            .I1(n2221), .I2(VCC_net), .I3(n44154), .O(n2288)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1503_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1503_15 (.CI(n44154), 
            .I0(n2221), .I1(VCC_net), .CO(n44155));
    SB_LUT4 dti_counter_2279_add_4_9_lut (.I0(n54547), .I1(n36544), .I2(dti_counter[7]), 
            .I3(n44447), .O(n48)) /* synthesis syn_instantiated=1 */ ;
    defparam dti_counter_2279_add_4_9_lut.LUT_INIT = 16'hE22E;
    SB_CARRY add_5094_10 (.CI(n43887), .I0(encoder0_position[9]), .I1(VCC_net), 
            .CO(n43888));
    SB_LUT4 dti_counter_2279_add_4_8_lut (.I0(n54548), .I1(n36544), .I2(dti_counter[6]), 
            .I3(n44446), .O(n49)) /* synthesis syn_instantiated=1 */ ;
    defparam dti_counter_2279_add_4_8_lut.LUT_INIT = 16'hE22E;
    SB_CARRY dti_counter_2279_add_4_8 (.CI(n44446), .I0(n36544), .I1(dti_counter[6]), 
            .CO(n44447));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1503_14_lut (.I0(GND_net), 
            .I1(n2222), .I2(VCC_net), .I3(n44153), .O(n2289)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1503_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1503_14 (.CI(n44153), 
            .I0(n2222), .I1(VCC_net), .CO(n44154));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1503_13_lut (.I0(GND_net), 
            .I1(n2223), .I2(VCC_net), .I3(n44152), .O(n2290)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1503_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1503_13 (.CI(n44152), 
            .I0(n2223), .I1(VCC_net), .CO(n44153));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1503_12_lut (.I0(GND_net), 
            .I1(n2224), .I2(VCC_net), .I3(n44151), .O(n2291)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1503_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 n10829_bdd_4_lut_40846 (.I0(n10829), .I1(n436), .I2(current[5]), 
            .I3(duty[23]), .O(n56676));
    defparam n10829_bdd_4_lut_40846.LUT_INIT = 16'he4aa;
    SB_LUT4 dti_counter_2279_add_4_7_lut (.I0(n54549), .I1(n36544), .I2(dti_counter[5]), 
            .I3(n44445), .O(n50)) /* synthesis syn_instantiated=1 */ ;
    defparam dti_counter_2279_add_4_7_lut.LUT_INIT = 16'hE22E;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1503_12 (.CI(n44151), 
            .I0(n2224), .I1(VCC_net), .CO(n44152));
    SB_LUT4 add_5094_9_lut (.I0(GND_net), .I1(encoder0_position[8]), .I2(VCC_net), 
            .I3(n43886), .O(encoder0_position_scaled_23__N_327[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5094_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY dti_counter_2279_add_4_7 (.CI(n44445), .I0(n36544), .I1(dti_counter[5]), 
            .CO(n44446));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i971_3_lut (.I0(n1424), .I1(n1491), 
            .I2(n1455), .I3(GND_net), .O(n1523));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i971_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 dti_counter_2279_add_4_6_lut (.I0(n54550), .I1(n36544), .I2(dti_counter[4]), 
            .I3(n44444), .O(n51)) /* synthesis syn_instantiated=1 */ ;
    defparam dti_counter_2279_add_4_6_lut.LUT_INIT = 16'hE22E;
    SB_CARRY dti_counter_2279_add_4_6 (.CI(n44444), .I0(n36544), .I1(dti_counter[4]), 
            .CO(n44445));
    SB_LUT4 dti_counter_2279_add_4_5_lut (.I0(n54551), .I1(n36544), .I2(dti_counter[3]), 
            .I3(n44443), .O(n52)) /* synthesis syn_instantiated=1 */ ;
    defparam dti_counter_2279_add_4_5_lut.LUT_INIT = 16'hE22E;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1503_11_lut (.I0(GND_net), 
            .I1(n2225), .I2(VCC_net), .I3(n44150), .O(n2292)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1503_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY dti_counter_2279_add_4_5 (.CI(n44443), .I0(n36544), .I1(dti_counter[3]), 
            .CO(n44444));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1503_11 (.CI(n44150), 
            .I0(n2225), .I1(VCC_net), .CO(n44151));
    SB_LUT4 i22664_2_lut_2_lut (.I0(duty[16]), .I1(n296), .I2(GND_net), 
            .I3(GND_net), .O(n4913));   // verilog/TinyFPGA_B.v(123[17] 125[11])
    defparam i22664_2_lut_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 dti_counter_2279_add_4_4_lut (.I0(n54552), .I1(n36544), .I2(dti_counter[2]), 
            .I3(n44442), .O(n53)) /* synthesis syn_instantiated=1 */ ;
    defparam dti_counter_2279_add_4_4_lut.LUT_INIT = 16'hE22E;
    SB_LUT4 n56676_bdd_4_lut (.I0(n56676), .I1(duty[5]), .I2(n265), .I3(duty[23]), 
            .O(pwm_setpoint_23__N_11[5]));
    defparam n56676_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_CARRY dti_counter_2279_add_4_4 (.CI(n44442), .I0(n36544), .I1(dti_counter[2]), 
            .CO(n44443));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1503_10_lut (.I0(GND_net), 
            .I1(n2226), .I2(VCC_net), .I3(n44149), .O(n2293)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1503_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5094_9 (.CI(n43886), .I0(encoder0_position[8]), .I1(VCC_net), 
            .CO(n43887));
    SB_LUT4 dti_counter_2279_add_4_3_lut (.I0(n54553), .I1(n36544), .I2(dti_counter[1]), 
            .I3(n44441), .O(n54)) /* synthesis syn_instantiated=1 */ ;
    defparam dti_counter_2279_add_4_3_lut.LUT_INIT = 16'hE22E;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1503_10 (.CI(n44149), 
            .I0(n2226), .I1(VCC_net), .CO(n44150));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1503_9_lut (.I0(GND_net), 
            .I1(n2227), .I2(VCC_net), .I3(n44148), .O(n2294)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1503_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY dti_counter_2279_add_4_3 (.CI(n44441), .I0(n36544), .I1(dti_counter[1]), 
            .CO(n44442));
    SB_LUT4 dti_counter_2279_add_4_2_lut (.I0(n54586), .I1(n2573), .I2(dti_counter[0]), 
            .I3(VCC_net), .O(n55)) /* synthesis syn_instantiated=1 */ ;
    defparam dti_counter_2279_add_4_2_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY dti_counter_2279_add_4_2 (.CI(VCC_net), .I0(n2573), .I1(dti_counter[0]), 
            .CO(n44441));
    SB_LUT4 add_2797_25_lut (.I0(n56458), .I1(n2_adj_5611), .I2(n1059), 
            .I3(n44440), .O(encoder0_position_scaled_23__N_51[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2797_25_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 add_5094_8_lut (.I0(GND_net), .I1(encoder0_position[7]), .I2(VCC_net), 
            .I3(n43885), .O(encoder0_position_scaled_23__N_327[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5094_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1503_9 (.CI(n44148), 
            .I0(n2227), .I1(VCC_net), .CO(n44149));
    SB_LUT4 add_2797_24_lut (.I0(n56444), .I1(n2_adj_5611), .I2(n1158), 
            .I3(n44439), .O(encoder0_position_scaled_23__N_51[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2797_24_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1038_rep_50_3_lut (.I0(n1523), 
            .I1(n1590), .I2(n1554_adj_5597), .I3(GND_net), .O(n1622));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1038_rep_50_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_5094_8 (.CI(n43885), .I0(encoder0_position[7]), .I1(VCC_net), 
            .CO(n43886));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1105_3_lut (.I0(n1622), 
            .I1(n1689), .I2(n1653), .I3(GND_net), .O(n1721));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1105_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_2797_24 (.CI(n44439), .I0(n2_adj_5611), .I1(n1158), .CO(n44440));
    SB_LUT4 add_2797_23_lut (.I0(n56430), .I1(n2_adj_5611), .I2(n1257), 
            .I3(n44438), .O(encoder0_position_scaled_23__N_51[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2797_23_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1503_8_lut (.I0(GND_net), 
            .I1(n2228), .I2(VCC_net), .I3(n44147), .O(n2295)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1503_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1503_8 (.CI(n44147), 
            .I0(n2228), .I1(VCC_net), .CO(n44148));
    SB_CARRY add_2797_23 (.CI(n44438), .I0(n2_adj_5611), .I1(n1257), .CO(n44439));
    SB_LUT4 add_2797_22_lut (.I0(n56415), .I1(n2_adj_5611), .I2(n1356), 
            .I3(n44437), .O(encoder0_position_scaled_23__N_51[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2797_22_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2797_22 (.CI(n44437), .I0(n2_adj_5611), .I1(n1356), .CO(n44438));
    SB_LUT4 add_2797_21_lut (.I0(n56399), .I1(n2_adj_5611), .I2(n1455), 
            .I3(n44436), .O(encoder0_position_scaled_23__N_51[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2797_21_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1503_7_lut (.I0(GND_net), 
            .I1(n2229), .I2(GND_net), .I3(n44146), .O(n2296)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1503_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2797_21 (.CI(n44436), .I0(n2_adj_5611), .I1(n1455), .CO(n44437));
    SB_LUT4 add_2797_20_lut (.I0(n56382), .I1(n2_adj_5611), .I2(n1554_adj_5597), 
            .I3(n44435), .O(encoder0_position_scaled_23__N_51[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2797_20_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2797_20 (.CI(n44435), .I0(n2_adj_5611), .I1(n1554_adj_5597), 
            .CO(n44436));
    SB_LUT4 add_2797_19_lut (.I0(n56364), .I1(n2_adj_5611), .I2(n1653), 
            .I3(n44434), .O(encoder0_position_scaled_23__N_51[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2797_19_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 add_5094_7_lut (.I0(GND_net), .I1(encoder0_position[6]), .I2(VCC_net), 
            .I3(n43884), .O(encoder0_position_scaled_23__N_327[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5094_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2797_19 (.CI(n44434), .I0(n2_adj_5611), .I1(n1653), .CO(n44435));
    SB_CARRY add_5094_7 (.CI(n43884), .I0(encoder0_position[6]), .I1(VCC_net), 
            .CO(n43885));
    SB_LUT4 add_2797_18_lut (.I0(n56328), .I1(n2_adj_5611), .I2(n1752), 
            .I3(n44433), .O(encoder0_position_scaled_23__N_51[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2797_18_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 i22481_1_lut_2_lut (.I0(n24553), .I1(dti), .I2(GND_net), .I3(GND_net), 
            .O(n2573));
    defparam i22481_1_lut_2_lut.LUT_INIT = 16'h7777;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1172_3_lut (.I0(n1721), 
            .I1(n1788), .I2(n1752), .I3(GND_net), .O(n1820));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1172_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1503_7 (.CI(n44146), 
            .I0(n2229), .I1(GND_net), .CO(n44147));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1503_6_lut (.I0(GND_net), 
            .I1(n2230), .I2(GND_net), .I3(n44145), .O(n2297)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1503_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1503_6 (.CI(n44145), 
            .I0(n2230), .I1(GND_net), .CO(n44146));
    SB_CARRY add_2797_18 (.CI(n44433), .I0(n2_adj_5611), .I1(n1752), .CO(n44434));
    SB_LUT4 add_2797_17_lut (.I0(n56323), .I1(n2_adj_5611), .I2(n1851), 
            .I3(n44432), .O(encoder0_position_scaled_23__N_51[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2797_17_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1239_3_lut (.I0(n1820), 
            .I1(n1887), .I2(n1851), .I3(GND_net), .O(n1919));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1239_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_2797_17 (.CI(n44432), .I0(n2_adj_5611), .I1(n1851), .CO(n44433));
    SB_LUT4 add_5094_6_lut (.I0(GND_net), .I1(encoder0_position[5]), .I2(VCC_net), 
            .I3(n43883), .O(encoder0_position_scaled_23__N_327[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5094_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1306_3_lut (.I0(n1919), 
            .I1(n1986), .I2(n1950), .I3(GND_net), .O(n2018));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1306_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_5094_6 (.CI(n43883), .I0(encoder0_position[5]), .I1(VCC_net), 
            .CO(n43884));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1503_5_lut (.I0(GND_net), 
            .I1(n2231), .I2(VCC_net), .I3(n44144), .O(n2298)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1503_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1503_5 (.CI(n44144), 
            .I0(n2231), .I1(VCC_net), .CO(n44145));
    SB_LUT4 add_2797_16_lut (.I0(n56302), .I1(n2_adj_5611), .I2(n1950), 
            .I3(n44431), .O(encoder0_position_scaled_23__N_51[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2797_16_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2797_16 (.CI(n44431), .I0(n2_adj_5611), .I1(n1950), .CO(n44432));
    SB_LUT4 add_5094_5_lut (.I0(GND_net), .I1(encoder0_position[4]), .I2(VCC_net), 
            .I3(n43882), .O(encoder0_position_scaled_23__N_327[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5094_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2797_15_lut (.I0(n56280), .I1(n2_adj_5611), .I2(n2049), 
            .I3(n44430), .O(encoder0_position_scaled_23__N_51[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2797_15_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1503_4_lut (.I0(GND_net), 
            .I1(n2232), .I2(GND_net), .I3(n44143), .O(n2299)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1503_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1503_4 (.CI(n44143), 
            .I0(n2232), .I1(GND_net), .CO(n44144));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1503_3_lut (.I0(GND_net), 
            .I1(n2233_adj_5599), .I2(VCC_net), .I3(n44142), .O(n2300)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1503_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5094_5 (.CI(n43882), .I0(encoder0_position[4]), .I1(VCC_net), 
            .CO(n43883));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1503_3 (.CI(n44142), 
            .I0(n2233_adj_5599), .I1(VCC_net), .CO(n44143));
    SB_LUT4 add_5094_4_lut (.I0(GND_net), .I1(encoder0_position[3]), .I2(VCC_net), 
            .I3(n43881), .O(encoder0_position_scaled_23__N_327[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5094_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5094_4 (.CI(n43881), .I0(encoder0_position[3]), .I1(VCC_net), 
            .CO(n43882));
    SB_CARRY add_2797_15 (.CI(n44430), .I0(n2_adj_5611), .I1(n2049), .CO(n44431));
    SB_LUT4 add_5094_3_lut (.I0(GND_net), .I1(encoder0_position[2]), .I2(VCC_net), 
            .I3(n43880), .O(encoder0_position_scaled_23__N_327[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5094_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2797_14_lut (.I0(n56237), .I1(n2_adj_5611), .I2(n2148), 
            .I3(n44429), .O(encoder0_position_scaled_23__N_51[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2797_14_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2797_14 (.CI(n44429), .I0(n2_adj_5611), .I1(n2148), .CO(n44430));
    SB_CARRY add_5094_3 (.CI(n43880), .I0(encoder0_position[2]), .I1(VCC_net), 
            .CO(n43881));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1503_2_lut (.I0(GND_net), 
            .I1(n533), .I2(GND_net), .I3(VCC_net), .O(n2301)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1503_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5094_2_lut (.I0(GND_net), .I1(encoder0_position[1]), .I2(VCC_net), 
            .I3(n43879), .O(encoder0_position_scaled_23__N_327[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5094_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5094_2 (.CI(n43879), .I0(encoder0_position[1]), .I1(VCC_net), 
            .CO(n43880));
    SB_LUT4 add_2797_13_lut (.I0(n56233), .I1(n2_adj_5611), .I2(n2247), 
            .I3(n44428), .O(encoder0_position_scaled_23__N_51[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2797_13_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2797_13 (.CI(n44428), .I0(n2_adj_5611), .I1(n2247), .CO(n44429));
    SB_CARRY add_5094_1 (.CI(GND_net), .I0(encoder0_position[0]), .I1(encoder0_position[0]), 
            .CO(n43879));
    SB_LUT4 add_2797_12_lut (.I0(n56200), .I1(n2_adj_5611), .I2(n2346), 
            .I3(n44427), .O(encoder0_position_scaled_23__N_51[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2797_12_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1503_2 (.CI(VCC_net), 
            .I0(n533), .I1(GND_net), .CO(n44142));
    SB_CARRY add_2797_12 (.CI(n44427), .I0(n2_adj_5611), .I1(n2346), .CO(n44428));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1436_21_lut (.I0(n56237), 
            .I1(n2115), .I2(VCC_net), .I3(n44141), .O(n2214)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1436_21_lut.LUT_INIT = 16'h8228;
    SB_LUT4 add_2797_11_lut (.I0(n56171), .I1(n2_adj_5611), .I2(n2445), 
            .I3(n44426), .O(encoder0_position_scaled_23__N_51[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2797_11_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2797_11 (.CI(n44426), .I0(n2_adj_5611), .I1(n2445), .CO(n44427));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1436_20_lut (.I0(GND_net), 
            .I1(n2116), .I2(VCC_net), .I3(n44140), .O(n2183)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1436_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2797_10_lut (.I0(n56142), .I1(n2_adj_5611), .I2(n2544), 
            .I3(n44425), .O(encoder0_position_scaled_23__N_51[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2797_10_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1436_20 (.CI(n44140), 
            .I0(n2116), .I1(VCC_net), .CO(n44141));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1436_19_lut (.I0(GND_net), 
            .I1(n2117), .I2(VCC_net), .I3(n44139), .O(n2184)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1436_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1436_19 (.CI(n44139), 
            .I0(n2117), .I1(VCC_net), .CO(n44140));
    SB_CARRY add_2797_10 (.CI(n44425), .I0(n2_adj_5611), .I1(n2544), .CO(n44426));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1436_18_lut (.I0(GND_net), 
            .I1(n2118), .I2(VCC_net), .I3(n44138), .O(n2185)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1436_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1373_3_lut (.I0(n2018), 
            .I1(n2085), .I2(n2049), .I3(GND_net), .O(n2117));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1373_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_2797_9_lut (.I0(n56115), .I1(n2_adj_5611), .I2(n2643), 
            .I3(n44424), .O(encoder0_position_scaled_23__N_51[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2797_9_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2797_9 (.CI(n44424), .I0(n2_adj_5611), .I1(n2643), .CO(n44425));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1436_18 (.CI(n44138), 
            .I0(n2118), .I1(VCC_net), .CO(n44139));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1436_17_lut (.I0(GND_net), 
            .I1(n2119), .I2(VCC_net), .I3(n44137), .O(n2186)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1436_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1436_17 (.CI(n44137), 
            .I0(n2119), .I1(VCC_net), .CO(n44138));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1436_16_lut (.I0(GND_net), 
            .I1(n2120), .I2(VCC_net), .I3(n44136), .O(n2187)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1436_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2797_8_lut (.I0(n56086), .I1(n2_adj_5611), .I2(n2742), 
            .I3(n44423), .O(encoder0_position_scaled_23__N_51[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2797_8_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2797_8 (.CI(n44423), .I0(n2_adj_5611), .I1(n2742), .CO(n44424));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1436_16 (.CI(n44136), 
            .I0(n2120), .I1(VCC_net), .CO(n44137));
    SB_LUT4 add_2797_7_lut (.I0(n56056), .I1(n2_adj_5611), .I2(n2841), 
            .I3(n44422), .O(encoder0_position_scaled_23__N_51[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2797_7_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2797_7 (.CI(n44422), .I0(n2_adj_5611), .I1(n2841), .CO(n44423));
    SB_LUT4 add_2797_6_lut (.I0(n56025), .I1(n2_adj_5611), .I2(n2940), 
            .I3(n44421), .O(encoder0_position_scaled_23__N_51[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2797_6_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2797_6 (.CI(n44421), .I0(n2_adj_5611), .I1(n2940), .CO(n44422));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1436_15_lut (.I0(GND_net), 
            .I1(n2121), .I2(VCC_net), .I3(n44135), .O(n2188)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1436_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1436_15 (.CI(n44135), 
            .I0(n2121), .I1(VCC_net), .CO(n44136));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1436_14_lut (.I0(GND_net), 
            .I1(n2122), .I2(VCC_net), .I3(n44134), .O(n2189)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1436_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1436_14 (.CI(n44134), 
            .I0(n2122), .I1(VCC_net), .CO(n44135));
    SB_LUT4 add_2797_5_lut (.I0(n56595), .I1(n2_adj_5611), .I2(n3039), 
            .I3(n44420), .O(encoder0_position_scaled_23__N_51[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2797_5_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2797_5 (.CI(n44420), .I0(n2_adj_5611), .I1(n3039), .CO(n44421));
    SB_LUT4 add_2797_4_lut (.I0(n56561), .I1(n2_adj_5611), .I2(n3138), 
            .I3(n44419), .O(encoder0_position_scaled_23__N_51[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2797_4_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1436_13_lut (.I0(GND_net), 
            .I1(n2123), .I2(VCC_net), .I3(n44133), .O(n2190)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1436_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2797_4 (.CI(n44419), .I0(n2_adj_5611), .I1(n3138), .CO(n44420));
    SB_LUT4 add_2797_3_lut (.I0(n56498), .I1(n2_adj_5611), .I2(n3237), 
            .I3(n44418), .O(encoder0_position_scaled_23__N_51[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2797_3_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1436_13 (.CI(n44133), 
            .I0(n2123), .I1(VCC_net), .CO(n44134));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1436_12_lut (.I0(GND_net), 
            .I1(n2124), .I2(VCC_net), .I3(n44132), .O(n2191)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1436_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1436_12 (.CI(n44132), 
            .I0(n2124), .I1(VCC_net), .CO(n44133));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1436_11_lut (.I0(GND_net), 
            .I1(n2125), .I2(VCC_net), .I3(n44131), .O(n2192)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1436_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2797_3 (.CI(n44418), .I0(n2_adj_5611), .I1(n3237), .CO(n44419));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1436_11 (.CI(n44131), 
            .I0(n2125), .I1(VCC_net), .CO(n44132));
    SB_LUT4 add_2797_2_lut (.I0(n56490), .I1(n2_adj_5611), .I2(n37482), 
            .I3(VCC_net), .O(encoder0_position_scaled_23__N_51[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2797_2_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1436_10_lut (.I0(GND_net), 
            .I1(n2126), .I2(VCC_net), .I3(n44130), .O(n2193)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1436_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2797_2 (.CI(VCC_net), .I0(n2_adj_5611), .I1(n37482), 
            .CO(n44418));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1436_10 (.CI(n44130), 
            .I0(n2126), .I1(VCC_net), .CO(n44131));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_2173_33_lut (.I0(n56498), 
            .I1(n3204), .I2(VCC_net), .I3(n44417), .O(n53025)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_2173_33_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_2173_32_lut (.I0(GND_net), 
            .I1(n3205), .I2(VCC_net), .I3(n44416), .O(n3272)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_2173_32_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_2173_32 (.CI(n44416), 
            .I0(n3205), .I1(VCC_net), .CO(n44417));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1436_9_lut (.I0(GND_net), 
            .I1(n2127), .I2(VCC_net), .I3(n44129), .O(n2194)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1436_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_2173_31_lut (.I0(GND_net), 
            .I1(n3206), .I2(VCC_net), .I3(n44415), .O(n3273)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_2173_31_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_2173_31 (.CI(n44415), 
            .I0(n3206), .I1(VCC_net), .CO(n44416));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_2173_30_lut (.I0(GND_net), 
            .I1(n3207), .I2(VCC_net), .I3(n44414), .O(n3274)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_2173_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_2173_30 (.CI(n44414), 
            .I0(n3207), .I1(VCC_net), .CO(n44415));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_2173_29_lut (.I0(GND_net), 
            .I1(n3208), .I2(VCC_net), .I3(n44413), .O(n3275)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_2173_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1436_9 (.CI(n44129), 
            .I0(n2127), .I1(VCC_net), .CO(n44130));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_2173_29 (.CI(n44413), 
            .I0(n3208), .I1(VCC_net), .CO(n44414));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1436_8_lut (.I0(GND_net), 
            .I1(n2128), .I2(VCC_net), .I3(n44128), .O(n2195)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1436_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1436_8 (.CI(n44128), 
            .I0(n2128), .I1(VCC_net), .CO(n44129));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1436_7_lut (.I0(GND_net), 
            .I1(n2129), .I2(GND_net), .I3(n44127), .O(n2196)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1436_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_2173_28_lut (.I0(GND_net), 
            .I1(n3209), .I2(VCC_net), .I3(n44412), .O(n3276)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_2173_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1436_7 (.CI(n44127), 
            .I0(n2129), .I1(GND_net), .CO(n44128));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1436_6_lut (.I0(GND_net), 
            .I1(n2130), .I2(GND_net), .I3(n44126), .O(n2197)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1436_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_2173_28 (.CI(n44412), 
            .I0(n3209), .I1(VCC_net), .CO(n44413));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i844_3_lut (.I0(n1233), .I1(n1300), 
            .I2(n1257), .I3(GND_net), .O(n1332));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i844_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1436_6 (.CI(n44126), 
            .I0(n2130), .I1(GND_net), .CO(n44127));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1436_5_lut (.I0(GND_net), 
            .I1(n2131), .I2(VCC_net), .I3(n44125), .O(n2198)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1436_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_2173_27_lut (.I0(GND_net), 
            .I1(n3210), .I2(VCC_net), .I3(n44411), .O(n3277)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_2173_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1436_5 (.CI(n44125), 
            .I0(n2131), .I1(VCC_net), .CO(n44126));
    SB_LUT4 add_261_5_lut (.I0(current[3]), .I1(duty[6]), .I2(n56614), 
            .I3(n43560), .O(n267)) /* synthesis syn_instantiated=1 */ ;
    defparam add_261_5_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_2173_27 (.CI(n44411), 
            .I0(n3210), .I1(VCC_net), .CO(n44412));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_2173_26_lut (.I0(GND_net), 
            .I1(n3211), .I2(VCC_net), .I3(n44410), .O(n3278)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_2173_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1436_4_lut (.I0(GND_net), 
            .I1(n2132), .I2(GND_net), .I3(n44124), .O(n2199)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1436_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_2173_26 (.CI(n44410), 
            .I0(n3211), .I1(VCC_net), .CO(n44411));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_2173_25_lut (.I0(GND_net), 
            .I1(n3212), .I2(VCC_net), .I3(n44409), .O(n3279)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_2173_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1436_4 (.CI(n44124), 
            .I0(n2132), .I1(GND_net), .CO(n44125));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1436_3_lut (.I0(GND_net), 
            .I1(n2133), .I2(VCC_net), .I3(n44123), .O(n2200)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1436_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1436_3 (.CI(n44123), 
            .I0(n2133), .I1(VCC_net), .CO(n44124));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1436_2_lut (.I0(GND_net), 
            .I1(n532), .I2(GND_net), .I3(VCC_net), .O(n2201)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1436_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_2173_25 (.CI(n44409), 
            .I0(n3212), .I1(VCC_net), .CO(n44410));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1436_2 (.CI(VCC_net), 
            .I0(n532), .I1(GND_net), .CO(n44123));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1369_20_lut (.I0(n56280), 
            .I1(n2016), .I2(VCC_net), .I3(n44122), .O(n2115)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1369_20_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_2173_24_lut (.I0(GND_net), 
            .I1(n3213), .I2(VCC_net), .I3(n44408), .O(n3280)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_2173_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_2173_24 (.CI(n44408), 
            .I0(n3213), .I1(VCC_net), .CO(n44409));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_2173_23_lut (.I0(GND_net), 
            .I1(n3214), .I2(VCC_net), .I3(n44407), .O(n3281)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_2173_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1369_19_lut (.I0(GND_net), 
            .I1(n2017), .I2(VCC_net), .I3(n44121), .O(n2084)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1369_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1369_19 (.CI(n44121), 
            .I0(n2017), .I1(VCC_net), .CO(n44122));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_2173_23 (.CI(n44407), 
            .I0(n3214), .I1(VCC_net), .CO(n44408));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_2173_22_lut (.I0(GND_net), 
            .I1(n3215), .I2(VCC_net), .I3(n44406), .O(n3282)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_2173_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1369_18_lut (.I0(GND_net), 
            .I1(n2018), .I2(VCC_net), .I3(n44120), .O(n2085)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1369_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1369_18 (.CI(n44120), 
            .I0(n2018), .I1(VCC_net), .CO(n44121));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_2173_22 (.CI(n44406), 
            .I0(n3215), .I1(VCC_net), .CO(n44407));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_2173_21_lut (.I0(GND_net), 
            .I1(n3216), .I2(VCC_net), .I3(n44405), .O(n3283)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_2173_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1369_17_lut (.I0(GND_net), 
            .I1(n2019), .I2(VCC_net), .I3(n44119), .O(n2086)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1369_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1369_17 (.CI(n44119), 
            .I0(n2019), .I1(VCC_net), .CO(n44120));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1369_16_lut (.I0(GND_net), 
            .I1(n2020), .I2(VCC_net), .I3(n44118), .O(n2087)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1369_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_261_5 (.CI(n43560), .I0(duty[6]), .I1(n56614), .CO(n43561));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_2173_21 (.CI(n44405), 
            .I0(n3216), .I1(VCC_net), .CO(n44406));
    SB_LUT4 add_261_4_lut (.I0(current[2]), .I1(duty[5]), .I2(n56614), 
            .I3(n43559), .O(n268)) /* synthesis syn_instantiated=1 */ ;
    defparam add_261_4_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_2173_20_lut (.I0(GND_net), 
            .I1(n3217), .I2(VCC_net), .I3(n44404), .O(n3284)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_2173_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1369_16 (.CI(n44118), 
            .I0(n2020), .I1(VCC_net), .CO(n44119));
    SB_LUT4 add_263_3_lut (.I0(GND_net), .I1(encoder1_position[4]), .I2(GND_net), 
            .I3(n43535), .O(encoder1_position_scaled_23__N_75[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_263_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i40340_1_lut (.I0(n2445), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n56171));
    defparam i40340_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_2173_20 (.CI(n44404), 
            .I0(n3217), .I1(VCC_net), .CO(n44405));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1369_15_lut (.I0(GND_net), 
            .I1(n2021), .I2(VCC_net), .I3(n44117), .O(n2088)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1369_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_263_3 (.CI(n43535), .I0(encoder1_position[4]), .I1(GND_net), 
            .CO(n43536));
    SB_LUT4 i40497_1_lut (.I0(n1752), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n56328));
    defparam i40497_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_2173_19_lut (.I0(GND_net), 
            .I1(n3218), .I2(VCC_net), .I3(n44403), .O(n3285)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_2173_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_2173_19 (.CI(n44403), 
            .I0(n3218), .I1(VCC_net), .CO(n44404));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1369_15 (.CI(n44117), 
            .I0(n2021), .I1(VCC_net), .CO(n44118));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_2173_18_lut (.I0(GND_net), 
            .I1(n3219), .I2(VCC_net), .I3(n44402), .O(n3286)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_2173_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1369_14_lut (.I0(GND_net), 
            .I1(n2022), .I2(VCC_net), .I3(n44116), .O(n2089)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1369_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1369_14 (.CI(n44116), 
            .I0(n2022), .I1(VCC_net), .CO(n44117));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1369_13_lut (.I0(GND_net), 
            .I1(n2023), .I2(VCC_net), .I3(n44115), .O(n2090)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1369_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_2173_18 (.CI(n44402), 
            .I0(n3219), .I1(VCC_net), .CO(n44403));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_2173_17_lut (.I0(GND_net), 
            .I1(n3220), .I2(VCC_net), .I3(n44401), .O(n3287)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_2173_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_2173_17 (.CI(n44401), 
            .I0(n3220), .I1(VCC_net), .CO(n44402));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1369_13 (.CI(n44115), 
            .I0(n2023), .I1(VCC_net), .CO(n44116));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1369_12_lut (.I0(GND_net), 
            .I1(n2024), .I2(VCC_net), .I3(n44114), .O(n2091_adj_5598)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1369_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_2173_16_lut (.I0(GND_net), 
            .I1(n3221), .I2(VCC_net), .I3(n44400), .O(n3288)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_2173_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_2173_16 (.CI(n44400), 
            .I0(n3221), .I1(VCC_net), .CO(n44401));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_2173_15_lut (.I0(GND_net), 
            .I1(n3222), .I2(VCC_net), .I3(n44399), .O(n3289)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_2173_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i40406_1_lut (.I0(n2148), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n56237));
    defparam i40406_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1369_12 (.CI(n44114), 
            .I0(n2024), .I1(VCC_net), .CO(n44115));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1369_11_lut (.I0(GND_net), 
            .I1(n2025), .I2(VCC_net), .I3(n44113), .O(n2092)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1369_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1369_11 (.CI(n44113), 
            .I0(n2025), .I1(VCC_net), .CO(n44114));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1369_10_lut (.I0(GND_net), 
            .I1(n2026), .I2(VCC_net), .I3(n44112), .O(n2093)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1369_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_261_4 (.CI(n43559), .I0(duty[5]), .I1(n56614), .CO(n43560));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_2173_15 (.CI(n44399), 
            .I0(n3222), .I1(VCC_net), .CO(n44400));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_2173_14_lut (.I0(GND_net), 
            .I1(n3223), .I2(VCC_net), .I3(n44398), .O(n3290)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_2173_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1369_10 (.CI(n44112), 
            .I0(n2026), .I1(VCC_net), .CO(n44113));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_2173_14 (.CI(n44398), 
            .I0(n3223), .I1(VCC_net), .CO(n44399));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_2173_13_lut (.I0(GND_net), 
            .I1(n3224), .I2(VCC_net), .I3(n44397), .O(n3291)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_2173_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_2173_13 (.CI(n44397), 
            .I0(n3224), .I1(VCC_net), .CO(n44398));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1369_9_lut (.I0(GND_net), 
            .I1(n2027), .I2(VCC_net), .I3(n44111), .O(n2094)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1369_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_281_i5_4_lut (.I0(encoder1_position_scaled[4]), .I1(displacement[4]), 
            .I2(n15), .I3(n15_adj_5471), .O(motor_state_23__N_123[4]));   // verilog/TinyFPGA_B.v(284[5] 286[10])
    defparam mux_281_i5_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 add_261_3_lut (.I0(current[1]), .I1(duty[4]), .I2(n56614), 
            .I3(n43558), .O(n269)) /* synthesis syn_instantiated=1 */ ;
    defparam add_261_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1369_9 (.CI(n44111), 
            .I0(n2027), .I1(VCC_net), .CO(n44112));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1369_8_lut (.I0(GND_net), 
            .I1(n2028), .I2(VCC_net), .I3(n44110), .O(n2095)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1369_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_2173_12_lut (.I0(GND_net), 
            .I1(n3225), .I2(VCC_net), .I3(n44396), .O(n3292)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_2173_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1369_8 (.CI(n44110), 
            .I0(n2028), .I1(VCC_net), .CO(n44111));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_2173_12 (.CI(n44396), 
            .I0(n3225), .I1(VCC_net), .CO(n44397));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_2173_11_lut (.I0(GND_net), 
            .I1(n3226), .I2(VCC_net), .I3(n44395), .O(n3293)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_2173_11_lut.LUT_INIT = 16'hC33C;
    SB_DFFESS commutation_state_i0 (.Q(commutation_state[0]), .C(clk16MHz), 
            .E(n6_adj_5656), .D(commutation_state_7__N_264[0]), .S(commutation_state_7__N_272));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_2173_11 (.CI(n44395), 
            .I0(n3226), .I1(VCC_net), .CO(n44396));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1369_7_lut (.I0(GND_net), 
            .I1(n2029), .I2(GND_net), .I3(n44109), .O(n2096)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1369_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_2173_10_lut (.I0(GND_net), 
            .I1(n3227), .I2(VCC_net), .I3(n44394), .O(n3294)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_2173_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1369_7 (.CI(n44109), 
            .I0(n2029), .I1(GND_net), .CO(n44110));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1369_6_lut (.I0(GND_net), 
            .I1(n2030), .I2(GND_net), .I3(n44108), .O(n2097)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1369_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_2173_10 (.CI(n44394), 
            .I0(n3227), .I1(VCC_net), .CO(n44395));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1369_6 (.CI(n44108), 
            .I0(n2030), .I1(GND_net), .CO(n44109));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1369_5_lut (.I0(GND_net), 
            .I1(n2031), .I2(VCC_net), .I3(n44107), .O(n2098)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1369_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1369_5 (.CI(n44107), 
            .I0(n2031), .I1(VCC_net), .CO(n44108));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_2173_9_lut (.I0(GND_net), 
            .I1(n3228), .I2(VCC_net), .I3(n44393), .O(n3295)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_2173_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_2173_9 (.CI(n44393), 
            .I0(n3228), .I1(VCC_net), .CO(n44394));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_2173_8_lut (.I0(GND_net), 
            .I1(n3229), .I2(GND_net), .I3(n44392), .O(n3296)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_2173_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1369_4_lut (.I0(GND_net), 
            .I1(n2032), .I2(GND_net), .I3(n44106), .O(n2099)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1369_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_2173_8 (.CI(n44392), 
            .I0(n3229), .I1(GND_net), .CO(n44393));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1369_4 (.CI(n44106), 
            .I0(n2032), .I1(GND_net), .CO(n44107));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1369_3_lut (.I0(GND_net), 
            .I1(n2033), .I2(VCC_net), .I3(n44105), .O(n2100)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1369_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1369_3 (.CI(n44105), 
            .I0(n2033), .I1(VCC_net), .CO(n44106));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1369_2_lut (.I0(GND_net), 
            .I1(n531), .I2(GND_net), .I3(VCC_net), .O(n2101)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1369_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1369_2 (.CI(VCC_net), 
            .I0(n531), .I1(GND_net), .CO(n44105));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_2173_7_lut (.I0(n3298), 
            .I1(n3230), .I2(GND_net), .I3(n44391), .O(n54589)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_2173_7_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1302_19_lut (.I0(n56302), 
            .I1(n1917), .I2(VCC_net), .I3(n44104), .O(n2016)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1302_19_lut.LUT_INIT = 16'h8228;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_2173_7 (.CI(n44391), 
            .I0(n3230), .I1(GND_net), .CO(n44392));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1302_18_lut (.I0(GND_net), 
            .I1(n1918), .I2(VCC_net), .I3(n44103), .O(n1985)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1302_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_2173_6_lut (.I0(GND_net), 
            .I1(n3231), .I2(VCC_net), .I3(n44390), .O(n3298)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_2173_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_2173_6 (.CI(n44390), 
            .I0(n3231), .I1(VCC_net), .CO(n44391));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_2173_5_lut (.I0(GND_net), 
            .I1(n3232), .I2(GND_net), .I3(n44389), .O(n3299)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_2173_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1302_18 (.CI(n44103), 
            .I0(n1918), .I1(VCC_net), .CO(n44104));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1302_17_lut (.I0(GND_net), 
            .I1(n1919), .I2(VCC_net), .I3(n44102), .O(n1986)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1302_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1302_17 (.CI(n44102), 
            .I0(n1919), .I1(VCC_net), .CO(n44103));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1302_16_lut (.I0(GND_net), 
            .I1(n1920), .I2(VCC_net), .I3(n44101), .O(n1987)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1302_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_2173_5 (.CI(n44389), 
            .I0(n3232), .I1(GND_net), .CO(n44390));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_2173_4_lut (.I0(GND_net), 
            .I1(n3233), .I2(VCC_net), .I3(n44388), .O(n3300)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_2173_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1302_16 (.CI(n44101), 
            .I0(n1920), .I1(VCC_net), .CO(n44102));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1302_15_lut (.I0(GND_net), 
            .I1(n1921), .I2(VCC_net), .I3(n44100), .O(n1988)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1302_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i39315_3_lut_4_lut (.I0(n2247), .I1(n2148), .I2(n2125), .I3(n53094), 
            .O(n2323));
    defparam i39315_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_2173_4 (.CI(n44388), 
            .I0(n3233), .I1(VCC_net), .CO(n44389));
    SB_CARRY add_261_3 (.CI(n43558), .I0(duty[4]), .I1(n56614), .CO(n43559));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_2173_3_lut (.I0(GND_net), 
            .I1(n543), .I2(GND_net), .I3(n44387), .O(n3301)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_2173_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1302_15 (.CI(n44100), 
            .I0(n1921), .I1(VCC_net), .CO(n44101));
    SB_LUT4 add_261_2_lut (.I0(GND_net), .I1(duty[3]), .I2(n211), .I3(GND_net), 
            .O(n2091)) /* synthesis syn_instantiated=1 */ ;
    defparam add_261_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1302_14_lut (.I0(GND_net), 
            .I1(n1922), .I2(VCC_net), .I3(n44099), .O(n1989)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1302_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_2173_3 (.CI(n44387), 
            .I0(n543), .I1(GND_net), .CO(n44388));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_2173_2 (.CI(VCC_net), 
            .I0(n544), .I1(VCC_net), .CO(n44387));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1302_14 (.CI(n44099), 
            .I0(n1922), .I1(VCC_net), .CO(n44100));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_2106_31_lut (.I0(n56561), 
            .I1(n3105), .I2(VCC_net), .I3(n44386), .O(n3204)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_2106_31_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_2106_30_lut (.I0(GND_net), 
            .I1(n3106), .I2(VCC_net), .I3(n44385), .O(n3173)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_2106_30_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1302_13_lut (.I0(GND_net), 
            .I1(n1923), .I2(VCC_net), .I3(n44098), .O(n1990)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1302_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_2106_30 (.CI(n44385), 
            .I0(n3106), .I1(VCC_net), .CO(n44386));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1302_13 (.CI(n44098), 
            .I0(n1923), .I1(VCC_net), .CO(n44099));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_2106_29_lut (.I0(GND_net), 
            .I1(n3107), .I2(VCC_net), .I3(n44384), .O(n3174)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_2106_29_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1302_12_lut (.I0(GND_net), 
            .I1(n1924), .I2(VCC_net), .I3(n44097), .O(n1991)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1302_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1302_12 (.CI(n44097), 
            .I0(n1924), .I1(VCC_net), .CO(n44098));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_2106_29 (.CI(n44384), 
            .I0(n3107), .I1(VCC_net), .CO(n44385));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_2106_28_lut (.I0(GND_net), 
            .I1(n3108), .I2(VCC_net), .I3(n44383), .O(n3175)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_2106_28_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1302_11_lut (.I0(GND_net), 
            .I1(n1925), .I2(VCC_net), .I3(n44096), .O(n1992)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1302_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1302_11 (.CI(n44096), 
            .I0(n1925), .I1(VCC_net), .CO(n44097));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1302_10_lut (.I0(GND_net), 
            .I1(n1926), .I2(VCC_net), .I3(n44095), .O(n1993)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1302_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_2106_28 (.CI(n44383), 
            .I0(n3108), .I1(VCC_net), .CO(n44384));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1302_10 (.CI(n44095), 
            .I0(n1926), .I1(VCC_net), .CO(n44096));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1302_9_lut (.I0(GND_net), 
            .I1(n1927), .I2(VCC_net), .I3(n44094), .O(n1994)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1302_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_2106_27_lut (.I0(GND_net), 
            .I1(n3109), .I2(VCC_net), .I3(n44382), .O(n3176)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_2106_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1302_9 (.CI(n44094), 
            .I0(n1927), .I1(VCC_net), .CO(n44095));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_2106_27 (.CI(n44382), 
            .I0(n3109), .I1(VCC_net), .CO(n44383));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_2106_26_lut (.I0(GND_net), 
            .I1(n3110), .I2(VCC_net), .I3(n44381), .O(n3177)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_2106_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_2106_26 (.CI(n44381), 
            .I0(n3110), .I1(VCC_net), .CO(n44382));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1302_8_lut (.I0(GND_net), 
            .I1(n1928), .I2(VCC_net), .I3(n44093), .O(n1995)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1302_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1302_8 (.CI(n44093), 
            .I0(n1928), .I1(VCC_net), .CO(n44094));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_2106_25_lut (.I0(GND_net), 
            .I1(n3111), .I2(VCC_net), .I3(n44380), .O(n3178)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_2106_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1302_7_lut (.I0(GND_net), 
            .I1(n1929), .I2(GND_net), .I3(n44092), .O(n1996)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1302_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_2106_25 (.CI(n44380), 
            .I0(n3111), .I1(VCC_net), .CO(n44381));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1302_7 (.CI(n44092), 
            .I0(n1929), .I1(GND_net), .CO(n44093));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_2106_24_lut (.I0(GND_net), 
            .I1(n3112), .I2(VCC_net), .I3(n44379), .O(n3179)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_2106_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_2106_24 (.CI(n44379), 
            .I0(n3112), .I1(VCC_net), .CO(n44380));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1302_6_lut (.I0(GND_net), 
            .I1(n1930), .I2(GND_net), .I3(n44091), .O(n1997)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1302_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1302_6 (.CI(n44091), 
            .I0(n1930), .I1(GND_net), .CO(n44092));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_2106_23_lut (.I0(GND_net), 
            .I1(n3113), .I2(VCC_net), .I3(n44378), .O(n3180)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_2106_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_2106_23 (.CI(n44378), 
            .I0(n3113), .I1(VCC_net), .CO(n44379));
    SB_CARRY add_263_10 (.CI(n43542), .I0(encoder1_position[11]), .I1(GND_net), 
            .CO(n43543));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1302_5_lut (.I0(GND_net), 
            .I1(n1931), .I2(VCC_net), .I3(n44090), .O(n1998)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1302_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_2106_22_lut (.I0(GND_net), 
            .I1(n3114), .I2(VCC_net), .I3(n44377), .O(n3181)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_2106_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_261_2 (.CI(GND_net), .I0(duty[3]), .I1(n211), .CO(n43558));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_2106_22 (.CI(n44377), 
            .I0(n3114), .I1(VCC_net), .CO(n44378));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1302_5 (.CI(n44090), 
            .I0(n1931), .I1(VCC_net), .CO(n44091));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_2106_21_lut (.I0(GND_net), 
            .I1(n3115), .I2(VCC_net), .I3(n44376), .O(n3182)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_2106_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_2106_21 (.CI(n44376), 
            .I0(n3115), .I1(VCC_net), .CO(n44377));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1302_4_lut (.I0(GND_net), 
            .I1(n1932), .I2(GND_net), .I3(n44089), .O(n1999)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1302_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1302_4 (.CI(n44089), 
            .I0(n1932), .I1(GND_net), .CO(n44090));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1302_3_lut (.I0(GND_net), 
            .I1(n1933), .I2(VCC_net), .I3(n44088), .O(n2000)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1302_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1302_3 (.CI(n44088), 
            .I0(n1933), .I1(VCC_net), .CO(n44089));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1302_2_lut (.I0(GND_net), 
            .I1(n530), .I2(GND_net), .I3(VCC_net), .O(n2001)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1302_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_2106_20_lut (.I0(GND_net), 
            .I1(n3116), .I2(VCC_net), .I3(n44375), .O(n3183)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_2106_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_2106_20 (.CI(n44375), 
            .I0(n3116), .I1(VCC_net), .CO(n44376));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_2106_19_lut (.I0(GND_net), 
            .I1(n3117), .I2(VCC_net), .I3(n44374), .O(n3184)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_2106_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_2106_19 (.CI(n44374), 
            .I0(n3117), .I1(VCC_net), .CO(n44375));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1302_2 (.CI(VCC_net), 
            .I0(n530), .I1(GND_net), .CO(n44088));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1235_18_lut (.I0(n56323), 
            .I1(n1818), .I2(VCC_net), .I3(n44087), .O(n1917)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1235_18_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1235_17_lut (.I0(GND_net), 
            .I1(n1819), .I2(VCC_net), .I3(n44086), .O(n1886)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1235_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_2106_18_lut (.I0(GND_net), 
            .I1(n3118), .I2(VCC_net), .I3(n44373), .O(n3185)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_2106_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_2106_18 (.CI(n44373), 
            .I0(n3118), .I1(VCC_net), .CO(n44374));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1235_17 (.CI(n44086), 
            .I0(n1819), .I1(VCC_net), .CO(n44087));
    SB_LUT4 add_263_2_lut (.I0(GND_net), .I1(encoder1_position[3]), .I2(encoder1_position_scaled_23__N_359), 
            .I3(GND_net), .O(encoder1_position_scaled_23__N_75[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_263_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_263_9_lut (.I0(GND_net), .I1(encoder1_position[10]), .I2(GND_net), 
            .I3(n43541), .O(encoder1_position_scaled_23__N_75[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_263_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_263_25_lut (.I0(GND_net), .I1(encoder1_position[26]), .I2(GND_net), 
            .I3(n43557), .O(encoder1_position_scaled_23__N_75[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_263_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_2106_17_lut (.I0(GND_net), 
            .I1(n3119), .I2(VCC_net), .I3(n44372), .O(n3186)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_2106_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_263_24_lut (.I0(GND_net), .I1(encoder1_position[25]), .I2(GND_net), 
            .I3(n43556), .O(encoder1_position_scaled_23__N_75[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_263_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_2106_17 (.CI(n44372), 
            .I0(n3119), .I1(VCC_net), .CO(n44373));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_2106_16_lut (.I0(GND_net), 
            .I1(n3120), .I2(VCC_net), .I3(n44371), .O(n3187)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_2106_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_263_9 (.CI(n43541), .I0(encoder1_position[10]), .I1(GND_net), 
            .CO(n43542));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1235_16_lut (.I0(GND_net), 
            .I1(n1820), .I2(VCC_net), .I3(n44085), .O(n1887)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1235_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1235_16 (.CI(n44085), 
            .I0(n1820), .I1(VCC_net), .CO(n44086));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1235_15_lut (.I0(GND_net), 
            .I1(n1821), .I2(VCC_net), .I3(n44084), .O(n1888)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1235_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1235_15 (.CI(n44084), 
            .I0(n1821), .I1(VCC_net), .CO(n44085));
    SB_CARRY add_263_24 (.CI(n43556), .I0(encoder1_position[25]), .I1(GND_net), 
            .CO(n43557));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1235_14_lut (.I0(GND_net), 
            .I1(n1822), .I2(VCC_net), .I3(n44083), .O(n1889)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1235_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_263_23_lut (.I0(GND_net), .I1(encoder1_position[24]), .I2(GND_net), 
            .I3(n43555), .O(encoder1_position_scaled_23__N_75[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_263_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_263_23 (.CI(n43555), .I0(encoder1_position[24]), .I1(GND_net), 
            .CO(n43556));
    SB_LUT4 mux_281_i6_4_lut (.I0(encoder1_position_scaled[5]), .I1(displacement[5]), 
            .I2(n15), .I3(n15_adj_5471), .O(motor_state_23__N_123[5]));   // verilog/TinyFPGA_B.v(284[5] 286[10])
    defparam mux_281_i6_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 add_263_22_lut (.I0(GND_net), .I1(encoder1_position[23]), .I2(GND_net), 
            .I3(n43554), .O(encoder1_position_scaled_23__N_75[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_263_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_263_22 (.CI(n43554), .I0(encoder1_position[23]), .I1(GND_net), 
            .CO(n43555));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_2106_16 (.CI(n44371), 
            .I0(n3120), .I1(VCC_net), .CO(n44372));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_2106_15_lut (.I0(GND_net), 
            .I1(n3121), .I2(VCC_net), .I3(n44370), .O(n3188)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_2106_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_2106_15 (.CI(n44370), 
            .I0(n3121), .I1(VCC_net), .CO(n44371));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_2106_14_lut (.I0(GND_net), 
            .I1(n3122), .I2(VCC_net), .I3(n44369), .O(n3189)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_2106_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_2106_14 (.CI(n44369), 
            .I0(n3122), .I1(VCC_net), .CO(n44370));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1235_14 (.CI(n44083), 
            .I0(n1822), .I1(VCC_net), .CO(n44084));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_2106_13_lut (.I0(GND_net), 
            .I1(n3123), .I2(VCC_net), .I3(n44368), .O(n3190)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_2106_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1235_13_lut (.I0(GND_net), 
            .I1(n1823), .I2(VCC_net), .I3(n44082), .O(n1890)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1235_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_2106_13 (.CI(n44368), 
            .I0(n3123), .I1(VCC_net), .CO(n44369));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1235_13 (.CI(n44082), 
            .I0(n1823), .I1(VCC_net), .CO(n44083));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_2106_12_lut (.I0(GND_net), 
            .I1(n3124), .I2(VCC_net), .I3(n44367), .O(n3191)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_2106_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i40402_1_lut (.I0(n2247), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n56233));
    defparam i40402_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1235_12_lut (.I0(GND_net), 
            .I1(n1824), .I2(VCC_net), .I3(n44081), .O(n1891)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1235_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1235_12 (.CI(n44081), 
            .I0(n1824), .I1(VCC_net), .CO(n44082));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1235_11_lut (.I0(GND_net), 
            .I1(n1825), .I2(VCC_net), .I3(n44080), .O(n1892)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1235_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_2106_12 (.CI(n44367), 
            .I0(n3124), .I1(VCC_net), .CO(n44368));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1235_11 (.CI(n44080), 
            .I0(n1825), .I1(VCC_net), .CO(n44081));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_2106_11_lut (.I0(GND_net), 
            .I1(n3125), .I2(VCC_net), .I3(n44366), .O(n3192)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_2106_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_2106_11 (.CI(n44366), 
            .I0(n3125), .I1(VCC_net), .CO(n44367));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1235_10_lut (.I0(GND_net), 
            .I1(n1826), .I2(VCC_net), .I3(n44079), .O(n1893)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1235_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_2106_10_lut (.I0(GND_net), 
            .I1(n3126), .I2(VCC_net), .I3(n44365), .O(n3193)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_2106_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1235_10 (.CI(n44079), 
            .I0(n1826), .I1(VCC_net), .CO(n44080));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_2106_10 (.CI(n44365), 
            .I0(n3126), .I1(VCC_net), .CO(n44366));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1235_9_lut (.I0(GND_net), 
            .I1(n1827), .I2(VCC_net), .I3(n44078), .O(n1894)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1235_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1235_9 (.CI(n44078), 
            .I0(n1827), .I1(VCC_net), .CO(n44079));
    SB_LUT4 n10829_bdd_4_lut_40836 (.I0(n10829), .I1(n437), .I2(current[4]), 
            .I3(duty[23]), .O(n56658));
    defparam n10829_bdd_4_lut_40836.LUT_INIT = 16'he4aa;
    SB_LUT4 add_261_23_lut (.I0(current[15]), .I1(duty[23]), .I2(n56614), 
            .I3(n43578), .O(n249)) /* synthesis syn_instantiated=1 */ ;
    defparam add_261_23_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 n56658_bdd_4_lut (.I0(n56658), .I1(duty[4]), .I2(n266), .I3(duty[23]), 
            .O(pwm_setpoint_23__N_11[4]));
    defparam n56658_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_2106_9_lut (.I0(GND_net), 
            .I1(n3127), .I2(VCC_net), .I3(n44364), .O(n3194)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_2106_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_2106_9 (.CI(n44364), 
            .I0(n3127), .I1(VCC_net), .CO(n44365));
    SB_LUT4 n10829_bdd_4_lut_40821 (.I0(n10829), .I1(n438), .I2(current[3]), 
            .I3(duty[23]), .O(n56652));
    defparam n10829_bdd_4_lut_40821.LUT_INIT = 16'he4aa;
    SB_LUT4 n56652_bdd_4_lut (.I0(n56652), .I1(duty[3]), .I2(n267), .I3(duty[23]), 
            .O(pwm_setpoint_23__N_11[3]));
    defparam n56652_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_2106_8_lut (.I0(GND_net), 
            .I1(n3128), .I2(VCC_net), .I3(n44363), .O(n3195)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_2106_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_2106_8 (.CI(n44363), 
            .I0(n3128), .I1(VCC_net), .CO(n44364));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1235_8_lut (.I0(GND_net), 
            .I1(n1828), .I2(VCC_net), .I3(n44077), .O(n1895)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1235_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_2106_7_lut (.I0(GND_net), 
            .I1(n3129), .I2(GND_net), .I3(n44362), .O(n3196)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_2106_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1235_8 (.CI(n44077), 
            .I0(n1828), .I1(VCC_net), .CO(n44078));
    SB_DFFESR GLA_211 (.Q(INLA_c_0), .C(clk16MHz), .E(n28672), .D(GLA_N_495), 
            .R(n29145));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_2106_7 (.CI(n44362), 
            .I0(n3129), .I1(GND_net), .CO(n44363));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1235_7_lut (.I0(GND_net), 
            .I1(n1829), .I2(GND_net), .I3(n44076), .O(n1896)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1235_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_2106_6_lut (.I0(GND_net), 
            .I1(n3130), .I2(GND_net), .I3(n44361), .O(n3197)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_2106_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1235_7 (.CI(n44076), 
            .I0(n1829), .I1(GND_net), .CO(n44077));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_2106_6 (.CI(n44361), 
            .I0(n3130), .I1(GND_net), .CO(n44362));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_2106_5_lut (.I0(GND_net), 
            .I1(n3131), .I2(VCC_net), .I3(n44360), .O(n3198)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_2106_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_2106_5 (.CI(n44360), 
            .I0(n3131), .I1(VCC_net), .CO(n44361));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1235_6_lut (.I0(GND_net), 
            .I1(n1830), .I2(GND_net), .I3(n44075), .O(n1897)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1235_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i911_3_lut (.I0(n1332), .I1(n1399), 
            .I2(n1356), .I3(GND_net), .O(n1431));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i911_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1235_6 (.CI(n44075), 
            .I0(n1830), .I1(GND_net), .CO(n44076));
    SB_LUT4 add_261_22_lut (.I0(current[15]), .I1(duty[23]), .I2(n56614), 
            .I3(n43577), .O(n250)) /* synthesis syn_instantiated=1 */ ;
    defparam add_261_22_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_2106_4_lut (.I0(GND_net), 
            .I1(n3132), .I2(GND_net), .I3(n44359), .O(n3199)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_2106_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_2106_4 (.CI(n44359), 
            .I0(n3132), .I1(GND_net), .CO(n44360));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_2106_3_lut (.I0(GND_net), 
            .I1(n3133), .I2(VCC_net), .I3(n44358), .O(n3200)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_2106_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1235_5_lut (.I0(GND_net), 
            .I1(n1831), .I2(VCC_net), .I3(n44074), .O(n1898)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1235_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_2106_3 (.CI(n44358), 
            .I0(n3133), .I1(VCC_net), .CO(n44359));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_2106_2_lut (.I0(GND_net), 
            .I1(n542), .I2(GND_net), .I3(VCC_net), .O(n3201)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_2106_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_2106_2 (.CI(VCC_net), 
            .I0(n542), .I1(GND_net), .CO(n44358));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_2039_30_lut (.I0(n56595), 
            .I1(n3006), .I2(VCC_net), .I3(n44357), .O(n3105)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_2039_30_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_2039_29_lut (.I0(GND_net), 
            .I1(n3007), .I2(VCC_net), .I3(n44356), .O(n3074)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_2039_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_2039_29 (.CI(n44356), 
            .I0(n3007), .I1(VCC_net), .CO(n44357));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_2039_28_lut (.I0(GND_net), 
            .I1(n3008), .I2(VCC_net), .I3(n44355), .O(n3075)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_2039_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_2039_28 (.CI(n44355), 
            .I0(n3008), .I1(VCC_net), .CO(n44356));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_2039_27_lut (.I0(GND_net), 
            .I1(n3009), .I2(VCC_net), .I3(n44354), .O(n3076)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_2039_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_2039_27 (.CI(n44354), 
            .I0(n3009), .I1(VCC_net), .CO(n44355));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1235_5 (.CI(n44074), 
            .I0(n1831), .I1(VCC_net), .CO(n44075));
    SB_LUT4 mux_281_i7_4_lut (.I0(encoder1_position_scaled[6]), .I1(displacement[6]), 
            .I2(n15), .I3(n15_adj_5471), .O(motor_state_23__N_123[6]));   // verilog/TinyFPGA_B.v(284[5] 286[10])
    defparam mux_281_i7_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1235_4_lut (.I0(GND_net), 
            .I1(n1832), .I2(GND_net), .I3(n44073), .O(n1899)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1235_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1235_4 (.CI(n44073), 
            .I0(n1832), .I1(GND_net), .CO(n44074));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1235_3_lut (.I0(GND_net), 
            .I1(n1833), .I2(VCC_net), .I3(n44072), .O(n1900)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1235_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1235_3 (.CI(n44072), 
            .I0(n1833), .I1(VCC_net), .CO(n44073));
    SB_CARRY add_261_22 (.CI(n43577), .I0(duty[23]), .I1(n56614), .CO(n43578));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_2039_26_lut (.I0(GND_net), 
            .I1(n3010), .I2(VCC_net), .I3(n44353), .O(n3077)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_2039_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_2039_26 (.CI(n44353), 
            .I0(n3010), .I1(VCC_net), .CO(n44354));
    SB_LUT4 add_261_21_lut (.I0(current[15]), .I1(duty[22]), .I2(n56614), 
            .I3(n43576), .O(n251)) /* synthesis syn_instantiated=1 */ ;
    defparam add_261_21_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_2039_25_lut (.I0(GND_net), 
            .I1(n3011), .I2(VCC_net), .I3(n44352), .O(n3078)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_2039_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_2039_25 (.CI(n44352), 
            .I0(n3011), .I1(VCC_net), .CO(n44353));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_2039_24_lut (.I0(GND_net), 
            .I1(n3012), .I2(VCC_net), .I3(n44351), .O(n3079)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_2039_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_2039_24 (.CI(n44351), 
            .I0(n3012), .I1(VCC_net), .CO(n44352));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1235_2_lut (.I0(GND_net), 
            .I1(n529), .I2(GND_net), .I3(VCC_net), .O(n1901)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1235_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1235_2 (.CI(VCC_net), 
            .I0(n529), .I1(GND_net), .CO(n44072));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1168_17_lut (.I0(n56328), 
            .I1(n1719), .I2(VCC_net), .I3(n44071), .O(n1818)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1168_17_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_2039_23_lut (.I0(GND_net), 
            .I1(n3013), .I2(VCC_net), .I3(n44350), .O(n3080)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_2039_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_2039_23 (.CI(n44350), 
            .I0(n3013), .I1(VCC_net), .CO(n44351));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_2039_22_lut (.I0(GND_net), 
            .I1(n3014), .I2(VCC_net), .I3(n44349), .O(n3081)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_2039_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_2039_22 (.CI(n44349), 
            .I0(n3014), .I1(VCC_net), .CO(n44350));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_2039_21_lut (.I0(GND_net), 
            .I1(n3015), .I2(VCC_net), .I3(n44348), .O(n3082)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_2039_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_2039_21 (.CI(n44348), 
            .I0(n3015), .I1(VCC_net), .CO(n44349));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1168_16_lut (.I0(GND_net), 
            .I1(n1720), .I2(VCC_net), .I3(n44070), .O(n1787)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1168_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_261_21 (.CI(n43576), .I0(duty[22]), .I1(n56614), .CO(n43577));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1168_16 (.CI(n44070), 
            .I0(n1720), .I1(VCC_net), .CO(n44071));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_2039_20_lut (.I0(GND_net), 
            .I1(n3016), .I2(VCC_net), .I3(n44347), .O(n3083)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_2039_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1168_15_lut (.I0(GND_net), 
            .I1(n1721), .I2(VCC_net), .I3(n44069), .O(n1788)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1168_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_2039_20 (.CI(n44347), 
            .I0(n3016), .I1(VCC_net), .CO(n44348));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_2039_19_lut (.I0(GND_net), 
            .I1(n3017), .I2(VCC_net), .I3(n44346), .O(n3084)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_2039_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_2039_19 (.CI(n44346), 
            .I0(n3017), .I1(VCC_net), .CO(n44347));
    SB_LUT4 add_263_8_lut (.I0(GND_net), .I1(encoder1_position[9]), .I2(GND_net), 
            .I3(n43540), .O(encoder1_position_scaled_23__N_75[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_263_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_2039_18_lut (.I0(GND_net), 
            .I1(n3018), .I2(VCC_net), .I3(n44345), .O(n3085)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_2039_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_2039_18 (.CI(n44345), 
            .I0(n3018), .I1(VCC_net), .CO(n44346));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1168_15 (.CI(n44069), 
            .I0(n1721), .I1(VCC_net), .CO(n44070));
    SB_LUT4 i15830_3_lut (.I0(\PID_CONTROLLER.integral [6]), .I1(\PID_CONTROLLER.integral_23__N_3996 [6]), 
            .I2(control_update), .I3(GND_net), .O(n29910));   // verilog/motorControl.v(41[14] 61[8])
    defparam i15830_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_2039_17_lut (.I0(GND_net), 
            .I1(n3019), .I2(VCC_net), .I3(n44344), .O(n3086)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_2039_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15831_3_lut (.I0(\PID_CONTROLLER.integral [5]), .I1(\PID_CONTROLLER.integral_23__N_3996 [5]), 
            .I2(control_update), .I3(GND_net), .O(n29911));   // verilog/motorControl.v(41[14] 61[8])
    defparam i15831_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_261_20_lut (.I0(current[15]), .I1(duty[21]), .I2(n56614), 
            .I3(n43575), .O(n252)) /* synthesis syn_instantiated=1 */ ;
    defparam add_261_20_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 add_263_21_lut (.I0(GND_net), .I1(encoder1_position[22]), .I2(GND_net), 
            .I3(n43553), .O(encoder1_position_scaled_23__N_75[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_263_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_263_21 (.CI(n43553), .I0(encoder1_position[22]), .I1(GND_net), 
            .CO(n43554));
    SB_CARRY add_261_20 (.CI(n43575), .I0(duty[21]), .I1(n56614), .CO(n43576));
    SB_LUT4 add_263_20_lut (.I0(GND_net), .I1(encoder1_position[21]), .I2(GND_net), 
            .I3(n43552), .O(encoder1_position_scaled_23__N_75[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_263_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_263_20 (.CI(n43552), .I0(encoder1_position[21]), .I1(GND_net), 
            .CO(n43553));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_2039_17 (.CI(n44344), 
            .I0(n3019), .I1(VCC_net), .CO(n44345));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1168_14_lut (.I0(GND_net), 
            .I1(n1722), .I2(VCC_net), .I3(n44068), .O(n1789)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1168_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1168_14 (.CI(n44068), 
            .I0(n1722), .I1(VCC_net), .CO(n44069));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1168_13_lut (.I0(GND_net), 
            .I1(n1723), .I2(VCC_net), .I3(n44067), .O(n1790)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1168_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_2039_16_lut (.I0(GND_net), 
            .I1(n3020), .I2(VCC_net), .I3(n44343), .O(n3087)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_2039_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_263_19_lut (.I0(GND_net), .I1(encoder1_position[20]), .I2(GND_net), 
            .I3(n43551), .O(encoder1_position_scaled_23__N_75[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_263_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_2039_16 (.CI(n44343), 
            .I0(n3020), .I1(VCC_net), .CO(n44344));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1168_13 (.CI(n44067), 
            .I0(n1723), .I1(VCC_net), .CO(n44068));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_2039_15_lut (.I0(GND_net), 
            .I1(n3021), .I2(VCC_net), .I3(n44342), .O(n3088)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_2039_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15832_3_lut (.I0(\PID_CONTROLLER.integral [4]), .I1(\PID_CONTROLLER.integral_23__N_3996 [4]), 
            .I2(control_update), .I3(GND_net), .O(n29912));   // verilog/motorControl.v(41[14] 61[8])
    defparam i15832_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1168_12_lut (.I0(GND_net), 
            .I1(n1724), .I2(VCC_net), .I3(n44066), .O(n1791)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1168_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1168_12 (.CI(n44066), 
            .I0(n1724), .I1(VCC_net), .CO(n44067));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1168_11_lut (.I0(GND_net), 
            .I1(n1725), .I2(VCC_net), .I3(n44065), .O(n1792)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1168_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1168_11 (.CI(n44065), 
            .I0(n1725), .I1(VCC_net), .CO(n44066));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_2039_15 (.CI(n44342), 
            .I0(n3021), .I1(VCC_net), .CO(n44343));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_2039_14_lut (.I0(GND_net), 
            .I1(n3022), .I2(VCC_net), .I3(n44341), .O(n3089)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_2039_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_261_19_lut (.I0(current[15]), .I1(duty[20]), .I2(n56614), 
            .I3(n43574), .O(n253)) /* synthesis syn_instantiated=1 */ ;
    defparam add_261_19_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1168_10_lut (.I0(GND_net), 
            .I1(n1726), .I2(VCC_net), .I3(n44064), .O(n1793)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1168_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_2039_14 (.CI(n44341), 
            .I0(n3022), .I1(VCC_net), .CO(n44342));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1168_10 (.CI(n44064), 
            .I0(n1726), .I1(VCC_net), .CO(n44065));
    SB_LUT4 i15833_3_lut (.I0(\PID_CONTROLLER.integral [3]), .I1(\PID_CONTROLLER.integral_23__N_3996 [3]), 
            .I2(control_update), .I3(GND_net), .O(n29913));   // verilog/motorControl.v(41[14] 61[8])
    defparam i15833_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_2039_13_lut (.I0(GND_net), 
            .I1(n3023), .I2(VCC_net), .I3(n44340), .O(n3090)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_2039_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_2039_13 (.CI(n44340), 
            .I0(n3023), .I1(VCC_net), .CO(n44341));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_2039_12_lut (.I0(GND_net), 
            .I1(n3024), .I2(VCC_net), .I3(n44339), .O(n3091)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_2039_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_2039_12 (.CI(n44339), 
            .I0(n3024), .I1(VCC_net), .CO(n44340));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1168_9_lut (.I0(GND_net), 
            .I1(n1727), .I2(VCC_net), .I3(n44063), .O(n1794)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1168_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_2039_11_lut (.I0(GND_net), 
            .I1(n3025), .I2(VCC_net), .I3(n44338), .O(n3092)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_2039_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_2039_11 (.CI(n44338), 
            .I0(n3025), .I1(VCC_net), .CO(n44339));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1168_9 (.CI(n44063), 
            .I0(n1727), .I1(VCC_net), .CO(n44064));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_2039_10_lut (.I0(GND_net), 
            .I1(n3026), .I2(VCC_net), .I3(n44337), .O(n3093)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_2039_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_2039_10 (.CI(n44337), 
            .I0(n3026), .I1(VCC_net), .CO(n44338));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_2039_9_lut (.I0(GND_net), 
            .I1(n3027), .I2(VCC_net), .I3(n44336), .O(n3094)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_2039_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1168_8_lut (.I0(GND_net), 
            .I1(n1728), .I2(VCC_net), .I3(n44062), .O(n1795)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1168_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_2039_9 (.CI(n44336), 
            .I0(n3027), .I1(VCC_net), .CO(n44337));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_2039_8_lut (.I0(GND_net), 
            .I1(n3028), .I2(VCC_net), .I3(n44335), .O(n3095)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_2039_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1168_8 (.CI(n44062), 
            .I0(n1728), .I1(VCC_net), .CO(n44063));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1168_7_lut (.I0(GND_net), 
            .I1(n1729), .I2(GND_net), .I3(n44061), .O(n1796)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1168_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1168_7 (.CI(n44061), 
            .I0(n1729), .I1(GND_net), .CO(n44062));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1168_6_lut (.I0(GND_net), 
            .I1(n1730), .I2(GND_net), .I3(n44060), .O(n1797)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1168_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_2039_8 (.CI(n44335), 
            .I0(n3028), .I1(VCC_net), .CO(n44336));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1168_6 (.CI(n44060), 
            .I0(n1730), .I1(GND_net), .CO(n44061));
    SB_LUT4 i15834_3_lut (.I0(\PID_CONTROLLER.integral [2]), .I1(\PID_CONTROLLER.integral_23__N_3996 [2]), 
            .I2(control_update), .I3(GND_net), .O(n29914));   // verilog/motorControl.v(41[14] 61[8])
    defparam i15834_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_2039_7_lut (.I0(GND_net), 
            .I1(n3029), .I2(GND_net), .I3(n44334), .O(n3096)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_2039_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_2039_7 (.CI(n44334), 
            .I0(n3029), .I1(GND_net), .CO(n44335));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_2039_6_lut (.I0(GND_net), 
            .I1(n3030), .I2(GND_net), .I3(n44333), .O(n3097)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_2039_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_2039_6 (.CI(n44333), 
            .I0(n3030), .I1(GND_net), .CO(n44334));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_2039_5_lut (.I0(GND_net), 
            .I1(n3031), .I2(VCC_net), .I3(n44332), .O(n3098)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_2039_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1168_5_lut (.I0(GND_net), 
            .I1(n1731), .I2(VCC_net), .I3(n44059), .O(n1798)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1168_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1168_5 (.CI(n44059), 
            .I0(n1731), .I1(VCC_net), .CO(n44060));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1168_4_lut (.I0(GND_net), 
            .I1(n1732), .I2(GND_net), .I3(n44058), .O(n1799)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1168_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1168_4 (.CI(n44058), 
            .I0(n1732), .I1(GND_net), .CO(n44059));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_2039_5 (.CI(n44332), 
            .I0(n3031), .I1(VCC_net), .CO(n44333));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1168_3_lut (.I0(GND_net), 
            .I1(n1733), .I2(VCC_net), .I3(n44057), .O(n1800)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1168_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_21_add_3_26_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_setpoint_23__N_263), 
            .I3(n43664), .O(n356)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_2039_4_lut (.I0(GND_net), 
            .I1(n3032), .I2(GND_net), .I3(n44331), .O(n3099)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_2039_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_2039_4 (.CI(n44331), 
            .I0(n3032), .I1(GND_net), .CO(n44332));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_2039_3_lut (.I0(GND_net), 
            .I1(n3033), .I2(VCC_net), .I3(n44330), .O(n3100)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_2039_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_2039_3 (.CI(n44330), 
            .I0(n3033), .I1(VCC_net), .CO(n44331));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_2039_2_lut (.I0(GND_net), 
            .I1(n541), .I2(GND_net), .I3(VCC_net), .O(n3101)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_2039_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_33_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n2_adj_5611), .I3(n44696), .O(n2_adj_5497)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_33_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1168_3 (.CI(n44057), 
            .I0(n1733), .I1(VCC_net), .CO(n44058));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_2039_2 (.CI(VCC_net), 
            .I0(n541), .I1(GND_net), .CO(n44330));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1168_2_lut (.I0(GND_net), 
            .I1(n942), .I2(GND_net), .I3(VCC_net), .O(n1801)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1168_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_21_add_3_25_lut (.I0(n4748), .I1(GND_net), .I2(pwm_setpoint_23__N_263), 
            .I3(n43663), .O(n4884)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_25_lut.LUT_INIT = 16'h8228;
    SB_CARRY unary_minus_21_add_3_25 (.CI(n43663), .I0(GND_net), .I1(pwm_setpoint_23__N_263), 
            .CO(n43664));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1972_29_lut (.I0(n56025), 
            .I1(n2907), .I2(VCC_net), .I3(n44329), .O(n3006)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1972_29_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1972_28_lut (.I0(GND_net), 
            .I1(n2908), .I2(VCC_net), .I3(n44328), .O(n2975)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1972_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1972_28 (.CI(n44328), 
            .I0(n2908), .I1(VCC_net), .CO(n44329));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1972_27_lut (.I0(GND_net), 
            .I1(n2909), .I2(VCC_net), .I3(n44327), .O(n2976)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1972_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1168_2 (.CI(VCC_net), 
            .I0(n942), .I1(GND_net), .CO(n44057));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1101_16_lut (.I0(n56364), 
            .I1(n1620), .I2(VCC_net), .I3(n44056), .O(n1719)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1101_16_lut.LUT_INIT = 16'h8228;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1972_27 (.CI(n44327), 
            .I0(n2909), .I1(VCC_net), .CO(n44328));
    SB_CARRY add_261_19 (.CI(n43574), .I0(duty[20]), .I1(n56614), .CO(n43575));
    SB_LUT4 unary_minus_21_add_3_24_lut (.I0(n4748), .I1(GND_net), .I2(n3), 
            .I3(n43662), .O(n4885)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_24_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1972_26_lut (.I0(GND_net), 
            .I1(n2910), .I2(VCC_net), .I3(n44326), .O(n2977)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1972_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_32_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n3_adj_5612), .I3(n44695), .O(n3_adj_5496)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_32_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1972_26 (.CI(n44326), 
            .I0(n2910), .I1(VCC_net), .CO(n44327));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1972_25_lut (.I0(GND_net), 
            .I1(n2911), .I2(VCC_net), .I3(n44325), .O(n2978)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1972_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_32 (.CI(n44695), 
            .I0(GND_net), .I1(n3_adj_5612), .CO(n44696));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1972_25 (.CI(n44325), 
            .I0(n2911), .I1(VCC_net), .CO(n44326));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1972_24_lut (.I0(GND_net), 
            .I1(n2912), .I2(VCC_net), .I3(n44324), .O(n2979)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1972_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1101_15_lut (.I0(GND_net), 
            .I1(n1621), .I2(VCC_net), .I3(n44055), .O(n1688)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1101_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_31_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n4_adj_5613), .I3(n44694), .O(n4_adj_5495)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_31_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1972_24 (.CI(n44324), 
            .I0(n2912), .I1(VCC_net), .CO(n44325));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1972_23_lut (.I0(GND_net), 
            .I1(n2913), .I2(VCC_net), .I3(n44323), .O(n2980)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1972_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1972_23 (.CI(n44323), 
            .I0(n2913), .I1(VCC_net), .CO(n44324));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1101_15 (.CI(n44055), 
            .I0(n1621), .I1(VCC_net), .CO(n44056));
    SB_CARRY encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_31 (.CI(n44694), 
            .I0(GND_net), .I1(n4_adj_5613), .CO(n44695));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1101_14_lut (.I0(GND_net), 
            .I1(n1622), .I2(VCC_net), .I3(n44054), .O(n1689)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1101_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1101_14 (.CI(n44054), 
            .I0(n1622), .I1(VCC_net), .CO(n44055));
    SB_CARRY unary_minus_21_add_3_24 (.CI(n43662), .I0(GND_net), .I1(n3), 
            .CO(n43663));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1972_22_lut (.I0(GND_net), 
            .I1(n2914), .I2(VCC_net), .I3(n44322), .O(n2981)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1972_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_30_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n5_adj_5614), .I3(n44693), .O(n5_adj_5494)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1972_22 (.CI(n44322), 
            .I0(n2914), .I1(VCC_net), .CO(n44323));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1972_21_lut (.I0(GND_net), 
            .I1(n2915), .I2(VCC_net), .I3(n44321), .O(n2982)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1972_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1101_13_lut (.I0(GND_net), 
            .I1(n1623), .I2(VCC_net), .I3(n44053), .O(n1690)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1101_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1101_13 (.CI(n44053), 
            .I0(n1623), .I1(VCC_net), .CO(n44054));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1972_21 (.CI(n44321), 
            .I0(n2915), .I1(VCC_net), .CO(n44322));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1101_12_lut (.I0(GND_net), 
            .I1(n1624), .I2(VCC_net), .I3(n44052), .O(n1691)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1101_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1972_20_lut (.I0(GND_net), 
            .I1(n2916), .I2(VCC_net), .I3(n44320), .O(n2983)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1972_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_30 (.CI(n44693), 
            .I0(GND_net), .I1(n5_adj_5614), .CO(n44694));
    SB_LUT4 add_261_18_lut (.I0(current[15]), .I1(duty[19]), .I2(n56614), 
            .I3(n43573), .O(n254)) /* synthesis syn_instantiated=1 */ ;
    defparam add_261_18_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY add_261_18 (.CI(n43573), .I0(duty[19]), .I1(n56614), .CO(n43574));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_29_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n6_adj_5615), .I3(n44692), .O(n6_adj_5493)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1972_20 (.CI(n44320), 
            .I0(n2916), .I1(VCC_net), .CO(n44321));
    SB_LUT4 unary_minus_21_add_3_23_lut (.I0(n4748), .I1(GND_net), .I2(n4_adj_5446), 
            .I3(n43661), .O(n4886)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_23_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1972_19_lut (.I0(GND_net), 
            .I1(n2917), .I2(VCC_net), .I3(n44319), .O(n2984)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1972_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1972_19 (.CI(n44319), 
            .I0(n2917), .I1(VCC_net), .CO(n44320));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1101_12 (.CI(n44052), 
            .I0(n1624), .I1(VCC_net), .CO(n44053));
    SB_CARRY unary_minus_21_add_3_23 (.CI(n43661), .I0(GND_net), .I1(n4_adj_5446), 
            .CO(n43662));
    SB_CARRY encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_29 (.CI(n44692), 
            .I0(GND_net), .I1(n6_adj_5615), .CO(n44693));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1972_18_lut (.I0(GND_net), 
            .I1(n2918), .I2(VCC_net), .I3(n44318), .O(n2985)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1972_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_21_add_3_22_lut (.I0(n4748), .I1(GND_net), .I2(n5_adj_5447), 
            .I3(n43660), .O(n4887)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_22_lut.LUT_INIT = 16'h8228;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1972_18 (.CI(n44318), 
            .I0(n2918), .I1(VCC_net), .CO(n44319));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_28_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n7_adj_5616), .I3(n44691), .O(n7_adj_5492)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_28_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1972_17_lut (.I0(GND_net), 
            .I1(n2919), .I2(VCC_net), .I3(n44317), .O(n2986)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1972_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_28 (.CI(n44691), 
            .I0(GND_net), .I1(n7_adj_5616), .CO(n44692));
    SB_CARRY unary_minus_21_add_3_22 (.CI(n43660), .I0(GND_net), .I1(n5_adj_5447), 
            .CO(n43661));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_27_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n8_adj_5617), .I3(n44690), .O(n8_adj_5491)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1972_17 (.CI(n44317), 
            .I0(n2919), .I1(VCC_net), .CO(n44318));
    SB_LUT4 unary_minus_21_add_3_21_lut (.I0(n4748), .I1(GND_net), .I2(n6_adj_5448), 
            .I3(n43659), .O(n4888)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_21_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1101_11_lut (.I0(GND_net), 
            .I1(n1625), .I2(VCC_net), .I3(n44051), .O(n1692)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1101_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1972_16_lut (.I0(GND_net), 
            .I1(n2920), .I2(VCC_net), .I3(n44316), .O(n2987)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1972_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_261_17_lut (.I0(current[15]), .I1(duty[18]), .I2(n56614), 
            .I3(n43572), .O(n255)) /* synthesis syn_instantiated=1 */ ;
    defparam add_261_17_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY add_261_17 (.CI(n43572), .I0(duty[18]), .I1(n56614), .CO(n43573));
    SB_CARRY unary_minus_21_add_3_21 (.CI(n43659), .I0(GND_net), .I1(n6_adj_5448), 
            .CO(n43660));
    SB_LUT4 unary_minus_21_add_3_20_lut (.I0(n4748), .I1(GND_net), .I2(n7_adj_5449), 
            .I3(n43658), .O(n4889)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_20_lut.LUT_INIT = 16'h8228;
    SB_CARRY encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_27 (.CI(n44690), 
            .I0(GND_net), .I1(n8_adj_5617), .CO(n44691));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1972_16 (.CI(n44316), 
            .I0(n2920), .I1(VCC_net), .CO(n44317));
    SB_CARRY unary_minus_21_add_3_20 (.CI(n43658), .I0(GND_net), .I1(n7_adj_5449), 
            .CO(n43659));
    SB_CARRY add_263_19 (.CI(n43551), .I0(encoder1_position[20]), .I1(GND_net), 
            .CO(n43552));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1972_15_lut (.I0(GND_net), 
            .I1(n2921), .I2(VCC_net), .I3(n44315), .O(n2988)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1972_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1972_15 (.CI(n44315), 
            .I0(n2921), .I1(VCC_net), .CO(n44316));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1972_14_lut (.I0(GND_net), 
            .I1(n2922), .I2(VCC_net), .I3(n44314), .O(n2989)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1972_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1101_11 (.CI(n44051), 
            .I0(n1625), .I1(VCC_net), .CO(n44052));
    SB_LUT4 LessThan_17_i6_3_lut_3_lut (.I0(current_limit[2]), .I1(current_limit[3]), 
            .I2(current[3]), .I3(GND_net), .O(n6_adj_5587));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam LessThan_17_i6_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 unary_minus_21_add_3_19_lut (.I0(n4748), .I1(GND_net), .I2(n8_adj_5450), 
            .I3(n43657), .O(n4890)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_19_lut.LUT_INIT = 16'h8228;
    SB_CARRY unary_minus_21_add_3_19 (.CI(n43657), .I0(GND_net), .I1(n8_adj_5450), 
            .CO(n43658));
    SB_CARRY add_263_8 (.CI(n43540), .I0(encoder1_position[9]), .I1(GND_net), 
            .CO(n43541));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1972_14 (.CI(n44314), 
            .I0(n2922), .I1(VCC_net), .CO(n44315));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_26_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n9_adj_5618), .I3(n44689), .O(n9_adj_5490)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_26 (.CI(n44689), 
            .I0(GND_net), .I1(n9_adj_5618), .CO(n44690));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1101_10_lut (.I0(GND_net), 
            .I1(n1626), .I2(VCC_net), .I3(n44050), .O(n1693)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1101_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_281_i8_4_lut (.I0(encoder1_position_scaled[7]), .I1(displacement[7]), 
            .I2(n15), .I3(n15_adj_5471), .O(motor_state_23__N_123[7]));   // verilog/TinyFPGA_B.v(284[5] 286[10])
    defparam mux_281_i8_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1972_13_lut (.I0(GND_net), 
            .I1(n2923), .I2(VCC_net), .I3(n44313), .O(n2990)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1972_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i10_1_lut_adj_1868 (.I0(duty[23]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(pwm_setpoint_23__N_263));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i10_1_lut_adj_1868.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1972_13 (.CI(n44313), 
            .I0(n2923), .I1(VCC_net), .CO(n44314));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_25_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n10_adj_5619), .I3(n44688), .O(n10_adj_5489)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_25 (.CI(n44688), 
            .I0(GND_net), .I1(n10_adj_5619), .CO(n44689));
    SB_LUT4 unary_minus_21_add_3_18_lut (.I0(n4748), .I1(GND_net), .I2(n9), 
            .I3(n43656), .O(n4891)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_18_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1972_12_lut (.I0(GND_net), 
            .I1(n2924), .I2(VCC_net), .I3(n44312), .O(n2991)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1972_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1972_12 (.CI(n44312), 
            .I0(n2924), .I1(VCC_net), .CO(n44313));
    SB_CARRY unary_minus_21_add_3_18 (.CI(n43656), .I0(GND_net), .I1(n9), 
            .CO(n43657));
    SB_LUT4 add_263_18_lut (.I0(GND_net), .I1(encoder1_position[19]), .I2(GND_net), 
            .I3(n43550), .O(encoder1_position_scaled_23__N_75[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_263_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_21_add_3_17_lut (.I0(n4748), .I1(GND_net), .I2(n10_adj_5451), 
            .I3(n43655), .O(n4892)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_17_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_263_2 (.CI(GND_net), .I0(encoder1_position[3]), .I1(encoder1_position_scaled_23__N_359), 
            .CO(n43535));
    SB_CARRY unary_minus_21_add_3_17 (.CI(n43655), .I0(GND_net), .I1(n10_adj_5451), 
            .CO(n43656));
    SB_LUT4 unary_minus_21_add_3_16_lut (.I0(n4748), .I1(GND_net), .I2(n11), 
            .I3(n43654), .O(n4893)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_16_lut.LUT_INIT = 16'h8228;
    SB_CARRY unary_minus_21_add_3_16 (.CI(n43654), .I0(GND_net), .I1(n11), 
            .CO(n43655));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1972_11_lut (.I0(GND_net), 
            .I1(n2925), .I2(VCC_net), .I3(n44311), .O(n2992)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1972_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_21_add_3_15_lut (.I0(n4748), .I1(GND_net), .I2(n12), 
            .I3(n43653), .O(n4894)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_15_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_24_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n11_adj_5620), .I3(n44687), .O(n11_adj_5488)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_263_18 (.CI(n43550), .I0(encoder1_position[19]), .I1(GND_net), 
            .CO(n43551));
    SB_LUT4 add_263_7_lut (.I0(GND_net), .I1(encoder1_position[8]), .I2(GND_net), 
            .I3(n43539), .O(encoder1_position_scaled_23__N_75[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_263_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_24 (.CI(n44687), 
            .I0(GND_net), .I1(n11_adj_5620), .CO(n44688));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1101_10 (.CI(n44050), 
            .I0(n1626), .I1(VCC_net), .CO(n44051));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1972_11 (.CI(n44311), 
            .I0(n2925), .I1(VCC_net), .CO(n44312));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1101_9_lut (.I0(GND_net), 
            .I1(n1627), .I2(VCC_net), .I3(n44049), .O(n1694)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1101_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_23_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n12_adj_5621), .I3(n44686), .O(n12_adj_5487)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_21_add_3_15 (.CI(n43653), .I0(GND_net), .I1(n12), 
            .CO(n43654));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1101_9 (.CI(n44049), 
            .I0(n1627), .I1(VCC_net), .CO(n44050));
    SB_CARRY encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_23 (.CI(n44686), 
            .I0(GND_net), .I1(n12_adj_5621), .CO(n44687));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1972_10_lut (.I0(GND_net), 
            .I1(n2926), .I2(VCC_net), .I3(n44310), .O(n2993)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1972_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1972_10 (.CI(n44310), 
            .I0(n2926), .I1(VCC_net), .CO(n44311));
    SB_LUT4 unary_minus_21_add_3_14_lut (.I0(n4748), .I1(GND_net), .I2(n13), 
            .I3(n43652), .O(n4895)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_14_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_22_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n13_adj_5622), .I3(n44685), .O(n13_adj_5486)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1101_8_lut (.I0(GND_net), 
            .I1(n1628), .I2(VCC_net), .I3(n44048), .O(n1695)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1101_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_263_17_lut (.I0(GND_net), .I1(encoder1_position[18]), .I2(GND_net), 
            .I3(n43549), .O(encoder1_position_scaled_23__N_75[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_263_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1101_8 (.CI(n44048), 
            .I0(n1628), .I1(VCC_net), .CO(n44049));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1101_7_lut (.I0(GND_net), 
            .I1(n1629), .I2(GND_net), .I3(n44047), .O(n1696)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1101_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_22 (.CI(n44685), 
            .I0(GND_net), .I1(n13_adj_5622), .CO(n44686));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_21_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n14_adj_5623), .I3(n44684), .O(n14_adj_5485)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_21_add_3_14 (.CI(n43652), .I0(GND_net), .I1(n13), 
            .CO(n43653));
    SB_DFFESR GLB_213 (.Q(INLB_c_0), .C(clk16MHz), .E(n28672), .D(GLB_N_509), 
            .R(n29145));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1972_9_lut (.I0(GND_net), 
            .I1(n2927), .I2(VCC_net), .I3(n44309), .O(n2994)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1972_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1972_9 (.CI(n44309), 
            .I0(n2927), .I1(VCC_net), .CO(n44310));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1972_8_lut (.I0(GND_net), 
            .I1(n2928), .I2(VCC_net), .I3(n44308), .O(n2995)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1972_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_263_17 (.CI(n43549), .I0(encoder1_position[18]), .I1(GND_net), 
            .CO(n43550));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1972_8 (.CI(n44308), 
            .I0(n2928), .I1(VCC_net), .CO(n44309));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1972_7_lut (.I0(GND_net), 
            .I1(n2929), .I2(GND_net), .I3(n44307), .O(n2996)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1972_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1972_7 (.CI(n44307), 
            .I0(n2929), .I1(GND_net), .CO(n44308));
    SB_LUT4 unary_minus_21_add_3_13_lut (.I0(n4748), .I1(GND_net), .I2(n14), 
            .I3(n43651), .O(n4896)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_13_lut.LUT_INIT = 16'h8228;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1101_7 (.CI(n44047), 
            .I0(n1629), .I1(GND_net), .CO(n44048));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1101_6_lut (.I0(GND_net), 
            .I1(n1630), .I2(GND_net), .I3(n44046), .O(n1697)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1101_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_21 (.CI(n44684), 
            .I0(GND_net), .I1(n14_adj_5623), .CO(n44685));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1972_6_lut (.I0(GND_net), 
            .I1(n2930), .I2(GND_net), .I3(n44306), .O(n2997)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1972_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1101_6 (.CI(n44046), 
            .I0(n1630), .I1(GND_net), .CO(n44047));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1101_5_lut (.I0(GND_net), 
            .I1(n1631), .I2(VCC_net), .I3(n44045), .O(n1698)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1101_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_21_add_3_13 (.CI(n43651), .I0(GND_net), .I1(n14), 
            .CO(n43652));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_20_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n15_adj_5624), .I3(n44683), .O(n15_adj_5484)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_21_add_3_12_lut (.I0(n4748), .I1(GND_net), .I2(n15_adj_5452), 
            .I3(n43650), .O(n4897)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_12_lut.LUT_INIT = 16'h8228;
    SB_CARRY encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_20 (.CI(n44683), 
            .I0(GND_net), .I1(n15_adj_5624), .CO(n44684));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1101_5 (.CI(n44045), 
            .I0(n1631), .I1(VCC_net), .CO(n44046));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1972_6 (.CI(n44306), 
            .I0(n2930), .I1(GND_net), .CO(n44307));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_19_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n16_adj_5625), .I3(n44682), .O(n16_adj_5483)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_263_16_lut (.I0(GND_net), .I1(encoder1_position[17]), .I2(GND_net), 
            .I3(n43548), .O(encoder1_position_scaled_23__N_75[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_263_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1972_5_lut (.I0(GND_net), 
            .I1(n2931), .I2(VCC_net), .I3(n44305), .O(n2998)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1972_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1101_4_lut (.I0(GND_net), 
            .I1(n1632), .I2(GND_net), .I3(n44044), .O(n1699)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1101_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1972_5 (.CI(n44305), 
            .I0(n2931), .I1(VCC_net), .CO(n44306));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1101_4 (.CI(n44044), 
            .I0(n1632), .I1(GND_net), .CO(n44045));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1101_3_lut (.I0(GND_net), 
            .I1(n1633), .I2(VCC_net), .I3(n44043), .O(n1700)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1101_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_21_add_3_12 (.CI(n43650), .I0(GND_net), .I1(n15_adj_5452), 
            .CO(n43651));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1101_3 (.CI(n44043), 
            .I0(n1633), .I1(VCC_net), .CO(n44044));
    SB_CARRY encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_19 (.CI(n44682), 
            .I0(GND_net), .I1(n16_adj_5625), .CO(n44683));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_18_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n17_adj_5626), .I3(n44681), .O(n17_adj_5482)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15842_3_lut (.I0(PWMLimit[19]), .I1(\data_in_frame[8] [3]), 
            .I2(n50654), .I3(GND_net), .O(n29922));   // verilog/coms.v(128[12] 303[6])
    defparam i15842_3_lut.LUT_INIT = 16'hacac;
    SB_DFFESR GLC_215 (.Q(INLC_c_0), .C(clk16MHz), .E(n28672), .D(GLC_N_523), 
            .R(n29145));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    SB_LUT4 i22675_2_lut (.I0(duty[5]), .I1(n296), .I2(GND_net), .I3(GND_net), 
            .O(n4924));   // verilog/TinyFPGA_B.v(123[17] 125[11])
    defparam i22675_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1101_2_lut (.I0(GND_net), 
            .I1(n941), .I2(GND_net), .I3(VCC_net), .O(n1701)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1101_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1972_4_lut (.I0(GND_net), 
            .I1(n2932), .I2(GND_net), .I3(n44304), .O(n2999)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1972_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1972_4 (.CI(n44304), 
            .I0(n2932), .I1(GND_net), .CO(n44305));
    SB_CARRY encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_18 (.CI(n44681), 
            .I0(GND_net), .I1(n17_adj_5626), .CO(n44682));
    SB_LUT4 i39173_2_lut_4_lut (.I0(current[8]), .I1(current_limit[8]), 
            .I2(current[4]), .I3(current_limit[4]), .O(n55003));
    defparam i39173_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1972_3_lut (.I0(GND_net), 
            .I1(n2933), .I2(VCC_net), .I3(n44303), .O(n3000)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1972_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1178_3_lut (.I0(n1727), 
            .I1(n1794), .I2(n1752), .I3(GND_net), .O(n1826));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1178_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1972_3 (.CI(n44303), 
            .I0(n2933), .I1(VCC_net), .CO(n44304));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_17_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n18_adj_5627), .I3(n44680), .O(n18_adj_5481)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1972_2_lut (.I0(GND_net), 
            .I1(n540), .I2(GND_net), .I3(VCC_net), .O(n3001)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1972_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1972_2 (.CI(VCC_net), 
            .I0(n540), .I1(GND_net), .CO(n44303));
    SB_CARRY encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_17 (.CI(n44680), 
            .I0(GND_net), .I1(n18_adj_5627), .CO(n44681));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1905_28_lut (.I0(n56056), 
            .I1(n2808), .I2(VCC_net), .I3(n44302), .O(n2907)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1905_28_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_16_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n19_adj_5628), .I3(n44679), .O(n19_adj_5480)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1101_2 (.CI(VCC_net), 
            .I0(n941), .I1(GND_net), .CO(n44043));
    SB_CARRY encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_16 (.CI(n44679), 
            .I0(GND_net), .I1(n19_adj_5628), .CO(n44680));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_15_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n20_adj_5629), .I3(n44678), .O(n20_adj_5479)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_15 (.CI(n44678), 
            .I0(GND_net), .I1(n20_adj_5629), .CO(n44679));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1905_27_lut (.I0(GND_net), 
            .I1(n2809), .I2(VCC_net), .I3(n44301), .O(n2876)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1905_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1905_27 (.CI(n44301), 
            .I0(n2809), .I1(VCC_net), .CO(n44302));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1905_26_lut (.I0(GND_net), 
            .I1(n2810), .I2(VCC_net), .I3(n44300), .O(n2877)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1905_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_14_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n21_adj_5630), .I3(n44677), .O(n21_adj_5478)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_14 (.CI(n44677), 
            .I0(GND_net), .I1(n21_adj_5630), .CO(n44678));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_13_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n22_adj_5631), .I3(n44676), .O(n22_adj_5477)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1034_15_lut (.I0(n56382), 
            .I1(n1521), .I2(VCC_net), .I3(n44042), .O(n1620)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1034_15_lut.LUT_INIT = 16'h8228;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1905_26 (.CI(n44300), 
            .I0(n2810), .I1(VCC_net), .CO(n44301));
    SB_LUT4 unary_minus_21_add_3_11_lut (.I0(n4748), .I1(GND_net), .I2(n16), 
            .I3(n43649), .O(n4898)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_11_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1905_25_lut (.I0(GND_net), 
            .I1(n2811), .I2(VCC_net), .I3(n44299), .O(n2878)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1905_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_13 (.CI(n44676), 
            .I0(GND_net), .I1(n22_adj_5631), .CO(n44677));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1034_14_lut (.I0(GND_net), 
            .I1(n1522), .I2(VCC_net), .I3(n44041), .O(n1589)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1034_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_21_add_3_11 (.CI(n43649), .I0(GND_net), .I1(n16), 
            .CO(n43650));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1034_14 (.CI(n44041), 
            .I0(n1522), .I1(VCC_net), .CO(n44042));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1905_25 (.CI(n44299), 
            .I0(n2811), .I1(VCC_net), .CO(n44300));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_12_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n23_adj_5632), .I3(n44675), .O(n23_adj_5476)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1905_24_lut (.I0(GND_net), 
            .I1(n2812), .I2(VCC_net), .I3(n44298), .O(n2879)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1905_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1905_24 (.CI(n44298), 
            .I0(n2812), .I1(VCC_net), .CO(n44299));
    SB_LUT4 unary_minus_21_add_3_10_lut (.I0(n4748), .I1(GND_net), .I2(n17), 
            .I3(n43648), .O(n4899)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_10_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1905_23_lut (.I0(GND_net), 
            .I1(n2813), .I2(VCC_net), .I3(n44297), .O(n2880)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1905_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1905_23 (.CI(n44297), 
            .I0(n2813), .I1(VCC_net), .CO(n44298));
    SB_CARRY unary_minus_21_add_3_10 (.CI(n43648), .I0(GND_net), .I1(n17), 
            .CO(n43649));
    SB_LUT4 unary_minus_21_add_3_9_lut (.I0(n4748), .I1(GND_net), .I2(n18), 
            .I3(n43647), .O(n4900)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_9_lut.LUT_INIT = 16'h8228;
    SB_LUT4 LessThan_17_i8_3_lut_3_lut (.I0(current_limit[4]), .I1(current_limit[8]), 
            .I2(current[8]), .I3(GND_net), .O(n8_adj_5585));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam LessThan_17_i8_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_CARRY unary_minus_21_add_3_9 (.CI(n43647), .I0(GND_net), .I1(n18), 
            .CO(n43648));
    SB_CARRY add_263_16 (.CI(n43548), .I0(encoder1_position[17]), .I1(GND_net), 
            .CO(n43549));
    SB_LUT4 unary_minus_21_add_3_8_lut (.I0(n4748), .I1(GND_net), .I2(n19), 
            .I3(n43646), .O(n4901)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_8_lut.LUT_INIT = 16'h8228;
    SB_LUT4 add_1039_25_lut (.I0(GND_net), .I1(n4883), .I2(n4906), .I3(n43794), 
            .O(n418)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1039_25_lut.LUT_INIT = 16'hC33C;
    SB_DFF commutation_state_i1 (.Q(commutation_state[1]), .C(clk16MHz), 
           .D(n48778));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    SB_CARRY unary_minus_21_add_3_8 (.CI(n43646), .I0(GND_net), .I1(n19), 
            .CO(n43647));
    SB_LUT4 add_263_15_lut (.I0(GND_net), .I1(encoder1_position[16]), .I2(GND_net), 
            .I3(n43547), .O(encoder1_position_scaled_23__N_75[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_263_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_21_add_3_7_lut (.I0(n4748), .I1(GND_net), .I2(n20), 
            .I3(n43645), .O(n4902)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_7_lut.LUT_INIT = 16'h8228;
    SB_LUT4 add_1039_24_lut (.I0(GND_net), .I1(n4883), .I2(n4907), .I3(n43793), 
            .O(n419)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1039_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_12 (.CI(n44675), 
            .I0(GND_net), .I1(n23_adj_5632), .CO(n44676));
    SB_CARRY add_263_15 (.CI(n43547), .I0(encoder1_position[16]), .I1(GND_net), 
            .CO(n43548));
    SB_CARRY add_1039_24 (.CI(n43793), .I0(n4883), .I1(n4907), .CO(n43794));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1905_22_lut (.I0(GND_net), 
            .I1(n2814), .I2(VCC_net), .I3(n44296), .O(n2881)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1905_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1905_22 (.CI(n44296), 
            .I0(n2814), .I1(VCC_net), .CO(n44297));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1905_21_lut (.I0(GND_net), 
            .I1(n2815), .I2(VCC_net), .I3(n44295), .O(n2882)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1905_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_11_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n24_adj_5633), .I3(n44674), .O(n24_adj_5475)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_11 (.CI(n44674), 
            .I0(GND_net), .I1(n24_adj_5633), .CO(n44675));
    SB_LUT4 add_1039_23_lut (.I0(GND_net), .I1(n4883), .I2(n4908), .I3(n43792), 
            .O(n420)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1039_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_21_add_3_7 (.CI(n43645), .I0(GND_net), .I1(n20), 
            .CO(n43646));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1177_3_lut (.I0(n1726), 
            .I1(n1793), .I2(n1752), .I3(GND_net), .O(n1825));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1177_3_lut.LUT_INIT = 16'hacac;
    SB_DFF commutation_state_i2 (.Q(commutation_state[2]), .C(clk16MHz), 
           .D(n49779));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    SB_DFF ID_i0_i1 (.Q(ID[1]), .C(clk16MHz), .D(n29821));   // verilog/TinyFPGA_B.v(368[10] 396[6])
    SB_DFF ID_i0_i2 (.Q(ID[2]), .C(clk16MHz), .D(n29820));   // verilog/TinyFPGA_B.v(368[10] 396[6])
    SB_DFF ID_i0_i3 (.Q(ID[3]), .C(clk16MHz), .D(n29819));   // verilog/TinyFPGA_B.v(368[10] 396[6])
    SB_DFF ID_i0_i4 (.Q(ID[4]), .C(clk16MHz), .D(n29818));   // verilog/TinyFPGA_B.v(368[10] 396[6])
    SB_DFF ID_i0_i5 (.Q(ID[5]), .C(clk16MHz), .D(n29817));   // verilog/TinyFPGA_B.v(368[10] 396[6])
    SB_DFF ID_i0_i6 (.Q(ID[6]), .C(clk16MHz), .D(n29816));   // verilog/TinyFPGA_B.v(368[10] 396[6])
    SB_DFF ID_i0_i7 (.Q(ID[7]), .C(clk16MHz), .D(n29815));   // verilog/TinyFPGA_B.v(368[10] 396[6])
    SB_LUT4 LessThan_17_i15_2_lut (.I0(current[7]), .I1(current_limit[7]), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_5562));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam LessThan_17_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i40784_1_lut_4_lut (.I0(current[15]), .I1(duty[23]), .I2(n51078), 
            .I3(n51081), .O(n56614));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i40784_1_lut_4_lut.LUT_INIT = 16'h4c5d;
    SB_LUT4 i22674_2_lut (.I0(duty[6]), .I1(n296), .I2(GND_net), .I3(GND_net), 
            .O(n4923));   // verilog/TinyFPGA_B.v(123[17] 125[11])
    defparam i22674_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1034_13_lut (.I0(GND_net), 
            .I1(n1523), .I2(VCC_net), .I3(n44040), .O(n1590)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1034_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1905_21 (.CI(n44295), 
            .I0(n2815), .I1(VCC_net), .CO(n44296));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_10_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n25_adj_5634), .I3(n44673), .O(n25_adj_5474)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1034_13 (.CI(n44040), 
            .I0(n1523), .I1(VCC_net), .CO(n44041));
    SB_CARRY add_1039_23 (.CI(n43792), .I0(n4883), .I1(n4908), .CO(n43793));
    SB_LUT4 i22673_2_lut (.I0(duty[7]), .I1(n296), .I2(GND_net), .I3(GND_net), 
            .O(n4922));   // verilog/TinyFPGA_B.v(123[17] 125[11])
    defparam i22673_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 add_1039_22_lut (.I0(GND_net), .I1(n4884), .I2(n4909), .I3(n43791), 
            .O(n421)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1039_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_281_i9_4_lut (.I0(encoder1_position_scaled[8]), .I1(displacement[8]), 
            .I2(n15), .I3(n15_adj_5471), .O(motor_state_23__N_123[8]));   // verilog/TinyFPGA_B.v(284[5] 286[10])
    defparam mux_281_i9_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 unary_minus_21_add_3_6_lut (.I0(n4748), .I1(GND_net), .I2(n21), 
            .I3(n43644), .O(n4903)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_6_lut.LUT_INIT = 16'h8228;
    SB_CARRY encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_10 (.CI(n44673), 
            .I0(GND_net), .I1(n25_adj_5634), .CO(n44674));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_9_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n26_adj_5635), .I3(n44672), .O(n26)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1905_20_lut (.I0(GND_net), 
            .I1(n2816), .I2(VCC_net), .I3(n44294), .O(n2883)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1905_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1034_12_lut (.I0(GND_net), 
            .I1(n1524), .I2(VCC_net), .I3(n44039), .O(n1591)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1034_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1034_12 (.CI(n44039), 
            .I0(n1524), .I1(VCC_net), .CO(n44040));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1905_20 (.CI(n44294), 
            .I0(n2816), .I1(VCC_net), .CO(n44295));
    SB_CARRY unary_minus_21_add_3_6 (.CI(n43644), .I0(GND_net), .I1(n21), 
            .CO(n43645));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1034_11_lut (.I0(GND_net), 
            .I1(n1525), .I2(VCC_net), .I3(n44038), .O(n1592)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1034_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_4_lut (.I0(current[15]), .I1(duty[23]), .I2(n51078), 
            .I3(n51081), .O(n209));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i1_4_lut_4_lut.LUT_INIT = 16'hb3a2;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1034_11 (.CI(n44038), 
            .I0(n1525), .I1(VCC_net), .CO(n44039));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1034_10_lut (.I0(GND_net), 
            .I1(n1526), .I2(VCC_net), .I3(n44037), .O(n1593)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1034_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 n10829_bdd_4_lut_40816 (.I0(n10829), .I1(n439), .I2(current[2]), 
            .I3(duty[23]), .O(n56628));
    defparam n10829_bdd_4_lut_40816.LUT_INIT = 16'he4aa;
    SB_LUT4 unary_minus_21_add_3_5_lut (.I0(n296), .I1(GND_net), .I2(n22), 
            .I3(n43643), .O(n4904)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_5_lut.LUT_INIT = 16'hebbe;
    SB_CARRY add_1039_22 (.CI(n43791), .I0(n4884), .I1(n4909), .CO(n43792));
    SB_CARRY encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_9 (.CI(n44672), 
            .I0(GND_net), .I1(n26_adj_5635), .CO(n44673));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1034_10 (.CI(n44037), 
            .I0(n1526), .I1(VCC_net), .CO(n44038));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1905_19_lut (.I0(GND_net), 
            .I1(n2817), .I2(VCC_net), .I3(n44293), .O(n2884)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1905_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder1_position_scaled_23__I_4_4_lut (.I0(encoder1_position[0]), 
            .I1(encoder1_position[31]), .I2(encoder1_position[1]), .I3(encoder1_position[2]), 
            .O(encoder1_position_scaled_23__N_359));   // verilog/TinyFPGA_B.v(323[33:52])
    defparam encoder1_position_scaled_23__I_4_4_lut.LUT_INIT = 16'hccc8;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_8_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n27_adj_5636), .I3(n44671), .O(n27)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_1039_21_lut (.I0(GND_net), .I1(n4885), .I2(n4910), .I3(n43790), 
            .O(n422)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1039_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1905_19 (.CI(n44293), 
            .I0(n2817), .I1(VCC_net), .CO(n44294));
    SB_CARRY unary_minus_21_add_3_5 (.CI(n43643), .I0(GND_net), .I1(n22), 
            .CO(n43644));
    SB_CARRY add_263_7 (.CI(n43539), .I0(encoder1_position[8]), .I1(GND_net), 
            .CO(n43540));
    SB_LUT4 add_263_6_lut (.I0(GND_net), .I1(encoder1_position[7]), .I2(GND_net), 
            .I3(n43538), .O(encoder1_position_scaled_23__N_75[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_263_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1905_18_lut (.I0(GND_net), 
            .I1(n2818), .I2(VCC_net), .I3(n44292), .O(n2885)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1905_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_8 (.CI(n44671), 
            .I0(GND_net), .I1(n27_adj_5636), .CO(n44672));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1905_18 (.CI(n44292), 
            .I0(n2818), .I1(VCC_net), .CO(n44293));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_7_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n28_adj_5637), .I3(n44670), .O(n28)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_7 (.CI(n44670), 
            .I0(GND_net), .I1(n28_adj_5637), .CO(n44671));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1034_9_lut (.I0(GND_net), 
            .I1(n1527), .I2(VCC_net), .I3(n44036), .O(n1594)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1034_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i40492_1_lut (.I0(n1851), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n56323));
    defparam i40492_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1034_9 (.CI(n44036), 
            .I0(n1527), .I1(VCC_net), .CO(n44037));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1034_8_lut (.I0(GND_net), 
            .I1(n1528), .I2(VCC_net), .I3(n44035), .O(n1595)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1034_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1039_21 (.CI(n43790), .I0(n4885), .I1(n4910), .CO(n43791));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_6_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n29_adj_5638), .I3(n44669), .O(n29)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1905_17_lut (.I0(GND_net), 
            .I1(n2819), .I2(VCC_net), .I3(n44291), .O(n2886)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1905_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1905_17 (.CI(n44291), 
            .I0(n2819), .I1(VCC_net), .CO(n44292));
    SB_LUT4 unary_minus_21_add_3_4_lut (.I0(n379), .I1(GND_net), .I2(n23), 
            .I3(n43642), .O(n4_adj_5444)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_4_lut.LUT_INIT = 16'hebbe;
    SB_CARRY encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_6 (.CI(n44669), 
            .I0(GND_net), .I1(n29_adj_5638), .CO(n44670));
    SB_CARRY unary_minus_21_add_3_4 (.CI(n43642), .I0(GND_net), .I1(n23), 
            .CO(n43643));
    SB_DFF \ID_READOUT_FSM.state__i1  (.Q(\ID_READOUT_FSM.state [1]), .C(clk16MHz), 
           .D(n48068));   // verilog/TinyFPGA_B.v(368[10] 396[6])
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1905_16_lut (.I0(GND_net), 
            .I1(n2820), .I2(VCC_net), .I3(n44290), .O(n2887)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1905_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_5_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n30_adj_5639), .I3(n44668), .O(n30)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_5 (.CI(n44668), 
            .I0(GND_net), .I1(n30_adj_5639), .CO(n44669));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1034_8 (.CI(n44035), 
            .I0(n1528), .I1(VCC_net), .CO(n44036));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_4_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n31_adj_5640), .I3(n44667), .O(n31)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1905_16 (.CI(n44290), 
            .I0(n2820), .I1(VCC_net), .CO(n44291));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1905_15_lut (.I0(GND_net), 
            .I1(n2821), .I2(VCC_net), .I3(n44289), .O(n2888)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1905_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1034_7_lut (.I0(GND_net), 
            .I1(n1529), .I2(GND_net), .I3(n44034), .O(n1596)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1034_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1034_7 (.CI(n44034), 
            .I0(n1529), .I1(GND_net), .CO(n44035));
    SB_CARRY encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_4 (.CI(n44667), 
            .I0(GND_net), .I1(n31_adj_5640), .CO(n44668));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1905_15 (.CI(n44289), 
            .I0(n2821), .I1(VCC_net), .CO(n44290));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1905_14_lut (.I0(GND_net), 
            .I1(n2822), .I2(VCC_net), .I3(n44288), .O(n2889)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1905_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1905_14 (.CI(n44288), 
            .I0(n2822), .I1(VCC_net), .CO(n44289));
    SB_LUT4 add_1039_20_lut (.I0(GND_net), .I1(n4886), .I2(n4911), .I3(n43789), 
            .O(n423)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1039_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_3_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n32_adj_5641), .I3(n44666), .O(n32)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1034_6_lut (.I0(GND_net), 
            .I1(n1530), .I2(GND_net), .I3(n44033), .O(n1597)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1034_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1905_13_lut (.I0(GND_net), 
            .I1(n2823), .I2(VCC_net), .I3(n44287), .O(n2890)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1905_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1034_6 (.CI(n44033), 
            .I0(n1530), .I1(GND_net), .CO(n44034));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_mux_3_i7_3_lut (.I0(encoder0_position_scaled_23__N_327[6]), 
            .I1(n27), .I2(encoder0_position_scaled_23__N_327[31]), .I3(GND_net), 
            .O(n538));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_mux_3_i7_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_17_i19_2_lut (.I0(current[9]), .I1(current_limit[9]), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_5559));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam LessThan_17_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1797_3_lut (.I0(n537), .I1(n2701), 
            .I2(n2643), .I3(GND_net), .O(n2733));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1797_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1034_5_lut (.I0(GND_net), 
            .I1(n1531), .I2(VCC_net), .I3(n44032), .O(n1598)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1034_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1905_13 (.CI(n44287), 
            .I0(n2823), .I1(VCC_net), .CO(n44288));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1905_12_lut (.I0(GND_net), 
            .I1(n2824), .I2(VCC_net), .I3(n44286), .O(n2891)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1905_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1905_12 (.CI(n44286), 
            .I0(n2824), .I1(VCC_net), .CO(n44287));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1034_5 (.CI(n44032), 
            .I0(n1531), .I1(VCC_net), .CO(n44033));
    SB_CARRY encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_3 (.CI(n44666), 
            .I0(GND_net), .I1(n32_adj_5641), .CO(n44667));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1034_4_lut (.I0(GND_net), 
            .I1(n1532_adj_5595), .I2(GND_net), .I3(n44031), .O(n1599)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1034_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_2_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n33_adj_5642), .I3(VCC_net), .O(n33)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_21_add_3_3_lut (.I0(GND_net), .I1(GND_net), .I2(n24), 
            .I3(n43641), .O(n379)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1034_4 (.CI(n44031), 
            .I0(n1532_adj_5595), .I1(GND_net), .CO(n44032));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1034_3_lut (.I0(GND_net), 
            .I1(n1533_adj_5596), .I2(VCC_net), .I3(n44030), .O(n1600)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1034_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1034_3 (.CI(n44030), 
            .I0(n1533_adj_5596), .I1(VCC_net), .CO(n44031));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1905_11_lut (.I0(GND_net), 
            .I1(n2825), .I2(VCC_net), .I3(n44285), .O(n2892)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1905_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1034_2_lut (.I0(GND_net), 
            .I1(n415), .I2(GND_net), .I3(VCC_net), .O(n1601)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1034_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1039_20 (.CI(n43789), .I0(n4886), .I1(n4911), .CO(n43790));
    SB_LUT4 add_263_14_lut (.I0(GND_net), .I1(encoder1_position[15]), .I2(GND_net), 
            .I3(n43546), .O(encoder1_position_scaled_23__N_75[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_263_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_2 (.CI(VCC_net), 
            .I0(GND_net), .I1(n33_adj_5642), .CO(n44666));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1905_11 (.CI(n44285), 
            .I0(n2825), .I1(VCC_net), .CO(n44286));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1034_2 (.CI(VCC_net), 
            .I0(n415), .I1(GND_net), .CO(n44030));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1905_10_lut (.I0(GND_net), 
            .I1(n2826), .I2(VCC_net), .I3(n44284), .O(n2893)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1905_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1905_10 (.CI(n44284), 
            .I0(n2826), .I1(VCC_net), .CO(n44285));
    SB_LUT4 i38792_2_lut_4_lut (.I0(duty[8]), .I1(n338), .I2(duty[4]), 
            .I3(n342), .O(n54622));
    defparam i38792_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 LessThan_11_i6_3_lut_3_lut (.I0(duty[2]), .I1(duty[3]), .I2(current[3]), 
            .I3(GND_net), .O(n6_adj_5580));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i6_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 mux_281_i10_4_lut (.I0(encoder1_position_scaled[9]), .I1(displacement[9]), 
            .I2(n15), .I3(n15_adj_5471), .O(motor_state_23__N_123[9]));   // verilog/TinyFPGA_B.v(284[5] 286[10])
    defparam mux_281_i10_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i39157_2_lut_4_lut (.I0(current[8]), .I1(duty[8]), .I2(current[4]), 
            .I3(duty[4]), .O(n54987));
    defparam i39157_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1905_9_lut (.I0(GND_net), 
            .I1(n2827), .I2(VCC_net), .I3(n44283), .O(n2894)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1905_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1905_9 (.CI(n44283), 
            .I0(n2827), .I1(VCC_net), .CO(n44284));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_967_14_lut (.I0(n56399), 
            .I1(n1422), .I2(VCC_net), .I3(n44029), .O(n1521)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_967_14_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1905_8_lut (.I0(GND_net), 
            .I1(n2828), .I2(VCC_net), .I3(n44282), .O(n2895)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1905_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_21_add_3_3 (.CI(n43641), .I0(GND_net), .I1(n24), 
            .CO(n43642));
    SB_CARRY add_263_6 (.CI(n43538), .I0(encoder1_position[7]), .I1(GND_net), 
            .CO(n43539));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1796_3_lut (.I0(n2633), 
            .I1(n2700), .I2(n2643), .I3(GND_net), .O(n2732));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1796_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_1039_19_lut (.I0(GND_net), .I1(n4887), .I2(n4912), .I3(n43788), 
            .O(n424)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1039_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_11_i8_3_lut_3_lut (.I0(duty[4]), .I1(duty[8]), .I2(current[8]), 
            .I3(GND_net), .O(n8_adj_5578));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i8_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1905_8 (.CI(n44282), 
            .I0(n2828), .I1(VCC_net), .CO(n44283));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_967_13_lut (.I0(GND_net), 
            .I1(n1423), .I2(VCC_net), .I3(n44028), .O(n1490)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_967_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1905_7_lut (.I0(GND_net), 
            .I1(n2829), .I2(GND_net), .I3(n44281), .O(n2896)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1905_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_21_add_3_2_lut (.I0(n4_adj_5444), .I1(GND_net), 
            .I2(n25), .I3(VCC_net), .O(n54531)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_2_lut.LUT_INIT = 16'hebbe;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1905_7 (.CI(n44281), 
            .I0(n2829), .I1(GND_net), .CO(n44282));
    SB_CARRY add_263_14 (.CI(n43546), .I0(encoder1_position[15]), .I1(GND_net), 
            .CO(n43547));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_967_13 (.CI(n44028), 
            .I0(n1423), .I1(VCC_net), .CO(n44029));
    SB_CARRY unary_minus_21_add_3_2 (.CI(VCC_net), .I0(GND_net), .I1(n25), 
            .CO(n43641));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1905_6_lut (.I0(GND_net), 
            .I1(n2830), .I2(GND_net), .I3(n44280), .O(n2897)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1905_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_967_12_lut (.I0(GND_net), 
            .I1(n1424), .I2(VCC_net), .I3(n44027), .O(n1491)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_967_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_967_12 (.CI(n44027), 
            .I0(n1424), .I1(VCC_net), .CO(n44028));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_967_11_lut (.I0(GND_net), 
            .I1(n1425), .I2(VCC_net), .I3(n44026), .O(n1492)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_967_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1905_6 (.CI(n44280), 
            .I0(n2830), .I1(GND_net), .CO(n44281));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1905_5_lut (.I0(GND_net), 
            .I1(n2831), .I2(VCC_net), .I3(n44279), .O(n2898)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1905_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1905_5 (.CI(n44279), 
            .I0(n2831), .I1(VCC_net), .CO(n44280));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_967_11 (.CI(n44026), 
            .I0(n1425), .I1(VCC_net), .CO(n44027));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1905_4_lut (.I0(GND_net), 
            .I1(n2832), .I2(GND_net), .I3(n44278), .O(n2899)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1905_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1905_4 (.CI(n44278), 
            .I0(n2832), .I1(GND_net), .CO(n44279));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_967_10_lut (.I0(GND_net), 
            .I1(n1426), .I2(VCC_net), .I3(n44025), .O(n1493)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_967_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_967_10 (.CI(n44025), 
            .I0(n1426), .I1(VCC_net), .CO(n44026));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1905_3_lut (.I0(GND_net), 
            .I1(n2833), .I2(VCC_net), .I3(n44277), .O(n2900)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1905_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1905_3 (.CI(n44277), 
            .I0(n2833), .I1(VCC_net), .CO(n44278));
    \quadrature_decoder(1)_U0  quad_counter0 (.n2269(clk16MHz), .b_prev(b_prev), 
            .GND_net(GND_net), .a_new({a_new[1], Open_0}), .position_31__N_4108(position_31__N_4108), 
            .ENCODER0_B_N_keep(ENCODER0_B_N), .ENCODER0_A_N_keep(ENCODER0_A_N), 
            .encoder0_position({encoder0_position}), .n29501(n29501), .n2233(n2233), 
            .VCC_net(VCC_net)) /* synthesis lattice_noprune=1 */ ;   // verilog/TinyFPGA_B.v(302[49] 308[6])
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1905_2_lut (.I0(GND_net), 
            .I1(n539), .I2(GND_net), .I3(VCC_net), .O(n2901)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1905_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_967_9_lut (.I0(GND_net), 
            .I1(n1427), .I2(VCC_net), .I3(n44024), .O(n1494)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_967_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1905_2 (.CI(VCC_net), 
            .I0(n539), .I1(GND_net), .CO(n44277));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_967_9 (.CI(n44024), 
            .I0(n1427), .I1(VCC_net), .CO(n44025));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1838_27_lut (.I0(GND_net), 
            .I1(n2709), .I2(VCC_net), .I3(n44276), .O(n2776)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1838_27_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1838_26_lut (.I0(GND_net), 
            .I1(n2710), .I2(VCC_net), .I3(n44275), .O(n2777)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1838_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_967_8_lut (.I0(GND_net), 
            .I1(n1428), .I2(VCC_net), .I3(n44023), .O(n1495)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_967_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1795_3_lut (.I0(n2632), 
            .I1(n2699), .I2(n2643), .I3(GND_net), .O(n2731));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1795_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_967_8 (.CI(n44023), 
            .I0(n1428), .I1(VCC_net), .CO(n44024));
    SB_CARRY add_1039_19 (.CI(n43788), .I0(n4887), .I1(n4912), .CO(n43789));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1838_26 (.CI(n44275), 
            .I0(n2710), .I1(VCC_net), .CO(n44276));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1838_25_lut (.I0(GND_net), 
            .I1(n2711), .I2(VCC_net), .I3(n44274), .O(n2778)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1838_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_1039_18_lut (.I0(GND_net), .I1(n4888), .I2(n4913), .I3(n43787), 
            .O(n425)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1039_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_967_7_lut (.I0(GND_net), 
            .I1(n1429), .I2(GND_net), .I3(n44022), .O(n1496)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_967_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_175_33_lut (.I0(GND_net), .I1(delay_counter[31]), .I2(GND_net), 
            .I3(n43640), .O(n1532)) /* synthesis syn_instantiated=1 */ ;
    defparam add_175_33_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_967_7 (.CI(n44022), 
            .I0(n1429), .I1(GND_net), .CO(n44023));
    SB_DFF pwm_setpoint_i0 (.Q(pwm_setpoint[0]), .C(clk16MHz), .D(pwm_setpoint_23__N_11[0]));   // verilog/TinyFPGA_B.v(103[9] 129[5])
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_967_6_lut (.I0(GND_net), 
            .I1(n1430), .I2(GND_net), .I3(n44021), .O(n1497)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_967_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_281_i11_4_lut (.I0(encoder1_position_scaled[10]), .I1(displacement[10]), 
            .I2(n15), .I3(n15_adj_5471), .O(motor_state_23__N_123[10]));   // verilog/TinyFPGA_B.v(284[5] 286[10])
    defparam mux_281_i11_4_lut.LUT_INIT = 16'h0aca;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1838_25 (.CI(n44274), 
            .I0(n2711), .I1(VCC_net), .CO(n44275));
    SB_CARRY add_1039_18 (.CI(n43787), .I0(n4888), .I1(n4913), .CO(n43788));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_967_6 (.CI(n44021), 
            .I0(n1430), .I1(GND_net), .CO(n44022));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_967_5_lut (.I0(GND_net), 
            .I1(n1431), .I2(VCC_net), .I3(n44020), .O(n1498)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_967_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_175_32_lut (.I0(GND_net), .I1(delay_counter[30]), .I2(GND_net), 
            .I3(n43639), .O(n1533)) /* synthesis syn_instantiated=1 */ ;
    defparam add_175_32_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_175_32 (.CI(n43639), .I0(delay_counter[30]), .I1(GND_net), 
            .CO(n43640));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1838_24_lut (.I0(GND_net), 
            .I1(n2712), .I2(VCC_net), .I3(n44273), .O(n2779)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1838_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_175_31_lut (.I0(GND_net), .I1(delay_counter[29]), .I2(GND_net), 
            .I3(n43638), .O(n1534)) /* synthesis syn_instantiated=1 */ ;
    defparam add_175_31_lut.LUT_INIT = 16'hC33C;
    SB_DFF ID_i0_i0 (.Q(ID[0]), .C(clk16MHz), .D(n29352));   // verilog/TinyFPGA_B.v(368[10] 396[6])
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1838_24 (.CI(n44273), 
            .I0(n2712), .I1(VCC_net), .CO(n44274));
    SB_LUT4 i22672_2_lut (.I0(duty[8]), .I1(n296), .I2(GND_net), .I3(GND_net), 
            .O(n4921));   // verilog/TinyFPGA_B.v(123[17] 125[11])
    defparam i22672_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 mux_281_i12_4_lut (.I0(encoder1_position_scaled[11]), .I1(displacement[11]), 
            .I2(n15), .I3(n15_adj_5471), .O(motor_state_23__N_123[11]));   // verilog/TinyFPGA_B.v(284[5] 286[10])
    defparam mux_281_i12_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1794_3_lut (.I0(n2631), 
            .I1(n2698), .I2(n2643), .I3(GND_net), .O(n2730));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1794_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1793_3_lut (.I0(n2630), 
            .I1(n2697), .I2(n2643), .I3(GND_net), .O(n2729));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1793_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1241_3_lut (.I0(n1822), 
            .I1(n1889), .I2(n1851), .I3(GND_net), .O(n1921));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1241_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_281_i13_4_lut (.I0(encoder1_position_scaled[12]), .I1(displacement[12]), 
            .I2(n15), .I3(n15_adj_5471), .O(motor_state_23__N_123[12]));   // verilog/TinyFPGA_B.v(284[5] 286[10])
    defparam mux_281_i13_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1792_3_lut (.I0(n2629), 
            .I1(n2696), .I2(n2643), .I3(GND_net), .O(n2728));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1792_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1791_3_lut (.I0(n2628), 
            .I1(n2695), .I2(n2643), .I3(GND_net), .O(n2727));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1791_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1790_3_lut (.I0(n2627), 
            .I1(n2694), .I2(n2643), .I3(GND_net), .O(n2726));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1790_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i22671_2_lut (.I0(duty[9]), .I1(n296), .I2(GND_net), .I3(GND_net), 
            .O(n4920));   // verilog/TinyFPGA_B.v(123[17] 125[11])
    defparam i22671_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 mux_281_i14_4_lut (.I0(encoder1_position_scaled[13]), .I1(displacement[13]), 
            .I2(n15), .I3(n15_adj_5471), .O(motor_state_23__N_123[13]));   // verilog/TinyFPGA_B.v(284[5] 286[10])
    defparam mux_281_i14_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1789_3_lut (.I0(n2626), 
            .I1(n2693), .I2(n2643), .I3(GND_net), .O(n2725));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1789_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1788_3_lut (.I0(n2625), 
            .I1(n2692), .I2(n2643), .I3(GND_net), .O(n2724));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1788_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i22670_2_lut (.I0(duty[10]), .I1(n296), .I2(GND_net), .I3(GND_net), 
            .O(n4919));   // verilog/TinyFPGA_B.v(123[17] 125[11])
    defparam i22670_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1787_3_lut (.I0(n2624), 
            .I1(n2691), .I2(n2643), .I3(GND_net), .O(n2723));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1787_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15273_3_lut (.I0(\data_out_frame[11] [6]), .I1(encoder1_position_scaled[6]), 
            .I2(n24210), .I3(GND_net), .O(n29353));   // verilog/coms.v(128[12] 303[6])
    defparam i15273_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_281_i15_4_lut (.I0(encoder1_position_scaled[14]), .I1(displacement[14]), 
            .I2(n15), .I3(n15_adj_5471), .O(motor_state_23__N_123[14]));   // verilog/TinyFPGA_B.v(284[5] 286[10])
    defparam mux_281_i15_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1786_3_lut (.I0(n2623), 
            .I1(n2690), .I2(n2643), .I3(GND_net), .O(n2722));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1786_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_281_i16_4_lut (.I0(encoder1_position_scaled[15]), .I1(displacement[15]), 
            .I2(n15), .I3(n15_adj_5471), .O(motor_state_23__N_123[15]));   // verilog/TinyFPGA_B.v(284[5] 286[10])
    defparam mux_281_i16_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1785_3_lut (.I0(n2622), 
            .I1(n2689), .I2(n2643), .I3(GND_net), .O(n2721));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1785_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1784_3_lut (.I0(n2621), 
            .I1(n2688), .I2(n2643), .I3(GND_net), .O(n2720));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1784_3_lut.LUT_INIT = 16'hacac;
    pll32MHz pll32MHz_inst (.GND_net(GND_net), .clk16MHz(clk16MHz), .VCC_net(VCC_net), 
            .clk32MHz(clk32MHz)) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(34[10] 38[2])
    SB_LUT4 LessThan_11_i15_2_lut (.I0(current[7]), .I1(duty[7]), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_5567));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_11_i13_2_lut (.I0(current[6]), .I1(duty[6]), .I2(GND_net), 
            .I3(GND_net), .O(n13_adj_5568));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i14_4_lut (.I0(duty[0]), .I1(duty[23]), .I2(duty[1]), .I3(duty[2]), 
            .O(n211));   // verilog/TinyFPGA_B.v(111[25:31])
    defparam i14_4_lut.LUT_INIT = 16'hccc8;
    SB_LUT4 LessThan_11_i19_2_lut (.I0(current[9]), .I1(duty[9]), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_5564));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_11_i17_2_lut (.I0(current[8]), .I1(duty[8]), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_5565));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mux_281_i17_4_lut (.I0(encoder1_position_scaled[16]), .I1(displacement[16]), 
            .I2(n15), .I3(n15_adj_5471), .O(motor_state_23__N_123[16]));   // verilog/TinyFPGA_B.v(284[5] 286[10])
    defparam mux_281_i17_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_281_i18_4_lut (.I0(encoder1_position_scaled[17]), .I1(displacement[17]), 
            .I2(n15), .I3(n15_adj_5471), .O(motor_state_23__N_123[17]));   // verilog/TinyFPGA_B.v(284[5] 286[10])
    defparam mux_281_i18_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 LessThan_11_i7_2_lut (.I0(current[3]), .I1(duty[3]), .I2(GND_net), 
            .I3(GND_net), .O(n7_adj_5579));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i7_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i5577_3_lut_4_lut_4_lut (.I0(commutation_state[2]), .I1(commutation_state[1]), 
            .I2(dir), .I3(commutation_state[0]), .O(GHA_N_478));   // verilog/TinyFPGA_B.v(179[7] 198[15])
    defparam i5577_3_lut_4_lut_4_lut.LUT_INIT = 16'h12c2;
    SB_LUT4 LessThan_11_i9_2_lut (.I0(current[4]), .I1(duty[4]), .I2(GND_net), 
            .I3(GND_net), .O(n9_adj_5570));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_11_i11_2_lut (.I0(current[5]), .I1(duty[5]), .I2(GND_net), 
            .I3(GND_net), .O(n11_adj_5569));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i5579_3_lut_4_lut_4_lut (.I0(commutation_state[2]), .I1(commutation_state[1]), 
            .I2(dir), .I3(commutation_state[0]), .O(GLA_N_495));   // verilog/TinyFPGA_B.v(179[7] 198[15])
    defparam i5579_3_lut_4_lut_4_lut.LUT_INIT = 16'h212c;
    SB_LUT4 LessThan_11_i5_2_lut (.I0(current[2]), .I1(duty[2]), .I2(GND_net), 
            .I3(GND_net), .O(n5_adj_5581));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i5_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i39165_4_lut (.I0(n11_adj_5569), .I1(n9_adj_5570), .I2(n7_adj_5579), 
            .I3(n5_adj_5581), .O(n54995));
    defparam i39165_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 LessThan_11_i16_3_lut (.I0(n8_adj_5578), .I1(duty[9]), .I2(n19_adj_5564), 
            .I3(GND_net), .O(n16_adj_5566));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_11_i4_4_lut (.I0(duty[0]), .I1(duty[1]), .I2(current[1]), 
            .I3(current[0]), .O(n4_adj_5590));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i4_4_lut.LUT_INIT = 16'h0c8e;
    SB_LUT4 LessThan_20_i15_2_lut (.I0(duty[7]), .I1(n339), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_5536));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam LessThan_20_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_20_i13_2_lut (.I0(duty[6]), .I1(n340), .I2(GND_net), 
            .I3(GND_net), .O(n13_adj_5537));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam LessThan_20_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mux_281_i19_4_lut (.I0(encoder1_position_scaled[18]), .I1(displacement[18]), 
            .I2(n15), .I3(n15_adj_5471), .O(motor_state_23__N_123[18]));   // verilog/TinyFPGA_B.v(284[5] 286[10])
    defparam mux_281_i19_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 LessThan_20_i19_2_lut (.I0(duty[9]), .I1(n337), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_5533));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam LessThan_20_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i39791_3_lut (.I0(n4_adj_5590), .I1(duty[5]), .I2(n11_adj_5569), 
            .I3(GND_net), .O(n55622));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i39791_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5581_3_lut_4_lut_4_lut (.I0(commutation_state[2]), .I1(commutation_state[1]), 
            .I2(dir), .I3(commutation_state[0]), .O(GHB_N_500));
    defparam i5581_3_lut_4_lut_4_lut.LUT_INIT = 16'hc121;
    SB_LUT4 i39792_3_lut (.I0(n55622), .I1(duty[6]), .I2(n13_adj_5568), 
            .I3(GND_net), .O(n55623));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i39792_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_20_i17_2_lut (.I0(duty[8]), .I1(n338), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_5534));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam LessThan_20_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i5583_3_lut_4_lut_4_lut (.I0(commutation_state[2]), .I1(commutation_state[1]), 
            .I2(dir), .I3(commutation_state[0]), .O(GLB_N_509));
    defparam i5583_3_lut_4_lut_4_lut.LUT_INIT = 16'h1c12;
    SB_LUT4 LessThan_20_i7_2_lut (.I0(duty[3]), .I1(n343), .I2(GND_net), 
            .I3(GND_net), .O(n7_adj_5541));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam LessThan_20_i7_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_20_i9_2_lut (.I0(duty[4]), .I1(n342), .I2(GND_net), 
            .I3(GND_net), .O(n9_adj_5539));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam LessThan_20_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mux_281_i20_4_lut (.I0(encoder1_position_scaled[19]), .I1(displacement[19]), 
            .I2(n15), .I3(n15_adj_5471), .O(motor_state_23__N_123[19]));   // verilog/TinyFPGA_B.v(284[5] 286[10])
    defparam mux_281_i20_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 LessThan_20_i11_2_lut (.I0(duty[5]), .I1(n341), .I2(GND_net), 
            .I3(GND_net), .O(n11_adj_5538));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam LessThan_20_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_20_i5_2_lut (.I0(duty[2]), .I1(n344), .I2(GND_net), 
            .I3(GND_net), .O(n5_adj_5543));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam LessThan_20_i5_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i39159_4_lut (.I0(n17_adj_5565), .I1(n15_adj_5567), .I2(n13_adj_5568), 
            .I3(n54995), .O(n54989));
    defparam i39159_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i39947_4_lut (.I0(n16_adj_5566), .I1(n6_adj_5580), .I2(n19_adj_5564), 
            .I3(n54987), .O(n55778));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i39947_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i38830_4_lut (.I0(n11_adj_5538), .I1(n9_adj_5539), .I2(n7_adj_5541), 
            .I3(n5_adj_5543), .O(n54660));
    defparam i38830_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 LessThan_20_i8_3_lut (.I0(n342), .I1(n338), .I2(n17_adj_5534), 
            .I3(GND_net), .O(n8_adj_5540));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam LessThan_20_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i39310_3_lut (.I0(n55623), .I1(duty[7]), .I2(n15_adj_5567), 
            .I3(GND_net), .O(n55141));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i39310_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_4_lut (.I0(\ID_READOUT_FSM.state [0]), .I1(\ID_READOUT_FSM.state [1]), 
            .I2(n27093), .I3(n1650), .O(n7974));   // verilog/TinyFPGA_B.v(386[7:11])
    defparam i1_2_lut_3_lut_4_lut.LUT_INIT = 16'h0400;
    SB_LUT4 i40031_4_lut (.I0(n55141), .I1(n55778), .I2(n19_adj_5564), 
            .I3(n54989), .O(n55862));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i40031_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i40032_3_lut (.I0(n55862), .I1(duty[10]), .I2(current[10]), 
            .I3(GND_net), .O(n55863));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i40032_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i1_3_lut_3_lut (.I0(\ID_READOUT_FSM.state [0]), .I1(\ID_READOUT_FSM.state [1]), 
            .I2(n27093), .I3(GND_net), .O(n7593));   // verilog/TinyFPGA_B.v(386[7:11])
    defparam i1_3_lut_3_lut.LUT_INIT = 16'h1515;
    SB_LUT4 i22377_2_lut_3_lut_4_lut (.I0(\ID_READOUT_FSM.state [0]), .I1(\ID_READOUT_FSM.state [1]), 
            .I2(n27093), .I3(n1650), .O(n36436));   // verilog/TinyFPGA_B.v(386[7:11])
    defparam i22377_2_lut_3_lut_4_lut.LUT_INIT = 16'hbfbb;
    SB_LUT4 LessThan_20_i6_3_lut (.I0(n344), .I1(n343), .I2(n7_adj_5541), 
            .I3(GND_net), .O(n6_adj_5542));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam LessThan_20_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut (.I0(\ID_READOUT_FSM.state [0]), .I1(\ID_READOUT_FSM.state [1]), 
            .I2(n27093), .I3(GND_net), .O(n27094));   // verilog/TinyFPGA_B.v(386[7:11])
    defparam i1_2_lut_3_lut.LUT_INIT = 16'hfbfb;
    SB_LUT4 LessThan_20_i16_3_lut (.I0(n8_adj_5540), .I1(n337), .I2(n19_adj_5533), 
            .I3(GND_net), .O(n16_adj_5535));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam LessThan_20_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i37269_3_lut (.I0(duty[17]), .I1(duty[19]), .I2(n330), .I3(GND_net), 
            .O(n53032));
    defparam i37269_3_lut.LUT_INIT = 16'h7e7e;
    SB_LUT4 mux_281_i21_4_lut (.I0(encoder1_position_scaled[20]), .I1(displacement[20]), 
            .I2(n15), .I3(n15_adj_5471), .O(motor_state_23__N_123[20]));   // verilog/TinyFPGA_B.v(284[5] 286[10])
    defparam mux_281_i21_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i22711_2_lut_2_lut (.I0(n296), .I1(n356), .I2(GND_net), .I3(GND_net), 
            .O(n4883));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam i22711_2_lut_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i39998_3_lut (.I0(n55863), .I1(duty[11]), .I2(current[11]), 
            .I3(GND_net), .O(n24_adj_5563));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i39998_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i3_4_lut_adj_1869 (.I0(duty[14]), .I1(n24_adj_5563), .I2(duty[12]), 
            .I3(duty[13]), .O(n50822));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i3_4_lut_adj_1869.LUT_INIT = 16'hfffe;
    SB_LUT4 i3_4_lut_adj_1870 (.I0(duty[14]), .I1(n24_adj_5563), .I2(duty[12]), 
            .I3(duty[13]), .O(n50825));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i3_4_lut_adj_1870.LUT_INIT = 16'h8000;
    SB_LUT4 i1_4_lut_adj_1871 (.I0(duty[15]), .I1(current[15]), .I2(n50825), 
            .I3(n50822), .O(n32_adj_5525));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i1_4_lut_adj_1871.LUT_INIT = 16'hb3a2;
    SB_LUT4 i40471_1_lut (.I0(n1950), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n56302));
    defparam i40471_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_281_i22_4_lut (.I0(encoder1_position_scaled[21]), .I1(displacement[21]), 
            .I2(n15), .I3(n15_adj_5471), .O(motor_state_23__N_123[21]));   // verilog/TinyFPGA_B.v(284[5] 286[10])
    defparam mux_281_i22_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i37273_3_lut (.I0(duty[21]), .I1(duty[15]), .I2(n330), .I3(GND_net), 
            .O(n53036));
    defparam i37273_3_lut.LUT_INIT = 16'h7e7e;
    SB_LUT4 i37303_4_lut (.I0(duty[20]), .I1(n53032), .I2(duty[22]), .I3(n330), 
            .O(n53069));
    defparam i37303_4_lut.LUT_INIT = 16'hdffe;
    SB_LUT4 i3_4_lut_adj_1872 (.I0(duty[18]), .I1(n32_adj_5525), .I2(duty[16]), 
            .I3(duty[17]), .O(n50886));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i3_4_lut_adj_1872.LUT_INIT = 16'hfffe;
    SB_LUT4 i3_4_lut_adj_1873 (.I0(duty[18]), .I1(n32_adj_5525), .I2(duty[16]), 
            .I3(duty[17]), .O(n50888));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i3_4_lut_adj_1873.LUT_INIT = 16'h8000;
    SB_LUT4 LessThan_20_i4_3_lut (.I0(n54539), .I1(n345), .I2(duty[1]), 
            .I3(GND_net), .O(n4_adj_5544));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam LessThan_20_i4_3_lut.LUT_INIT = 16'h8e8e;
    motorControl control (.\Kp[14] (Kp[14]), .GND_net(GND_net), .\Kp[0] (Kp[0]), 
            .\Kp[2] (Kp[2]), .\Kp[11] (Kp[11]), .\Kp[12] (Kp[12]), .\Kp[3] (Kp[3]), 
            .\Kp[4] (Kp[4]), .\Kp[5] (Kp[5]), .\Ki[12] (Ki[12]), .\PID_CONTROLLER.integral_23__N_3996 ({\PID_CONTROLLER.integral_23__N_3996 }), 
            .\Kp[13] (Kp[13]), .\Ki[7] (Ki[7]), .\Ki[8] (Ki[8]), .\Kp[6] (Kp[6]), 
            .\Ki[13] (Ki[13]), .\Ki[14] (Ki[14]), .\Ki[9] (Ki[9]), .\Kp[15] (Kp[15]), 
            .\Kp[7] (Kp[7]), .\Kp[8] (Kp[8]), .\Ki[15] (Ki[15]), .control_update(control_update), 
            .duty({duty}), .clk16MHz(clk16MHz), .\Kp[9] (Kp[9]), .\Kp[10] (Kp[10]), 
            .IntegralLimit({IntegralLimit}), .\Ki[1] (Ki[1]), .\Ki[0] (Ki[0]), 
            .\Kp[1] (Kp[1]), .\Ki[2] (Ki[2]), .\Ki[3] (Ki[3]), .\Ki[4] (Ki[4]), 
            .\Ki[5] (Ki[5]), .\Ki[6] (Ki[6]), .\Ki[10] (Ki[10]), .\Ki[11] (Ki[11]), 
            .PWMLimit({PWMLimit}), .n363(n363), .n32464(n32464), .deadband({deadband}), 
            .VCC_net(VCC_net), .\PID_CONTROLLER.integral ({\PID_CONTROLLER.integral }), 
            .n29381(n29381), .setpoint({setpoint}), .motor_state({motor_state}), 
            .n29915(n29915), .n29914(n29914), .n29913(n29913), .n29912(n29912), 
            .n29911(n29911), .n29910(n29910), .n29909(n29909), .n29908(n29908), 
            .n29907(n29907), .n29906(n29906), .n29905(n29905), .n29904(n29904), 
            .n29903(n29903), .n29902(n29902), .n29901(n29901), .n29900(n29900), 
            .n29899(n29899), .n29898(n29898), .n29897(n29897), .n29896(n29896), 
            .n29895(n29895), .n29894(n29894), .n29893(n29893)) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(288[16] 300[4])
    SB_LUT4 i39863_3_lut (.I0(n4_adj_5544), .I1(n341), .I2(n11_adj_5538), 
            .I3(GND_net), .O(n55694));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam i39863_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i39864_3_lut (.I0(n55694), .I1(n340), .I2(n13_adj_5537), .I3(GND_net), 
            .O(n55695));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam i39864_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1874 (.I0(duty[19]), .I1(current[15]), .I2(n50888), 
            .I3(n50886), .O(n40));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i1_4_lut_adj_1874.LUT_INIT = 16'hb3a2;
    SB_LUT4 i15274_3_lut (.I0(\neo_pixel_transmitter.t0 [0]), .I1(timer[0]), 
            .I2(n47790), .I3(GND_net), .O(n29354));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15274_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i38794_4_lut (.I0(n17_adj_5534), .I1(n15_adj_5536), .I2(n13_adj_5537), 
            .I3(n54660), .O(n54624));
    defparam i38794_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i3_4_lut_adj_1875 (.I0(duty[22]), .I1(n40), .I2(duty[20]), 
            .I3(duty[21]), .O(n51081));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i3_4_lut_adj_1875.LUT_INIT = 16'hfffe;
    SB_LUT4 i39975_4_lut (.I0(n16_adj_5535), .I1(n6_adj_5542), .I2(n19_adj_5533), 
            .I3(n54622), .O(n55806));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam i39975_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i39738_3_lut (.I0(n55695), .I1(n339), .I2(n15_adj_5536), .I3(GND_net), 
            .O(n55569));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam i39738_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i40053_4_lut (.I0(n55569), .I1(n55806), .I2(n19_adj_5533), 
            .I3(n54624), .O(n55884));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam i40053_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i40054_3_lut (.I0(n55884), .I1(n336), .I2(duty[10]), .I3(GND_net), 
            .O(n55885));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam i40054_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i40038_3_lut (.I0(n55885), .I1(n335), .I2(duty[11]), .I3(GND_net), 
            .O(n55869));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam i40038_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i39992_3_lut (.I0(n55869), .I1(n334), .I2(duty[12]), .I3(GND_net), 
            .O(n55823));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam i39992_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i7_4_lut_adj_1876 (.I0(duty[18]), .I1(n55823), .I2(n330), 
            .I3(duty[23]), .O(n20_adj_5466));
    defparam i7_4_lut_adj_1876.LUT_INIT = 16'h2100;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i568_3_lut_4_lut (.I0(n861), 
            .I1(encoder0_position_scaled_23__N_327[31]), .I2(n53127), .I3(n49749), 
            .O(n928));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i568_3_lut_4_lut.LUT_INIT = 16'hf4b0;
    SB_LUT4 i11_4_lut (.I0(n330), .I1(n53069), .I2(n53036), .I3(duty[13]), 
            .O(n24_adj_5465));
    defparam i11_4_lut.LUT_INIT = 16'h0200;
    SB_LUT4 i3_4_lut_adj_1877 (.I0(duty[22]), .I1(n40), .I2(duty[20]), 
            .I3(duty[21]), .O(n51078));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i3_4_lut_adj_1877.LUT_INIT = 16'h8000;
    SB_LUT4 i38941_4_lut (.I0(duty[16]), .I1(n20_adj_5466), .I2(duty[14]), 
            .I3(n330), .O(n54594));
    defparam i38941_4_lut.LUT_INIT = 16'h8004;
    SB_LUT4 i14_4_lut_adj_1878 (.I0(n54594), .I1(pwm_setpoint_23__N_263), 
            .I2(n296), .I3(n24_adj_5465), .O(n10829));
    defparam i14_4_lut_adj_1878.LUT_INIT = 16'hcac0;
    SB_LUT4 LessThan_17_i5_2_lut (.I0(current[2]), .I1(current_limit[2]), 
            .I2(GND_net), .I3(GND_net), .O(n5_adj_5588));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam LessThan_17_i5_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i572_3_lut_4_lut (.I0(n861), 
            .I1(encoder0_position_scaled_23__N_327[31]), .I2(n53125), .I3(n49757), 
            .O(n932));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i572_3_lut_4_lut.LUT_INIT = 16'hf4b0;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_mux_3_i28_3_lut (.I0(encoder0_position_scaled_23__N_327[27]), 
            .I1(n6_adj_5493), .I2(encoder0_position_scaled_23__N_327[31]), 
            .I3(GND_net), .O(n625));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_mux_3_i28_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_adj_1879 (.I0(n2_adj_5497), .I1(n3_adj_5496), 
            .I2(encoder0_position_scaled_23__N_327[31]), .I3(GND_net), .O(n51996));
    defparam i1_2_lut_3_lut_adj_1879.LUT_INIT = 16'h8080;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_mux_3_i29_3_lut (.I0(encoder0_position_scaled_23__N_327[28]), 
            .I1(n5_adj_5494), .I2(encoder0_position_scaled_23__N_327[31]), 
            .I3(GND_net), .O(n516));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_mux_3_i29_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34000_2_lut_3_lut (.I0(n2_adj_5497), .I1(n3_adj_5496), .I2(n5_adj_5643), 
            .I3(GND_net), .O(n49748));
    defparam i34000_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i39179_4_lut (.I0(n11_adj_5583), .I1(n9_adj_5584), .I2(n7_adj_5586), 
            .I3(n5_adj_5588), .O(n55009));
    defparam i39179_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_mux_3_i30_3_lut (.I0(encoder0_position_scaled_23__N_327[29]), 
            .I1(n4_adj_5495), .I2(encoder0_position_scaled_23__N_327[31]), 
            .I3(GND_net), .O(n623));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_mux_3_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i22367_2_lut (.I0(pwm_out), .I1(GHC), .I2(GND_net), .I3(GND_net), 
            .O(INHC_c_0));   // verilog/TinyFPGA_B.v(91[16:31])
    defparam i22367_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i22366_2_lut (.I0(pwm_out), .I1(GHB), .I2(GND_net), .I3(GND_net), 
            .O(INHB_c_0));   // verilog/TinyFPGA_B.v(89[16:31])
    defparam i22366_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i22365_2_lut (.I0(pwm_out), .I1(GHA), .I2(GND_net), .I3(GND_net), 
            .O(INHA_c_0));   // verilog/TinyFPGA_B.v(87[16:31])
    defparam i22365_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_mux_3_i31_3_lut (.I0(encoder0_position_scaled_23__N_327[30]), 
            .I1(n3_adj_5496), .I2(encoder0_position_scaled_23__N_327[31]), 
            .I3(GND_net), .O(n622));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_mux_3_i31_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n56628_bdd_4_lut (.I0(n56628), .I1(duty[2]), .I2(n268), .I3(duty[23]), 
            .O(pwm_setpoint_23__N_11[2]));
    defparam n56628_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i12_3_lut_4_lut (.I0(r_SM_Main[1]), .I1(r_SM_Main[2]), .I2(n28753), 
            .I3(rx_data_ready), .O(n48522));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i12_3_lut_4_lut.LUT_INIT = 16'h2f20;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1880 (.I0(r_SM_Main[1]), .I1(r_SM_Main[2]), 
            .I2(r_SM_Main[0]), .I3(r_SM_Main_2__N_3777[2]), .O(n48878));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i1_2_lut_3_lut_4_lut_adj_1880.LUT_INIT = 16'h2000;
    SB_LUT4 i13_3_lut_4_lut_4_lut (.I0(r_SM_Main[1]), .I1(r_SM_Main[2]), 
            .I2(r_SM_Main[0]), .I3(r_SM_Main_2__N_3777[2]), .O(n28753));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i13_3_lut_4_lut_4_lut.LUT_INIT = 16'h2505;
    SB_LUT4 i22657_2_lut_2_lut (.I0(duty[23]), .I1(n296), .I2(GND_net), 
            .I3(GND_net), .O(n4906));   // verilog/TinyFPGA_B.v(123[17] 125[11])
    defparam i22657_2_lut_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1783_3_lut (.I0(n2620), 
            .I1(n2687), .I2(n2643), .I3(GND_net), .O(n2719));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1783_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i22658_2_lut_2_lut (.I0(duty[22]), .I1(n296), .I2(GND_net), 
            .I3(GND_net), .O(n4907));   // verilog/TinyFPGA_B.v(123[17] 125[11])
    defparam i22658_2_lut_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1782_3_lut (.I0(n2619), 
            .I1(n2686), .I2(n2643), .I3(GND_net), .O(n2718));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1782_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 LessThan_17_i16_3_lut (.I0(n8_adj_5585), .I1(current_limit[9]), 
            .I2(n19_adj_5559), .I3(GND_net), .O(n16_adj_5561));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam LessThan_17_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_17_i4_4_lut (.I0(current_limit[0]), .I1(current_limit[1]), 
            .I2(current[1]), .I3(current[0]), .O(n4_adj_5589));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam LessThan_17_i4_4_lut.LUT_INIT = 16'h0c8e;
    SB_LUT4 i40584_1_lut (.I0(n1356), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n56415));
    defparam i40584_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i22669_2_lut (.I0(duty[11]), .I1(n296), .I2(GND_net), .I3(GND_net), 
            .O(n4918));   // verilog/TinyFPGA_B.v(123[17] 125[11])
    defparam i22669_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i39793_3_lut (.I0(n4_adj_5589), .I1(current_limit[5]), .I2(n11_adj_5583), 
            .I3(GND_net), .O(n55624));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam i39793_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1781_3_lut (.I0(n2618), 
            .I1(n2685), .I2(n2643), .I3(GND_net), .O(n2717));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1781_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1780_3_lut (.I0(n2617), 
            .I1(n2684), .I2(n2643), .I3(GND_net), .O(n2716));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1780_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i39794_3_lut (.I0(n55624), .I1(current_limit[6]), .I2(n13_adj_5582), 
            .I3(GND_net), .O(n55625));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam i39794_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i39175_4_lut (.I0(n17_adj_5560), .I1(n15_adj_5562), .I2(n13_adj_5582), 
            .I3(n55009), .O(n55005));
    defparam i39175_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1779_3_lut (.I0(n2616), 
            .I1(n2683), .I2(n2643), .I3(GND_net), .O(n2715));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1779_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15438_3_lut (.I0(Kp[4]), .I1(\data_in_frame[3] [4]), .I2(n50654), 
            .I3(GND_net), .O(n29518));   // verilog/coms.v(128[12] 303[6])
    defparam i15438_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i39951_4_lut (.I0(n16_adj_5561), .I1(n6_adj_5587), .I2(n19_adj_5559), 
            .I3(n55003), .O(n55782));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam i39951_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i39306_3_lut (.I0(n55625), .I1(current_limit[7]), .I2(n15_adj_5562), 
            .I3(GND_net), .O(n55137));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam i39306_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i40033_4_lut (.I0(n55137), .I1(n55782), .I2(n19_adj_5559), 
            .I3(n55005), .O(n55864));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam i40033_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i40034_3_lut (.I0(n55864), .I1(current_limit[10]), .I2(current[10]), 
            .I3(GND_net), .O(n55865));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam i40034_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i39996_3_lut (.I0(n55865), .I1(current_limit[11]), .I2(current[11]), 
            .I3(GND_net), .O(n24_adj_5558));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam i39996_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i22659_2_lut_2_lut (.I0(duty[21]), .I1(n296), .I2(GND_net), 
            .I3(GND_net), .O(n4908));   // verilog/TinyFPGA_B.v(123[17] 125[11])
    defparam i22659_2_lut_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i16_4_lut_4_lut (.I0(state_adj_5736[0]), .I1(n54609), .I2(n7354), 
            .I3(n10), .O(n8_adj_5654));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i16_4_lut_4_lut.LUT_INIT = 16'h3a7a;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1308_3_lut (.I0(n1921), 
            .I1(n1988), .I2(n1950), .I3(GND_net), .O(n2020));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1308_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15749_4_lut_4_lut (.I0(state[0]), .I1(state[1]), .I2(n28778), 
            .I3(state_3__N_639[1]), .O(n29829));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15749_4_lut_4_lut.LUT_INIT = 16'hfc7c;
    SB_LUT4 i1_4_lut_adj_1881 (.I0(current_limit[13]), .I1(n24_adj_5558), 
            .I2(current_limit[14]), .I3(current_limit[12]), .O(n50829));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam i1_4_lut_adj_1881.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1882 (.I0(current_limit[13]), .I1(n24_adj_5558), 
            .I2(current_limit[14]), .I3(current_limit[12]), .O(n50836));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam i1_4_lut_adj_1882.LUT_INIT = 16'h8000;
    SB_LUT4 i1_4_lut_adj_1883 (.I0(current[15]), .I1(current_limit[15]), 
            .I2(n50836), .I3(n50829), .O(n296));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam i1_4_lut_adj_1883.LUT_INIT = 16'hb3a2;
    SB_LUT4 i15843_3_lut (.I0(PWMLimit[18]), .I1(\data_in_frame[8] [2]), 
            .I2(n50654), .I3(GND_net), .O(n29923));   // verilog/coms.v(128[12] 303[6])
    defparam i15843_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i22665_2_lut (.I0(duty[15]), .I1(n296), .I2(GND_net), .I3(GND_net), 
            .O(n4914));   // verilog/TinyFPGA_B.v(123[17] 125[11])
    defparam i22665_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i22668_2_lut (.I0(duty[12]), .I1(n296), .I2(GND_net), .I3(GND_net), 
            .O(n4917));   // verilog/TinyFPGA_B.v(123[17] 125[11])
    defparam i22668_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i22667_2_lut (.I0(duty[13]), .I1(n296), .I2(GND_net), .I3(GND_net), 
            .O(n4916));   // verilog/TinyFPGA_B.v(123[17] 125[11])
    defparam i22667_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i22666_2_lut (.I0(duty[14]), .I1(n296), .I2(GND_net), .I3(GND_net), 
            .O(n4915));   // verilog/TinyFPGA_B.v(123[17] 125[11])
    defparam i22666_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1708_3_lut (.I0(n2513), 
            .I1(n2580), .I2(n2544), .I3(GND_net), .O(n2612));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1708_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1707_3_lut (.I0(n2512), 
            .I1(n2579), .I2(n2544), .I3(GND_net), .O(n2611));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1707_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1710_3_lut (.I0(n2515), 
            .I1(n2582), .I2(n2544), .I3(GND_net), .O(n2614));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1710_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1709_3_lut (.I0(n2514), 
            .I1(n2581), .I2(n2544), .I3(GND_net), .O(n2613));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1709_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1713_3_lut (.I0(n2518), 
            .I1(n2585), .I2(n2544), .I3(GND_net), .O(n2617));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1713_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1712_3_lut (.I0(n2517), 
            .I1(n2584), .I2(n2544), .I3(GND_net), .O(n2616));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1712_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1726_3_lut (.I0(n2531), 
            .I1(n2598), .I2(n2544), .I3(GND_net), .O(n2630));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1726_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1725_3_lut (.I0(n2530), 
            .I1(n2597), .I2(n2544), .I3(GND_net), .O(n2629));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1725_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1719_3_lut (.I0(n2524), 
            .I1(n2591), .I2(n2544), .I3(GND_net), .O(n2623));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1719_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1723_3_lut (.I0(n2528), 
            .I1(n2595), .I2(n2544), .I3(GND_net), .O(n2627));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1723_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1721_3_lut (.I0(n2526), 
            .I1(n2593), .I2(n2544), .I3(GND_net), .O(n2625));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1721_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1715_3_lut (.I0(n2520), 
            .I1(n2587), .I2(n2544), .I3(GND_net), .O(n2619));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1715_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1729_3_lut (.I0(n536), .I1(n2601), 
            .I2(n2544), .I3(GND_net), .O(n2633));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1729_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1728_3_lut (.I0(n2533), 
            .I1(n2600), .I2(n2544), .I3(GND_net), .O(n2632));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1728_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1727_3_lut (.I0(n2532), 
            .I1(n2599), .I2(n2544), .I3(GND_net), .O(n2631));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1727_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_mux_3_i8_3_lut (.I0(encoder0_position_scaled_23__N_327[7]), 
            .I1(n26), .I2(encoder0_position_scaled_23__N_327[31]), .I3(GND_net), 
            .O(n537));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_mux_3_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1722_3_lut (.I0(n2527), 
            .I1(n2594), .I2(n2544), .I3(GND_net), .O(n2626));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1722_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1724_3_lut (.I0(n2529), 
            .I1(n2596), .I2(n2544), .I3(GND_net), .O(n2628));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1724_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1720_3_lut (.I0(n2525), 
            .I1(n2592), .I2(n2544), .I3(GND_net), .O(n2624));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1720_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1716_3_lut (.I0(n2521), 
            .I1(n2588), .I2(n2544), .I3(GND_net), .O(n2620));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1716_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1714_3_lut (.I0(n2519), 
            .I1(n2586), .I2(n2544), .I3(GND_net), .O(n2618));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1714_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1641_3_lut (.I0(n2414), 
            .I1(n2481), .I2(n2445), .I3(GND_net), .O(n2513));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1641_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 n10829_bdd_4_lut_40798 (.I0(n10829), .I1(n440), .I2(current[1]), 
            .I3(duty[23]), .O(n56622));
    defparam n10829_bdd_4_lut_40798.LUT_INIT = 16'he4aa;
    SB_LUT4 n56622_bdd_4_lut (.I0(n56622), .I1(duty[1]), .I2(n269), .I3(duty[23]), 
            .O(pwm_setpoint_23__N_11[1]));
    defparam n56622_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1640_3_lut (.I0(n2413), 
            .I1(n2480), .I2(n2445), .I3(GND_net), .O(n2512));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1640_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1644_3_lut (.I0(n2417), 
            .I1(n2484), .I2(n2445), .I3(GND_net), .O(n2516));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1644_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1643_3_lut (.I0(n2416), 
            .I1(n2483), .I2(n2445), .I3(GND_net), .O(n2515));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1643_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1642_3_lut (.I0(n2415), 
            .I1(n2482), .I2(n2445), .I3(GND_net), .O(n2514));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1642_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1649_3_lut (.I0(n2422), 
            .I1(n2489), .I2(n2445), .I3(GND_net), .O(n2521));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1649_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1648_3_lut (.I0(n2421), 
            .I1(n2488), .I2(n2445), .I3(GND_net), .O(n2520));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1648_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1647_3_lut (.I0(n2420), 
            .I1(n2487), .I2(n2445), .I3(GND_net), .O(n2519));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1647_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1661_3_lut (.I0(n535), .I1(n2501), 
            .I2(n2445), .I3(GND_net), .O(n2533));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1661_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1660_3_lut (.I0(n2433), 
            .I1(n2500), .I2(n2445), .I3(GND_net), .O(n2532));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1660_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_mux_3_i9_3_lut (.I0(encoder0_position_scaled_23__N_327[8]), 
            .I1(n25_adj_5474), .I2(encoder0_position_scaled_23__N_327[31]), 
            .I3(GND_net), .O(n536));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_mux_3_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1646_3_lut (.I0(n2419), 
            .I1(n2486), .I2(n2445), .I3(GND_net), .O(n2518));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1646_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1645_3_lut (.I0(n2418), 
            .I1(n2485), .I2(n2445), .I3(GND_net), .O(n2517));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1645_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1650_3_lut (.I0(n2423), 
            .I1(n2490), .I2(n2445), .I3(GND_net), .O(n2522));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1650_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i39843_3_lut (.I0(n2228), .I1(n2295), .I2(n2247), .I3(GND_net), 
            .O(n2327));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam i39843_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i39844_3_lut (.I0(n2327), .I1(n2394), .I2(n2346), .I3(GND_net), 
            .O(n2426));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam i39844_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i39760_3_lut (.I0(n2426), .I1(n2493), .I2(n2445), .I3(GND_net), 
            .O(n2525));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam i39760_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1652_3_lut (.I0(n2425), 
            .I1(n2492), .I2(n2445), .I3(GND_net), .O(n2524));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1652_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1659_3_lut (.I0(n2432), 
            .I1(n2499), .I2(n2445), .I3(GND_net), .O(n2531));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1659_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1658_3_lut (.I0(n2431), 
            .I1(n2498), .I2(n2445), .I3(GND_net), .O(n2530));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1658_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1657_3_lut (.I0(n2430), 
            .I1(n2497), .I2(n2445), .I3(GND_net), .O(n2529));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1657_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1655_3_lut (.I0(n2428), 
            .I1(n2495), .I2(n2445), .I3(GND_net), .O(n2527));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1655_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1656_3_lut (.I0(n2429), 
            .I1(n2496), .I2(n2445), .I3(GND_net), .O(n2528));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1656_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1654_3_lut (.I0(n2427), 
            .I1(n2494), .I2(n2445), .I3(GND_net), .O(n2526));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1654_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i39845_3_lut (.I0(n2226), .I1(n2293), .I2(n2247), .I3(GND_net), 
            .O(n2325));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam i39845_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i39846_3_lut (.I0(n2325), .I1(n2392), .I2(n2346), .I3(GND_net), 
            .O(n2424));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam i39846_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i39758_3_lut (.I0(n2424), .I1(n2491), .I2(n2445), .I3(GND_net), 
            .O(n2523));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam i39758_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1884 (.I0(n2523), .I1(n2526), .I2(n2528), .I3(n2527), 
            .O(n51792));
    defparam i1_4_lut_adj_1884.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1885 (.I0(n2524), .I1(n51792), .I2(n2525), .I3(n2522), 
            .O(n51794));
    defparam i1_4_lut_adj_1885.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i905_3_lut (.I0(n1326), .I1(n1393), 
            .I2(n1356), .I3(GND_net), .O(n1425));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i905_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i23226_3_lut (.I0(n536), .I1(n2532), .I2(n2533), .I3(GND_net), 
            .O(n37316));
    defparam i23226_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i1_4_lut_adj_1886 (.I0(n2519), .I1(n2520), .I2(n51794), .I3(n2521), 
            .O(n51800));
    defparam i1_4_lut_adj_1886.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1887 (.I0(n2529), .I1(n37316), .I2(n2530), .I3(n2531), 
            .O(n50075));
    defparam i1_4_lut_adj_1887.LUT_INIT = 16'ha080;
    SB_LUT4 i1_4_lut_adj_1888 (.I0(n2517), .I1(n2518), .I2(n50075), .I3(n51800), 
            .O(n51806));
    defparam i1_4_lut_adj_1888.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1889 (.I0(n2514), .I1(n2515), .I2(n2516), .I3(n51806), 
            .O(n51812));
    defparam i1_4_lut_adj_1889.LUT_INIT = 16'hfffe;
    SB_LUT4 i40315_4_lut (.I0(n2512), .I1(n2511), .I2(n2513), .I3(n51812), 
            .O(n2544));
    defparam i40315_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1590_3_lut (.I0(n2331), 
            .I1(n2398), .I2(n2346), .I3(GND_net), .O(n2430));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1590_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1589_3_lut (.I0(n2330), 
            .I1(n2397), .I2(n2346), .I3(GND_net), .O(n2429));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1589_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1580_3_lut (.I0(n2321), 
            .I1(n2388), .I2(n2346), .I3(GND_net), .O(n2420));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1580_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1579_3_lut (.I0(n2320), 
            .I1(n2387), .I2(n2346), .I3(GND_net), .O(n2419));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1579_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1506_3_lut (.I0(n2215), 
            .I1(n2282), .I2(n2247), .I3(GND_net), .O(n2314));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1506_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1507_3_lut (.I0(n2216), 
            .I1(n2283), .I2(n2247), .I3(GND_net), .O(n2315));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1507_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1574_3_lut (.I0(n2315), 
            .I1(n2382), .I2(n2346), .I3(GND_net), .O(n2414));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1574_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1573_3_lut (.I0(n2314), 
            .I1(n2381), .I2(n2346), .I3(GND_net), .O(n2413));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1573_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1577_3_lut (.I0(n2318), 
            .I1(n2385), .I2(n2346), .I3(GND_net), .O(n2417));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1577_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1576_3_lut (.I0(n2317), 
            .I1(n2384), .I2(n2346), .I3(GND_net), .O(n2416));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1576_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1575_3_lut (.I0(n2316), 
            .I1(n2383), .I2(n2346), .I3(GND_net), .O(n2415));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1575_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1578_3_lut (.I0(n2319), 
            .I1(n2386), .I2(n2346), .I3(GND_net), .O(n2418));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1578_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1593_3_lut (.I0(n534), .I1(n2401), 
            .I2(n2346), .I3(GND_net), .O(n2433));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1593_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1592_3_lut (.I0(n2333), 
            .I1(n2400), .I2(n2346), .I3(GND_net), .O(n2432));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1592_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1591_3_lut (.I0(n2332), 
            .I1(n2399), .I2(n2346), .I3(GND_net), .O(n2431));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1591_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_mux_3_i10_3_lut (.I0(encoder0_position_scaled_23__N_327[9]), 
            .I1(n24_adj_5475), .I2(encoder0_position_scaled_23__N_327[31]), 
            .I3(GND_net), .O(n535));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_mux_3_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1585_3_lut (.I0(n2326), 
            .I1(n2393), .I2(n2346), .I3(GND_net), .O(n2425));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1585_3_lut.LUT_INIT = 16'hacac;
    EEPROM eeprom (.\state[3] (state_adj_5736[3]), .n6(n6), .GND_net(GND_net), 
           .clk16MHz(clk16MHz), .read(read), .\state[0] (state_adj_5705[0]), 
           .enable_slow_N_4393(enable_slow_N_4393), .n6271({n6272}), .\state[1] (state_adj_5705[1]), 
           .n48526(n48526), .VCC_net(VCC_net), .n48558(n48558), .n29393(n29393), 
           .rw(rw), .n48670(n48670), .data_ready(data_ready), .n36659(n36659), 
           .n49838(n49838), .n49919(n49919), .\state_7__N_4290[0] (state_7__N_4290[0]), 
           .n4(n4_adj_5555), .n4_adj_18(n4), .n36542(n36542), .n7354(n7354), 
           .\state[2] (state_adj_5736[2]), .n26(n26_adj_5575), .\state_7__N_4306[3] (state_7__N_4306[3]), 
           .n7936(n7936), .scl_enable(scl_enable), .\saved_addr[0] (saved_addr[0]), 
           .\state[0]_adj_19 (state_adj_5736[0]), .n29452(n29452), .sda_enable(sda_enable), 
           .n29364(n29364), .data({data}), .n29363(n29363), .n29362(n29362), 
           .n29361(n29361), .n29360(n29360), .n29359(n29359), .n29358(n29358), 
           .n10(n10), .n10_adj_20(n10_adj_5610), .n8(n8_adj_5654), .n29835(n29835), 
           .n54609(n54609), .n27243(n27243), .n27238(n27238), .scl(scl), 
           .sda_out(sda_out)) /* synthesis syn_noprune=1, syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(398[10] 409[6])
    SB_LUT4 i39316_3_lut (.I0(n2323), .I1(n2390), .I2(n2346), .I3(GND_net), 
            .O(n2422));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam i39316_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1587_3_lut (.I0(n2328), 
            .I1(n2395), .I2(n2346), .I3(GND_net), .O(n2427));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1587_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1583_3_lut (.I0(n2324), 
            .I1(n2391), .I2(n2346), .I3(GND_net), .O(n2423));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1583_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1588_3_lut (.I0(n2329), 
            .I1(n2396), .I2(n2346), .I3(GND_net), .O(n2428));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1588_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i2_2_lut_3_lut (.I0(hall1), .I1(hall3), .I2(hall2), .I3(GND_net), 
            .O(commutation_state_7__N_272));   // verilog/TinyFPGA_B.v(166[7:32])
    defparam i2_2_lut_3_lut.LUT_INIT = 16'h0404;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1581_3_lut (.I0(n2322), 
            .I1(n2389), .I2(n2346), .I3(GND_net), .O(n2421));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1581_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 n10829_bdd_4_lut_40793 (.I0(n10829), .I1(n441), .I2(current[0]), 
            .I3(duty[23]), .O(n56616));
    defparam n10829_bdd_4_lut_40793.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_4_lut_adj_1890 (.I0(n2423), .I1(n2427), .I2(n2422), .I3(n2425), 
            .O(n52084));
    defparam i1_4_lut_adj_1890.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1891 (.I0(n2426), .I1(n2421), .I2(n2428), .I3(n2424), 
            .O(n52086));
    defparam i1_4_lut_adj_1891.LUT_INIT = 16'hfffe;
    SB_LUT4 i23296_4_lut (.I0(n535), .I1(n2431), .I2(n2432), .I3(n2433), 
            .O(n37386));
    defparam i23296_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 i1_4_lut_adj_1892 (.I0(n2419), .I1(n2420), .I2(n52086), .I3(n52084), 
            .O(n52092));
    defparam i1_4_lut_adj_1892.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_adj_1893 (.I0(n2429), .I1(n2430), .I2(GND_net), .I3(GND_net), 
            .O(n52278));
    defparam i1_2_lut_adj_1893.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut_adj_1894 (.I0(n2418), .I1(n52278), .I2(n52092), .I3(n37386), 
            .O(n52096));
    defparam i1_4_lut_adj_1894.LUT_INIT = 16'hfefa;
    SB_LUT4 i1_4_lut_adj_1895 (.I0(n2415), .I1(n2416), .I2(n2417), .I3(n52096), 
            .O(n52102));
    defparam i1_4_lut_adj_1895.LUT_INIT = 16'hfffe;
    SB_LUT4 i40344_4_lut (.I0(n2413), .I1(n2412), .I2(n2414), .I3(n52102), 
            .O(n2445));
    defparam i40344_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i979_3_lut (.I0(n1432), .I1(n1499), 
            .I2(n1455), .I3(GND_net), .O(n1531));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i979_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1046_3_lut (.I0(n1531), 
            .I1(n1598), .I2(n1554_adj_5597), .I3(GND_net), .O(n1630));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1046_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1113_3_lut (.I0(n1630), 
            .I1(n1697), .I2(n1653), .I3(GND_net), .O(n1729));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1113_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1180_rep_44_3_lut (.I0(n1729), 
            .I1(n1796), .I2(n1752), .I3(GND_net), .O(n1828));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1180_rep_44_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1247_3_lut (.I0(n1828), 
            .I1(n1895), .I2(n1851), .I3(GND_net), .O(n1927));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1247_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1314_3_lut (.I0(n1927), 
            .I1(n1994), .I2(n1950), .I3(GND_net), .O(n2026));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1314_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1381_rep_36_3_lut (.I0(n2026), 
            .I1(n2093), .I2(n2049), .I3(GND_net), .O(n2125));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1381_rep_36_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1448_rep_27_3_lut (.I0(n2192), 
            .I1(n2291), .I2(n2247), .I3(GND_net), .O(n53094));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1448_rep_27_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1510_3_lut (.I0(n2219), 
            .I1(n2286), .I2(n2247), .I3(GND_net), .O(n2318));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1510_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1509_3_lut (.I0(n2218), 
            .I1(n2285), .I2(n2247), .I3(GND_net), .O(n2317));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1509_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1508_3_lut (.I0(n2217), 
            .I1(n2284), .I2(n2247), .I3(GND_net), .O(n2316));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1508_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_mux_3_i15_3_lut (.I0(encoder0_position_scaled_23__N_327[14]), 
            .I1(n19_adj_5480), .I2(encoder0_position_scaled_23__N_327[31]), 
            .I3(GND_net), .O(n530));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_mux_3_i15_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1321_3_lut (.I0(n530), .I1(n2001), 
            .I2(n1950), .I3(GND_net), .O(n2033));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1321_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1388_3_lut (.I0(n2033), 
            .I1(n2100), .I2(n2049), .I3(GND_net), .O(n2132));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1388_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_mux_3_i16_3_lut (.I0(encoder0_position_scaled_23__N_327[15]), 
            .I1(n18_adj_5481), .I2(encoder0_position_scaled_23__N_327[31]), 
            .I3(GND_net), .O(n529));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_mux_3_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1253_3_lut (.I0(n529), .I1(n1901), 
            .I2(n1851), .I3(GND_net), .O(n1933));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1253_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1320_3_lut (.I0(n1933), 
            .I1(n2000), .I2(n1950), .I3(GND_net), .O(n2032));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1320_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1387_3_lut (.I0(n2032), 
            .I1(n2099), .I2(n2049), .I3(GND_net), .O(n2131));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1387_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1454_3_lut (.I0(n2131), 
            .I1(n2198), .I2(n2148), .I3(GND_net), .O(n2230));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1454_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1455_3_lut (.I0(n2132), 
            .I1(n2199), .I2(n2148), .I3(GND_net), .O(n2231));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1455_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1522_3_lut (.I0(n2231), 
            .I1(n2298), .I2(n2247), .I3(GND_net), .O(n2330));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1522_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1521_3_lut (.I0(n2230), 
            .I1(n2297), .I2(n2247), .I3(GND_net), .O(n2329));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1521_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_mux_3_i14_3_lut (.I0(encoder0_position_scaled_23__N_327[13]), 
            .I1(n20_adj_5479), .I2(encoder0_position_scaled_23__N_327[31]), 
            .I3(GND_net), .O(n531));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_mux_3_i14_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1389_3_lut (.I0(n531), .I1(n2101), 
            .I2(n2049), .I3(GND_net), .O(n2133));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1389_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_mux_3_i13_3_lut (.I0(encoder0_position_scaled_23__N_327[12]), 
            .I1(n21_adj_5478), .I2(encoder0_position_scaled_23__N_327[31]), 
            .I3(GND_net), .O(n532));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_mux_3_i13_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1457_3_lut (.I0(n532), .I1(n2201), 
            .I2(n2148), .I3(GND_net), .O(n2233_adj_5599));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1457_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_mux_3_i12_3_lut (.I0(encoder0_position_scaled_23__N_327[11]), 
            .I1(n22_adj_5477), .I2(encoder0_position_scaled_23__N_327[31]), 
            .I3(GND_net), .O(n533));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_mux_3_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1456_3_lut (.I0(n2133), 
            .I1(n2200), .I2(n2148), .I3(GND_net), .O(n2232));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1456_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1525_3_lut (.I0(n533), .I1(n2301), 
            .I2(n2247), .I3(GND_net), .O(n2333));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1525_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i40627_1_lut (.I0(n1059), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n56458));
    defparam i40627_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_unary_minus_2_inv_0_i32_1_lut (.I0(encoder0_position_scaled_23__N_327[31]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n2_adj_5611));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_unary_minus_2_inv_0_i32_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1524_3_lut (.I0(n2233_adj_5599), 
            .I1(n2300), .I2(n2247), .I3(GND_net), .O(n2332));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1524_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1523_3_lut (.I0(n2232), 
            .I1(n2299), .I2(n2247), .I3(GND_net), .O(n2331));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1523_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_mux_3_i11_3_lut (.I0(encoder0_position_scaled_23__N_327[10]), 
            .I1(n23_adj_5476), .I2(encoder0_position_scaled_23__N_327[31]), 
            .I3(GND_net), .O(n534));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_mux_3_i11_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i908_3_lut (.I0(n1329), .I1(n1396), 
            .I2(n1356), .I3(GND_net), .O(n1428));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i908_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15845_3_lut (.I0(PWMLimit[16]), .I1(\data_in_frame[8] [0]), 
            .I2(n50654), .I3(GND_net), .O(n29925));   // verilog/coms.v(128[12] 303[6])
    defparam i15845_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i34010_3_lut (.I0(encoder0_position_scaled_23__N_327[26]), .I1(n49757), 
            .I2(encoder0_position_scaled_23__N_327[31]), .I3(GND_net), .O(n833));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam i34010_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i975_3_lut (.I0(n1428), .I1(n1495), 
            .I2(n1455), .I3(GND_net), .O(n1527));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i975_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1042_3_lut (.I0(n1527), 
            .I1(n1594), .I2(n1554_adj_5597), .I3(GND_net), .O(n1626));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1042_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1109_3_lut (.I0(n1626), 
            .I1(n1693), .I2(n1653), .I3(GND_net), .O(n1725));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1109_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1176_3_lut (.I0(n1725), 
            .I1(n1792), .I2(n1752), .I3(GND_net), .O(n1824));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1176_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15339_3_lut (.I0(\data_out_frame[7] [4]), .I1(encoder0_position_scaled[12]), 
            .I2(n24210), .I3(GND_net), .O(n29419));   // verilog/coms.v(128[12] 303[6])
    defparam i15339_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1243_3_lut (.I0(n1824), 
            .I1(n1891), .I2(n1851), .I3(GND_net), .O(n1923));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1243_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15340_3_lut (.I0(\data_out_frame[7] [3]), .I1(encoder0_position_scaled[11]), 
            .I2(n24210), .I3(GND_net), .O(n29420));   // verilog/coms.v(128[12] 303[6])
    defparam i15340_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15341_3_lut (.I0(\data_out_frame[7] [2]), .I1(encoder0_position_scaled[10]), 
            .I2(n24210), .I3(GND_net), .O(n29421));   // verilog/coms.v(128[12] 303[6])
    defparam i15341_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15342_3_lut (.I0(\data_out_frame[7] [1]), .I1(encoder0_position_scaled[9]), 
            .I2(n24210), .I3(GND_net), .O(n29422));   // verilog/coms.v(128[12] 303[6])
    defparam i15342_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15343_3_lut (.I0(\data_out_frame[7] [0]), .I1(encoder0_position_scaled[8]), 
            .I2(n24210), .I3(GND_net), .O(n29423));   // verilog/coms.v(128[12] 303[6])
    defparam i15343_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15344_3_lut (.I0(\data_out_frame[6] [7]), .I1(encoder0_position_scaled[23]), 
            .I2(n24210), .I3(GND_net), .O(n29424));   // verilog/coms.v(128[12] 303[6])
    defparam i15344_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1310_3_lut (.I0(n1923), 
            .I1(n1990), .I2(n1950), .I3(GND_net), .O(n2022));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1310_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15345_3_lut (.I0(\data_out_frame[6] [6]), .I1(encoder0_position_scaled[22]), 
            .I2(n24210), .I3(GND_net), .O(n29425));   // verilog/coms.v(128[12] 303[6])
    defparam i15345_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15346_3_lut (.I0(\data_out_frame[6] [5]), .I1(encoder0_position_scaled[21]), 
            .I2(n24210), .I3(GND_net), .O(n29426));   // verilog/coms.v(128[12] 303[6])
    defparam i15346_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15347_3_lut (.I0(\data_out_frame[6] [4]), .I1(encoder0_position_scaled[20]), 
            .I2(n24210), .I3(GND_net), .O(n29427));   // verilog/coms.v(128[12] 303[6])
    defparam i15347_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1377_3_lut (.I0(n2022), 
            .I1(n2089), .I2(n2049), .I3(GND_net), .O(n2121));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1377_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1444_3_lut (.I0(n2121), 
            .I1(n2188), .I2(n2148), .I3(GND_net), .O(n2220));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1444_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1511_3_lut (.I0(n2220), 
            .I1(n2287), .I2(n2247), .I3(GND_net), .O(n2319));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1511_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_mux_3_i17_3_lut (.I0(encoder0_position_scaled_23__N_327[16]), 
            .I1(n17_adj_5482), .I2(encoder0_position_scaled_23__N_327[31]), 
            .I3(GND_net), .O(n942));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_mux_3_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15348_3_lut (.I0(\data_out_frame[6] [3]), .I1(encoder0_position_scaled[19]), 
            .I2(n24210), .I3(GND_net), .O(n29428));   // verilog/coms.v(128[12] 303[6])
    defparam i15348_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1185_3_lut (.I0(n942), .I1(n1801), 
            .I2(n1752), .I3(GND_net), .O(n1833));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1185_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1252_3_lut (.I0(n1833), 
            .I1(n1900), .I2(n1851), .I3(GND_net), .O(n1932));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1252_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15349_3_lut (.I0(\data_out_frame[6] [2]), .I1(encoder0_position_scaled[18]), 
            .I2(n24210), .I3(GND_net), .O(n29429));   // verilog/coms.v(128[12] 303[6])
    defparam i15349_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1319_3_lut (.I0(n1932), 
            .I1(n1999), .I2(n1950), .I3(GND_net), .O(n2031));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1319_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1386_3_lut (.I0(n2031), 
            .I1(n2098), .I2(n2049), .I3(GND_net), .O(n2130));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1386_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i913_3_lut (.I0(n413), .I1(n1401), 
            .I2(n1356), .I3(GND_net), .O(n1433));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i913_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i980_3_lut (.I0(n1433), .I1(n1500), 
            .I2(n1455), .I3(GND_net), .O(n1532_adj_5595));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i980_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15350_3_lut (.I0(\data_out_frame[6] [1]), .I1(encoder0_position_scaled[17]), 
            .I2(n24210), .I3(GND_net), .O(n29430));   // verilog/coms.v(128[12] 303[6])
    defparam i15350_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15351_3_lut (.I0(\data_out_frame[6] [0]), .I1(encoder0_position_scaled[16]), 
            .I2(n24210), .I3(GND_net), .O(n29431));   // verilog/coms.v(128[12] 303[6])
    defparam i15351_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15352_3_lut (.I0(\data_out_frame[5] [7]), .I1(control_mode[7]), 
            .I2(n24210), .I3(GND_net), .O(n29432));   // verilog/coms.v(128[12] 303[6])
    defparam i15352_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15353_3_lut (.I0(\data_out_frame[5] [6]), .I1(control_mode[6]), 
            .I2(n24210), .I3(GND_net), .O(n29433));   // verilog/coms.v(128[12] 303[6])
    defparam i15353_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1047_3_lut (.I0(n1532_adj_5595), 
            .I1(n1599), .I2(n1554_adj_5597), .I3(GND_net), .O(n1631));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1047_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15354_3_lut (.I0(\data_out_frame[5] [5]), .I1(control_mode[5]), 
            .I2(n24210), .I3(GND_net), .O(n29434));   // verilog/coms.v(128[12] 303[6])
    defparam i15354_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1114_3_lut (.I0(n1631), 
            .I1(n1698), .I2(n1653), .I3(GND_net), .O(n1730));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1114_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1181_3_lut (.I0(n1730), 
            .I1(n1797), .I2(n1752), .I3(GND_net), .O(n1829));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1181_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15355_3_lut (.I0(\data_out_frame[5] [4]), .I1(control_mode[4]), 
            .I2(n24210), .I3(GND_net), .O(n29435));   // verilog/coms.v(128[12] 303[6])
    defparam i15355_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i22660_2_lut_2_lut (.I0(duty[20]), .I1(n296), .I2(GND_net), 
            .I3(GND_net), .O(n4909));   // verilog/TinyFPGA_B.v(123[17] 125[11])
    defparam i22660_2_lut_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i15356_3_lut (.I0(\data_out_frame[5] [3]), .I1(control_mode[3]), 
            .I2(n24210), .I3(GND_net), .O(n29436));   // verilog/coms.v(128[12] 303[6])
    defparam i15356_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15357_3_lut (.I0(\data_out_frame[5] [2]), .I1(control_mode[2]), 
            .I2(n24210), .I3(GND_net), .O(n29437));   // verilog/coms.v(128[12] 303[6])
    defparam i15357_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15358_3_lut (.I0(\data_out_frame[5] [1]), .I1(control_mode[1]), 
            .I2(n24210), .I3(GND_net), .O(n29438));   // verilog/coms.v(128[12] 303[6])
    defparam i15358_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1248_3_lut (.I0(n1829), 
            .I1(n1896), .I2(n1851), .I3(GND_net), .O(n1928));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1248_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1315_3_lut (.I0(n1928), 
            .I1(n1995), .I2(n1950), .I3(GND_net), .O(n2027));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1315_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15359_3_lut (.I0(\data_out_frame[5] [0]), .I1(control_mode[0]), 
            .I2(n24210), .I3(GND_net), .O(n29439));   // verilog/coms.v(128[12] 303[6])
    defparam i15359_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15360_3_lut (.I0(\data_out_frame[4] [7]), .I1(ID[7]), .I2(n24210), 
            .I3(GND_net), .O(n29440));   // verilog/coms.v(128[12] 303[6])
    defparam i15360_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15361_3_lut (.I0(\data_out_frame[4] [6]), .I1(ID[6]), .I2(n24210), 
            .I3(GND_net), .O(n29441));   // verilog/coms.v(128[12] 303[6])
    defparam i15361_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1382_3_lut (.I0(n2027), 
            .I1(n2094), .I2(n2049), .I3(GND_net), .O(n2126));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1382_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1449_3_lut (.I0(n2126), 
            .I1(n2193), .I2(n2148), .I3(GND_net), .O(n2225));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1449_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1453_3_lut (.I0(n2130), 
            .I1(n2197), .I2(n2148), .I3(GND_net), .O(n2229));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1453_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15362_3_lut (.I0(\data_out_frame[4] [5]), .I1(ID[5]), .I2(n24210), 
            .I3(GND_net), .O(n29442));   // verilog/coms.v(128[12] 303[6])
    defparam i15362_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1516_3_lut (.I0(n2225), 
            .I1(n2292), .I2(n2247), .I3(GND_net), .O(n2324));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1516_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1520_3_lut (.I0(n2229), 
            .I1(n2296), .I2(n2247), .I3(GND_net), .O(n2328));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1520_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15363_3_lut (.I0(\data_out_frame[4] [4]), .I1(ID[4]), .I2(n24210), 
            .I3(GND_net), .O(n29443));   // verilog/coms.v(128[12] 303[6])
    defparam i15363_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15364_3_lut (.I0(\data_out_frame[4] [3]), .I1(ID[3]), .I2(n24210), 
            .I3(GND_net), .O(n29444));   // verilog/coms.v(128[12] 303[6])
    defparam i15364_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15365_3_lut (.I0(\data_out_frame[4] [2]), .I1(ID[2]), .I2(n24210), 
            .I3(GND_net), .O(n29445));   // verilog/coms.v(128[12] 303[6])
    defparam i15365_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15366_3_lut (.I0(\data_out_frame[4] [1]), .I1(ID[1]), .I2(n24210), 
            .I3(GND_net), .O(n29446));   // verilog/coms.v(128[12] 303[6])
    defparam i15366_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i978_3_lut (.I0(n1431), .I1(n1498), 
            .I2(n1455), .I3(GND_net), .O(n1530));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i978_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1045_3_lut (.I0(n1530), 
            .I1(n1597), .I2(n1554_adj_5597), .I3(GND_net), .O(n1629));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1045_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1112_3_lut (.I0(n1629), 
            .I1(n1696), .I2(n1653), .I3(GND_net), .O(n1728));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1112_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1179_rep_45_3_lut (.I0(n1728), 
            .I1(n1795), .I2(n1752), .I3(GND_net), .O(n1827));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1179_rep_45_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1246_3_lut (.I0(n1827), 
            .I1(n1894), .I2(n1851), .I3(GND_net), .O(n1926));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1246_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i38982_2_lut_4_lut (.I0(commutation_state[0]), .I1(n4_adj_5607), 
            .I2(commutation_state_prev[0]), .I3(dti_counter[0]), .O(n54586));   // verilog/TinyFPGA_B.v(146[7:48])
    defparam i38982_2_lut_4_lut.LUT_INIT = 16'h2100;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1313_3_lut (.I0(n1926), 
            .I1(n1993), .I2(n1950), .I3(GND_net), .O(n2025));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1313_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1380_3_lut (.I0(n2025), 
            .I1(n2092), .I2(n2049), .I3(GND_net), .O(n2124));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1380_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i910_3_lut (.I0(n1331), .I1(n1398), 
            .I2(n1356), .I3(GND_net), .O(n1430));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i910_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i977_3_lut (.I0(n1430), .I1(n1497), 
            .I2(n1455), .I3(GND_net), .O(n1529));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i977_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1044_3_lut (.I0(n1529), 
            .I1(n1596), .I2(n1554_adj_5597), .I3(GND_net), .O(n1628));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1044_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i38917_2_lut_4_lut (.I0(commutation_state[0]), .I1(n4_adj_5607), 
            .I2(commutation_state_prev[0]), .I3(dti_counter[1]), .O(n54553));   // verilog/TinyFPGA_B.v(146[7:48])
    defparam i38917_2_lut_4_lut.LUT_INIT = 16'h2100;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1111_3_lut (.I0(n1628), 
            .I1(n1695), .I2(n1653), .I3(GND_net), .O(n1727));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1111_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i39618_3_lut (.I0(n1826), .I1(n1893), .I2(n1851), .I3(GND_net), 
            .O(n1925));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam i39618_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i38988_2_lut_4_lut (.I0(commutation_state[0]), .I1(n4_adj_5607), 
            .I2(commutation_state_prev[0]), .I3(dti_counter[2]), .O(n54552));   // verilog/TinyFPGA_B.v(146[7:48])
    defparam i38988_2_lut_4_lut.LUT_INIT = 16'h2100;
    SB_LUT4 i38986_2_lut_4_lut (.I0(commutation_state[0]), .I1(n4_adj_5607), 
            .I2(commutation_state_prev[0]), .I3(dti_counter[3]), .O(n54551));   // verilog/TinyFPGA_B.v(146[7:48])
    defparam i38986_2_lut_4_lut.LUT_INIT = 16'h2100;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1312_3_lut (.I0(n1925), 
            .I1(n1992), .I2(n1950), .I3(GND_net), .O(n2024));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1312_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1379_3_lut (.I0(n2024), 
            .I1(n2091_adj_5598), .I2(n2049), .I3(GND_net), .O(n2123));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1379_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1446_3_lut (.I0(n2123), 
            .I1(n2190), .I2(n2148), .I3(GND_net), .O(n2222));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1446_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i38985_2_lut_4_lut (.I0(commutation_state[0]), .I1(n4_adj_5607), 
            .I2(commutation_state_prev[0]), .I3(dti_counter[4]), .O(n54550));   // verilog/TinyFPGA_B.v(146[7:48])
    defparam i38985_2_lut_4_lut.LUT_INIT = 16'h2100;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i909_3_lut (.I0(n1330), .I1(n1397), 
            .I2(n1356), .I3(GND_net), .O(n1429));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i909_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i976_3_lut (.I0(n1429), .I1(n1496), 
            .I2(n1455), .I3(GND_net), .O(n1528));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i976_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1043_3_lut (.I0(n1528), 
            .I1(n1595), .I2(n1554_adj_5597), .I3(GND_net), .O(n1627));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1043_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1110_3_lut (.I0(n1627), 
            .I1(n1694), .I2(n1653), .I3(GND_net), .O(n1726));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1110_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i39616_3_lut (.I0(n1825), .I1(n1892), .I2(n1851), .I3(GND_net), 
            .O(n1924));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam i39616_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1311_3_lut (.I0(n1924), 
            .I1(n1991), .I2(n1950), .I3(GND_net), .O(n2023));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1311_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i38984_2_lut_4_lut (.I0(commutation_state[0]), .I1(n4_adj_5607), 
            .I2(commutation_state_prev[0]), .I3(dti_counter[5]), .O(n54549));   // verilog/TinyFPGA_B.v(146[7:48])
    defparam i38984_2_lut_4_lut.LUT_INIT = 16'h2100;
    SB_LUT4 i15367_3_lut (.I0(\data_out_frame[4] [0]), .I1(ID[0]), .I2(n24210), 
            .I3(GND_net), .O(n29447));   // verilog/coms.v(128[12] 303[6])
    defparam i15367_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15368_3_lut (.I0(\data_in[3] [7]), .I1(rx_data[7]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n29448));   // verilog/coms.v(128[12] 303[6])
    defparam i15368_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15369_3_lut (.I0(\data_in[3] [6]), .I1(rx_data[6]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n29449));   // verilog/coms.v(128[12] 303[6])
    defparam i15369_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15370_3_lut (.I0(\data_in[3] [5]), .I1(rx_data[5]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n29450));   // verilog/coms.v(128[12] 303[6])
    defparam i15370_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1378_3_lut (.I0(n2023), 
            .I1(n2090), .I2(n2049), .I3(GND_net), .O(n2122));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1378_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i38946_2_lut_4_lut (.I0(commutation_state[0]), .I1(n4_adj_5607), 
            .I2(commutation_state_prev[0]), .I3(dti_counter[6]), .O(n54548));   // verilog/TinyFPGA_B.v(146[7:48])
    defparam i38946_2_lut_4_lut.LUT_INIT = 16'h2100;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1445_3_lut (.I0(n2122), 
            .I1(n2189), .I2(n2148), .I3(GND_net), .O(n2221));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1445_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1447_3_lut (.I0(n2124), 
            .I1(n2191), .I2(n2148), .I3(GND_net), .O(n2223));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1447_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1514_3_lut (.I0(n2223), 
            .I1(n2290), .I2(n2247), .I3(GND_net), .O(n2322));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1514_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1513_3_lut (.I0(n2222), 
            .I1(n2289), .I2(n2247), .I3(GND_net), .O(n2321));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1513_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1512_3_lut (.I0(n2221), 
            .I1(n2288), .I2(n2247), .I3(GND_net), .O(n2320));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1512_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_mux_3_i18_3_lut (.I0(encoder0_position_scaled_23__N_327[17]), 
            .I1(n16_adj_5483), .I2(encoder0_position_scaled_23__N_327[31]), 
            .I3(GND_net), .O(n941));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_mux_3_i18_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1117_3_lut (.I0(n941), .I1(n1701), 
            .I2(n1653), .I3(GND_net), .O(n1733));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1117_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i38925_2_lut_4_lut (.I0(commutation_state[0]), .I1(n4_adj_5607), 
            .I2(commutation_state_prev[0]), .I3(dti_counter[7]), .O(n54547));   // verilog/TinyFPGA_B.v(146[7:48])
    defparam i38925_2_lut_4_lut.LUT_INIT = 16'h2100;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1448_3_lut (.I0(n2125), 
            .I1(n2192), .I2(n2148), .I3(GND_net), .O(n2224));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1448_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut (.I0(commutation_state[0]), .I1(n4_adj_5607), 
            .I2(commutation_state_prev[0]), .I3(dti_N_527), .O(n28648));   // verilog/TinyFPGA_B.v(146[7:48])
    defparam i1_2_lut_4_lut.LUT_INIT = 16'hdeff;
    SB_LUT4 i15846_3_lut (.I0(PWMLimit[15]), .I1(\data_in_frame[9] [7]), 
            .I2(n50654), .I3(GND_net), .O(n29926));   // verilog/coms.v(128[12] 303[6])
    defparam i15846_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1184_3_lut (.I0(n1733), 
            .I1(n1800), .I2(n1752), .I3(GND_net), .O(n1832));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1184_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15371_3_lut (.I0(\data_in[3] [4]), .I1(rx_data[4]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n29451));   // verilog/coms.v(128[12] 303[6])
    defparam i15371_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1251_3_lut (.I0(n1832), 
            .I1(n1899), .I2(n1851), .I3(GND_net), .O(n1931));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1251_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1318_3_lut (.I0(n1931), 
            .I1(n1998), .I2(n1950), .I3(GND_net), .O(n2030));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1318_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15372_4_lut (.I0(saved_addr[0]), .I1(rw), .I2(state_7__N_4290[0]), 
            .I3(enable_slow_N_4393), .O(n29452));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i15372_4_lut.LUT_INIT = 16'haaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1385_3_lut (.I0(n2030), 
            .I1(n2097), .I2(n2049), .I3(GND_net), .O(n2129));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1385_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1452_rep_32_3_lut (.I0(n2129), 
            .I1(n2196), .I2(n2148), .I3(GND_net), .O(n2228));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1452_rep_32_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15373_3_lut (.I0(\data_in[3] [3]), .I1(rx_data[3]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n29453));   // verilog/coms.v(128[12] 303[6])
    defparam i15373_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15374_3_lut (.I0(\data_in[3] [2]), .I1(rx_data[2]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n29454));   // verilog/coms.v(128[12] 303[6])
    defparam i15374_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_mux_3_i19_3_lut (.I0(encoder0_position_scaled_23__N_327[18]), 
            .I1(n15_adj_5484), .I2(encoder0_position_scaled_23__N_327[31]), 
            .I3(GND_net), .O(n415));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_mux_3_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1049_3_lut (.I0(n415), .I1(n1601), 
            .I2(n1554_adj_5597), .I3(GND_net), .O(n1633));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1049_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1116_3_lut (.I0(n1633), 
            .I1(n1700), .I2(n1653), .I3(GND_net), .O(n1732));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1116_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1183_3_lut (.I0(n1732), 
            .I1(n1799), .I2(n1752), .I3(GND_net), .O(n1831));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1183_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1250_3_lut (.I0(n1831), 
            .I1(n1898), .I2(n1851), .I3(GND_net), .O(n1930));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1250_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1317_3_lut (.I0(n1930), 
            .I1(n1997), .I2(n1950), .I3(GND_net), .O(n2029));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1317_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1384_3_lut (.I0(n2029), 
            .I1(n2096), .I2(n2049), .I3(GND_net), .O(n2128));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1384_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1451_3_lut (.I0(n2128), 
            .I1(n2195), .I2(n2148), .I3(GND_net), .O(n2227));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1451_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15375_3_lut (.I0(\data_in[3] [1]), .I1(rx_data[1]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n29455));   // verilog/coms.v(128[12] 303[6])
    defparam i15375_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15376_3_lut (.I0(\data_in[3] [0]), .I1(rx_data[0]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n29456));   // verilog/coms.v(128[12] 303[6])
    defparam i15376_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15380_3_lut (.I0(\data_in[2] [7]), .I1(\data_in[3] [7]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n29460));   // verilog/coms.v(128[12] 303[6])
    defparam i15380_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15381_3_lut (.I0(\data_in[2] [6]), .I1(\data_in[3] [6]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n29461));   // verilog/coms.v(128[12] 303[6])
    defparam i15381_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_mux_3_i20_3_lut (.I0(encoder0_position_scaled_23__N_327[19]), 
            .I1(n14_adj_5485), .I2(encoder0_position_scaled_23__N_327[31]), 
            .I3(GND_net), .O(n414));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_mux_3_i20_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i981_rep_51_3_lut (.I0(n414), 
            .I1(n1501), .I2(n1455), .I3(GND_net), .O(n1533_adj_5596));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i981_rep_51_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1048_3_lut (.I0(n1533_adj_5596), 
            .I1(n1600), .I2(n1554_adj_5597), .I3(GND_net), .O(n1632));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1048_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15382_3_lut (.I0(\data_in[2] [5]), .I1(\data_in[3] [5]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n29462));   // verilog/coms.v(128[12] 303[6])
    defparam i15382_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1115_3_lut (.I0(n1632), 
            .I1(n1699), .I2(n1653), .I3(GND_net), .O(n1731));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1115_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1182_3_lut (.I0(n1731), 
            .I1(n1798), .I2(n1752), .I3(GND_net), .O(n1830));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1182_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15383_3_lut (.I0(\data_in[2] [4]), .I1(\data_in[3] [4]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n29463));   // verilog/coms.v(128[12] 303[6])
    defparam i15383_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1249_3_lut (.I0(n1830), 
            .I1(n1897), .I2(n1851), .I3(GND_net), .O(n1929));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1249_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15384_3_lut (.I0(\data_in[2] [3]), .I1(\data_in[3] [3]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n29464));   // verilog/coms.v(128[12] 303[6])
    defparam i15384_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1316_3_lut (.I0(n1929), 
            .I1(n1996), .I2(n1950), .I3(GND_net), .O(n2028));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1316_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1383_3_lut (.I0(n2028), 
            .I1(n2095), .I2(n2049), .I3(GND_net), .O(n2127));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1383_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i906_3_lut (.I0(n1327), .I1(n1394), 
            .I2(n1356), .I3(GND_net), .O(n1426));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i906_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i22480_2_lut (.I0(n24553), .I1(dti), .I2(GND_net), .I3(GND_net), 
            .O(n36544));
    defparam i22480_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i15385_3_lut (.I0(\data_in[2] [2]), .I1(\data_in[3] [2]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n29465));   // verilog/coms.v(128[12] 303[6])
    defparam i15385_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15386_3_lut (.I0(\data_in[2] [1]), .I1(\data_in[3] [1]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n29466));   // verilog/coms.v(128[12] 303[6])
    defparam i15386_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15387_3_lut (.I0(\data_in[2] [0]), .I1(\data_in[3] [0]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n29467));   // verilog/coms.v(128[12] 303[6])
    defparam i15387_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15847_3_lut (.I0(PWMLimit[14]), .I1(\data_in_frame[9] [6]), 
            .I2(n50654), .I3(GND_net), .O(n29927));   // verilog/coms.v(128[12] 303[6])
    defparam i15847_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15388_3_lut (.I0(\data_in[1] [7]), .I1(\data_in[2] [7]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n29468));   // verilog/coms.v(128[12] 303[6])
    defparam i15388_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i22661_2_lut_2_lut (.I0(duty[19]), .I1(n296), .I2(GND_net), 
            .I3(GND_net), .O(n4910));   // verilog/TinyFPGA_B.v(123[17] 125[11])
    defparam i22661_2_lut_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i34002_3_lut (.I0(encoder0_position_scaled_23__N_327[30]), .I1(n49749), 
            .I2(encoder0_position_scaled_23__N_327[31]), .I3(GND_net), .O(n829));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam i34002_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5047_2_lut (.I0(n2_adj_5497), .I1(encoder0_position_scaled_23__N_327[31]), 
            .I2(GND_net), .I3(GND_net), .O(n621));
    defparam i5047_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i500_4_lut (.I0(n621), .I1(n8581), 
            .I2(n51996), .I3(n5_adj_5643), .O(n828));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i500_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i15389_3_lut (.I0(\data_in[1] [6]), .I1(\data_in[2] [6]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n29469));   // verilog/coms.v(128[12] 303[6])
    defparam i15389_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5585_3_lut_4_lut (.I0(commutation_state[2]), .I1(commutation_state[1]), 
            .I2(commutation_state[0]), .I3(dir), .O(GHC_N_514));   // verilog/TinyFPGA_B.v(200[7] 219[14])
    defparam i5585_3_lut_4_lut.LUT_INIT = 16'h21cc;
    SB_LUT4 i5587_3_lut_4_lut (.I0(commutation_state[2]), .I1(commutation_state[1]), 
            .I2(commutation_state[0]), .I3(dir), .O(GLC_N_523));   // verilog/TinyFPGA_B.v(200[7] 219[14])
    defparam i5587_3_lut_4_lut.LUT_INIT = 16'hcc21;
    SB_LUT4 mux_276_i1_3_lut_4_lut (.I0(n27100), .I1(control_mode[1]), .I2(motor_state_23__N_123[0]), 
            .I3(encoder0_position_scaled[0]), .O(motor_state[0]));   // verilog/TinyFPGA_B.v(283[5:22])
    defparam mux_276_i1_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 i15390_3_lut (.I0(\data_in[1] [5]), .I1(\data_in[2] [5]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n29470));   // verilog/coms.v(128[12] 303[6])
    defparam i15390_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_276_i2_3_lut_4_lut (.I0(n27100), .I1(control_mode[1]), .I2(motor_state_23__N_123[1]), 
            .I3(encoder0_position_scaled[1]), .O(motor_state[1]));   // verilog/TinyFPGA_B.v(283[5:22])
    defparam mux_276_i2_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 mux_276_i3_3_lut_4_lut (.I0(n27100), .I1(control_mode[1]), .I2(motor_state_23__N_123[2]), 
            .I3(encoder0_position_scaled[2]), .O(motor_state[2]));   // verilog/TinyFPGA_B.v(283[5:22])
    defparam mux_276_i3_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 mux_276_i4_3_lut_4_lut (.I0(n27100), .I1(control_mode[1]), .I2(motor_state_23__N_123[3]), 
            .I3(encoder0_position_scaled[3]), .O(motor_state[3]));   // verilog/TinyFPGA_B.v(283[5:22])
    defparam mux_276_i4_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 i22662_2_lut_2_lut (.I0(duty[18]), .I1(n296), .I2(GND_net), 
            .I3(GND_net), .O(n4911));   // verilog/TinyFPGA_B.v(123[17] 125[11])
    defparam i22662_2_lut_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i1_2_lut_4_lut_adj_1896 (.I0(control_mode[0]), .I1(n52298), 
            .I2(control_mode[7]), .I3(control_mode[5]), .O(n27100));   // verilog/TinyFPGA_B.v(285[5:22])
    defparam i1_2_lut_4_lut_adj_1896.LUT_INIT = 16'hfffe;
    SB_LUT4 i34031_4_lut_4_lut_4_lut (.I0(hall1), .I1(commutation_state[2]), 
            .I2(hall2), .I3(hall3), .O(n49779));
    defparam i34031_4_lut_4_lut_4_lut.LUT_INIT = 16'hd504;
    SB_LUT4 mux_276_i5_3_lut_4_lut (.I0(n27100), .I1(control_mode[1]), .I2(motor_state_23__N_123[4]), 
            .I3(encoder0_position_scaled[4]), .O(motor_state[4]));   // verilog/TinyFPGA_B.v(283[5:22])
    defparam mux_276_i5_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 mux_276_i6_3_lut_4_lut (.I0(n27100), .I1(control_mode[1]), .I2(motor_state_23__N_123[5]), 
            .I3(encoder0_position_scaled[5]), .O(motor_state[5]));   // verilog/TinyFPGA_B.v(283[5:22])
    defparam mux_276_i6_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 mux_276_i7_3_lut_4_lut (.I0(n27100), .I1(control_mode[1]), .I2(motor_state_23__N_123[6]), 
            .I3(encoder0_position_scaled[6]), .O(motor_state[6]));   // verilog/TinyFPGA_B.v(283[5:22])
    defparam mux_276_i7_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 i15391_3_lut (.I0(\data_in[1] [4]), .I1(\data_in[2] [4]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n29471));   // verilog/coms.v(128[12] 303[6])
    defparam i15391_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_17_i9_2_lut (.I0(current[4]), .I1(current_limit[4]), 
            .I2(GND_net), .I3(GND_net), .O(n9_adj_5584));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam LessThan_17_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_17_i7_2_lut (.I0(current[3]), .I1(current_limit[3]), 
            .I2(GND_net), .I3(GND_net), .O(n7_adj_5586));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam LessThan_17_i7_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mux_276_i8_3_lut_4_lut (.I0(n27100), .I1(control_mode[1]), .I2(motor_state_23__N_123[7]), 
            .I3(encoder0_position_scaled[7]), .O(motor_state[7]));   // verilog/TinyFPGA_B.v(283[5:22])
    defparam mux_276_i8_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 LessThan_17_i11_2_lut (.I0(current[5]), .I1(current_limit[5]), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_5583));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam LessThan_17_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mux_276_i9_3_lut_4_lut (.I0(n27100), .I1(control_mode[1]), .I2(motor_state_23__N_123[8]), 
            .I3(encoder0_position_scaled[8]), .O(motor_state[8]));   // verilog/TinyFPGA_B.v(283[5:22])
    defparam mux_276_i9_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 LessThan_17_i13_2_lut (.I0(current[6]), .I1(current_limit[6]), 
            .I2(GND_net), .I3(GND_net), .O(n13_adj_5582));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam LessThan_17_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mux_276_i10_3_lut_4_lut (.I0(n27100), .I1(control_mode[1]), 
            .I2(motor_state_23__N_123[9]), .I3(encoder0_position_scaled[9]), 
            .O(motor_state[9]));   // verilog/TinyFPGA_B.v(283[5:22])
    defparam mux_276_i10_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 mux_276_i11_3_lut_4_lut (.I0(n27100), .I1(control_mode[1]), 
            .I2(motor_state_23__N_123[10]), .I3(encoder0_position_scaled[10]), 
            .O(motor_state[10]));   // verilog/TinyFPGA_B.v(283[5:22])
    defparam mux_276_i11_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 mux_276_i12_3_lut_4_lut (.I0(n27100), .I1(control_mode[1]), 
            .I2(motor_state_23__N_123[11]), .I3(encoder0_position_scaled[11]), 
            .O(motor_state[11]));   // verilog/TinyFPGA_B.v(283[5:22])
    defparam mux_276_i12_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 LessThan_17_i17_2_lut (.I0(current[8]), .I1(current_limit[8]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_5560));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam LessThan_17_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mux_276_i13_3_lut_4_lut (.I0(n27100), .I1(control_mode[1]), 
            .I2(motor_state_23__N_123[12]), .I3(encoder0_position_scaled[12]), 
            .O(motor_state[12]));   // verilog/TinyFPGA_B.v(283[5:22])
    defparam mux_276_i13_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 mux_276_i14_3_lut_4_lut (.I0(n27100), .I1(control_mode[1]), 
            .I2(motor_state_23__N_123[13]), .I3(encoder0_position_scaled[13]), 
            .O(motor_state[13]));   // verilog/TinyFPGA_B.v(283[5:22])
    defparam mux_276_i14_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    \quadrature_decoder(1)  quad_counter1 (.encoder1_position({encoder1_position}), 
            .GND_net(GND_net), .b_prev(b_prev_adj_5527), .a_new({a_new_adj_5692[1], 
            Open_1}), .position_31__N_4108(position_31__N_4108_adj_5528), 
            .VCC_net(VCC_net), .ENCODER1_B_N_keep(ENCODER1_B_N), .n2269(clk16MHz), 
            .ENCODER1_A_N_keep(ENCODER1_A_N), .n29500(n29500), .n2274(n2274)) /* synthesis lattice_noprune=1 */ ;   // verilog/TinyFPGA_B.v(310[49] 316[6])
    SB_LUT4 mux_276_i15_3_lut_4_lut (.I0(n27100), .I1(control_mode[1]), 
            .I2(motor_state_23__N_123[14]), .I3(encoder0_position_scaled[14]), 
            .O(motor_state[14]));   // verilog/TinyFPGA_B.v(283[5:22])
    defparam mux_276_i15_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 mux_276_i16_3_lut_4_lut (.I0(n27100), .I1(control_mode[1]), 
            .I2(motor_state_23__N_123[15]), .I3(encoder0_position_scaled[15]), 
            .O(motor_state[15]));   // verilog/TinyFPGA_B.v(283[5:22])
    defparam mux_276_i16_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 mux_15_i1_3_lut (.I0(current[0]), .I1(n2091), .I2(n209), .I3(GND_net), 
            .O(n270));   // verilog/TinyFPGA_B.v(112[16] 114[10])
    defparam mux_15_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_276_i17_3_lut_4_lut (.I0(n27100), .I1(control_mode[1]), 
            .I2(motor_state_23__N_123[16]), .I3(encoder0_position_scaled[16]), 
            .O(motor_state[16]));   // verilog/TinyFPGA_B.v(283[5:22])
    defparam mux_276_i17_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 mux_276_i18_3_lut_4_lut (.I0(n27100), .I1(control_mode[1]), 
            .I2(motor_state_23__N_123[17]), .I3(encoder0_position_scaled[17]), 
            .O(motor_state[17]));   // verilog/TinyFPGA_B.v(283[5:22])
    defparam mux_276_i18_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 mux_276_i19_3_lut_4_lut (.I0(n27100), .I1(control_mode[1]), 
            .I2(motor_state_23__N_123[18]), .I3(encoder0_position_scaled[18]), 
            .O(motor_state[18]));   // verilog/TinyFPGA_B.v(283[5:22])
    defparam mux_276_i19_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 mux_276_i20_3_lut_4_lut (.I0(n27100), .I1(control_mode[1]), 
            .I2(motor_state_23__N_123[19]), .I3(encoder0_position_scaled[19]), 
            .O(motor_state[19]));   // verilog/TinyFPGA_B.v(283[5:22])
    defparam mux_276_i20_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 mux_276_i21_3_lut_4_lut (.I0(n27100), .I1(control_mode[1]), 
            .I2(motor_state_23__N_123[20]), .I3(encoder0_position_scaled[20]), 
            .O(motor_state[20]));   // verilog/TinyFPGA_B.v(283[5:22])
    defparam mux_276_i21_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 i15421_3_lut_4_lut (.I0(n2233), .I1(b_prev), .I2(a_new[1]), 
            .I3(position_31__N_4108), .O(n29501));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    defparam i15421_3_lut_4_lut.LUT_INIT = 16'h3caa;
    SB_LUT4 i15444_3_lut (.I0(deadband[21]), .I1(\data_in_frame[14] [5]), 
            .I2(n50654), .I3(GND_net), .O(n29524));   // verilog/coms.v(128[12] 303[6])
    defparam i15444_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15420_3_lut_4_lut (.I0(n2274), .I1(b_prev_adj_5527), .I2(a_new_adj_5692[1]), 
            .I3(position_31__N_4108_adj_5528), .O(n29500));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    defparam i15420_3_lut_4_lut.LUT_INIT = 16'h3caa;
    SB_LUT4 i15445_3_lut (.I0(deadband[20]), .I1(\data_in_frame[14] [4]), 
            .I2(n50654), .I3(GND_net), .O(n29525));   // verilog/coms.v(128[12] 303[6])
    defparam i15445_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15446_3_lut (.I0(deadband[19]), .I1(\data_in_frame[14] [3]), 
            .I2(n50654), .I3(GND_net), .O(n29526));   // verilog/coms.v(128[12] 303[6])
    defparam i15446_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15447_3_lut (.I0(deadband[18]), .I1(\data_in_frame[14] [2]), 
            .I2(n50654), .I3(GND_net), .O(n29527));   // verilog/coms.v(128[12] 303[6])
    defparam i15447_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_276_i22_3_lut_4_lut (.I0(n27100), .I1(control_mode[1]), 
            .I2(motor_state_23__N_123[21]), .I3(encoder0_position_scaled[21]), 
            .O(motor_state[21]));   // verilog/TinyFPGA_B.v(283[5:22])
    defparam mux_276_i22_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 i15448_4_lut (.I0(r_Rx_Data), .I1(rx_data[6]), .I2(n36556), 
            .I3(n27208), .O(n29528));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i15448_4_lut.LUT_INIT = 16'hccac;
    SB_LUT4 i15449_3_lut (.I0(deadband[17]), .I1(\data_in_frame[14] [1]), 
            .I2(n50654), .I3(GND_net), .O(n29529));   // verilog/coms.v(128[12] 303[6])
    defparam i15449_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15272_3_lut (.I0(ID[0]), .I1(data[0]), .I2(n51509), .I3(GND_net), 
            .O(n29352));   // verilog/TinyFPGA_B.v(368[10] 396[6])
    defparam i15272_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15450_3_lut (.I0(deadband[16]), .I1(\data_in_frame[14] [0]), 
            .I2(n50654), .I3(GND_net), .O(n29530));   // verilog/coms.v(128[12] 303[6])
    defparam i15450_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i3_4_lut_4_lut (.I0(r_SM_Main_adj_5723[2]), .I1(r_SM_Main_adj_5723[0]), 
            .I2(r_SM_Main_adj_5723[1]), .I3(r_SM_Main_2__N_3848[1]), .O(n57032));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i3_4_lut_4_lut.LUT_INIT = 16'h4000;
    SB_LUT4 i15392_3_lut (.I0(\data_in[1] [3]), .I1(\data_in[2] [3]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n29472));   // verilog/coms.v(128[12] 303[6])
    defparam i15392_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_276_i23_3_lut_4_lut (.I0(n27100), .I1(control_mode[1]), 
            .I2(motor_state_23__N_123[22]), .I3(encoder0_position_scaled[22]), 
            .O(motor_state[22]));   // verilog/TinyFPGA_B.v(283[5:22])
    defparam mux_276_i23_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 i15451_3_lut (.I0(deadband[15]), .I1(\data_in_frame[15] [7]), 
            .I2(n50654), .I3(GND_net), .O(n29531));   // verilog/coms.v(128[12] 303[6])
    defparam i15451_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15452_3_lut (.I0(deadband[14]), .I1(\data_in_frame[15] [6]), 
            .I2(n50654), .I3(GND_net), .O(n29532));   // verilog/coms.v(128[12] 303[6])
    defparam i15452_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_276_i24_3_lut_4_lut (.I0(n27100), .I1(control_mode[1]), 
            .I2(motor_state_23__N_123[23]), .I3(encoder0_position_scaled[23]), 
            .O(motor_state[23]));   // verilog/TinyFPGA_B.v(283[5:22])
    defparam mux_276_i24_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 i15453_3_lut (.I0(deadband[13]), .I1(\data_in_frame[15] [5]), 
            .I2(n50654), .I3(GND_net), .O(n29533));   // verilog/coms.v(128[12] 303[6])
    defparam i15453_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 n56616_bdd_4_lut (.I0(n56616), .I1(duty[0]), .I2(n270), .I3(duty[23]), 
            .O(pwm_setpoint_23__N_11[0]));
    defparam n56616_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i15454_3_lut (.I0(deadband[12]), .I1(\data_in_frame[15] [4]), 
            .I2(n50654), .I3(GND_net), .O(n29534));   // verilog/coms.v(128[12] 303[6])
    defparam i15454_3_lut.LUT_INIT = 16'hacac;
    coms neopxl_color_23__I_0 (.n29523(n29523), .deadband({deadband}), .clk16MHz(clk16MHz), 
         .n29522(n29522), .n29521(n29521), .\Kp[1] (Kp[1]), .n29520(n29520), 
         .\Kp[2] (Kp[2]), .n29519(n29519), .\Kp[3] (Kp[3]), .n29518(n29518), 
         .\Kp[4] (Kp[4]), .GND_net(GND_net), .\data_in_frame[3] ({\data_in_frame[3] }), 
         .n63(n63), .n3303(n3303), .n27219(n27219), .n48947(n48947), 
         .n48957(n48957), .\data_out_frame[16] ({\data_out_frame[16] }), 
         .\data_out_frame[17] ({\data_out_frame[17] }), .\data_out_frame[18] ({\data_out_frame[18] }), 
         .\data_out_frame[19] ({\data_out_frame[19] }), .n27218(n27218), 
         .\FRAME_MATCHER.state[3] (\FRAME_MATCHER.state [3]), .\data_out_frame[22] ({\data_out_frame[22] }), 
         .\data_out_frame[23] ({\data_out_frame[23] }), .\data_out_frame[20] ({\data_out_frame[20] }), 
         .\data_out_frame[21] ({\data_out_frame[21] }), .\data_in_frame[2] ({\data_in_frame[2] }), 
         .rx_data_ready(rx_data_ready), .n22875(n22875), .\data_out_frame[6] ({\data_out_frame[6] }), 
         .\data_out_frame[7] ({\data_out_frame[7] }), .\data_out_frame[4] ({\data_out_frame[4] }), 
         .\data_out_frame[5] ({\data_out_frame[5] }), .n29516(n29516), .\Kp[5] (Kp[5]), 
         .\data_in_frame[4] ({\data_in_frame[4] }), .\data_in_frame[5] ({\data_in_frame[5] }), 
         .PWMLimit({PWMLimit}), .n50654(n50654), .\data_in[0] ({\data_in[0] }), 
         .\data_in[1] ({\data_in[1] }), .\data_in[2] ({\data_in[2] }), .\data_in[3] ({\data_in[3] }), 
         .n29515(n29515), .\Kp[6] (Kp[6]), .n63_adj_6(n63_adj_5605), .n29514(n29514), 
         .\Kp[7] (Kp[7]), .rx_data({rx_data}), .n122(n122), .n8(n8_adj_5609), 
         .n7(n7_adj_5608), .\data_in_frame[1] ({\data_in_frame[1] }), .\data_in_frame[8] ({\data_in_frame[8] [7], 
         Open_2, Open_3, Open_4, \data_in_frame[8] [3], Open_5, Open_6, 
         \data_in_frame[8] [0]}), .ID({ID}), .\data_out_frame[8] ({\data_out_frame[8] }), 
         .\data_out_frame[9] ({\data_out_frame[9] }), .\data_out_frame[10] ({\data_out_frame[10] }), 
         .\data_out_frame[11] ({\data_out_frame[11] }), .\data_out_frame[14] ({\data_out_frame[14] }), 
         .\data_out_frame[15] ({\data_out_frame[15] }), .\data_out_frame[12] ({\data_out_frame[12] }), 
         .\data_out_frame[13] ({\data_out_frame[13] }), .tx_active(tx_active), 
         .\data_in_frame[13] ({\data_in_frame[13] }), .\data_in_frame[15] ({\data_in_frame[15] }), 
         .\FRAME_MATCHER.state[0] (\FRAME_MATCHER.state [0]), .n29513(n29513), 
         .\Kp[8] (Kp[8]), .n29512(n29512), .\Kp[9] (Kp[9]), .setpoint({setpoint}), 
         .n19602(n19602), .\data_in_frame[8][2] (\data_in_frame[8] [2]), 
         .n29511(n29511), .\Kp[10] (Kp[10]), .\data_in_frame[9] ({\data_in_frame[9] }), 
         .n29510(n29510), .\Kp[11] (Kp[11]), .n29509(n29509), .\Kp[12] (Kp[12]), 
         .\data_in_frame[10][2] (\data_in_frame[10] [2]), .n29508(n29508), 
         .\Kp[13] (Kp[13]), .n29507(n29507), .\Kp[14] (Kp[14]), .n363(n363), 
         .n32464(n32464), .\data_in_frame[12] ({\data_in_frame[12] }), .\data_in_frame[10][1] (\data_in_frame[10] [1]), 
         .n29506(n29506), .\Kp[15] (Kp[15]), .\data_in_frame[16] ({\data_in_frame[16] }), 
         .n29505(n29505), .\Ki[1] (Ki[1]), .n29504(n29504), .\Ki[2] (Ki[2]), 
         .n29503(n29503), .\Ki[3] (Ki[3]), .n29502(n29502), .\Ki[4] (Ki[4]), 
         .n29499(n29499), .\Ki[5] (Ki[5]), .n29498(n29498), .\Ki[6] (Ki[6]), 
         .n29497(n29497), .\Ki[7] (Ki[7]), .n29496(n29496), .\Ki[8] (Ki[8]), 
         .n29495(n29495), .\Ki[9] (Ki[9]), .n29494(n29494), .\Ki[10] (Ki[10]), 
         .n29493(n29493), .\Ki[11] (Ki[11]), .n29492(n29492), .\Ki[12] (Ki[12]), 
         .n29491(n29491), .\Ki[13] (Ki[13]), .n29490(n29490), .\Ki[14] (Ki[14]), 
         .n29486(n29486), .\Ki[15] (Ki[15]), .n29485(n29485), .n29484(n29484), 
         .n29483(n29483), .n29482(n29482), .n29481(n29481), .n29480(n29480), 
         .n29479(n29479), .n29478(n29478), .n29477(n29477), .n29476(n29476), 
         .\data_in_frame[14] ({\data_in_frame[14] }), .n29472(n29472), .n4(n4_adj_5472), 
         .n29471(n29471), .\data_in_frame[8][6] (\data_in_frame[8] [6]), 
         .\data_in_frame[11] ({\data_in_frame[11] }), .n29470(n29470), .n29469(n29469), 
         .DE_c(DE_c), .n29468(n29468), .n29467(n29467), .n29466(n29466), 
         .n29465(n29465), .n29464(n29464), .n29463(n29463), .n29462(n29462), 
         .n29461(n29461), .n29460(n29460), .n29456(n29456), .n29455(n29455), 
         .n29454(n29454), .n29453(n29453), .n29451(n29451), .\data_out_frame[25] ({\data_out_frame[25] }), 
         .n29450(n29450), .\data_in_frame[21] ({\data_in_frame[21] }), .\data_in_frame[20] ({\data_in_frame[20] }), 
         .n29449(n29449), .n29448(n29448), .n29447(n29447), .n29446(n29446), 
         .n29445(n29445), .n29444(n29444), .n29443(n29443), .n29442(n29442), 
         .n29441(n29441), .n29440(n29440), .n29439(n29439), .n29438(n29438), 
         .n29437(n29437), .n29436(n29436), .n29435(n29435), .n29434(n29434), 
         .n29433(n29433), .n29432(n29432), .n29431(n29431), .n29430(n29430), 
         .n29429(n29429), .n29428(n29428), .n29427(n29427), .n29426(n29426), 
         .n29425(n29425), .n29424(n29424), .n29423(n29423), .n29422(n29422), 
         .n29421(n29421), .n29420(n29420), .n29419(n29419), .\data_out_frame[24] ({\data_out_frame[24] }), 
         .\data_in_frame[8][4] (\data_in_frame[8] [4]), .\data_in_frame[8][5] (\data_in_frame[8] [5]), 
         .n29418(n29418), .n30058(n30058), .n30057(n30057), .n30056(n30056), 
         .n30055(n30055), .n30054(n30054), .n30053(n30053), .n30052(n30052), 
         .n30051(n30051), .n30050(n30050), .n30049(n30049), .n30048(n30048), 
         .n30047(n30047), .n30046(n30046), .n30045(n30045), .n30044(n30044), 
         .n30043(n30043), .n30042(n30042), .n30041(n30041), .n30040(n30040), 
         .n30039(n30039), .n30038(n30038), .n30037(n30037), .n30036(n30036), 
         .n30035(n30035), .n30034(n30034), .n30033(n30033), .n30032(n30032), 
         .n30031(n30031), .n30030(n30030), .n30029(n30029), .n30028(n30028), 
         .n30027(n30027), .n30026(n30026), .n30025(n30025), .n30024(n30024), 
         .n30023(n30023), .n30022(n30022), .n30021(n30021), .n30020(n30020), 
         .n30019(n30019), .n30018(n30018), .n30017(n30017), .n30016(n30016), 
         .n30015(n30015), .n30014(n30014), .n30013(n30013), .n30012(n30012), 
         .n30011(n30011), .n30010(n30010), .n30009(n30009), .n30008(n30008), 
         .n30007(n30007), .n30006(n30006), .n30005(n30005), .n30004(n30004), 
         .n30003(n30003), .n30002(n30002), .n30001(n30001), .n30000(n30000), 
         .n29999(n29999), .n29998(n29998), .n29997(n29997), .n29996(n29996), 
         .n29995(n29995), .n29994(n29994), .n29993(n29993), .n29992(n29992), 
         .n29991(n29991), .n29990(n29990), .n29989(n29989), .n29988(n29988), 
         .n29987(n29987), .n29986(n29986), .n29985(n29985), .n29984(n29984), 
         .n29983(n29983), .n29982(n29982), .n29981(n29981), .n29980(n29980), 
         .n29979(n29979), .n29978(n29978), .n29977(n29977), .n29976(n29976), 
         .n29417(n29417), .n29416(n29416), .n29415(n29415), .n29414(n29414), 
         .n29412(n29412), .n29411(n29411), .n29410(n29410), .n29408(n29408), 
         .n29406(n29406), .n29405(n29405), .n29404(n29404), .n29403(n29403), 
         .n29402(n29402), .n29401(n29401), .n29400(n29400), .n29397(n29397), 
         .n29396(n29396), .n29395(n29395), .n29394(n29394), .LED_c(LED_c), 
         .n29975(n29975), .n29974(n29974), .n29973(n29973), .n29972(n29972), 
         .n29971(n29971), .n29970(n29970), .n29969(n29969), .n29968(n29968), 
         .n29967(n29967), .n29962(n29962), .control_mode({control_mode}), 
         .n29961(n29961), .n29960(n29960), .n29959(n29959), .n29958(n29958), 
         .n29957(n29957), .n29956(n29956), .n29955(n29955), .current_limit({current_limit}), 
         .n29954(n29954), .n29953(n29953), .n29952(n29952), .n29951(n29951), 
         .n29950(n29950), .n29949(n29949), .n29948(n29948), .n29947(n29947), 
         .n29946(n29946), .n29945(n29945), .n29944(n29944), .n29943(n29943), 
         .n29942(n29942), .n29941(n29941), .n29940(n29940), .n29939(n29939), 
         .n29390(n29390), .n29938(n29938), .n29389(n29389), .n29937(n29937), 
         .n29936(n29936), .n29935(n29935), .n29934(n29934), .n29388(n29388), 
         .n29387(n29387), .n29386(n29386), .n29385(n29385), .n29384(n29384), 
         .n29383(n29383), .n29382(n29382), .n29380(n29380), .n29379(n29379), 
         .n29378(n29378), .n50741(n50741), .n29375(n29375), .n29374(n29374), 
         .neopxl_color({neopxl_color}), .n29371(n29371), .n29370(n29370), 
         .\Ki[0] (Ki[0]), .n29369(n29369), .\Kp[0] (Kp[0]), .n29368(n29368), 
         .IntegralLimit({IntegralLimit}), .n29933(n29933), .n29932(n29932), 
         .n29931(n29931), .n29930(n29930), .n29929(n29929), .n29928(n29928), 
         .n29927(n29927), .n29926(n29926), .n6(n6_adj_5645), .n29925(n29925), 
         .n29923(n29923), .n29922(n29922), .n29356(n29356), .n29355(n29355), 
         .n29921(n29921), .n29920(n29920), .n29919(n29919), .n29918(n29918), 
         .n57033(n57033), .n29353(n29353), .n29874(n29874), .n29873(n29873), 
         .n29872(n29872), .n29870(n29870), .n29868(n29868), .n29867(n29867), 
         .n29866(n29866), .n29865(n29865), .n29864(n29864), .n29863(n29863), 
         .n29862(n29862), .n29861(n29861), .n29834(n29834), .n29833(n29833), 
         .n29832(n29832), .n29831(n29831), .n29830(n29830), .n29827(n29827), 
         .n29826(n29826), .n29825(n29825), .n29824(n29824), .\data_in_frame[10][3] (\data_in_frame[10] [3]), 
         .\data_in_frame[10][4] (\data_in_frame[10] [4]), .\data_in_frame[10][5] (\data_in_frame[10] [5]), 
         .\data_in_frame[10][6] (\data_in_frame[10] [6]), .\data_in_frame[10][7] (\data_in_frame[10] [7]), 
         .n29571(n29571), .n29570(n29570), .n29569(n29569), .n29568(n29568), 
         .n29567(n29567), .n29566(n29566), .n29565(n29565), .n29564(n29564), 
         .n29563(n29563), .n29562(n29562), .n29561(n29561), .n29560(n29560), 
         .n29559(n29559), .n29558(n29558), .n29557(n29557), .n29556(n29556), 
         .n29555(n29555), .n29554(n29554), .n29553(n29553), .n29552(n29552), 
         .n29551(n29551), .n29550(n29550), .n29549(n29549), .n29546(n29546), 
         .n29545(n29545), .n29544(n29544), .n29543(n29543), .n29542(n29542), 
         .n29541(n29541), .n29540(n29540), .n29539(n29539), .n29538(n29538), 
         .n29537(n29537), .n29536(n29536), .n29534(n29534), .n29533(n29533), 
         .n29532(n29532), .n29531(n29531), .n29530(n29530), .n29529(n29529), 
         .n29527(n29527), .n29526(n29526), .n29525(n29525), .n29524(n29524), 
         .n24210(n24210), .\state[0] (state_adj_5736[0]), .\state[2] (state_adj_5736[2]), 
         .\state[3] (state_adj_5736[3]), .n7936(n7936), .\FRAME_MATCHER.state_31__N_3007[2] (\FRAME_MATCHER.state_31__N_3007 [2]), 
         .n28848(n28848), .n29280(n29280), .r_SM_Main({r_SM_Main_adj_5723}), 
         .\r_SM_Main_2__N_3848[1] (r_SM_Main_2__N_3848[1]), .\r_Bit_Index[0] (r_Bit_Index_adj_5725[0]), 
         .VCC_net(VCC_net), .tx_o(tx_o), .n19728(n19728), .n29842(n29842), 
         .n29413(n29413), .n57032(n57032), .n4_adj_7(n4_adj_5644), .tx_enable(tx_enable), 
         .r_SM_Main_adj_15({r_SM_Main}), .\r_SM_Main_2__N_3777[2] (r_SM_Main_2__N_3777[2]), 
         .r_Rx_Data(r_Rx_Data), .n28852(n28852), .n29282(n29282), .RX_N_10(RX_N_10), 
         .\r_Bit_Index[0]_adj_11 (r_Bit_Index[0]), .n4_adj_12(n4_adj_5443), 
         .n36556(n36556), .n4_adj_13(n4_adj_5469), .n4_adj_14(n4_adj_5445), 
         .n29845(n29845), .n48522(n48522), .n48878(n48878), .n29880(n29880), 
         .n29878(n29878), .n29877(n29877), .n29871(n29871), .n29860(n29860), 
         .n29849(n29849), .n29759(n29759), .n29528(n29528), .n27208(n27208), 
         .n27203(n27203)) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(254[8] 278[4])
    SB_LUT4 i15456_3_lut (.I0(deadband[11]), .I1(\data_in_frame[15] [3]), 
            .I2(n50654), .I3(GND_net), .O(n29536));   // verilog/coms.v(128[12] 303[6])
    defparam i15456_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15457_3_lut (.I0(deadband[10]), .I1(\data_in_frame[15] [2]), 
            .I2(n50654), .I3(GND_net), .O(n29537));   // verilog/coms.v(128[12] 303[6])
    defparam i15457_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15458_3_lut (.I0(deadband[9]), .I1(\data_in_frame[15] [1]), 
            .I2(n50654), .I3(GND_net), .O(n29538));   // verilog/coms.v(128[12] 303[6])
    defparam i15458_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15459_3_lut (.I0(deadband[8]), .I1(\data_in_frame[15] [0]), 
            .I2(n50654), .I3(GND_net), .O(n29539));   // verilog/coms.v(128[12] 303[6])
    defparam i15459_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15460_3_lut (.I0(deadband[7]), .I1(\data_in_frame[16] [7]), 
            .I2(n50654), .I3(GND_net), .O(n29540));   // verilog/coms.v(128[12] 303[6])
    defparam i15460_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i22663_2_lut_2_lut (.I0(duty[17]), .I1(n296), .I2(GND_net), 
            .I3(GND_net), .O(n4912));   // verilog/TinyFPGA_B.v(123[17] 125[11])
    defparam i22663_2_lut_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i15461_3_lut (.I0(deadband[6]), .I1(\data_in_frame[16] [6]), 
            .I2(n50654), .I3(GND_net), .O(n29541));   // verilog/coms.v(128[12] 303[6])
    defparam i15461_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15462_3_lut (.I0(deadband[5]), .I1(\data_in_frame[16] [5]), 
            .I2(n50654), .I3(GND_net), .O(n29542));   // verilog/coms.v(128[12] 303[6])
    defparam i15462_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15463_3_lut (.I0(deadband[4]), .I1(\data_in_frame[16] [4]), 
            .I2(n50654), .I3(GND_net), .O(n29543));   // verilog/coms.v(128[12] 303[6])
    defparam i15463_3_lut.LUT_INIT = 16'hacac;
    pwm PWM (.pwm_out(pwm_out), .clk32MHz(clk32MHz), .GND_net(GND_net), 
        .VCC_net(VCC_net), .pwm_setpoint({pwm_setpoint})) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(96[6] 101[3])
    SB_LUT4 i15464_3_lut (.I0(deadband[3]), .I1(\data_in_frame[16] [3]), 
            .I2(n50654), .I3(GND_net), .O(n29544));   // verilog/coms.v(128[12] 303[6])
    defparam i15464_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15465_3_lut (.I0(deadband[2]), .I1(\data_in_frame[16] [2]), 
            .I2(n50654), .I3(GND_net), .O(n29545));   // verilog/coms.v(128[12] 303[6])
    defparam i15465_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15466_3_lut (.I0(deadband[1]), .I1(\data_in_frame[16] [1]), 
            .I2(n50654), .I3(GND_net), .O(n29546));   // verilog/coms.v(128[12] 303[6])
    defparam i15466_3_lut.LUT_INIT = 16'hacac;
    TLI4970 tli (.\state[0] (state_adj_5713[0]), .GND_net(GND_net), .\data[12] (data_adj_5711[12]), 
            .n5(n5_adj_5557), .\state[1] (state_adj_5713[1]), .\data[15] (data_adj_5711[15]), 
            .n28729(n28729), .clk16MHz(clk16MHz), .VCC_net(VCC_net), .n15(n15_adj_5470), 
            .n5_adj_1(n5), .n36554(n36554), .n36528(n36528), .n6(n6_adj_5523), 
            .n30067(n30067), .n30066(n30066), .\data[11] (data_adj_5711[11]), 
            .n30059(n30059), .\data[10] (data_adj_5711[10]), .n29407(n29407), 
            .n9(n9_adj_5601), .clk_out(clk_out), .n29398(n29398), .CS_c(CS_c), 
            .n29391(n29391), .\current[0] (current[0]), .\current[15] (current[15]), 
            .n7(n7_adj_5577), .n29916(n29916), .\data[9] (data_adj_5711[9]), 
            .n29892(n29892), .\data[8] (data_adj_5711[8]), .n29891(n29891), 
            .\current[1] (current[1]), .n29890(n29890), .\current[2] (current[2]), 
            .n29889(n29889), .\current[3] (current[3]), .n29888(n29888), 
            .\current[4] (current[4]), .n29887(n29887), .\current[5] (current[5]), 
            .n29886(n29886), .\current[6] (current[6]), .n29885(n29885), 
            .\current[7] (current[7]), .n29884(n29884), .\current[8] (current[8]), 
            .n29883(n29883), .\current[9] (current[9]), .n29882(n29882), 
            .\current[10] (current[10]), .n29881(n29881), .\current[11] (current[11]), 
            .n29879(n29879), .\data[7] (data_adj_5711[7]), .n29876(n29876), 
            .\data[6] (data_adj_5711[6]), .n29869(n29869), .\data[5] (data_adj_5711[5]), 
            .n29850(n29850), .\data[0] (data_adj_5711[0]), .n29839(n29839), 
            .\data[4] (data_adj_5711[4]), .n29838(n29838), .\data[3] (data_adj_5711[3]), 
            .n29823(n29823), .\data[2] (data_adj_5711[2]), .n29758(n29758), 
            .\data[1] (data_adj_5711[1]), .CS_CLK_c(CS_CLK_c), .n27258(n27258), 
            .n27271(n27271), .n27232(n27232), .n27198(n27198), .n6_adj_2(n6_adj_5556), 
            .n5_adj_3(n5_adj_5524), .n27264(n27264), .state_7__N_4499(state_7__N_4499)) /* synthesis syn_noprune=1, syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(411[11] 417[4])
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1777_3_lut (.I0(n2614), 
            .I1(n2681), .I2(n2643), .I3(GND_net), .O(n2713));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1777_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15469_3_lut (.I0(IntegralLimit[23]), .I1(\data_in_frame[11] [7]), 
            .I2(n50654), .I3(GND_net), .O(n29549));   // verilog/coms.v(128[12] 303[6])
    defparam i15469_3_lut.LUT_INIT = 16'hacac;
    
endmodule
//
// Verilog Description of module \neopixel(CLOCK_SPEED_HZ=16000000) 
//

module \neopixel(CLOCK_SPEED_HZ=16000000)  (clk16MHz, \state[0] , \state[1] , 
            GND_net, \neo_pixel_transmitter.t0 , n28778, \state_3__N_639[1] , 
            neopxl_color, timer, VCC_net, LED_c, n29354, n29829, 
            n29814, n29813, n29812, n29811, n29810, n29809, n29808, 
            n29807, n29806, n29805, n29804, n29803, n29802, n29801, 
            n29800, n29799, n29798, n29797, n29796, n29795, n29794, 
            n29793, n29792, n29791, n29790, n29789, n29788, n29785, 
            n29784, n29783, n29782, NEOPXL_c, n47790) /* synthesis syn_module_defined=1 */ ;
    input clk16MHz;
    output \state[0] ;
    output \state[1] ;
    input GND_net;
    output [31:0]\neo_pixel_transmitter.t0 ;
    output n28778;
    output \state_3__N_639[1] ;
    input [23:0]neopxl_color;
    output [31:0]timer;
    input VCC_net;
    input LED_c;
    input n29354;
    input n29829;
    input n29814;
    input n29813;
    input n29812;
    input n29811;
    input n29810;
    input n29809;
    input n29808;
    input n29807;
    input n29806;
    input n29805;
    input n29804;
    input n29803;
    input n29802;
    input n29801;
    input n29800;
    input n29799;
    input n29798;
    input n29797;
    input n29796;
    input n29795;
    input n29794;
    input n29793;
    input n29792;
    input n29791;
    input n29790;
    input n29789;
    input n29788;
    input n29785;
    input n29784;
    input n29783;
    input n29782;
    output NEOPXL_c;
    output n47790;
    
    wire clk16MHz /* synthesis SET_AS_NETWORK=clk16MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    
    wire \neo_pixel_transmitter.done_N_847 , n56981, \neo_pixel_transmitter.done , 
        start_N_838, n7, start, n45295, n49822, n55119, n54536, 
        n37356, n27111, n49937, n55120, n49955, \neo_pixel_transmitter.done_N_853 ;
    wire [31:0]bit_ctr;   // verilog/neopixel.v(18[12:19])
    wire [31:0]color_bit_N_833;
    wire [31:0]n133;
    
    wire n7792, n29197;
    wire [31:0]n1;
    
    wire n51332, n49892, n27251, n56643, n56949, n55504, n37163, 
        n45911, n56853, n55564, n56793, n54600;
    wire [3:0]state_3__N_639;
    
    wire n53312, n53313, n53304, n53303, n56946;
    wire [31:0]n133_adj_5442;
    
    wire n53210, n53211, n56850, n53205, n53204, n44509, n44508, 
        n44507, n44506, n44505, n44504, n44503, n44502, n44501, 
        n27299, n43609, n52818, n44500, n44499, n44498, n43608, 
        n52816, n43607, n52814, n44497, n44496, n44495, n44494, 
        n43606, n52812, n44493, n44492, n44491, n44490, n44489, 
        n44488, n44487, n44486, n43605, n52810, n43604, n52808, 
        n44485, n44484, n44483, n44482, n44481, n43603, n52806, 
        n44480, n44479, n44478, n44477, n43602, n52804, n44476, 
        n56790, n44475, n29172, n44474, n44473, n44472, n44471, 
        n44470, n44469, n44468, n30, n48, n46, n47, n44467, 
        n44466, n44465, n45, n44, n43, n54, n49, n44464, n44463, 
        n2586, n44462, n44461, n44460, n44459, n44458, n44457, 
        n44456, n44455, n44454, n43601, n52802, n54532, n6_adj_5437, 
        n44453, n44452, n44451, n44450, n54542, n44449, n43600, 
        n52800, n44448, n43599, n52798, n43598, n52796, n43597, 
        n52794, n43596, n52792, n43595, n52790, n43594, n52788, 
        n43593, n52786, n43592, n52784, n43591, n52782, n43590;
    wire [31:0]one_wire_N_790;
    
    wire n43589, n43588, n43587, n43586, n43585, n43584, n43583, 
        n43582, n43581, n43580, n43579, n56640, n51489, n49935, 
        n7_adj_5439, n52822, n52828, n54545, n49746, n49818, n48982, 
        n103, n16_adj_5440, n6_adj_5441;
    
    SB_DFFE \neo_pixel_transmitter.done_104  (.Q(\neo_pixel_transmitter.done ), 
            .C(clk16MHz), .E(n56981), .D(\neo_pixel_transmitter.done_N_847 ));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFE start_103 (.Q(start), .C(clk16MHz), .E(n7), .D(start_N_838));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 i39606_4_lut (.I0(n45295), .I1(n49822), .I2(\neo_pixel_transmitter.done ), 
            .I3(\state[0] ), .O(n55119));
    defparam i39606_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i53_4_lut (.I0(n54536), .I1(n37356), .I2(\state[1] ), .I3(n27111), 
            .O(n49937));
    defparam i53_4_lut.LUT_INIT = 16'hcfca;
    SB_LUT4 i52_4_lut (.I0(n49937), .I1(n55120), .I2(\state[0] ), .I3(\neo_pixel_transmitter.done ), 
            .O(n49955));
    defparam i52_4_lut.LUT_INIT = 16'h3335;
    SB_LUT4 i3_1_lut (.I0(\neo_pixel_transmitter.done ), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(\neo_pixel_transmitter.done_N_853 ));   // verilog/neopixel.v(35[12] 117[6])
    defparam i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_2_lut (.I0(bit_ctr[1]), .I1(bit_ctr[0]), .I2(GND_net), 
            .I3(GND_net), .O(color_bit_N_833[1]));
    defparam i1_2_lut.LUT_INIT = 16'h6666;
    SB_DFFESR bit_ctr_2281__i0 (.Q(bit_ctr[0]), .C(clk16MHz), .E(n7792), 
            .D(n133[0]), .R(n29197));   // verilog/neopixel.v(69[23:32])
    SB_DFFESR bit_ctr_2281__i1 (.Q(bit_ctr[1]), .C(clk16MHz), .E(n7792), 
            .D(n133[1]), .R(n29197));   // verilog/neopixel.v(69[23:32])
    SB_DFFESR bit_ctr_2281__i2 (.Q(bit_ctr[2]), .C(clk16MHz), .E(n7792), 
            .D(n133[2]), .R(n29197));   // verilog/neopixel.v(69[23:32])
    SB_DFFESR bit_ctr_2281__i3 (.Q(bit_ctr[3]), .C(clk16MHz), .E(n7792), 
            .D(n133[3]), .R(n29197));   // verilog/neopixel.v(69[23:32])
    SB_DFFESR bit_ctr_2281__i4 (.Q(bit_ctr[4]), .C(clk16MHz), .E(n7792), 
            .D(n133[4]), .R(n29197));   // verilog/neopixel.v(69[23:32])
    SB_DFFESR bit_ctr_2281__i5 (.Q(bit_ctr[5]), .C(clk16MHz), .E(n7792), 
            .D(n133[5]), .R(n29197));   // verilog/neopixel.v(69[23:32])
    SB_DFFESR bit_ctr_2281__i6 (.Q(bit_ctr[6]), .C(clk16MHz), .E(n7792), 
            .D(n133[6]), .R(n29197));   // verilog/neopixel.v(69[23:32])
    SB_DFFESR bit_ctr_2281__i7 (.Q(bit_ctr[7]), .C(clk16MHz), .E(n7792), 
            .D(n133[7]), .R(n29197));   // verilog/neopixel.v(69[23:32])
    SB_DFFESR bit_ctr_2281__i8 (.Q(bit_ctr[8]), .C(clk16MHz), .E(n7792), 
            .D(n133[8]), .R(n29197));   // verilog/neopixel.v(69[23:32])
    SB_DFFESR bit_ctr_2281__i9 (.Q(bit_ctr[9]), .C(clk16MHz), .E(n7792), 
            .D(n133[9]), .R(n29197));   // verilog/neopixel.v(69[23:32])
    SB_DFFESR bit_ctr_2281__i10 (.Q(bit_ctr[10]), .C(clk16MHz), .E(n7792), 
            .D(n133[10]), .R(n29197));   // verilog/neopixel.v(69[23:32])
    SB_DFFESR bit_ctr_2281__i11 (.Q(bit_ctr[11]), .C(clk16MHz), .E(n7792), 
            .D(n133[11]), .R(n29197));   // verilog/neopixel.v(69[23:32])
    SB_DFFESR bit_ctr_2281__i12 (.Q(bit_ctr[12]), .C(clk16MHz), .E(n7792), 
            .D(n133[12]), .R(n29197));   // verilog/neopixel.v(69[23:32])
    SB_DFFESR bit_ctr_2281__i13 (.Q(bit_ctr[13]), .C(clk16MHz), .E(n7792), 
            .D(n133[13]), .R(n29197));   // verilog/neopixel.v(69[23:32])
    SB_DFFESR bit_ctr_2281__i14 (.Q(bit_ctr[14]), .C(clk16MHz), .E(n7792), 
            .D(n133[14]), .R(n29197));   // verilog/neopixel.v(69[23:32])
    SB_DFFESR bit_ctr_2281__i15 (.Q(bit_ctr[15]), .C(clk16MHz), .E(n7792), 
            .D(n133[15]), .R(n29197));   // verilog/neopixel.v(69[23:32])
    SB_DFFESR bit_ctr_2281__i16 (.Q(bit_ctr[16]), .C(clk16MHz), .E(n7792), 
            .D(n133[16]), .R(n29197));   // verilog/neopixel.v(69[23:32])
    SB_DFFESR bit_ctr_2281__i17 (.Q(bit_ctr[17]), .C(clk16MHz), .E(n7792), 
            .D(n133[17]), .R(n29197));   // verilog/neopixel.v(69[23:32])
    SB_DFFESR bit_ctr_2281__i18 (.Q(bit_ctr[18]), .C(clk16MHz), .E(n7792), 
            .D(n133[18]), .R(n29197));   // verilog/neopixel.v(69[23:32])
    SB_DFFESR bit_ctr_2281__i19 (.Q(bit_ctr[19]), .C(clk16MHz), .E(n7792), 
            .D(n133[19]), .R(n29197));   // verilog/neopixel.v(69[23:32])
    SB_DFFESR bit_ctr_2281__i20 (.Q(bit_ctr[20]), .C(clk16MHz), .E(n7792), 
            .D(n133[20]), .R(n29197));   // verilog/neopixel.v(69[23:32])
    SB_DFFESR bit_ctr_2281__i21 (.Q(bit_ctr[21]), .C(clk16MHz), .E(n7792), 
            .D(n133[21]), .R(n29197));   // verilog/neopixel.v(69[23:32])
    SB_DFFESR bit_ctr_2281__i22 (.Q(bit_ctr[22]), .C(clk16MHz), .E(n7792), 
            .D(n133[22]), .R(n29197));   // verilog/neopixel.v(69[23:32])
    SB_DFFESR bit_ctr_2281__i23 (.Q(bit_ctr[23]), .C(clk16MHz), .E(n7792), 
            .D(n133[23]), .R(n29197));   // verilog/neopixel.v(69[23:32])
    SB_DFFESR bit_ctr_2281__i24 (.Q(bit_ctr[24]), .C(clk16MHz), .E(n7792), 
            .D(n133[24]), .R(n29197));   // verilog/neopixel.v(69[23:32])
    SB_DFFESR bit_ctr_2281__i25 (.Q(bit_ctr[25]), .C(clk16MHz), .E(n7792), 
            .D(n133[25]), .R(n29197));   // verilog/neopixel.v(69[23:32])
    SB_DFFESR bit_ctr_2281__i26 (.Q(bit_ctr[26]), .C(clk16MHz), .E(n7792), 
            .D(n133[26]), .R(n29197));   // verilog/neopixel.v(69[23:32])
    SB_DFFESR bit_ctr_2281__i27 (.Q(bit_ctr[27]), .C(clk16MHz), .E(n7792), 
            .D(n133[27]), .R(n29197));   // verilog/neopixel.v(69[23:32])
    SB_DFFESR bit_ctr_2281__i28 (.Q(bit_ctr[28]), .C(clk16MHz), .E(n7792), 
            .D(n133[28]), .R(n29197));   // verilog/neopixel.v(69[23:32])
    SB_DFFESR bit_ctr_2281__i29 (.Q(bit_ctr[29]), .C(clk16MHz), .E(n7792), 
            .D(n133[29]), .R(n29197));   // verilog/neopixel.v(69[23:32])
    SB_DFFESR bit_ctr_2281__i30 (.Q(bit_ctr[30]), .C(clk16MHz), .E(n7792), 
            .D(n133[30]), .R(n29197));   // verilog/neopixel.v(69[23:32])
    SB_DFFESR bit_ctr_2281__i31 (.Q(bit_ctr[31]), .C(clk16MHz), .E(n7792), 
            .D(n133[31]), .R(n29197));   // verilog/neopixel.v(69[23:32])
    SB_LUT4 sub_14_inv_0_i11_1_lut (.I0(\neo_pixel_transmitter.t0 [10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[10]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i12_1_lut (.I0(\neo_pixel_transmitter.t0 [11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[11]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i13_1_lut (.I0(\neo_pixel_transmitter.t0 [12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[12]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i14_1_lut (.I0(\neo_pixel_transmitter.t0 [13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[13]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i15_1_lut (.I0(\neo_pixel_transmitter.t0 [14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[14]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i16_1_lut (.I0(\neo_pixel_transmitter.t0 [15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[15]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i17_1_lut (.I0(\neo_pixel_transmitter.t0 [16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[16]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i18_1_lut (.I0(\neo_pixel_transmitter.t0 [17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[17]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_4_lut (.I0(\state[1] ), .I1(n37356), .I2(\state[0] ), .I3(\neo_pixel_transmitter.done ), 
            .O(n51332));
    defparam i1_4_lut.LUT_INIT = 16'hf5fd;
    SB_LUT4 i1_4_lut_adj_1702 (.I0(n51332), .I1(n49892), .I2(\state[1] ), 
            .I3(n27251), .O(n28778));
    defparam i1_4_lut_adj_1702.LUT_INIT = 16'ha0a8;
    SB_LUT4 i39673_3_lut (.I0(n56643), .I1(n56949), .I2(color_bit_N_833[2]), 
            .I3(GND_net), .O(n55504));
    defparam i39673_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_3_lut (.I0(bit_ctr[4]), .I1(bit_ctr[3]), .I2(n37163), .I3(GND_net), 
            .O(n45911));
    defparam i1_3_lut.LUT_INIT = 16'h6a6a;
    SB_LUT4 i39733_4_lut (.I0(n55504), .I1(n56853), .I2(bit_ctr[3]), .I3(n37163), 
            .O(n55564));   // verilog/neopixel.v(22[26:38])
    defparam i39733_4_lut.LUT_INIT = 16'hacca;
    SB_LUT4 i39030_3_lut (.I0(n56793), .I1(bit_ctr[3]), .I2(n37163), .I3(GND_net), 
            .O(n54600));
    defparam i39030_3_lut.LUT_INIT = 16'h2828;
    SB_LUT4 i22376_4_lut (.I0(n54600), .I1(\state_3__N_639[1] ), .I2(n55564), 
            .I3(n45911), .O(state_3__N_639[0]));   // verilog/neopixel.v(40[18] 45[12])
    defparam i22376_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 i37482_3_lut (.I0(neopxl_color[16]), .I1(neopxl_color[17]), 
            .I2(bit_ctr[0]), .I3(GND_net), .O(n53312));
    defparam i37482_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i37483_3_lut (.I0(neopxl_color[18]), .I1(neopxl_color[19]), 
            .I2(bit_ctr[0]), .I3(GND_net), .O(n53313));
    defparam i37483_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i37474_3_lut (.I0(neopxl_color[22]), .I1(neopxl_color[23]), 
            .I2(bit_ctr[0]), .I3(GND_net), .O(n53304));
    defparam i37474_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i37473_3_lut (.I0(neopxl_color[20]), .I1(neopxl_color[21]), 
            .I2(bit_ctr[0]), .I3(GND_net), .O(n53303));
    defparam i37473_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 sub_14_inv_0_i25_1_lut (.I0(\neo_pixel_transmitter.t0 [24]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[24]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i25_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 n56946_bdd_4_lut (.I0(n56946), .I1(neopxl_color[9]), .I2(neopxl_color[8]), 
            .I3(color_bit_N_833[1]), .O(n56949));
    defparam n56946_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 sub_14_inv_0_i26_1_lut (.I0(\neo_pixel_transmitter.t0 [25]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[25]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i26_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i27_1_lut (.I0(\neo_pixel_transmitter.t0 [26]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[26]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i27_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i28_1_lut (.I0(\neo_pixel_transmitter.t0 [27]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[27]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i28_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i19_1_lut (.I0(\neo_pixel_transmitter.t0 [18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[18]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_DFF timer_2280__i31 (.Q(timer[31]), .C(clk16MHz), .D(n133_adj_5442[31]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2280__i30 (.Q(timer[30]), .C(clk16MHz), .D(n133_adj_5442[30]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2280__i29 (.Q(timer[29]), .C(clk16MHz), .D(n133_adj_5442[29]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2280__i28 (.Q(timer[28]), .C(clk16MHz), .D(n133_adj_5442[28]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2280__i27 (.Q(timer[27]), .C(clk16MHz), .D(n133_adj_5442[27]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2280__i26 (.Q(timer[26]), .C(clk16MHz), .D(n133_adj_5442[26]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2280__i25 (.Q(timer[25]), .C(clk16MHz), .D(n133_adj_5442[25]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2280__i24 (.Q(timer[24]), .C(clk16MHz), .D(n133_adj_5442[24]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2280__i23 (.Q(timer[23]), .C(clk16MHz), .D(n133_adj_5442[23]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2280__i22 (.Q(timer[22]), .C(clk16MHz), .D(n133_adj_5442[22]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2280__i21 (.Q(timer[21]), .C(clk16MHz), .D(n133_adj_5442[21]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2280__i20 (.Q(timer[20]), .C(clk16MHz), .D(n133_adj_5442[20]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2280__i19 (.Q(timer[19]), .C(clk16MHz), .D(n133_adj_5442[19]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2280__i18 (.Q(timer[18]), .C(clk16MHz), .D(n133_adj_5442[18]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2280__i17 (.Q(timer[17]), .C(clk16MHz), .D(n133_adj_5442[17]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2280__i16 (.Q(timer[16]), .C(clk16MHz), .D(n133_adj_5442[16]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2280__i15 (.Q(timer[15]), .C(clk16MHz), .D(n133_adj_5442[15]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2280__i14 (.Q(timer[14]), .C(clk16MHz), .D(n133_adj_5442[14]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2280__i13 (.Q(timer[13]), .C(clk16MHz), .D(n133_adj_5442[13]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2280__i12 (.Q(timer[12]), .C(clk16MHz), .D(n133_adj_5442[12]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2280__i11 (.Q(timer[11]), .C(clk16MHz), .D(n133_adj_5442[11]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2280__i10 (.Q(timer[10]), .C(clk16MHz), .D(n133_adj_5442[10]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2280__i9 (.Q(timer[9]), .C(clk16MHz), .D(n133_adj_5442[9]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2280__i8 (.Q(timer[8]), .C(clk16MHz), .D(n133_adj_5442[8]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2280__i7 (.Q(timer[7]), .C(clk16MHz), .D(n133_adj_5442[7]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2280__i6 (.Q(timer[6]), .C(clk16MHz), .D(n133_adj_5442[6]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2280__i5 (.Q(timer[5]), .C(clk16MHz), .D(n133_adj_5442[5]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2280__i4 (.Q(timer[4]), .C(clk16MHz), .D(n133_adj_5442[4]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2280__i3 (.Q(timer[3]), .C(clk16MHz), .D(n133_adj_5442[3]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2280__i2 (.Q(timer[2]), .C(clk16MHz), .D(n133_adj_5442[2]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2280__i1 (.Q(timer[1]), .C(clk16MHz), .D(n133_adj_5442[1]));   // verilog/neopixel.v(12[12:21])
    SB_LUT4 sub_14_inv_0_i29_1_lut (.I0(\neo_pixel_transmitter.t0 [28]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[28]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i29_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 color_bit_N_833_1__bdd_4_lut (.I0(color_bit_N_833[1]), .I1(n53210), 
            .I2(n53211), .I3(color_bit_N_833[2]), .O(n56850));
    defparam color_bit_N_833_1__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n56850_bdd_4_lut (.I0(n56850), .I1(n53205), .I2(n53204), .I3(color_bit_N_833[2]), 
            .O(n56853));
    defparam n56850_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 sub_14_inv_0_i30_1_lut (.I0(\neo_pixel_transmitter.t0 [29]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[29]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i30_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i31_1_lut (.I0(\neo_pixel_transmitter.t0 [30]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[30]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i31_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 bit_ctr_2281_add_4_33_lut (.I0(GND_net), .I1(GND_net), .I2(bit_ctr[31]), 
            .I3(n44509), .O(n133[31])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_ctr_2281_add_4_33_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 bit_ctr_2281_add_4_32_lut (.I0(GND_net), .I1(GND_net), .I2(bit_ctr[30]), 
            .I3(n44508), .O(n133[30])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_ctr_2281_add_4_32_lut.LUT_INIT = 16'hC33C;
    SB_CARRY bit_ctr_2281_add_4_32 (.CI(n44508), .I0(GND_net), .I1(bit_ctr[30]), 
            .CO(n44509));
    SB_LUT4 bit_ctr_2281_add_4_31_lut (.I0(GND_net), .I1(GND_net), .I2(bit_ctr[29]), 
            .I3(n44507), .O(n133[29])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_ctr_2281_add_4_31_lut.LUT_INIT = 16'hC33C;
    SB_CARRY bit_ctr_2281_add_4_31 (.CI(n44507), .I0(GND_net), .I1(bit_ctr[29]), 
            .CO(n44508));
    SB_LUT4 bit_ctr_2281_add_4_30_lut (.I0(GND_net), .I1(GND_net), .I2(bit_ctr[28]), 
            .I3(n44506), .O(n133[28])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_ctr_2281_add_4_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY bit_ctr_2281_add_4_30 (.CI(n44506), .I0(GND_net), .I1(bit_ctr[28]), 
            .CO(n44507));
    SB_LUT4 bit_ctr_2281_add_4_29_lut (.I0(GND_net), .I1(GND_net), .I2(bit_ctr[27]), 
            .I3(n44505), .O(n133[27])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_ctr_2281_add_4_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY bit_ctr_2281_add_4_29 (.CI(n44505), .I0(GND_net), .I1(bit_ctr[27]), 
            .CO(n44506));
    SB_LUT4 bit_ctr_2281_add_4_28_lut (.I0(GND_net), .I1(GND_net), .I2(bit_ctr[26]), 
            .I3(n44504), .O(n133[26])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_ctr_2281_add_4_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY bit_ctr_2281_add_4_28 (.CI(n44504), .I0(GND_net), .I1(bit_ctr[26]), 
            .CO(n44505));
    SB_LUT4 bit_ctr_2281_add_4_27_lut (.I0(GND_net), .I1(GND_net), .I2(bit_ctr[25]), 
            .I3(n44503), .O(n133[25])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_ctr_2281_add_4_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY bit_ctr_2281_add_4_27 (.CI(n44503), .I0(GND_net), .I1(bit_ctr[25]), 
            .CO(n44504));
    SB_LUT4 bit_ctr_2281_add_4_26_lut (.I0(GND_net), .I1(GND_net), .I2(bit_ctr[24]), 
            .I3(n44502), .O(n133[24])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_ctr_2281_add_4_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY bit_ctr_2281_add_4_26 (.CI(n44502), .I0(GND_net), .I1(bit_ctr[24]), 
            .CO(n44503));
    SB_LUT4 bit_ctr_2281_add_4_25_lut (.I0(GND_net), .I1(GND_net), .I2(bit_ctr[23]), 
            .I3(n44501), .O(n133[23])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_ctr_2281_add_4_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY bit_ctr_2281_add_4_25 (.CI(n44501), .I0(GND_net), .I1(bit_ctr[23]), 
            .CO(n44502));
    SB_LUT4 sub_14_add_2_33_lut (.I0(n52818), .I1(timer[31]), .I2(n1[31]), 
            .I3(n43609), .O(n27299)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_33_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 bit_ctr_2281_add_4_24_lut (.I0(GND_net), .I1(GND_net), .I2(bit_ctr[22]), 
            .I3(n44500), .O(n133[22])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_ctr_2281_add_4_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY bit_ctr_2281_add_4_24 (.CI(n44500), .I0(GND_net), .I1(bit_ctr[22]), 
            .CO(n44501));
    SB_LUT4 bit_ctr_2281_add_4_23_lut (.I0(GND_net), .I1(GND_net), .I2(bit_ctr[21]), 
            .I3(n44499), .O(n133[21])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_ctr_2281_add_4_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY bit_ctr_2281_add_4_23 (.CI(n44499), .I0(GND_net), .I1(bit_ctr[21]), 
            .CO(n44500));
    SB_LUT4 bit_ctr_2281_add_4_22_lut (.I0(GND_net), .I1(GND_net), .I2(bit_ctr[20]), 
            .I3(n44498), .O(n133[20])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_ctr_2281_add_4_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_14_add_2_32_lut (.I0(n52816), .I1(timer[30]), .I2(n1[30]), 
            .I3(n43608), .O(n52818)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_32_lut.LUT_INIT = 16'hebbe;
    SB_CARRY bit_ctr_2281_add_4_22 (.CI(n44498), .I0(GND_net), .I1(bit_ctr[20]), 
            .CO(n44499));
    SB_CARRY sub_14_add_2_32 (.CI(n43608), .I0(timer[30]), .I1(n1[30]), 
            .CO(n43609));
    SB_LUT4 sub_14_add_2_31_lut (.I0(n52814), .I1(timer[29]), .I2(n1[29]), 
            .I3(n43607), .O(n52816)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_31_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 sub_14_inv_0_i32_1_lut (.I0(\neo_pixel_transmitter.t0 [31]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[31]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i32_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 bit_ctr_2281_add_4_21_lut (.I0(GND_net), .I1(GND_net), .I2(bit_ctr[19]), 
            .I3(n44497), .O(n133[19])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_ctr_2281_add_4_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY bit_ctr_2281_add_4_21 (.CI(n44497), .I0(GND_net), .I1(bit_ctr[19]), 
            .CO(n44498));
    SB_LUT4 bit_ctr_2281_add_4_20_lut (.I0(GND_net), .I1(GND_net), .I2(bit_ctr[18]), 
            .I3(n44496), .O(n133[18])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_ctr_2281_add_4_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY bit_ctr_2281_add_4_20 (.CI(n44496), .I0(GND_net), .I1(bit_ctr[18]), 
            .CO(n44497));
    SB_LUT4 bit_ctr_2281_add_4_19_lut (.I0(GND_net), .I1(GND_net), .I2(bit_ctr[17]), 
            .I3(n44495), .O(n133[17])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_ctr_2281_add_4_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY bit_ctr_2281_add_4_19 (.CI(n44495), .I0(GND_net), .I1(bit_ctr[17]), 
            .CO(n44496));
    SB_LUT4 bit_ctr_2281_add_4_18_lut (.I0(GND_net), .I1(GND_net), .I2(bit_ctr[16]), 
            .I3(n44494), .O(n133[16])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_ctr_2281_add_4_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY bit_ctr_2281_add_4_18 (.CI(n44494), .I0(GND_net), .I1(bit_ctr[16]), 
            .CO(n44495));
    SB_CARRY sub_14_add_2_31 (.CI(n43607), .I0(timer[29]), .I1(n1[29]), 
            .CO(n43608));
    SB_LUT4 sub_14_add_2_30_lut (.I0(n52812), .I1(timer[28]), .I2(n1[28]), 
            .I3(n43606), .O(n52814)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_30_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 bit_ctr_2281_add_4_17_lut (.I0(GND_net), .I1(GND_net), .I2(bit_ctr[15]), 
            .I3(n44493), .O(n133[15])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_ctr_2281_add_4_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY bit_ctr_2281_add_4_17 (.CI(n44493), .I0(GND_net), .I1(bit_ctr[15]), 
            .CO(n44494));
    SB_LUT4 bit_ctr_2281_add_4_16_lut (.I0(GND_net), .I1(GND_net), .I2(bit_ctr[14]), 
            .I3(n44492), .O(n133[14])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_ctr_2281_add_4_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY bit_ctr_2281_add_4_16 (.CI(n44492), .I0(GND_net), .I1(bit_ctr[14]), 
            .CO(n44493));
    SB_LUT4 bit_ctr_2281_add_4_15_lut (.I0(GND_net), .I1(GND_net), .I2(bit_ctr[13]), 
            .I3(n44491), .O(n133[13])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_ctr_2281_add_4_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY bit_ctr_2281_add_4_15 (.CI(n44491), .I0(GND_net), .I1(bit_ctr[13]), 
            .CO(n44492));
    SB_LUT4 bit_ctr_2281_add_4_14_lut (.I0(GND_net), .I1(GND_net), .I2(bit_ctr[12]), 
            .I3(n44490), .O(n133[12])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_ctr_2281_add_4_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_30 (.CI(n43606), .I0(timer[28]), .I1(n1[28]), 
            .CO(n43607));
    SB_CARRY bit_ctr_2281_add_4_14 (.CI(n44490), .I0(GND_net), .I1(bit_ctr[12]), 
            .CO(n44491));
    SB_LUT4 bit_ctr_2281_add_4_13_lut (.I0(GND_net), .I1(GND_net), .I2(bit_ctr[11]), 
            .I3(n44489), .O(n133[11])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_ctr_2281_add_4_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY bit_ctr_2281_add_4_13 (.CI(n44489), .I0(GND_net), .I1(bit_ctr[11]), 
            .CO(n44490));
    SB_LUT4 bit_ctr_2281_add_4_12_lut (.I0(GND_net), .I1(GND_net), .I2(bit_ctr[10]), 
            .I3(n44488), .O(n133[10])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_ctr_2281_add_4_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY bit_ctr_2281_add_4_12 (.CI(n44488), .I0(GND_net), .I1(bit_ctr[10]), 
            .CO(n44489));
    SB_LUT4 bit_ctr_2281_add_4_11_lut (.I0(GND_net), .I1(GND_net), .I2(bit_ctr[9]), 
            .I3(n44487), .O(n133[9])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_ctr_2281_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY bit_ctr_2281_add_4_11 (.CI(n44487), .I0(GND_net), .I1(bit_ctr[9]), 
            .CO(n44488));
    SB_LUT4 bit_ctr_2281_add_4_10_lut (.I0(GND_net), .I1(GND_net), .I2(bit_ctr[8]), 
            .I3(n44486), .O(n133[8])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_ctr_2281_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_14_add_2_29_lut (.I0(n52810), .I1(timer[27]), .I2(n1[27]), 
            .I3(n43605), .O(n52812)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_29_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_14_add_2_29 (.CI(n43605), .I0(timer[27]), .I1(n1[27]), 
            .CO(n43606));
    SB_LUT4 sub_14_add_2_28_lut (.I0(n52808), .I1(timer[26]), .I2(n1[26]), 
            .I3(n43604), .O(n52810)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_28_lut.LUT_INIT = 16'hebbe;
    SB_CARRY bit_ctr_2281_add_4_10 (.CI(n44486), .I0(GND_net), .I1(bit_ctr[8]), 
            .CO(n44487));
    SB_LUT4 bit_ctr_2281_add_4_9_lut (.I0(GND_net), .I1(GND_net), .I2(bit_ctr[7]), 
            .I3(n44485), .O(n133[7])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_ctr_2281_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY bit_ctr_2281_add_4_9 (.CI(n44485), .I0(GND_net), .I1(bit_ctr[7]), 
            .CO(n44486));
    SB_LUT4 bit_ctr_2281_add_4_8_lut (.I0(GND_net), .I1(GND_net), .I2(bit_ctr[6]), 
            .I3(n44484), .O(n133[6])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_ctr_2281_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY bit_ctr_2281_add_4_8 (.CI(n44484), .I0(GND_net), .I1(bit_ctr[6]), 
            .CO(n44485));
    SB_LUT4 bit_ctr_2281_add_4_7_lut (.I0(GND_net), .I1(GND_net), .I2(bit_ctr[5]), 
            .I3(n44483), .O(n133[5])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_ctr_2281_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY bit_ctr_2281_add_4_7 (.CI(n44483), .I0(GND_net), .I1(bit_ctr[5]), 
            .CO(n44484));
    SB_CARRY sub_14_add_2_28 (.CI(n43604), .I0(timer[26]), .I1(n1[26]), 
            .CO(n43605));
    SB_LUT4 bit_ctr_2281_add_4_6_lut (.I0(GND_net), .I1(GND_net), .I2(bit_ctr[4]), 
            .I3(n44482), .O(n133[4])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_ctr_2281_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY bit_ctr_2281_add_4_6 (.CI(n44482), .I0(GND_net), .I1(bit_ctr[4]), 
            .CO(n44483));
    SB_LUT4 bit_ctr_2281_add_4_5_lut (.I0(GND_net), .I1(GND_net), .I2(bit_ctr[3]), 
            .I3(n44481), .O(n133[3])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_ctr_2281_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_14_add_2_27_lut (.I0(n52806), .I1(timer[25]), .I2(n1[25]), 
            .I3(n43603), .O(n52808)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_27_lut.LUT_INIT = 16'hebbe;
    SB_CARRY bit_ctr_2281_add_4_5 (.CI(n44481), .I0(GND_net), .I1(bit_ctr[3]), 
            .CO(n44482));
    SB_CARRY sub_14_add_2_27 (.CI(n43603), .I0(timer[25]), .I1(n1[25]), 
            .CO(n43604));
    SB_LUT4 bit_ctr_2281_add_4_4_lut (.I0(GND_net), .I1(GND_net), .I2(bit_ctr[2]), 
            .I3(n44480), .O(n133[2])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_ctr_2281_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY bit_ctr_2281_add_4_4 (.CI(n44480), .I0(GND_net), .I1(bit_ctr[2]), 
            .CO(n44481));
    SB_DFF timer_2280__i0 (.Q(timer[0]), .C(clk16MHz), .D(n133_adj_5442[0]));   // verilog/neopixel.v(12[12:21])
    SB_LUT4 bit_ctr_2281_add_4_3_lut (.I0(GND_net), .I1(GND_net), .I2(bit_ctr[1]), 
            .I3(n44479), .O(n133[1])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_ctr_2281_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY bit_ctr_2281_add_4_3 (.CI(n44479), .I0(GND_net), .I1(bit_ctr[1]), 
            .CO(n44480));
    SB_LUT4 bit_ctr_2281_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(bit_ctr[0]), 
            .I3(VCC_net), .O(n133[0])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_ctr_2281_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY bit_ctr_2281_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(bit_ctr[0]), 
            .CO(n44479));
    SB_LUT4 timer_2280_add_4_33_lut (.I0(GND_net), .I1(GND_net), .I2(timer[31]), 
            .I3(n44478), .O(n133_adj_5442[31])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2280_add_4_33_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 timer_2280_add_4_32_lut (.I0(GND_net), .I1(GND_net), .I2(timer[30]), 
            .I3(n44477), .O(n133_adj_5442[30])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2280_add_4_32_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2280_add_4_32 (.CI(n44477), .I0(GND_net), .I1(timer[30]), 
            .CO(n44478));
    SB_LUT4 sub_14_add_2_26_lut (.I0(n52804), .I1(timer[24]), .I2(n1[24]), 
            .I3(n43602), .O(n52806)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_26_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 timer_2280_add_4_31_lut (.I0(GND_net), .I1(GND_net), .I2(timer[29]), 
            .I3(n44476), .O(n133_adj_5442[29])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2280_add_4_31_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2280_add_4_31 (.CI(n44476), .I0(GND_net), .I1(timer[29]), 
            .CO(n44477));
    SB_LUT4 color_bit_N_833_1__bdd_4_lut_40979 (.I0(color_bit_N_833[1]), .I1(n53303), 
            .I2(n53304), .I3(color_bit_N_833[2]), .O(n56790));
    defparam color_bit_N_833_1__bdd_4_lut_40979.LUT_INIT = 16'he4aa;
    SB_LUT4 n56790_bdd_4_lut (.I0(n56790), .I1(n53313), .I2(n53312), .I3(color_bit_N_833[2]), 
            .O(n56793));
    defparam n56790_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 timer_2280_add_4_30_lut (.I0(GND_net), .I1(GND_net), .I2(timer[28]), 
            .I3(n44475), .O(n133_adj_5442[28])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2280_add_4_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2280_add_4_30 (.CI(n44475), .I0(GND_net), .I1(timer[28]), 
            .CO(n44476));
    SB_CARRY sub_14_add_2_26 (.CI(n43602), .I0(timer[24]), .I1(n1[24]), 
            .CO(n43603));
    SB_DFFESS state_i0 (.Q(\state[0] ), .C(clk16MHz), .E(n28778), .D(state_3__N_639[0]), 
            .S(n29172));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 sub_14_inv_0_i20_1_lut (.I0(\neo_pixel_transmitter.t0 [19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[19]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 timer_2280_add_4_29_lut (.I0(GND_net), .I1(GND_net), .I2(timer[27]), 
            .I3(n44474), .O(n133_adj_5442[27])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2280_add_4_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2280_add_4_29 (.CI(n44474), .I0(GND_net), .I1(timer[27]), 
            .CO(n44475));
    SB_LUT4 timer_2280_add_4_28_lut (.I0(GND_net), .I1(GND_net), .I2(timer[26]), 
            .I3(n44473), .O(n133_adj_5442[26])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2280_add_4_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2280_add_4_28 (.CI(n44473), .I0(GND_net), .I1(timer[26]), 
            .CO(n44474));
    SB_LUT4 timer_2280_add_4_27_lut (.I0(GND_net), .I1(GND_net), .I2(timer[25]), 
            .I3(n44472), .O(n133_adj_5442[25])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2280_add_4_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2280_add_4_27 (.CI(n44472), .I0(GND_net), .I1(timer[25]), 
            .CO(n44473));
    SB_LUT4 timer_2280_add_4_26_lut (.I0(GND_net), .I1(GND_net), .I2(timer[24]), 
            .I3(n44471), .O(n133_adj_5442[24])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2280_add_4_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2280_add_4_26 (.CI(n44471), .I0(GND_net), .I1(timer[24]), 
            .CO(n44472));
    SB_LUT4 timer_2280_add_4_25_lut (.I0(GND_net), .I1(GND_net), .I2(timer[23]), 
            .I3(n44470), .O(n133_adj_5442[23])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2280_add_4_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2280_add_4_25 (.CI(n44470), .I0(GND_net), .I1(timer[23]), 
            .CO(n44471));
    SB_LUT4 timer_2280_add_4_24_lut (.I0(GND_net), .I1(GND_net), .I2(timer[22]), 
            .I3(n44469), .O(n133_adj_5442[22])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2280_add_4_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2280_add_4_24 (.CI(n44469), .I0(GND_net), .I1(timer[22]), 
            .CO(n44470));
    SB_LUT4 timer_2280_add_4_23_lut (.I0(GND_net), .I1(GND_net), .I2(timer[21]), 
            .I3(n44468), .O(n133_adj_5442[21])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2280_add_4_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2280_add_4_23 (.CI(n44468), .I0(GND_net), .I1(timer[21]), 
            .CO(n44469));
    SB_LUT4 i2_2_lut (.I0(bit_ctr[22]), .I1(bit_ctr[17]), .I2(GND_net), 
            .I3(GND_net), .O(n30));
    defparam i2_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i20_4_lut (.I0(bit_ctr[20]), .I1(bit_ctr[7]), .I2(bit_ctr[16]), 
            .I3(bit_ctr[30]), .O(n48));
    defparam i20_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i18_4_lut (.I0(bit_ctr[25]), .I1(bit_ctr[10]), .I2(bit_ctr[9]), 
            .I3(bit_ctr[27]), .O(n46));
    defparam i18_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i19_4_lut (.I0(bit_ctr[15]), .I1(bit_ctr[29]), .I2(bit_ctr[12]), 
            .I3(bit_ctr[23]), .O(n47));
    defparam i19_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 timer_2280_add_4_22_lut (.I0(GND_net), .I1(GND_net), .I2(timer[20]), 
            .I3(n44467), .O(n133_adj_5442[20])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2280_add_4_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2280_add_4_22 (.CI(n44467), .I0(GND_net), .I1(timer[20]), 
            .CO(n44468));
    SB_LUT4 timer_2280_add_4_21_lut (.I0(GND_net), .I1(GND_net), .I2(timer[19]), 
            .I3(n44466), .O(n133_adj_5442[19])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2280_add_4_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2280_add_4_21 (.CI(n44466), .I0(GND_net), .I1(timer[19]), 
            .CO(n44467));
    SB_LUT4 timer_2280_add_4_20_lut (.I0(GND_net), .I1(GND_net), .I2(timer[18]), 
            .I3(n44465), .O(n133_adj_5442[18])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2280_add_4_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i17_4_lut (.I0(bit_ctr[19]), .I1(bit_ctr[21]), .I2(bit_ctr[31]), 
            .I3(bit_ctr[14]), .O(n45));
    defparam i17_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut (.I0(bit_ctr[11]), .I1(bit_ctr[5]), .I2(bit_ctr[28]), 
            .I3(bit_ctr[6]), .O(n44));
    defparam i16_4_lut.LUT_INIT = 16'hfffe;
    SB_CARRY timer_2280_add_4_20 (.CI(n44465), .I0(GND_net), .I1(timer[18]), 
            .CO(n44466));
    SB_LUT4 i15_4_lut (.I0(bit_ctr[3]), .I1(n30), .I2(bit_ctr[13]), .I3(bit_ctr[4]), 
            .O(n43));
    defparam i15_4_lut.LUT_INIT = 16'hfefc;
    SB_LUT4 i26_4_lut (.I0(n45), .I1(n47), .I2(n46), .I3(n48), .O(n54));
    defparam i26_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i21_4_lut (.I0(bit_ctr[24]), .I1(bit_ctr[8]), .I2(bit_ctr[18]), 
            .I3(bit_ctr[26]), .O(n49));
    defparam i21_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 timer_2280_add_4_19_lut (.I0(GND_net), .I1(GND_net), .I2(timer[17]), 
            .I3(n44464), .O(n133_adj_5442[17])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2280_add_4_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2280_add_4_19 (.CI(n44464), .I0(GND_net), .I1(timer[17]), 
            .CO(n44465));
    SB_LUT4 timer_2280_add_4_18_lut (.I0(GND_net), .I1(GND_net), .I2(timer[16]), 
            .I3(n44463), .O(n133_adj_5442[16])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2280_add_4_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2280_add_4_18 (.CI(n44463), .I0(GND_net), .I1(timer[16]), 
            .CO(n44464));
    SB_LUT4 i27_4_lut (.I0(n49), .I1(n54), .I2(n43), .I3(n44), .O(\state_3__N_639[1] ));
    defparam i27_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i547_2_lut (.I0(LED_c), .I1(\state_3__N_639[1] ), .I2(GND_net), 
            .I3(GND_net), .O(n2586));   // verilog/neopixel.v(40[18] 45[12])
    defparam i547_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 timer_2280_add_4_17_lut (.I0(GND_net), .I1(GND_net), .I2(timer[15]), 
            .I3(n44462), .O(n133_adj_5442[15])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2280_add_4_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2280_add_4_17 (.CI(n44462), .I0(GND_net), .I1(timer[15]), 
            .CO(n44463));
    SB_LUT4 equal_704_i8_2_lut (.I0(\neo_pixel_transmitter.done ), .I1(start), 
            .I2(GND_net), .I3(GND_net), .O(n27251));
    defparam equal_704_i8_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 timer_2280_add_4_16_lut (.I0(GND_net), .I1(GND_net), .I2(timer[14]), 
            .I3(n44461), .O(n133_adj_5442[14])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2280_add_4_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2280_add_4_16 (.CI(n44461), .I0(GND_net), .I1(timer[14]), 
            .CO(n44462));
    SB_LUT4 timer_2280_add_4_15_lut (.I0(GND_net), .I1(GND_net), .I2(timer[13]), 
            .I3(n44460), .O(n133_adj_5442[13])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2280_add_4_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2280_add_4_15 (.CI(n44460), .I0(GND_net), .I1(timer[13]), 
            .CO(n44461));
    SB_LUT4 timer_2280_add_4_14_lut (.I0(GND_net), .I1(GND_net), .I2(timer[12]), 
            .I3(n44459), .O(n133_adj_5442[12])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2280_add_4_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2280_add_4_14 (.CI(n44459), .I0(GND_net), .I1(timer[12]), 
            .CO(n44460));
    SB_LUT4 timer_2280_add_4_13_lut (.I0(GND_net), .I1(GND_net), .I2(timer[11]), 
            .I3(n44458), .O(n133_adj_5442[11])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2280_add_4_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2280_add_4_13 (.CI(n44458), .I0(GND_net), .I1(timer[11]), 
            .CO(n44459));
    SB_LUT4 timer_2280_add_4_12_lut (.I0(GND_net), .I1(GND_net), .I2(timer[10]), 
            .I3(n44457), .O(n133_adj_5442[10])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2280_add_4_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2280_add_4_12 (.CI(n44457), .I0(GND_net), .I1(timer[10]), 
            .CO(n44458));
    SB_LUT4 timer_2280_add_4_11_lut (.I0(GND_net), .I1(GND_net), .I2(timer[9]), 
            .I3(n44456), .O(n133_adj_5442[9])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2280_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2280_add_4_11 (.CI(n44456), .I0(GND_net), .I1(timer[9]), 
            .CO(n44457));
    SB_LUT4 timer_2280_add_4_10_lut (.I0(GND_net), .I1(GND_net), .I2(timer[8]), 
            .I3(n44455), .O(n133_adj_5442[8])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2280_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2280_add_4_10 (.CI(n44455), .I0(GND_net), .I1(timer[8]), 
            .CO(n44456));
    SB_LUT4 timer_2280_add_4_9_lut (.I0(GND_net), .I1(GND_net), .I2(timer[7]), 
            .I3(n44454), .O(n133_adj_5442[7])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2280_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2280_add_4_9 (.CI(n44454), .I0(GND_net), .I1(timer[7]), 
            .CO(n44455));
    SB_LUT4 sub_14_add_2_25_lut (.I0(n52802), .I1(timer[23]), .I2(n1[23]), 
            .I3(n43601), .O(n52804)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_25_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 i3_4_lut (.I0(n54532), .I1(n6_adj_5437), .I2(n2586), .I3(\state[1] ), 
            .O(n29197));
    defparam i3_4_lut.LUT_INIT = 16'hc040;
    SB_LUT4 timer_2280_add_4_8_lut (.I0(GND_net), .I1(GND_net), .I2(timer[6]), 
            .I3(n44453), .O(n133_adj_5442[6])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2280_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2280_add_4_8 (.CI(n44453), .I0(GND_net), .I1(timer[6]), 
            .CO(n44454));
    SB_LUT4 timer_2280_add_4_7_lut (.I0(GND_net), .I1(GND_net), .I2(timer[5]), 
            .I3(n44452), .O(n133_adj_5442[5])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2280_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2280_add_4_7 (.CI(n44452), .I0(GND_net), .I1(timer[5]), 
            .CO(n44453));
    SB_LUT4 timer_2280_add_4_6_lut (.I0(GND_net), .I1(GND_net), .I2(timer[4]), 
            .I3(n44451), .O(n133_adj_5442[4])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2280_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2280_add_4_6 (.CI(n44451), .I0(GND_net), .I1(timer[4]), 
            .CO(n44452));
    SB_LUT4 timer_2280_add_4_5_lut (.I0(GND_net), .I1(GND_net), .I2(timer[3]), 
            .I3(n44450), .O(n133_adj_5442[3])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2280_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i26_4_lut_adj_1703 (.I0(n27251), .I1(n54542), .I2(\state[1] ), 
            .I3(n49892), .O(n7792));
    defparam i26_4_lut_adj_1703.LUT_INIT = 16'hc5c0;
    SB_CARRY timer_2280_add_4_5 (.CI(n44450), .I0(GND_net), .I1(timer[3]), 
            .CO(n44451));
    SB_LUT4 timer_2280_add_4_4_lut (.I0(GND_net), .I1(GND_net), .I2(timer[2]), 
            .I3(n44449), .O(n133_adj_5442[2])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2280_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_25 (.CI(n43601), .I0(timer[23]), .I1(n1[23]), 
            .CO(n43602));
    SB_LUT4 sub_14_add_2_24_lut (.I0(n52800), .I1(timer[22]), .I2(n1[22]), 
            .I3(n43600), .O(n52802)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_24_lut.LUT_INIT = 16'hebbe;
    SB_CARRY timer_2280_add_4_4 (.CI(n44449), .I0(GND_net), .I1(timer[2]), 
            .CO(n44450));
    SB_LUT4 timer_2280_add_4_3_lut (.I0(GND_net), .I1(GND_net), .I2(timer[1]), 
            .I3(n44448), .O(n133_adj_5442[1])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2280_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2280_add_4_3 (.CI(n44448), .I0(GND_net), .I1(timer[1]), 
            .CO(n44449));
    SB_LUT4 timer_2280_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(timer[0]), 
            .I3(VCC_net), .O(n133_adj_5442[0])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2280_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2280_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(timer[0]), 
            .CO(n44448));
    SB_CARRY sub_14_add_2_24 (.CI(n43600), .I0(timer[22]), .I1(n1[22]), 
            .CO(n43601));
    SB_LUT4 sub_14_add_2_23_lut (.I0(n52798), .I1(timer[21]), .I2(n1[21]), 
            .I3(n43599), .O(n52800)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_23_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_14_add_2_23 (.CI(n43599), .I0(timer[21]), .I1(n1[21]), 
            .CO(n43600));
    SB_LUT4 sub_14_add_2_22_lut (.I0(n52796), .I1(timer[20]), .I2(n1[20]), 
            .I3(n43598), .O(n52798)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_22_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_14_add_2_22 (.CI(n43598), .I0(timer[20]), .I1(n1[20]), 
            .CO(n43599));
    SB_LUT4 sub_14_add_2_21_lut (.I0(n52794), .I1(timer[19]), .I2(n1[19]), 
            .I3(n43597), .O(n52796)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_21_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_14_add_2_21 (.CI(n43597), .I0(timer[19]), .I1(n1[19]), 
            .CO(n43598));
    SB_LUT4 sub_14_add_2_20_lut (.I0(n52792), .I1(timer[18]), .I2(n1[18]), 
            .I3(n43596), .O(n52794)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_20_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_14_add_2_20 (.CI(n43596), .I0(timer[18]), .I1(n1[18]), 
            .CO(n43597));
    SB_LUT4 sub_14_add_2_19_lut (.I0(n52790), .I1(timer[17]), .I2(n1[17]), 
            .I3(n43595), .O(n52792)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_19_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_14_add_2_19 (.CI(n43595), .I0(timer[17]), .I1(n1[17]), 
            .CO(n43596));
    SB_LUT4 sub_14_add_2_18_lut (.I0(n52788), .I1(timer[16]), .I2(n1[16]), 
            .I3(n43594), .O(n52790)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_18_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_14_add_2_18 (.CI(n43594), .I0(timer[16]), .I1(n1[16]), 
            .CO(n43595));
    SB_LUT4 sub_14_add_2_17_lut (.I0(n52786), .I1(timer[15]), .I2(n1[15]), 
            .I3(n43593), .O(n52788)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_17_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_14_add_2_17 (.CI(n43593), .I0(timer[15]), .I1(n1[15]), 
            .CO(n43594));
    SB_LUT4 sub_14_add_2_16_lut (.I0(n52784), .I1(timer[14]), .I2(n1[14]), 
            .I3(n43592), .O(n52786)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_16_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_14_add_2_16 (.CI(n43592), .I0(timer[14]), .I1(n1[14]), 
            .CO(n43593));
    SB_LUT4 sub_14_add_2_15_lut (.I0(n52782), .I1(timer[13]), .I2(n1[13]), 
            .I3(n43591), .O(n52784)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_15_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_14_add_2_15 (.CI(n43591), .I0(timer[13]), .I1(n1[13]), 
            .CO(n43592));
    SB_LUT4 sub_14_add_2_14_lut (.I0(one_wire_N_790[11]), .I1(timer[12]), 
            .I2(n1[12]), .I3(n43590), .O(n52782)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_14_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_14_add_2_14 (.CI(n43590), .I0(timer[12]), .I1(n1[12]), 
            .CO(n43591));
    SB_LUT4 sub_14_add_2_13_lut (.I0(GND_net), .I1(timer[11]), .I2(n1[11]), 
            .I3(n43589), .O(one_wire_N_790[11])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_13 (.CI(n43589), .I0(timer[11]), .I1(n1[11]), 
            .CO(n43590));
    SB_LUT4 sub_14_add_2_12_lut (.I0(GND_net), .I1(timer[10]), .I2(n1[10]), 
            .I3(n43588), .O(one_wire_N_790[10])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_12 (.CI(n43588), .I0(timer[10]), .I1(n1[10]), 
            .CO(n43589));
    SB_DFF \neo_pixel_transmitter.t0_i0_i0  (.Q(\neo_pixel_transmitter.t0 [0]), 
           .C(clk16MHz), .D(n29354));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 sub_14_add_2_11_lut (.I0(GND_net), .I1(timer[9]), .I2(n1[9]), 
            .I3(n43587), .O(one_wire_N_790[9])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_11 (.CI(n43587), .I0(timer[9]), .I1(n1[9]), 
            .CO(n43588));
    SB_LUT4 sub_14_add_2_10_lut (.I0(GND_net), .I1(timer[8]), .I2(n1[8]), 
            .I3(n43586), .O(one_wire_N_790[8])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_10 (.CI(n43586), .I0(timer[8]), .I1(n1[8]), 
            .CO(n43587));
    SB_LUT4 sub_14_add_2_9_lut (.I0(GND_net), .I1(timer[7]), .I2(n1[7]), 
            .I3(n43585), .O(one_wire_N_790[7])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_9 (.CI(n43585), .I0(timer[7]), .I1(n1[7]), .CO(n43586));
    SB_LUT4 sub_14_add_2_8_lut (.I0(GND_net), .I1(timer[6]), .I2(n1[6]), 
            .I3(n43584), .O(one_wire_N_790[6])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_8 (.CI(n43584), .I0(timer[6]), .I1(n1[6]), .CO(n43585));
    SB_LUT4 sub_14_add_2_7_lut (.I0(GND_net), .I1(timer[5]), .I2(n1[5]), 
            .I3(n43583), .O(one_wire_N_790[5])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_7 (.CI(n43583), .I0(timer[5]), .I1(n1[5]), .CO(n43584));
    SB_LUT4 sub_14_add_2_6_lut (.I0(GND_net), .I1(timer[4]), .I2(n1[4]), 
            .I3(n43582), .O(one_wire_N_790[4])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_6 (.CI(n43582), .I0(timer[4]), .I1(n1[4]), .CO(n43583));
    SB_LUT4 sub_14_add_2_5_lut (.I0(GND_net), .I1(timer[3]), .I2(n1[3]), 
            .I3(n43581), .O(one_wire_N_790[3])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_5 (.CI(n43581), .I0(timer[3]), .I1(n1[3]), .CO(n43582));
    SB_LUT4 sub_14_add_2_4_lut (.I0(GND_net), .I1(timer[2]), .I2(n1[2]), 
            .I3(n43580), .O(one_wire_N_790[2])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_4 (.CI(n43580), .I0(timer[2]), .I1(n1[2]), .CO(n43581));
    SB_LUT4 sub_14_add_2_3_lut (.I0(GND_net), .I1(timer[1]), .I2(n1[1]), 
            .I3(n43579), .O(one_wire_N_790[1])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_3 (.CI(n43579), .I0(timer[1]), .I1(n1[1]), .CO(n43580));
    SB_CARRY sub_14_add_2_2 (.CI(VCC_net), .I0(timer[0]), .I1(n1[0]), 
            .CO(n43579));
    SB_LUT4 sub_14_inv_0_i21_1_lut (.I0(\neo_pixel_transmitter.t0 [20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[20]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i23080_2_lut_3_lut (.I0(bit_ctr[1]), .I1(bit_ctr[0]), .I2(bit_ctr[2]), 
            .I3(GND_net), .O(n37163));
    defparam i23080_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_2_lut_3_lut (.I0(bit_ctr[1]), .I1(bit_ctr[0]), .I2(bit_ctr[2]), 
            .I3(GND_net), .O(color_bit_N_833[2]));
    defparam i1_2_lut_3_lut.LUT_INIT = 16'h1e1e;
    SB_DFFE state_i1 (.Q(\state[1] ), .C(clk16MHz), .E(VCC_net), .D(n29829));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i1  (.Q(\neo_pixel_transmitter.t0 [1]), 
           .C(clk16MHz), .D(n29814));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i2  (.Q(\neo_pixel_transmitter.t0 [2]), 
           .C(clk16MHz), .D(n29813));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i3  (.Q(\neo_pixel_transmitter.t0 [3]), 
           .C(clk16MHz), .D(n29812));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i4  (.Q(\neo_pixel_transmitter.t0 [4]), 
           .C(clk16MHz), .D(n29811));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i5  (.Q(\neo_pixel_transmitter.t0 [5]), 
           .C(clk16MHz), .D(n29810));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i6  (.Q(\neo_pixel_transmitter.t0 [6]), 
           .C(clk16MHz), .D(n29809));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i7  (.Q(\neo_pixel_transmitter.t0 [7]), 
           .C(clk16MHz), .D(n29808));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i8  (.Q(\neo_pixel_transmitter.t0 [8]), 
           .C(clk16MHz), .D(n29807));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i9  (.Q(\neo_pixel_transmitter.t0 [9]), 
           .C(clk16MHz), .D(n29806));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i10  (.Q(\neo_pixel_transmitter.t0 [10]), 
           .C(clk16MHz), .D(n29805));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i11  (.Q(\neo_pixel_transmitter.t0 [11]), 
           .C(clk16MHz), .D(n29804));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i12  (.Q(\neo_pixel_transmitter.t0 [12]), 
           .C(clk16MHz), .D(n29803));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i13  (.Q(\neo_pixel_transmitter.t0 [13]), 
           .C(clk16MHz), .D(n29802));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i14  (.Q(\neo_pixel_transmitter.t0 [14]), 
           .C(clk16MHz), .D(n29801));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i15  (.Q(\neo_pixel_transmitter.t0 [15]), 
           .C(clk16MHz), .D(n29800));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i16  (.Q(\neo_pixel_transmitter.t0 [16]), 
           .C(clk16MHz), .D(n29799));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i17  (.Q(\neo_pixel_transmitter.t0 [17]), 
           .C(clk16MHz), .D(n29798));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i18  (.Q(\neo_pixel_transmitter.t0 [18]), 
           .C(clk16MHz), .D(n29797));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i19  (.Q(\neo_pixel_transmitter.t0 [19]), 
           .C(clk16MHz), .D(n29796));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i20  (.Q(\neo_pixel_transmitter.t0 [20]), 
           .C(clk16MHz), .D(n29795));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i21  (.Q(\neo_pixel_transmitter.t0 [21]), 
           .C(clk16MHz), .D(n29794));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i22  (.Q(\neo_pixel_transmitter.t0 [22]), 
           .C(clk16MHz), .D(n29793));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i23  (.Q(\neo_pixel_transmitter.t0 [23]), 
           .C(clk16MHz), .D(n29792));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i24  (.Q(\neo_pixel_transmitter.t0 [24]), 
           .C(clk16MHz), .D(n29791));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i25  (.Q(\neo_pixel_transmitter.t0 [25]), 
           .C(clk16MHz), .D(n29790));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i26  (.Q(\neo_pixel_transmitter.t0 [26]), 
           .C(clk16MHz), .D(n29789));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i27  (.Q(\neo_pixel_transmitter.t0 [27]), 
           .C(clk16MHz), .D(n29788));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i28  (.Q(\neo_pixel_transmitter.t0 [28]), 
           .C(clk16MHz), .D(n29785));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i29  (.Q(\neo_pixel_transmitter.t0 [29]), 
           .C(clk16MHz), .D(n29784));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i30  (.Q(\neo_pixel_transmitter.t0 [30]), 
           .C(clk16MHz), .D(n29783));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i31  (.Q(\neo_pixel_transmitter.t0 [31]), 
           .C(clk16MHz), .D(n29782));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 sub_14_inv_0_i1_1_lut (.I0(\neo_pixel_transmitter.t0 [0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[0]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i2_1_lut (.I0(\neo_pixel_transmitter.t0 [1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[1]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 n56640_bdd_4_lut_4_lut (.I0(color_bit_N_833[1]), .I1(neopxl_color[14]), 
            .I2(neopxl_color[15]), .I3(n56640), .O(n56643));   // verilog/neopixel.v(19[6:15])
    defparam n56640_bdd_4_lut_4_lut.LUT_INIT = 16'hf588;
    SB_LUT4 sub_14_inv_0_i3_1_lut (.I0(\neo_pixel_transmitter.t0 [2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[2]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i4_1_lut (.I0(\neo_pixel_transmitter.t0 [3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[3]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_DFFESR one_wire_108 (.Q(NEOPXL_c), .C(clk16MHz), .E(n49955), .D(\neo_pixel_transmitter.done_N_853 ), 
            .R(n51489));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 sub_14_inv_0_i5_1_lut (.I0(\neo_pixel_transmitter.t0 [4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[4]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 bit_ctr_0__bdd_4_lut_41057_4_lut_4_lut (.I0(bit_ctr[1]), .I1(bit_ctr[0]), 
            .I2(neopxl_color[13]), .I3(neopxl_color[12]), .O(n56640));   // verilog/neopixel.v(19[6:15])
    defparam bit_ctr_0__bdd_4_lut_41057_4_lut_4_lut.LUT_INIT = 16'hd5c4;
    SB_LUT4 sub_14_inv_0_i6_1_lut (.I0(\neo_pixel_transmitter.t0 [5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[5]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i37374_3_lut (.I0(neopxl_color[0]), .I1(neopxl_color[1]), .I2(bit_ctr[0]), 
            .I3(GND_net), .O(n53204));
    defparam i37374_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i37375_3_lut (.I0(neopxl_color[2]), .I1(neopxl_color[3]), .I2(bit_ctr[0]), 
            .I3(GND_net), .O(n53205));
    defparam i37375_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i37381_3_lut (.I0(neopxl_color[6]), .I1(neopxl_color[7]), .I2(bit_ctr[0]), 
            .I3(GND_net), .O(n53211));
    defparam i37381_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i37380_3_lut (.I0(neopxl_color[4]), .I1(neopxl_color[5]), .I2(bit_ctr[0]), 
            .I3(GND_net), .O(n53210));
    defparam i37380_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 sub_14_inv_0_i7_1_lut (.I0(\neo_pixel_transmitter.t0 [6]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[6]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i2_2_lut_3_lut (.I0(\state[0] ), .I1(\state[1] ), .I2(n7792), 
            .I3(GND_net), .O(n6_adj_5437));   // verilog/neopixel.v(36[4] 116[11])
    defparam i2_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 sub_14_inv_0_i8_1_lut (.I0(\neo_pixel_transmitter.t0 [7]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[7]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i15092_2_lut_3_lut (.I0(\state[0] ), .I1(\state[1] ), .I2(n28778), 
            .I3(GND_net), .O(n29172));   // verilog/neopixel.v(36[4] 116[11])
    defparam i15092_2_lut_3_lut.LUT_INIT = 16'h7070;
    SB_LUT4 sub_14_inv_0_i9_1_lut (.I0(\neo_pixel_transmitter.t0 [8]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[8]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i10_1_lut (.I0(\neo_pixel_transmitter.t0 [9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[9]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i34176_4_lut (.I0(n27111), .I1(n49822), .I2(n45295), .I3(\state[0] ), 
            .O(n49935));
    defparam i34176_4_lut.LUT_INIT = 16'hfaee;
    SB_LUT4 i20_4_lut_adj_1704 (.I0(\neo_pixel_transmitter.done ), .I1(\state[1] ), 
            .I2(start), .I3(n49935), .O(n7_adj_5439));
    defparam i20_4_lut_adj_1704.LUT_INIT = 16'hcecf;
    SB_LUT4 i1_4_lut_adj_1705 (.I0(n27251), .I1(n7_adj_5439), .I2(n49892), 
            .I3(\state[1] ), .O(n47790));
    defparam i1_4_lut_adj_1705.LUT_INIT = 16'hcc8c;
    SB_LUT4 i39017_2_lut_3_lut (.I0(LED_c), .I1(\state_3__N_639[1] ), .I2(\state[0] ), 
            .I3(GND_net), .O(n54542));
    defparam i39017_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i39009_3_lut_4_lut (.I0(n27111), .I1(\neo_pixel_transmitter.done ), 
            .I2(start), .I3(n49822), .O(n54532));
    defparam i39009_3_lut_4_lut.LUT_INIT = 16'hf3f7;
    SB_LUT4 i34070_2_lut (.I0(one_wire_N_790[3]), .I1(one_wire_N_790[2]), 
            .I2(GND_net), .I3(GND_net), .O(n49822));
    defparam i34070_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i2_3_lut (.I0(one_wire_N_790[3]), .I1(one_wire_N_790[2]), .I2(one_wire_N_790[1]), 
            .I3(GND_net), .O(n45295));
    defparam i2_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i1_2_lut_adj_1706 (.I0(one_wire_N_790[5]), .I1(one_wire_N_790[4]), 
            .I2(GND_net), .I3(GND_net), .O(n52822));   // verilog/neopixel.v(62[15:42])
    defparam i1_2_lut_adj_1706.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_1707 (.I0(one_wire_N_790[8]), .I1(one_wire_N_790[7]), 
            .I2(one_wire_N_790[6]), .I3(n52822), .O(n52828));   // verilog/neopixel.v(62[15:42])
    defparam i1_4_lut_adj_1707.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1708 (.I0(one_wire_N_790[10]), .I1(n27299), .I2(one_wire_N_790[9]), 
            .I3(n52828), .O(n27111));   // verilog/neopixel.v(62[15:42])
    defparam i1_4_lut_adj_1708.LUT_INIT = 16'hfffe;
    SB_LUT4 i34174_4_lut (.I0(n27111), .I1(n45295), .I2(n49822), .I3(\state[0] ), 
            .O(n49892));
    defparam i34174_4_lut.LUT_INIT = 16'hfaee;
    SB_LUT4 i23266_4_lut (.I0(one_wire_N_790[8]), .I1(n27299), .I2(one_wire_N_790[10]), 
            .I3(one_wire_N_790[9]), .O(n37356));
    defparam i23266_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 i39010_2_lut (.I0(\neo_pixel_transmitter.done ), .I1(\state[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n54545));
    defparam i39010_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i33998_3_lut (.I0(\neo_pixel_transmitter.done ), .I1(start), 
            .I2(n49892), .I3(GND_net), .O(n49746));
    defparam i33998_3_lut.LUT_INIT = 16'hecec;
    SB_LUT4 i15_4_lut_adj_1709 (.I0(n49746), .I1(n54545), .I2(\state[1] ), 
            .I3(n37356), .O(n7));
    defparam i15_4_lut_adj_1709.LUT_INIT = 16'h3a0a;
    SB_LUT4 i40650_2_lut (.I0(start), .I1(\state[1] ), .I2(GND_net), .I3(GND_net), 
            .O(start_N_838));   // verilog/neopixel.v(36[4] 116[11])
    defparam i40650_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 i34066_2_lut (.I0(start), .I1(\state[1] ), .I2(GND_net), .I3(GND_net), 
            .O(n49818));
    defparam i34066_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i40065_2_lut (.I0(\neo_pixel_transmitter.done ), .I1(\state[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n48982));
    defparam i40065_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1710 (.I0(one_wire_N_790[2]), .I1(n48982), .I2(one_wire_N_790[3]), 
            .I3(one_wire_N_790[1]), .O(n103));
    defparam i1_4_lut_adj_1710.LUT_INIT = 16'h4dcd;
    SB_LUT4 i6_4_lut (.I0(one_wire_N_790[7]), .I1(one_wire_N_790[9]), .I2(n49818), 
            .I3(n103), .O(n16_adj_5440));
    defparam i6_4_lut.LUT_INIT = 16'h0100;
    SB_LUT4 i1_4_lut_adj_1711 (.I0(one_wire_N_790[8]), .I1(one_wire_N_790[4]), 
            .I2(n16_adj_5440), .I3(n27299), .O(n6_adj_5441));
    defparam i1_4_lut_adj_1711.LUT_INIT = 16'hffef;
    SB_LUT4 i4_4_lut (.I0(one_wire_N_790[10]), .I1(one_wire_N_790[6]), .I2(one_wire_N_790[5]), 
            .I3(n6_adj_5441), .O(n56981));
    defparam i4_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 mux_1370_Mux_0_i3_3_lut (.I0(start), .I1(\neo_pixel_transmitter.done ), 
            .I2(\state[1] ), .I3(GND_net), .O(\neo_pixel_transmitter.done_N_847 ));   // verilog/neopixel.v(36[4] 116[11])
    defparam mux_1370_Mux_0_i3_3_lut.LUT_INIT = 16'hc1c1;
    SB_LUT4 sub_14_inv_0_i22_1_lut (.I0(\neo_pixel_transmitter.t0 [21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[21]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 bit_ctr_0__bdd_4_lut_4_lut (.I0(bit_ctr[0]), .I1(neopxl_color[10]), 
            .I2(neopxl_color[11]), .I3(bit_ctr[1]), .O(n56946));
    defparam bit_ctr_0__bdd_4_lut_4_lut.LUT_INIT = 16'heea0;
    SB_LUT4 sub_14_inv_0_i23_1_lut (.I0(\neo_pixel_transmitter.t0 [22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[22]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i24_1_lut (.I0(\neo_pixel_transmitter.t0 [23]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[23]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i39289_3_lut_4_lut (.I0(n27111), .I1(n55119), .I2(start), 
            .I3(\state[1] ), .O(n55120));
    defparam i39289_3_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i39012_2_lut_3_lut (.I0(one_wire_N_790[3]), .I1(one_wire_N_790[2]), 
            .I2(start), .I3(GND_net), .O(n54536));
    defparam i39012_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i3_4_lut_4_lut (.I0(n37356), .I1(\state[1] ), .I2(\state[0] ), 
            .I3(\neo_pixel_transmitter.done ), .O(n51489));
    defparam i3_4_lut_4_lut.LUT_INIT = 16'h0004;
    
endmodule
//
// Verilog Description of module \quadrature_decoder(1)_U0 
//

module \quadrature_decoder(1)_U0  (n2269, b_prev, GND_net, a_new, position_31__N_4108, 
            ENCODER0_B_N_keep, ENCODER0_A_N_keep, encoder0_position, n29501, 
            n2233, VCC_net) /* synthesis lattice_noprune=1 */ ;
    input n2269;
    output b_prev;
    input GND_net;
    output [1:0]a_new;
    output position_31__N_4108;
    input ENCODER0_B_N_keep;
    input ENCODER0_A_N_keep;
    output [31:0]encoder0_position;
    input n29501;
    output n2233;
    input VCC_net;
    
    
    wire n29517, a_prev;
    wire [1:0]b_new;   // vhdl/quadrature_decoder.vhd(40[9:14])
    
    wire position_31__N_4111, debounce_cnt, direction_N_4113;
    wire [1:0]a_new_c;   // vhdl/quadrature_decoder.vhd(39[9:14])
    
    wire a_prev_N_4116;
    wire [31:0]n133;
    
    wire n44594, n44593, n44592, n44591, n44590, n44589, n44588, 
        n44587, n44586, n44585, n44584, n44583, n44582, n44581, 
        n44580, n44579, n44578, n44577, n44576, n44575, n44574, 
        n44573, n44572, n44571, n44570, n44569, n44568, n44567, 
        n44566, n44565, n44564, n29535;
    
    SB_DFF a_prev_38 (.Q(a_prev), .C(n2269), .D(n29517));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_LUT4 b_prev_I_0_43_2_lut (.I0(b_prev), .I1(b_new[1]), .I2(GND_net), 
            .I3(GND_net), .O(position_31__N_4111));   // vhdl/quadrature_decoder.vhd(63[37:56])
    defparam b_prev_I_0_43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 debounce_cnt_I_0_4_lut (.I0(debounce_cnt), .I1(a_prev), .I2(position_31__N_4111), 
            .I3(a_new[1]), .O(position_31__N_4108));   // vhdl/quadrature_decoder.vhd(62[7] 63[64])
    defparam debounce_cnt_I_0_4_lut.LUT_INIT = 16'ha2a8;
    SB_LUT4 b_prev_I_0_45_2_lut (.I0(b_prev), .I1(a_new[1]), .I2(GND_net), 
            .I3(GND_net), .O(direction_N_4113));   // vhdl/quadrature_decoder.vhd(64[18:37])
    defparam b_prev_I_0_45_2_lut.LUT_INIT = 16'h9999;
    SB_DFF b_new_i0 (.Q(b_new[0]), .C(n2269), .D(ENCODER0_B_N_keep));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_DFF a_new_i0 (.Q(a_new_c[0]), .C(n2269), .D(ENCODER0_A_N_keep));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_DFF debounce_cnt_37 (.Q(debounce_cnt), .C(n2269), .D(a_prev_N_4116));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_LUT4 position_2284_add_4_33_lut (.I0(GND_net), .I1(direction_N_4113), 
            .I2(encoder0_position[31]), .I3(n44594), .O(n133[31])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2284_add_4_33_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 position_2284_add_4_32_lut (.I0(GND_net), .I1(direction_N_4113), 
            .I2(encoder0_position[30]), .I3(n44593), .O(n133[30])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2284_add_4_32_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2284_add_4_32 (.CI(n44593), .I0(direction_N_4113), 
            .I1(encoder0_position[30]), .CO(n44594));
    SB_LUT4 position_2284_add_4_31_lut (.I0(GND_net), .I1(direction_N_4113), 
            .I2(encoder0_position[29]), .I3(n44592), .O(n133[29])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2284_add_4_31_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2284_add_4_31 (.CI(n44592), .I0(direction_N_4113), 
            .I1(encoder0_position[29]), .CO(n44593));
    SB_LUT4 position_2284_add_4_30_lut (.I0(GND_net), .I1(direction_N_4113), 
            .I2(encoder0_position[28]), .I3(n44591), .O(n133[28])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2284_add_4_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2284_add_4_30 (.CI(n44591), .I0(direction_N_4113), 
            .I1(encoder0_position[28]), .CO(n44592));
    SB_LUT4 position_2284_add_4_29_lut (.I0(GND_net), .I1(direction_N_4113), 
            .I2(encoder0_position[27]), .I3(n44590), .O(n133[27])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2284_add_4_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2284_add_4_29 (.CI(n44590), .I0(direction_N_4113), 
            .I1(encoder0_position[27]), .CO(n44591));
    SB_LUT4 position_2284_add_4_28_lut (.I0(GND_net), .I1(direction_N_4113), 
            .I2(encoder0_position[26]), .I3(n44589), .O(n133[26])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2284_add_4_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2284_add_4_28 (.CI(n44589), .I0(direction_N_4113), 
            .I1(encoder0_position[26]), .CO(n44590));
    SB_LUT4 position_2284_add_4_27_lut (.I0(GND_net), .I1(direction_N_4113), 
            .I2(encoder0_position[25]), .I3(n44588), .O(n133[25])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2284_add_4_27_lut.LUT_INIT = 16'hC33C;
    SB_DFF direction_40 (.Q(n2233), .C(n2269), .D(n29501));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_CARRY position_2284_add_4_27 (.CI(n44588), .I0(direction_N_4113), 
            .I1(encoder0_position[25]), .CO(n44589));
    SB_LUT4 position_2284_add_4_26_lut (.I0(GND_net), .I1(direction_N_4113), 
            .I2(encoder0_position[24]), .I3(n44587), .O(n133[24])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2284_add_4_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2284_add_4_26 (.CI(n44587), .I0(direction_N_4113), 
            .I1(encoder0_position[24]), .CO(n44588));
    SB_LUT4 position_2284_add_4_25_lut (.I0(GND_net), .I1(direction_N_4113), 
            .I2(encoder0_position[23]), .I3(n44586), .O(n133[23])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2284_add_4_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2284_add_4_25 (.CI(n44586), .I0(direction_N_4113), 
            .I1(encoder0_position[23]), .CO(n44587));
    SB_LUT4 position_2284_add_4_24_lut (.I0(GND_net), .I1(direction_N_4113), 
            .I2(encoder0_position[22]), .I3(n44585), .O(n133[22])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2284_add_4_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2284_add_4_24 (.CI(n44585), .I0(direction_N_4113), 
            .I1(encoder0_position[22]), .CO(n44586));
    SB_LUT4 position_2284_add_4_23_lut (.I0(GND_net), .I1(direction_N_4113), 
            .I2(encoder0_position[21]), .I3(n44584), .O(n133[21])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2284_add_4_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2284_add_4_23 (.CI(n44584), .I0(direction_N_4113), 
            .I1(encoder0_position[21]), .CO(n44585));
    SB_LUT4 position_2284_add_4_22_lut (.I0(GND_net), .I1(direction_N_4113), 
            .I2(encoder0_position[20]), .I3(n44583), .O(n133[20])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2284_add_4_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2284_add_4_22 (.CI(n44583), .I0(direction_N_4113), 
            .I1(encoder0_position[20]), .CO(n44584));
    SB_LUT4 position_2284_add_4_21_lut (.I0(GND_net), .I1(direction_N_4113), 
            .I2(encoder0_position[19]), .I3(n44582), .O(n133[19])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2284_add_4_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2284_add_4_21 (.CI(n44582), .I0(direction_N_4113), 
            .I1(encoder0_position[19]), .CO(n44583));
    SB_LUT4 position_2284_add_4_20_lut (.I0(GND_net), .I1(direction_N_4113), 
            .I2(encoder0_position[18]), .I3(n44581), .O(n133[18])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2284_add_4_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2284_add_4_20 (.CI(n44581), .I0(direction_N_4113), 
            .I1(encoder0_position[18]), .CO(n44582));
    SB_LUT4 position_2284_add_4_19_lut (.I0(GND_net), .I1(direction_N_4113), 
            .I2(encoder0_position[17]), .I3(n44580), .O(n133[17])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2284_add_4_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2284_add_4_19 (.CI(n44580), .I0(direction_N_4113), 
            .I1(encoder0_position[17]), .CO(n44581));
    SB_LUT4 position_2284_add_4_18_lut (.I0(GND_net), .I1(direction_N_4113), 
            .I2(encoder0_position[16]), .I3(n44579), .O(n133[16])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2284_add_4_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2284_add_4_18 (.CI(n44579), .I0(direction_N_4113), 
            .I1(encoder0_position[16]), .CO(n44580));
    SB_LUT4 position_2284_add_4_17_lut (.I0(GND_net), .I1(direction_N_4113), 
            .I2(encoder0_position[15]), .I3(n44578), .O(n133[15])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2284_add_4_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2284_add_4_17 (.CI(n44578), .I0(direction_N_4113), 
            .I1(encoder0_position[15]), .CO(n44579));
    SB_LUT4 position_2284_add_4_16_lut (.I0(GND_net), .I1(direction_N_4113), 
            .I2(encoder0_position[14]), .I3(n44577), .O(n133[14])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2284_add_4_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2284_add_4_16 (.CI(n44577), .I0(direction_N_4113), 
            .I1(encoder0_position[14]), .CO(n44578));
    SB_LUT4 position_2284_add_4_15_lut (.I0(GND_net), .I1(direction_N_4113), 
            .I2(encoder0_position[13]), .I3(n44576), .O(n133[13])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2284_add_4_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2284_add_4_15 (.CI(n44576), .I0(direction_N_4113), 
            .I1(encoder0_position[13]), .CO(n44577));
    SB_LUT4 position_2284_add_4_14_lut (.I0(GND_net), .I1(direction_N_4113), 
            .I2(encoder0_position[12]), .I3(n44575), .O(n133[12])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2284_add_4_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2284_add_4_14 (.CI(n44575), .I0(direction_N_4113), 
            .I1(encoder0_position[12]), .CO(n44576));
    SB_LUT4 position_2284_add_4_13_lut (.I0(GND_net), .I1(direction_N_4113), 
            .I2(encoder0_position[11]), .I3(n44574), .O(n133[11])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2284_add_4_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2284_add_4_13 (.CI(n44574), .I0(direction_N_4113), 
            .I1(encoder0_position[11]), .CO(n44575));
    SB_LUT4 position_2284_add_4_12_lut (.I0(GND_net), .I1(direction_N_4113), 
            .I2(encoder0_position[10]), .I3(n44573), .O(n133[10])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2284_add_4_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2284_add_4_12 (.CI(n44573), .I0(direction_N_4113), 
            .I1(encoder0_position[10]), .CO(n44574));
    SB_LUT4 position_2284_add_4_11_lut (.I0(GND_net), .I1(direction_N_4113), 
            .I2(encoder0_position[9]), .I3(n44572), .O(n133[9])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2284_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2284_add_4_11 (.CI(n44572), .I0(direction_N_4113), 
            .I1(encoder0_position[9]), .CO(n44573));
    SB_LUT4 position_2284_add_4_10_lut (.I0(GND_net), .I1(direction_N_4113), 
            .I2(encoder0_position[8]), .I3(n44571), .O(n133[8])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2284_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2284_add_4_10 (.CI(n44571), .I0(direction_N_4113), 
            .I1(encoder0_position[8]), .CO(n44572));
    SB_LUT4 position_2284_add_4_9_lut (.I0(GND_net), .I1(direction_N_4113), 
            .I2(encoder0_position[7]), .I3(n44570), .O(n133[7])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2284_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2284_add_4_9 (.CI(n44570), .I0(direction_N_4113), 
            .I1(encoder0_position[7]), .CO(n44571));
    SB_LUT4 position_2284_add_4_8_lut (.I0(GND_net), .I1(direction_N_4113), 
            .I2(encoder0_position[6]), .I3(n44569), .O(n133[6])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2284_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2284_add_4_8 (.CI(n44569), .I0(direction_N_4113), 
            .I1(encoder0_position[6]), .CO(n44570));
    SB_LUT4 position_2284_add_4_7_lut (.I0(GND_net), .I1(direction_N_4113), 
            .I2(encoder0_position[5]), .I3(n44568), .O(n133[5])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2284_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2284_add_4_7 (.CI(n44568), .I0(direction_N_4113), 
            .I1(encoder0_position[5]), .CO(n44569));
    SB_LUT4 position_2284_add_4_6_lut (.I0(GND_net), .I1(direction_N_4113), 
            .I2(encoder0_position[4]), .I3(n44567), .O(n133[4])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2284_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2284_add_4_6 (.CI(n44567), .I0(direction_N_4113), 
            .I1(encoder0_position[4]), .CO(n44568));
    SB_LUT4 position_2284_add_4_5_lut (.I0(GND_net), .I1(direction_N_4113), 
            .I2(encoder0_position[3]), .I3(n44566), .O(n133[3])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2284_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2284_add_4_5 (.CI(n44566), .I0(direction_N_4113), 
            .I1(encoder0_position[3]), .CO(n44567));
    SB_LUT4 position_2284_add_4_4_lut (.I0(GND_net), .I1(direction_N_4113), 
            .I2(encoder0_position[2]), .I3(n44565), .O(n133[2])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2284_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2284_add_4_4 (.CI(n44565), .I0(direction_N_4113), 
            .I1(encoder0_position[2]), .CO(n44566));
    SB_LUT4 position_2284_add_4_3_lut (.I0(GND_net), .I1(direction_N_4113), 
            .I2(encoder0_position[1]), .I3(n44564), .O(n133[1])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2284_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2284_add_4_3 (.CI(n44564), .I0(direction_N_4113), 
            .I1(encoder0_position[1]), .CO(n44565));
    SB_LUT4 position_2284_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(encoder0_position[0]), 
            .I3(VCC_net), .O(n133[0])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2284_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2284_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(encoder0_position[0]), 
            .CO(n44564));
    SB_DFFE position_2284__i31 (.Q(encoder0_position[31]), .C(n2269), .E(position_31__N_4108), 
            .D(n133[31]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2284__i30 (.Q(encoder0_position[30]), .C(n2269), .E(position_31__N_4108), 
            .D(n133[30]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2284__i29 (.Q(encoder0_position[29]), .C(n2269), .E(position_31__N_4108), 
            .D(n133[29]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2284__i28 (.Q(encoder0_position[28]), .C(n2269), .E(position_31__N_4108), 
            .D(n133[28]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2284__i27 (.Q(encoder0_position[27]), .C(n2269), .E(position_31__N_4108), 
            .D(n133[27]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2284__i26 (.Q(encoder0_position[26]), .C(n2269), .E(position_31__N_4108), 
            .D(n133[26]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2284__i25 (.Q(encoder0_position[25]), .C(n2269), .E(position_31__N_4108), 
            .D(n133[25]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2284__i24 (.Q(encoder0_position[24]), .C(n2269), .E(position_31__N_4108), 
            .D(n133[24]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2284__i23 (.Q(encoder0_position[23]), .C(n2269), .E(position_31__N_4108), 
            .D(n133[23]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2284__i22 (.Q(encoder0_position[22]), .C(n2269), .E(position_31__N_4108), 
            .D(n133[22]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2284__i21 (.Q(encoder0_position[21]), .C(n2269), .E(position_31__N_4108), 
            .D(n133[21]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2284__i20 (.Q(encoder0_position[20]), .C(n2269), .E(position_31__N_4108), 
            .D(n133[20]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2284__i19 (.Q(encoder0_position[19]), .C(n2269), .E(position_31__N_4108), 
            .D(n133[19]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2284__i18 (.Q(encoder0_position[18]), .C(n2269), .E(position_31__N_4108), 
            .D(n133[18]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2284__i17 (.Q(encoder0_position[17]), .C(n2269), .E(position_31__N_4108), 
            .D(n133[17]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2284__i16 (.Q(encoder0_position[16]), .C(n2269), .E(position_31__N_4108), 
            .D(n133[16]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2284__i15 (.Q(encoder0_position[15]), .C(n2269), .E(position_31__N_4108), 
            .D(n133[15]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2284__i14 (.Q(encoder0_position[14]), .C(n2269), .E(position_31__N_4108), 
            .D(n133[14]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2284__i13 (.Q(encoder0_position[13]), .C(n2269), .E(position_31__N_4108), 
            .D(n133[13]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2284__i12 (.Q(encoder0_position[12]), .C(n2269), .E(position_31__N_4108), 
            .D(n133[12]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2284__i11 (.Q(encoder0_position[11]), .C(n2269), .E(position_31__N_4108), 
            .D(n133[11]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2284__i10 (.Q(encoder0_position[10]), .C(n2269), .E(position_31__N_4108), 
            .D(n133[10]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2284__i9 (.Q(encoder0_position[9]), .C(n2269), .E(position_31__N_4108), 
            .D(n133[9]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2284__i8 (.Q(encoder0_position[8]), .C(n2269), .E(position_31__N_4108), 
            .D(n133[8]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2284__i7 (.Q(encoder0_position[7]), .C(n2269), .E(position_31__N_4108), 
            .D(n133[7]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2284__i6 (.Q(encoder0_position[6]), .C(n2269), .E(position_31__N_4108), 
            .D(n133[6]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2284__i5 (.Q(encoder0_position[5]), .C(n2269), .E(position_31__N_4108), 
            .D(n133[5]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2284__i4 (.Q(encoder0_position[4]), .C(n2269), .E(position_31__N_4108), 
            .D(n133[4]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2284__i3 (.Q(encoder0_position[3]), .C(n2269), .E(position_31__N_4108), 
            .D(n133[3]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2284__i2 (.Q(encoder0_position[2]), .C(n2269), .E(position_31__N_4108), 
            .D(n133[2]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2284__i1 (.Q(encoder0_position[1]), .C(n2269), .E(position_31__N_4108), 
            .D(n133[1]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2284__i0 (.Q(encoder0_position[0]), .C(n2269), .E(position_31__N_4108), 
            .D(n133[0]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFF a_new_i1 (.Q(a_new[1]), .C(n2269), .D(a_new_c[0]));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_DFF b_new_i1 (.Q(b_new[1]), .C(n2269), .D(b_new[0]));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_LUT4 i15437_3_lut_4_lut (.I0(debounce_cnt), .I1(a_prev_N_4116), .I2(a_new[1]), 
            .I3(a_prev), .O(n29517));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    defparam i15437_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i15455_3_lut_4_lut (.I0(debounce_cnt), .I1(a_prev_N_4116), .I2(b_new[1]), 
            .I3(b_prev), .O(n29535));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    defparam i15455_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF b_prev_39 (.Q(b_prev), .C(n2269), .D(n29535));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_LUT4 i40078_4_lut (.I0(a_new_c[0]), .I1(b_new[0]), .I2(a_new[1]), 
            .I3(b_new[1]), .O(a_prev_N_4116));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    defparam i40078_4_lut.LUT_INIT = 16'h8421;
    
endmodule
//
// Verilog Description of module pll32MHz
//

module pll32MHz (GND_net, clk16MHz, VCC_net, clk32MHz) /* synthesis syn_module_defined=1 */ ;
    input GND_net;
    input clk16MHz;
    input VCC_net;
    output clk32MHz;
    
    wire clk16MHz /* synthesis SET_AS_NETWORK=clk16MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[16:24])
    
    SB_PLL40_CORE pll32MHz_inst (.REFERENCECLK(clk16MHz), .PLLOUTCORE(clk32MHz), 
            .BYPASS(GND_net), .RESETB(VCC_net)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=52, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=34, LSE_RLINE=38 */ ;   // verilog/TinyFPGA_B.v(34[10] 38[2])
    defparam pll32MHz_inst.FEEDBACK_PATH = "PHASE_AND_DELAY";
    defparam pll32MHz_inst.DELAY_ADJUSTMENT_MODE_FEEDBACK = "FIXED";
    defparam pll32MHz_inst.DELAY_ADJUSTMENT_MODE_RELATIVE = "FIXED";
    defparam pll32MHz_inst.SHIFTREG_DIV_MODE = 2'b00;
    defparam pll32MHz_inst.FDA_FEEDBACK = 4'b0000;
    defparam pll32MHz_inst.FDA_RELATIVE = 4'b0000;
    defparam pll32MHz_inst.PLLOUT_SELECT = "SHIFTREG_0deg";
    defparam pll32MHz_inst.DIVR = 4'b0000;
    defparam pll32MHz_inst.DIVF = 7'b0000001;
    defparam pll32MHz_inst.DIVQ = 3'b011;
    defparam pll32MHz_inst.FILTER_RANGE = 3'b001;
    defparam pll32MHz_inst.ENABLE_ICEGATE = 1'b0;
    defparam pll32MHz_inst.TEST_MODE = 1'b0;
    defparam pll32MHz_inst.EXTERNAL_DIVIDE_FACTOR = 1;
    
endmodule
//
// Verilog Description of module motorControl
//

module motorControl (\Kp[14] , GND_net, \Kp[0] , \Kp[2] , \Kp[11] , 
            \Kp[12] , \Kp[3] , \Kp[4] , \Kp[5] , \Ki[12] , \PID_CONTROLLER.integral_23__N_3996 , 
            \Kp[13] , \Ki[7] , \Ki[8] , \Kp[6] , \Ki[13] , \Ki[14] , 
            \Ki[9] , \Kp[15] , \Kp[7] , \Kp[8] , \Ki[15] , control_update, 
            duty, clk16MHz, \Kp[9] , \Kp[10] , IntegralLimit, \Ki[1] , 
            \Ki[0] , \Kp[1] , \Ki[2] , \Ki[3] , \Ki[4] , \Ki[5] , 
            \Ki[6] , \Ki[10] , \Ki[11] , PWMLimit, n363, n32464, 
            deadband, VCC_net, \PID_CONTROLLER.integral , n29381, setpoint, 
            motor_state, n29915, n29914, n29913, n29912, n29911, 
            n29910, n29909, n29908, n29907, n29906, n29905, n29904, 
            n29903, n29902, n29901, n29900, n29899, n29898, n29897, 
            n29896, n29895, n29894, n29893) /* synthesis syn_module_defined=1 */ ;
    input \Kp[14] ;
    input GND_net;
    input \Kp[0] ;
    input \Kp[2] ;
    input \Kp[11] ;
    input \Kp[12] ;
    input \Kp[3] ;
    input \Kp[4] ;
    input \Kp[5] ;
    input \Ki[12] ;
    output [23:0]\PID_CONTROLLER.integral_23__N_3996 ;
    input \Kp[13] ;
    input \Ki[7] ;
    input \Ki[8] ;
    input \Kp[6] ;
    input \Ki[13] ;
    input \Ki[14] ;
    input \Ki[9] ;
    input \Kp[15] ;
    input \Kp[7] ;
    input \Kp[8] ;
    input \Ki[15] ;
    output control_update;
    output [23:0]duty;
    input clk16MHz;
    input \Kp[9] ;
    input \Kp[10] ;
    input [23:0]IntegralLimit;
    input \Ki[1] ;
    input \Ki[0] ;
    input \Kp[1] ;
    input \Ki[2] ;
    input \Ki[3] ;
    input \Ki[4] ;
    input \Ki[5] ;
    input \Ki[6] ;
    input \Ki[10] ;
    input \Ki[11] ;
    input [23:0]PWMLimit;
    output n363;
    input n32464;
    input [23:0]deadband;
    input VCC_net;
    output [23:0]\PID_CONTROLLER.integral ;
    input n29381;
    input [23:0]setpoint;
    input [23:0]motor_state;
    input n29915;
    input n29914;
    input n29913;
    input n29912;
    input n29911;
    input n29910;
    input n29909;
    input n29908;
    input n29907;
    input n29906;
    input n29905;
    input n29904;
    input n29903;
    input n29902;
    input n29901;
    input n29900;
    input n29899;
    input n29898;
    input n29897;
    input n29896;
    input n29895;
    input n29894;
    input n29893;
    
    wire clk16MHz /* synthesis SET_AS_NETWORK=clk16MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    wire [23:0]n1;
    
    wire n1029, n44904;
    wire [20:0]n12422;
    
    wire n661, n44905, n44, n186, n828;
    wire [21:0]n11404;
    
    wire n588, n44903, n901, n259;
    wire [21:0]n11935;
    wire [20:0]n12905;
    
    wire n45150, n45033;
    wire [15:0]n16530;
    
    wire n165, n45034, n45104;
    wire [18:0]n14585;
    
    wire n1032, n45105;
    wire [16:0]n15953;
    
    wire n23, n92, n332, n515, n44902, n405, n442, n44901, n880, 
        n369, n44900;
    wire [7:0]n19026;
    wire [6:0]n19170;
    
    wire n630, n45032, n296, n44899, n557, n45031, n223, n44898;
    wire [19:0]n13786;
    
    wire n959, n45103, n150, n44897, n484, n45030, n8, n77, 
        n45151;
    wire [19:0]n13346;
    
    wire n44896, n886, n45102, n411, n45029, n44895, n44894, n45149, 
        n44893, n813, n45101, n338, n45028, n44892, n44891, n265, 
        n45027, n45148, n1102, n44890, n1029_adj_4864, n44889, n740, 
        n45100, n192, n45026, n956, n44888, n883, n44887, n50, 
        n119, n247, n810, n44886, n737, n44885, n45147, n45146, 
        n667, n45099;
    wire [14:0]n17041;
    
    wire n45025, n974, n594, n45098, n664, n44884, n1117, n45024, 
        n530, n150_adj_4866, n159, n223_adj_4867, n603, n478, n953, 
        n1026, n311, n676, n1105, n551, n624, n1099, n1047, 
        n29029, n29330, n29024, n29019, n29014, n29009, n29004, 
        n28999, n28994, n28989, n28984, n28979, n28974, n28969, 
        n28964, n28959, n28954, n28949, n28944, n28939, n28934, 
        n28929, n28924, n28919, n1120, n697, n770;
    wire [23:0]n130;
    wire [23:0]n182;
    
    wire n181;
    wire [23:0]n207;
    
    wire n155, n83, n14, n1044, n45023, n591, n44883, n95, n26, 
        n83_adj_4869, n14_adj_4870, n156, n1026_adj_4871, n168, n156_adj_4872, 
        n229, n302, n375, n448, n241, n521, n1099_adj_4873, n229_adj_4874, 
        n314, n594_adj_4875, n384, n387, n302_adj_4876, n667_adj_4877, 
        n740_adj_4878, n518, n44882, n460, n472, n813_adj_4879, 
        n533, n74, n886_adj_4880, n5, n959_adj_4881, n606, n466, 
        n232, n296_adj_4882, n320, n1032_adj_4883, n375_adj_4884, 
        n1105_adj_4885, n445, n44881, n971, n45022, n372, n44880, 
        n305, n898, n45021, n369_adj_4886, n1038, n539;
    wire [31:0]counter;   // verilog/motorControl.v(21[11:18])
    
    wire n8_adj_4887, n6, n12, n50419, n50978, n50560, n10, n10_adj_4888, 
        n9, n51315, counter_31__N_3995, n612, n1102_adj_4889, n679, 
        n545;
    wire [23:0]n1_adj_5401;
    
    wire n752, n448_adj_4890, n80, n685, n758, n831, n618, n1111, 
        n11, n825, n521_adj_4891, n153, n904, n226, n691, n299, 
        n44879, n977, n1050, n98, n29, n764, n171, n749, n244, 
        n822, n317, n837, n390, n463;
    wire [23:0]n356;
    wire [23:0]n436;
    
    wire n10860, n28918, n28923, n28928, n910, n28933, n28938, 
        n28943, n28948, n28953, n44878, n44877, n45097, n45020;
    wire [18:0]n14186;
    
    wire n44876, n44875, n45, n45096, n45019, n41, n43, n44874, 
        n39, n35, n37, n45018, n29_adj_4899, n31, n33, n44873, 
        n44872, n393, n28958, n28963, n27, n21, n19_adj_4901, 
        n17_adj_4902, n9_adj_4903, n54925, n44871, n45145, n45095, 
        n44870, n15_adj_4904, n13_adj_4905, n11_adj_4906, n54918, 
        n28968, n12_adj_4907, n28973, n28978, n45017, n44869, n44868, 
        n45016, n28983, n28988, n10_adj_4910, n28993, n30, n54935, 
        n55311, n55307, n25, n23_adj_4912, n55758, n55512, n44867, 
        n45015, n55802, n16_adj_4913, n44866, n28998, n29003, n29008, 
        n29013, n29018, n6_adj_4915, n55586, n55587, n29023, n8_adj_4916, 
        n44865, n24, n54904, n54902, n55462, n55183, n45094, n45014, 
        n457_adj_4917, n44864, n45013, n4, n45093, n45144, n44863, 
        n41_adj_4919, n39_adj_4920, n45_adj_4921, n45012, n55584, 
        n55585, n54914, n44862, n43_adj_4922, n29_adj_4923, n31_adj_4924, 
        n37_adj_4925, n44861, n23_adj_4926, n25_adj_4927, n54912, 
        n55776, n44860, n44859, n55185;
    wire [0:0]n11428;
    wire [0:0]n10897;
    
    wire n43771;
    wire [47:0]n257;
    wire [47:0]n306;
    
    wire n43770, n11_adj_4929, n55860, n55861, n13_adj_4930, n15_adj_4931, 
        n27_adj_4932, n33_adj_4933, n9_adj_4934, n17_adj_4935, n19_adj_4936, 
        n55831, n45092, n45011, n45143, n54906, n21_adj_4937, n44858, 
        n54712, n54704, n55716, n12_adj_4938, n55191, n55794, n43769, 
        n10_adj_4939, n30_adj_4940, n41_adj_4942, n54723, n55103;
    wire [9:0]n18746;
    wire [8:0]n18945;
    
    wire n44857, n442_adj_4943, n55099, n55688, n55422, n55788, 
        n16_adj_4944, n43_adj_4945, n6_adj_4946, n55656, n44856, n45_adj_4947, 
        n55657, n8_adj_4948;
    wire [13:0]n17490;
    
    wire n45010, n24_adj_4949, n54688, n54686, n55470, n37_adj_4950, 
        n55609, n4_adj_4951, n530_adj_4952, n39_adj_4953, n35_adj_4954, 
        n55668, n55669, n45009, n44855, n44854, n54700, n54698, 
        n55812, n55611, n55890, n55891, n55853, n54690, n29_adj_4956, 
        n44853, n28710, n55734, n147_adj_4958, n895, n40, n31_adj_4959, 
        n55736, n33_adj_4960, n409, n27_adj_4961;
    wire [17:0]n15306;
    
    wire n45091, n45008, n43768, n466_adj_4962, n21_adj_4963, n19_adj_4964, 
        n17_adj_4965, n9_adj_4966, n54890, n378_adj_4967, n39_adj_4968, 
        n41_adj_4969, n45_adj_4970, n968, n15_adj_4971, n13_adj_4972, 
        n11_adj_4973, n54883, n12_adj_4974, n43_adj_4975, n37_adj_4976, 
        n29_adj_4977, n31_adj_4978, n10_adj_4979, n23_adj_4980, n25_adj_4981, 
        n539_adj_4982, n30_adj_4983, n515_adj_4984, n35_adj_4985, n33_adj_4986, 
        n11_adj_4987, n13_adj_4988, n536, n15_adj_4989, n27_adj_4990, 
        n54900, n55267, n55263, n25_adj_4991, n23_adj_4992, n55752, 
        n9_adj_4993, n17_adj_4994, n19_adj_4995, n21_adj_4996, n54672, 
        n54666, n55494, n12_adj_4997, n55800, n16_adj_4998, n10_adj_4999, 
        n30_adj_5000, n54684, n55071, n55067, n55682, n55406, n55786, 
        n6_adj_5001, n55664, n16_adj_5002, n8_adj_5003, n24_adj_5004, 
        n55665, n54646, n6_adj_5005, n55580, n54644, n55472, n55581, 
        n8_adj_5006, n44852, n55615, n4_adj_5007, n55662, n55663, 
        n54658, n54656, n55814, n44851, n24_adj_5008, n55617, n55892, 
        n54868, n54866, n55464, n44850, n1041, n55893, n55851, 
        n55193, n54648, n55740, n45007, n45090, n1114, n40_adj_5009, 
        n55742, n55743, n125_adj_5010, n56, n612_adj_5011, n41_adj_5012, 
        n39_adj_5013, n45_adj_5014, n43_adj_5015, n37_adj_5016, n21_adj_5017, 
        n45006, n23_adj_5018, n25_adj_5019, n29_adj_5020, n44849, 
        n31_adj_5021, n4_adj_5022, n55578, n55579, n113, n54878, 
        n220, n54876, n55780, n55195, n55866;
    wire [17:0]n14946;
    
    wire n44848, n17_adj_5023, n43767, n55867, n19_adj_5024, n55825, 
        n9_adj_5025, n44847, n35_adj_5026, n953_adj_5027, n45142, 
        n33_adj_5028, n11_adj_5029, n13_adj_5030, n15_adj_5031, n27_adj_5032, 
        n451_adj_5033;
    wire [23:0]n382;
    
    wire n54761, n55144, n54870, n57142, n55123, n43766, n44846, 
        n57136, n755, n45005, n45089, n55718, n54757, n55138, 
        n57157, n55134, n55201, n55796, n57151, n16_adj_5035, n54725, 
        n44845, n603_adj_5036, n43765, n8_adj_5037, n24_adj_5039, 
        n682, n45004, n54765, n1108, n44844, n57150, n54763, n57178, 
        n55450, n1035, n44843, n43764, n880_adj_5041, n45141, n962, 
        n44842;
    wire [31:0]n28;
    
    wire n44563, n44562, n44561, n44560, n609, n45003, n44559, 
        n57175, n55142, n45088, n55570, n44558, n889, n44841, 
        n54748, n57140, n55440, n43763, n293, n44557, n536_adj_5049, 
        n45002, n1108_adj_5050, n45087, n43762, n463_adj_5051, n45001, 
        n816, n44840, n44556, n743, n44839, n44555, n44554, n57168, 
        n55692, n57131, n55820, n670, n44838, n44553, n390_adj_5058, 
        n45000, n1035_adj_5059, n45086, n44552, n597, n44837, n44551, 
        n524, n44836, n57128, n54835, n44550, n44549, n12_adj_5064, 
        n317_adj_5065, n44999, n10_adj_5066, n44548, n451_adj_5068, 
        n44835, n44547, n30_adj_5070, n44546, n378_adj_5072, n44834, 
        n54864, n55229, n44545, n44544, n305_adj_5074, n44833, n807, 
        n45140, n44543, n55225, n43761, n55746, n962_adj_5076, n45085, 
        n44542, n244_adj_5078, n44998, n171_adj_5079, n44997, n44541, 
        n232_adj_5081, n44832, n44540, n55478, n55798, n6_adj_5082, 
        n55566, n16_adj_5083, n43760, n159_adj_5085, n44831, n29_adj_5086, 
        n98_adj_5087, n44539, n8_adj_5088, n24_adj_5089, n54848, n116, 
        n47, n55567, n43759, n54780, n17_adj_5091, n86, n54777, 
        n55466, n55203, n12_adj_5092, n54560, n4_adj_5094, n55670, 
        n55671, n44538, n44537, n54735, n57163, n10_adj_5096, n30_adj_5097, 
        n54738, n685_adj_5098, n113_adj_5099, n55810, n55605, n55888, 
        n55889, n44536, n6_adj_5100, n44_adj_5101;
    wire [16:0]n15630;
    
    wire n44830, n44829, n44535, n524_adj_5102, n186_adj_5103, n259_adj_5104, 
        n44534, n55672, n44828, n43758, n55673, n54727, n189_adj_5105, 
        n332_adj_5106, n44533;
    wire [5:0]n19282;
    
    wire n560, n44996, n758_adj_5108, n1111_adj_5109, n44827, n57126, 
        n55468, n55603, n43757, n55855, n54729, n366_adj_5111, n55728, 
        n405_adj_5112, n478_adj_5113, n551_adj_5114, n40_adj_5115, n4_adj_5116, 
        n55562, n262, n55563, n54828, n54826, n55808, n609_adj_5117, 
        n198_adj_5118, n55205, n55886, n55887, n55857, n54782, n55722, 
        n335_adj_5121, n624_adj_5122, n597_adj_5123, n697_adj_5124, 
        n40_adj_5125, n55724, n55730, n588_adj_5126, n487, n44995, 
        n770_adj_5127, n52322, n47_adj_5128, n43756, n1038_adj_5129, 
        n44826, n965, n44825, n734, n45139, n408, n43755, n889_adj_5130, 
        n45084, n481, n414, n44994, n43754, n892, n44824, n43753, 
        n43752, n341_adj_5132, n44993, n819, n44823, n816_adj_5133, 
        n45083, n746, n44822, n673, n44821, n43751, n43750, n600, 
        n44820, n268, n44992, n43749, n527, n44819, n43748, n43747, 
        n743_adj_5136, n45082, n454_adj_5137, n44818, n43746, n43745, 
        n381, n44817, n195_adj_5138, n44991, n43744, n554, n661_adj_5139, 
        n45138, n670_adj_5140, n45081, n53, n122_adj_5141, n43743, 
        n308, n44816, n43742, n43741, n43740, n43739, n43738, 
        n43737, n235, n44815, n162_adj_5143, n44814, n439_adj_5144;
    wire [12:0]n17881;
    
    wire n1050_adj_5145, n44990, n43736, n74_adj_5146, n5_adj_5147, 
        n43735, n512, n977_adj_5148, n44989, n43734, n43733, n676_adj_5149, 
        n147_adj_5150, n43732, n20_adj_5151, n89, n43731, n831_adj_5152, 
        n627, n220_adj_5153, n80_adj_5154;
    wire [7:0]n19106;
    
    wire n700, n44813, n43730, n43729, n11_adj_5155, n904_adj_5156, 
        n44988, n43728, n44812, n44987, n44811, n43727, n43726, 
        n293_adj_5158, n749_adj_5159, n366_adj_5160, n585, n44810, 
        n44809;
    wire [9:0]n18626;
    wire [8:0]n18846;
    
    wire n43931, n45137, n43930, n45080, n43929, n44808, n439_adj_5161, 
        n822_adj_5162, n512_adj_5163, n44807, n153_adj_5164, n895_adj_5165, 
        n43928, n43927, n585_adj_5166, n226_adj_5167, n43926, n29028, 
        n44986, n658, n658_adj_5168, n43925, n968_adj_5169, n44806, 
        n43924, n43923, n45079, n44985;
    wire [23:0]n1_adj_5402;
    wire [15:0]n16242;
    
    wire n44805, n44804, n45078, n1041_adj_5173, n44984, n44803, 
        n731, n44802, n45136, n44983, n44801, n45077, n44982, 
        n44800, n28711, n45135, n804, n44981, n682_adj_5177, n44799, 
        n44798, n45134, n45076, n110_adj_5185, n41_adj_5186, n183_adj_5187, 
        n256, n877, n329, n44980, n45133, n45075, n1114_adj_5190, 
        n950, n402_adj_5192, n1023, n44797, n475, n44796, n45132, 
        n45074, n45131, n1096, n548, n299_adj_5196, n731_adj_5198, 
        n621, n44795, n694, n767, n840, n125_adj_5200, n44979, 
        n56_adj_5201, n37221, n457_adj_5202, n44794;
    wire [23:0]n1_adj_5403;
    
    wire n198_adj_5206, n384_adj_5207, n44793, n372_adj_5208, n271, 
        n174, n44978, n804_adj_5210, n8_adj_5212, n77_adj_5213, n32, 
        n101, n344_adj_5214, n17_adj_5215, n86_adj_5216, n311_adj_5217, 
        n44792;
    wire [11:0]n18218;
    
    wire n980, n44977, n238, n44791, n165_adj_5218, n44790, n45130, 
        n700_adj_5219, n45073, n907, n44976, n834, n44975, n755_adj_5221, 
        n23_adj_5222, n92_adj_5223, n627_adj_5224, n45072, n271_adj_5225;
    wire [14:0]n16786;
    
    wire n44789, n828_adj_5226, n1117_adj_5227, n44788, n45129, n45173, 
        n1044_adj_5229, n44787, n761, n44974, n971_adj_5231, n44786, 
        n554_adj_5232, n45071, n898_adj_5233, n44785, n688, n44973, 
        n825_adj_5235, n44784, n615, n44972, n752_adj_5236, n44783, 
        n417;
    wire [3:0]n19450;
    
    wire n6_adj_5237;
    wire [4:0]n19401;
    
    wire n204, n679_adj_5238, n44782, n606_adj_5239, n44781;
    wire [1:0]n19498;
    
    wire n481_adj_5240, n45070, n533_adj_5241, n44780, n542, n44971, 
        n460_adj_5242, n44779, n45128, n387_adj_5243, n44778, n469, 
        n44970, n314_adj_5244, n44777, n45172, n241_adj_5245, n44776, 
        n131_adj_5246, n62, n45127, n408_adj_5247, n45069, n45171, 
        n335_adj_5248, n45068, n396_adj_5249, n44969, n168_adj_5250, 
        n44775, n323, n44968, n26_adj_5251, n95_adj_5252;
    wire [6:0]n19233;
    
    wire n630_adj_5253, n44774, n250, n44967, n262_adj_5254, n45067, 
        n557_adj_5255, n44773, n484_adj_5256, n44772, n45126, n177, 
        n44966, n411_adj_5257, n44771, n338_adj_5258, n44770, n265_adj_5259, 
        n44769, n35_adj_5260, n104, n490, n52332, n52334, n189_adj_5261, 
        n45066, n192_adj_5262, n44768, n50_adj_5263, n119_adj_5264, 
        n210, n51074, n490_adj_5265, n44965;
    wire [13:0]n17266;
    
    wire n1120_adj_5266, n44767, n47_adj_5267, n116_adj_5268;
    wire [4:0]n19366;
    
    wire n417_adj_5269, n44964, n1047_adj_5270, n44766, n52338, n974_adj_5271, 
        n44765, n344_adj_5272, n44963, n901_adj_5273, n44764, n43305, 
        n44763, n52342, n44962, n44762, n43878, n43877, n43876, 
        n44761, n8_adj_5274, n45065, n43875, n45064, n43874, n44961, 
        n44760, n6_adj_5275, n4_adj_5276, n50980, n44759, n43873, 
        n43872;
    wire [10:0]n18505;
    
    wire n44960, n44758, n43871, n43870, n44757, n43869, n43868, 
        n44959, n44756, n44755, n44754, n43867, n45063, n44958, 
        n43866;
    wire [12:0]n17686;
    
    wire n44753, n44752, n44957, n107_adj_5277, n45170, n38, n45125, 
        n43865, n44751, n45062, n44956, n44750, n43864, n43863, 
        n44749, n44748, n43862, n43861, n180, n89_adj_5279, n20_adj_5280, 
        n43860, n44955, n45169, n45124, n44747, n43687, n445_adj_5283, 
        n45168, n44746, n162_adj_5284, n253, n326, n45061, n44745, 
        n43686, n44954, n45123, n45167, n877_adj_5287, n399_adj_5288, 
        n44953, n393_adj_5289, n44744, n45166, n956_adj_5290, n45122, 
        n326_adj_5291, n44952, n320_adj_5292, n44743, n247_adj_5293, 
        n44742, n174_adj_5294, n44741, n253_adj_5295, n44951, n43859, 
        n32_adj_5297, n101_adj_5298, n43685, n43858, n43684;
    wire [5:0]n19330;
    
    wire n560_adj_5300, n44740, n399_adj_5301, n487_adj_5302, n44739, 
        n43857, n43683, n43682, n883_adj_5304, n45121, n43856, n414_adj_5307, 
        n44738, n235_adj_5308, n180_adj_5309, n44950, n965_adj_5310, 
        n45060, n43681, n43680, n38_adj_5311, n107_adj_5312, n341_adj_5313, 
        n44737, n1096_adj_5314, n45165, n268_adj_5316, n44736, n892_adj_5317, 
        n45059, n810_adj_5318, n45120, n43679, n195_adj_5319, n44735, 
        n43678, n819_adj_5320, n45058, n840_adj_5321, n44949, n767_adj_5322, 
        n44948, n43855, n43677, n53_adj_5324, n122_adj_5325, n43854;
    wire [11:0]n18050;
    
    wire n980_adj_5327, n44734, n43676, n907_adj_5328, n44733, n694_adj_5329, 
        n44947, n834_adj_5330, n44732, n43853, n43675, n761_adj_5332, 
        n44731, n43852, n43851, n43674, n746_adj_5335, n45057, n621_adj_5336, 
        n44946, n688_adj_5337, n44730, n615_adj_5338, n44729, n43673, 
        n548_adj_5339, n44945, n542_adj_5340, n44728, n43850, n475_adj_5342, 
        n44944, n469_adj_5343, n44727, n43849, n43672, n396_adj_5345, 
        n44726, n737_adj_5347, n45119, n323_adj_5348, n44725, n43848, 
        n1023_adj_5350, n45164, n250_adj_5351, n44724, n664_adj_5352, 
        n45118, n673_adj_5353, n45056, n472_adj_5354, n402_adj_5355, 
        n44943, n177_adj_5356, n44723, n308_adj_5357, n43847, n43671, 
        n35_adj_5359, n104_adj_5360, n545_adj_5361, n600_adj_5362, n45055, 
        n110_adj_5363, n329_adj_5364, n44942;
    wire [10:0]n18362;
    
    wire n910_adj_5365, n44722, n527_adj_5366, n45054, n41_adj_5367, 
        n837_adj_5368, n44721, n256_adj_5369, n44941, n950_adj_5370, 
        n45163, n591_adj_5371, n45117, n43846, n764_adj_5373, n44720, 
        n691_adj_5374, n44719, n454_adj_5375, n45053, n43845, n518_adj_5377, 
        n45116, n43670, n381_adj_5378, n45052, n43844, n183_adj_5380, 
        n44940, n618_adj_5381, n44718, n44717, n44939, n44938, n45051, 
        n44716;
    wire [3:0]n19426;
    
    wire n6_adj_5382, n43669, n44937, n43843, n45050, n43842, n44715, 
        n45162, n43668, n44714, n44713, n43841, n45049, n45115, 
        n43840, n44936, n43839, n43838, n44712, n44935, n44711, 
        n44710, n43837, n43836, n43835, n43667, n43666, n43834, 
        n44709, n43833, n45161, n44708, n45114, n44707, n44934, 
        n43665, n44706, n44933, n44705, n43832, n43831, n45048, 
        n44932, n44704, n43830, n44703, n45160, n43829, n45113, 
        n45047, n43828, n44702, n44931, n43827, n43826, n44701, 
        n44930, n44700, n43825, n44929, n45046, n43824, n44699, 
        n43823, n44928, n44698, n44697, n43822, n43821, n43820, 
        n43819, n43818, n43817, n43816, n44927, n43815, n43814, 
        n43813, n44926, n43812, n45045, n43811, n43810, n45044, 
        n45159, n44925;
    wire [1:0]n19490;
    
    wire n43478;
    wire [2:0]n19466;
    
    wire n43280, n45112, n44924, n45043, n45111, n44923, n45042, 
        n4_adj_5384, n44922, n43362, n45158, n44921, n45041, n44920, 
        n44919, n44918, n45040, n45157, n45110, n45156, n44917, 
        n44916, n4_adj_5385, n6_adj_5386, n45109, n45155, n45154, 
        n45039, n62_adj_5387, n131_adj_5388, n204_adj_5389, n45108, 
        n45153, n44915, n45107, n44914, n45152, n45038, n44913, 
        n45037, n44912, n45106, n44911, n45036, n44910, n45035, 
        n44909, n44908, n44907, n238_adj_5390, n807_adj_5391, n44906, 
        n734_adj_5392, n43412;
    wire [2:0]n19481;
    
    wire n4_adj_5394, n43494, n4_adj_5395, n52300, n52304, n52302, 
        n52310, n4_adj_5397, n8_adj_5398;
    
    SB_LUT4 mult_16_i692_2_lut (.I0(\Kp[14] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n1029));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i692_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5070_10 (.CI(n44904), .I0(n12422[7]), .I1(n661), .CO(n44905));
    SB_LUT4 mult_16_i30_2_lut (.I0(\Kp[0] ), .I1(n1[14]), .I2(GND_net), 
            .I3(GND_net), .O(n44));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i30_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i126_2_lut (.I0(\Kp[2] ), .I1(n1[13]), .I2(GND_net), 
            .I3(GND_net), .O(n186));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i126_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i557_2_lut (.I0(\Kp[11] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n828));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i557_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5070_9_lut (.I0(GND_net), .I1(n12422[6]), .I2(n588), .I3(n44903), 
            .O(n11404[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5070_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i606_2_lut (.I0(\Kp[12] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n901));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i606_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i175_2_lut (.I0(\Kp[3] ), .I1(n1[13]), .I2(GND_net), 
            .I3(GND_net), .O(n259));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i175_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5070_9 (.CI(n44903), .I0(n12422[6]), .I1(n588), .CO(n44904));
    SB_LUT4 add_5093_22_lut (.I0(GND_net), .I1(n12905[19]), .I2(GND_net), 
            .I3(n45150), .O(n11935[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5093_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5284_3 (.CI(n45033), .I0(n16530[0]), .I1(n165), .CO(n45034));
    SB_CARRY add_5176_15 (.CI(n45104), .I0(n14585[12]), .I1(n1032), .CO(n45105));
    SB_LUT4 add_5284_2_lut (.I0(GND_net), .I1(n23), .I2(n92), .I3(GND_net), 
            .O(n15953[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5284_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i224_2_lut (.I0(\Kp[4] ), .I1(n1[13]), .I2(GND_net), 
            .I3(GND_net), .O(n332));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i224_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5070_8_lut (.I0(GND_net), .I1(n12422[5]), .I2(n515), .I3(n44902), 
            .O(n11404[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5070_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i273_2_lut (.I0(\Kp[5] ), .I1(n1[13]), .I2(GND_net), 
            .I3(GND_net), .O(n405));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i273_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5070_8 (.CI(n44902), .I0(n12422[5]), .I1(n515), .CO(n44903));
    SB_LUT4 add_5070_7_lut (.I0(GND_net), .I1(n12422[4]), .I2(n442), .I3(n44901), 
            .O(n11404[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5070_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_i592_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n880));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i592_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5070_7 (.CI(n44901), .I0(n12422[4]), .I1(n442), .CO(n44902));
    SB_CARRY add_5284_2 (.CI(GND_net), .I0(n23), .I1(n92), .CO(n45033));
    SB_LUT4 add_5070_6_lut (.I0(GND_net), .I1(n12422[3]), .I2(n369), .I3(n44900), 
            .O(n11404[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5070_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5492_9_lut (.I0(GND_net), .I1(n19170[6]), .I2(n630), .I3(n45032), 
            .O(n19026[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5492_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5070_6 (.CI(n44900), .I0(n12422[3]), .I1(n369), .CO(n44901));
    SB_LUT4 add_5070_5_lut (.I0(GND_net), .I1(n12422[2]), .I2(n296), .I3(n44899), 
            .O(n11404[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5070_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5492_8_lut (.I0(GND_net), .I1(n19170[5]), .I2(n557), .I3(n45031), 
            .O(n19026[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5492_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5070_5 (.CI(n44899), .I0(n12422[2]), .I1(n296), .CO(n44900));
    SB_LUT4 add_5070_4_lut (.I0(GND_net), .I1(n12422[1]), .I2(n223), .I3(n44898), 
            .O(n11404[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5070_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5176_14_lut (.I0(GND_net), .I1(n14585[11]), .I2(n959), 
            .I3(n45103), .O(n13786[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5176_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5492_8 (.CI(n45031), .I0(n19170[5]), .I1(n557), .CO(n45032));
    SB_CARRY add_5070_4 (.CI(n44898), .I0(n12422[1]), .I1(n223), .CO(n44899));
    SB_LUT4 add_5070_3_lut (.I0(GND_net), .I1(n12422[0]), .I2(n150), .I3(n44897), 
            .O(n11404[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5070_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5070_3 (.CI(n44897), .I0(n12422[0]), .I1(n150), .CO(n44898));
    SB_LUT4 add_5492_7_lut (.I0(GND_net), .I1(n19170[4]), .I2(n484), .I3(n45030), 
            .O(n19026[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5492_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5070_2_lut (.I0(GND_net), .I1(n8), .I2(n77), .I3(GND_net), 
            .O(n11404[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5070_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5492_7 (.CI(n45030), .I0(n19170[4]), .I1(n484), .CO(n45031));
    SB_CARRY add_5093_22 (.CI(n45150), .I0(n12905[19]), .I1(GND_net), 
            .CO(n45151));
    SB_CARRY add_5070_2 (.CI(GND_net), .I0(n8), .I1(n77), .CO(n44897));
    SB_LUT4 add_5115_22_lut (.I0(GND_net), .I1(n13346[19]), .I2(GND_net), 
            .I3(n44896), .O(n12422[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5115_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5176_14 (.CI(n45103), .I0(n14585[11]), .I1(n959), .CO(n45104));
    SB_LUT4 add_5176_13_lut (.I0(GND_net), .I1(n14585[10]), .I2(n886), 
            .I3(n45102), .O(n13786[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5176_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5492_6_lut (.I0(GND_net), .I1(n19170[3]), .I2(n411), .I3(n45029), 
            .O(n19026[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5492_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5115_21_lut (.I0(GND_net), .I1(n13346[18]), .I2(GND_net), 
            .I3(n44895), .O(n12422[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5115_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5115_21 (.CI(n44895), .I0(n13346[18]), .I1(GND_net), 
            .CO(n44896));
    SB_LUT4 add_5115_20_lut (.I0(GND_net), .I1(n13346[17]), .I2(GND_net), 
            .I3(n44894), .O(n12422[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5115_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5492_6 (.CI(n45029), .I0(n19170[3]), .I1(n411), .CO(n45030));
    SB_LUT4 add_5093_21_lut (.I0(GND_net), .I1(n12905[18]), .I2(GND_net), 
            .I3(n45149), .O(n11935[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5093_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5176_13 (.CI(n45102), .I0(n14585[10]), .I1(n886), .CO(n45103));
    SB_CARRY add_5115_20 (.CI(n44894), .I0(n13346[17]), .I1(GND_net), 
            .CO(n44895));
    SB_LUT4 add_5115_19_lut (.I0(GND_net), .I1(n13346[16]), .I2(GND_net), 
            .I3(n44893), .O(n12422[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5115_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5093_21 (.CI(n45149), .I0(n12905[18]), .I1(GND_net), 
            .CO(n45150));
    SB_LUT4 add_5176_12_lut (.I0(GND_net), .I1(n14585[9]), .I2(n813), 
            .I3(n45101), .O(n13786[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5176_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5492_5_lut (.I0(GND_net), .I1(n19170[2]), .I2(n338), .I3(n45028), 
            .O(n19026[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5492_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5115_19 (.CI(n44893), .I0(n13346[16]), .I1(GND_net), 
            .CO(n44894));
    SB_LUT4 add_5115_18_lut (.I0(GND_net), .I1(n13346[15]), .I2(GND_net), 
            .I3(n44892), .O(n12422[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5115_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5492_5 (.CI(n45028), .I0(n19170[2]), .I1(n338), .CO(n45029));
    SB_CARRY add_5115_18 (.CI(n44892), .I0(n13346[15]), .I1(GND_net), 
            .CO(n44893));
    SB_LUT4 add_5115_17_lut (.I0(GND_net), .I1(n13346[14]), .I2(GND_net), 
            .I3(n44891), .O(n12422[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5115_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5492_4_lut (.I0(GND_net), .I1(n19170[1]), .I2(n265), .I3(n45027), 
            .O(n19026[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5492_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5093_20_lut (.I0(GND_net), .I1(n12905[17]), .I2(GND_net), 
            .I3(n45148), .O(n11935[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5093_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5176_12 (.CI(n45101), .I0(n14585[9]), .I1(n813), .CO(n45102));
    SB_CARRY add_5115_17 (.CI(n44891), .I0(n13346[14]), .I1(GND_net), 
            .CO(n44892));
    SB_CARRY add_5492_4 (.CI(n45027), .I0(n19170[1]), .I1(n265), .CO(n45028));
    SB_LUT4 add_5115_16_lut (.I0(GND_net), .I1(n13346[13]), .I2(n1102), 
            .I3(n44890), .O(n12422[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5115_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5115_16 (.CI(n44890), .I0(n13346[13]), .I1(n1102), .CO(n44891));
    SB_LUT4 add_5115_15_lut (.I0(GND_net), .I1(n13346[12]), .I2(n1029_adj_4864), 
            .I3(n44889), .O(n12422[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5115_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5115_15 (.CI(n44889), .I0(n13346[12]), .I1(n1029_adj_4864), 
            .CO(n44890));
    SB_LUT4 add_5176_11_lut (.I0(GND_net), .I1(n14585[8]), .I2(n740), 
            .I3(n45100), .O(n13786[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5176_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5492_3_lut (.I0(GND_net), .I1(n19170[0]), .I2(n192), .I3(n45026), 
            .O(n19026[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5492_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5115_14_lut (.I0(GND_net), .I1(n13346[11]), .I2(n956), 
            .I3(n44888), .O(n12422[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5115_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5115_14 (.CI(n44888), .I0(n13346[11]), .I1(n956), .CO(n44889));
    SB_LUT4 add_5115_13_lut (.I0(GND_net), .I1(n13346[10]), .I2(n883), 
            .I3(n44887), .O(n12422[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5115_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5492_3 (.CI(n45026), .I0(n19170[0]), .I1(n192), .CO(n45027));
    SB_LUT4 add_5492_2_lut (.I0(GND_net), .I1(n50), .I2(n119), .I3(GND_net), 
            .O(n19026[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5492_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i167_2_lut (.I0(\Kp[3] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n247));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i167_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5115_13 (.CI(n44887), .I0(n13346[10]), .I1(n883), .CO(n44888));
    SB_LUT4 add_5115_12_lut (.I0(GND_net), .I1(n13346[9]), .I2(n810), 
            .I3(n44886), .O(n12422[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5115_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5492_2 (.CI(GND_net), .I0(n50), .I1(n119), .CO(n45026));
    SB_CARRY add_5115_12 (.CI(n44886), .I0(n13346[9]), .I1(n810), .CO(n44887));
    SB_CARRY add_5093_20 (.CI(n45148), .I0(n12905[17]), .I1(GND_net), 
            .CO(n45149));
    SB_LUT4 add_5115_11_lut (.I0(GND_net), .I1(n13346[8]), .I2(n737), 
            .I3(n44885), .O(n12422[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5115_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5115_11 (.CI(n44885), .I0(n13346[8]), .I1(n737), .CO(n44886));
    SB_CARRY add_5176_11 (.CI(n45100), .I0(n14585[8]), .I1(n740), .CO(n45101));
    SB_LUT4 add_5093_19_lut (.I0(GND_net), .I1(n12905[16]), .I2(GND_net), 
            .I3(n45147), .O(n11935[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5093_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5093_19 (.CI(n45147), .I0(n12905[16]), .I1(GND_net), 
            .CO(n45148));
    SB_LUT4 add_5093_18_lut (.I0(GND_net), .I1(n12905[15]), .I2(GND_net), 
            .I3(n45146), .O(n11935[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5093_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5176_10_lut (.I0(GND_net), .I1(n14585[7]), .I2(n667), 
            .I3(n45099), .O(n13786[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5176_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5176_10 (.CI(n45099), .I0(n14585[7]), .I1(n667), .CO(n45100));
    SB_LUT4 add_5316_17_lut (.I0(GND_net), .I1(n17041[14]), .I2(GND_net), 
            .I3(n45025), .O(n16530[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5316_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i655_2_lut (.I0(\Kp[13] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n974));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i655_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5176_9_lut (.I0(GND_net), .I1(n14585[6]), .I2(n594), .I3(n45098), 
            .O(n13786[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5176_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5115_10_lut (.I0(GND_net), .I1(n13346[7]), .I2(n664), 
            .I3(n44884), .O(n12422[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5115_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5115_10 (.CI(n44884), .I0(n13346[7]), .I1(n664), .CO(n44885));
    SB_LUT4 add_5316_16_lut (.I0(GND_net), .I1(n17041[13]), .I2(n1117), 
            .I3(n45024), .O(n16530[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5316_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5316_16 (.CI(n45024), .I0(n17041[13]), .I1(n1117), .CO(n45025));
    SB_LUT4 mult_17_i357_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n530));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i357_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i102_2_lut (.I0(\Kp[2] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n150_adj_4866));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i102_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i108_2_lut (.I0(\Kp[2] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n159));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i108_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i151_2_lut (.I0(\Kp[3] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n223_adj_4867));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i151_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i406_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n603));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i406_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i322_2_lut (.I0(\Kp[6] ), .I1(n1[13]), .I2(GND_net), 
            .I3(GND_net), .O(n478));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i322_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i641_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n953));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i641_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i690_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n1026));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i690_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i210_2_lut (.I0(\Kp[4] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n311));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i210_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i455_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n676));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i455_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i743_2_lut (.I0(\Kp[15] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n1105));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i743_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i371_2_lut (.I0(\Kp[7] ), .I1(n1[13]), .I2(GND_net), 
            .I3(GND_net), .O(n551));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i371_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i420_2_lut (.I0(\Kp[8] ), .I1(n1[13]), .I2(GND_net), 
            .I3(GND_net), .O(n624));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i420_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i739_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n1099));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i739_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i704_2_lut (.I0(\Kp[14] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n1047));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i704_2_lut.LUT_INIT = 16'h8888;
    SB_DFFESR result__i1 (.Q(duty[1]), .C(clk16MHz), .E(control_update), 
            .D(n29029), .R(n29330));   // verilog/motorControl.v(41[14] 61[8])
    SB_DFFESR result__i2 (.Q(duty[2]), .C(clk16MHz), .E(control_update), 
            .D(n29024), .R(n29330));   // verilog/motorControl.v(41[14] 61[8])
    SB_DFFESR result__i3 (.Q(duty[3]), .C(clk16MHz), .E(control_update), 
            .D(n29019), .R(n29330));   // verilog/motorControl.v(41[14] 61[8])
    SB_DFFESR result__i4 (.Q(duty[4]), .C(clk16MHz), .E(control_update), 
            .D(n29014), .R(n29330));   // verilog/motorControl.v(41[14] 61[8])
    SB_DFFESR result__i5 (.Q(duty[5]), .C(clk16MHz), .E(control_update), 
            .D(n29009), .R(n29330));   // verilog/motorControl.v(41[14] 61[8])
    SB_DFFESR result__i6 (.Q(duty[6]), .C(clk16MHz), .E(control_update), 
            .D(n29004), .R(n29330));   // verilog/motorControl.v(41[14] 61[8])
    SB_DFFESR result__i7 (.Q(duty[7]), .C(clk16MHz), .E(control_update), 
            .D(n28999), .R(n29330));   // verilog/motorControl.v(41[14] 61[8])
    SB_DFFESR result__i8 (.Q(duty[8]), .C(clk16MHz), .E(control_update), 
            .D(n28994), .R(n29330));   // verilog/motorControl.v(41[14] 61[8])
    SB_DFFESR result__i9 (.Q(duty[9]), .C(clk16MHz), .E(control_update), 
            .D(n28989), .R(n29330));   // verilog/motorControl.v(41[14] 61[8])
    SB_DFFESR result__i10 (.Q(duty[10]), .C(clk16MHz), .E(control_update), 
            .D(n28984), .R(n29330));   // verilog/motorControl.v(41[14] 61[8])
    SB_DFFESR result__i11 (.Q(duty[11]), .C(clk16MHz), .E(control_update), 
            .D(n28979), .R(n29330));   // verilog/motorControl.v(41[14] 61[8])
    SB_DFFESR result__i12 (.Q(duty[12]), .C(clk16MHz), .E(control_update), 
            .D(n28974), .R(n29330));   // verilog/motorControl.v(41[14] 61[8])
    SB_DFFESR result__i13 (.Q(duty[13]), .C(clk16MHz), .E(control_update), 
            .D(n28969), .R(n29330));   // verilog/motorControl.v(41[14] 61[8])
    SB_DFFESR result__i14 (.Q(duty[14]), .C(clk16MHz), .E(control_update), 
            .D(n28964), .R(n29330));   // verilog/motorControl.v(41[14] 61[8])
    SB_DFFESR result__i15 (.Q(duty[15]), .C(clk16MHz), .E(control_update), 
            .D(n28959), .R(n29330));   // verilog/motorControl.v(41[14] 61[8])
    SB_DFFESR result__i16 (.Q(duty[16]), .C(clk16MHz), .E(control_update), 
            .D(n28954), .R(n29330));   // verilog/motorControl.v(41[14] 61[8])
    SB_DFFESR result__i17 (.Q(duty[17]), .C(clk16MHz), .E(control_update), 
            .D(n28949), .R(n29330));   // verilog/motorControl.v(41[14] 61[8])
    SB_DFFESR result__i18 (.Q(duty[18]), .C(clk16MHz), .E(control_update), 
            .D(n28944), .R(n29330));   // verilog/motorControl.v(41[14] 61[8])
    SB_DFFESR result__i19 (.Q(duty[19]), .C(clk16MHz), .E(control_update), 
            .D(n28939), .R(n29330));   // verilog/motorControl.v(41[14] 61[8])
    SB_DFFESR result__i20 (.Q(duty[20]), .C(clk16MHz), .E(control_update), 
            .D(n28934), .R(n29330));   // verilog/motorControl.v(41[14] 61[8])
    SB_DFFESR result__i21 (.Q(duty[21]), .C(clk16MHz), .E(control_update), 
            .D(n28929), .R(n29330));   // verilog/motorControl.v(41[14] 61[8])
    SB_DFFESR result__i22 (.Q(duty[22]), .C(clk16MHz), .E(control_update), 
            .D(n28924), .R(n29330));   // verilog/motorControl.v(41[14] 61[8])
    SB_DFFESR result__i23 (.Q(duty[23]), .C(clk16MHz), .E(control_update), 
            .D(n28919), .R(n29330));   // verilog/motorControl.v(41[14] 61[8])
    SB_LUT4 mult_16_i753_2_lut (.I0(\Kp[15] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n1120));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i753_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i469_2_lut (.I0(\Kp[9] ), .I1(n1[13]), .I2(GND_net), 
            .I3(GND_net), .O(n697));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i469_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i518_2_lut (.I0(\Kp[10] ), .I1(n1[13]), .I2(GND_net), 
            .I3(GND_net), .O(n770));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i518_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_14_i5_3_lut (.I0(n130[4]), .I1(n182[4]), .I2(n181), .I3(GND_net), 
            .O(n207[4]));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_14_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_15_i5_3_lut (.I0(n207[4]), .I1(IntegralLimit[4]), .I2(n155), 
            .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3996 [4]));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_15_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_17_i57_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n83));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i57_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i10_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n14));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i10_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5316_15_lut (.I0(GND_net), .I1(n17041[12]), .I2(n1044), 
            .I3(n45023), .O(n16530[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5316_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5115_9_lut (.I0(GND_net), .I1(n13346[6]), .I2(n591), .I3(n44883), 
            .O(n12422[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5115_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i65_2_lut (.I0(\Kp[1] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n95));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i65_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i18_2_lut (.I0(\Kp[0] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n26));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i18_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i57_2_lut (.I0(\Kp[1] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n83_adj_4869));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i57_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i10_2_lut (.I0(\Kp[0] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n14_adj_4870));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i10_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i106_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n156));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i106_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i690_2_lut (.I0(\Kp[14] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n1026_adj_4871));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i690_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i114_2_lut (.I0(\Kp[2] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n168));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i114_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i106_2_lut (.I0(\Kp[2] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n156_adj_4872));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i106_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i155_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n229));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i155_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i204_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n302));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i204_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i253_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n375));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i253_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i302_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n448));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i302_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i163_2_lut (.I0(\Kp[3] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n241));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i163_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i351_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n521));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i351_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i739_2_lut (.I0(\Kp[15] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n1099_adj_4873));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i739_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i155_2_lut (.I0(\Kp[3] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n229_adj_4874));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i155_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i212_2_lut (.I0(\Kp[4] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n314));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i212_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i400_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n594_adj_4875));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i400_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i259_2_lut (.I0(\Kp[5] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n384));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i259_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i261_2_lut (.I0(\Kp[5] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n387));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i261_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i204_2_lut (.I0(\Kp[4] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n302_adj_4876));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i204_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5316_15 (.CI(n45023), .I0(n17041[12]), .I1(n1044), .CO(n45024));
    SB_CARRY add_5115_9 (.CI(n44883), .I0(n13346[6]), .I1(n591), .CO(n44884));
    SB_LUT4 mult_17_i449_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n667_adj_4877));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i449_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i498_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n740_adj_4878));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i498_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5115_8_lut (.I0(GND_net), .I1(n13346[5]), .I2(n518), .I3(n44882), 
            .O(n12422[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5115_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i310_2_lut (.I0(\Kp[6] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n460));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i310_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i318_2_lut (.I0(\Kp[6] ), .I1(n1[11]), .I2(GND_net), 
            .I3(GND_net), .O(n472));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i318_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i547_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n813_adj_4879));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i547_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i359_2_lut (.I0(\Kp[7] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n533));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i359_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i51_2_lut (.I0(\Kp[1] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n74));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i51_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i596_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n886_adj_4880));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i596_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i4_2_lut (.I0(\Kp[0] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n5));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i4_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i645_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n959_adj_4881));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i645_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i408_2_lut (.I0(\Kp[8] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n606));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i408_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i314_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n466));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i314_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i157_2_lut (.I0(\Kp[3] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n232));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i157_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i200_2_lut (.I0(\Kp[4] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n296_adj_4882));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i200_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i216_2_lut (.I0(\Kp[4] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n320));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i216_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i694_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n1032_adj_4883));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i694_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i253_2_lut (.I0(\Kp[5] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n375_adj_4884));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i253_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i743_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n1105_adj_4885));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i743_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5115_8 (.CI(n44882), .I0(n13346[5]), .I1(n518), .CO(n44883));
    SB_LUT4 add_5115_7_lut (.I0(GND_net), .I1(n13346[4]), .I2(n445), .I3(n44881), 
            .O(n12422[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5115_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5176_9 (.CI(n45098), .I0(n14585[6]), .I1(n594), .CO(n45099));
    SB_LUT4 add_5316_14_lut (.I0(GND_net), .I1(n17041[11]), .I2(n971), 
            .I3(n45022), .O(n16530[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5316_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5316_14 (.CI(n45022), .I0(n17041[11]), .I1(n971), .CO(n45023));
    SB_CARRY add_5115_7 (.CI(n44881), .I0(n13346[4]), .I1(n445), .CO(n44882));
    SB_LUT4 add_5115_6_lut (.I0(GND_net), .I1(n13346[3]), .I2(n372), .I3(n44880), 
            .O(n12422[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5115_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i206_2_lut (.I0(\Kp[4] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n305));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i206_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5316_13_lut (.I0(GND_net), .I1(n17041[10]), .I2(n898), 
            .I3(n45021), .O(n16530[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5316_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5115_6 (.CI(n44880), .I0(n13346[3]), .I1(n372), .CO(n44881));
    SB_LUT4 mult_16_i249_2_lut (.I0(\Kp[5] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n369_adj_4886));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i249_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i698_2_lut (.I0(\Kp[14] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n1038));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i698_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i363_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n539));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i363_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i3_3_lut (.I0(counter[19]), .I1(counter[29]), .I2(counter[28]), 
            .I3(GND_net), .O(n8_adj_4887));
    defparam i3_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_4_lut (.I0(counter[24]), .I1(counter[30]), .I2(n8_adj_4887), 
            .I3(counter[27]), .O(n6));
    defparam i1_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i5_4_lut (.I0(counter[4]), .I1(counter[6]), .I2(counter[1]), 
            .I3(counter[3]), .O(n12));
    defparam i5_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i6_4_lut (.I0(counter[5]), .I1(n12), .I2(counter[2]), .I3(counter[0]), 
            .O(n50419));
    defparam i6_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i4_4_lut (.I0(counter[16]), .I1(counter[14]), .I2(counter[20]), 
            .I3(n6), .O(n50978));
    defparam i4_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i3_4_lut (.I0(counter[23]), .I1(counter[15]), .I2(counter[26]), 
            .I3(counter[25]), .O(n50560));
    defparam i3_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i4_4_lut_adj_1677 (.I0(n50560), .I1(counter[17]), .I2(n50978), 
            .I3(counter[21]), .O(n10));
    defparam i4_4_lut_adj_1677.LUT_INIT = 16'hfffe;
    SB_LUT4 i4_4_lut_adj_1678 (.I0(counter[13]), .I1(counter[9]), .I2(counter[10]), 
            .I3(counter[11]), .O(n10_adj_4888));
    defparam i4_4_lut_adj_1678.LUT_INIT = 16'h8000;
    SB_LUT4 i3_4_lut_adj_1679 (.I0(counter[12]), .I1(n50419), .I2(counter[8]), 
            .I3(counter[7]), .O(n9));
    defparam i3_4_lut_adj_1679.LUT_INIT = 16'ha8a0;
    SB_LUT4 i5_3_lut (.I0(counter[22]), .I1(n10), .I2(counter[18]), .I3(GND_net), 
            .O(n51315));
    defparam i5_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i22597_4_lut (.I0(n51315), .I1(counter[31]), .I2(n9), .I3(n10_adj_4888), 
            .O(counter_31__N_3995));   // verilog/motorControl.v(26[8:41])
    defparam i22597_4_lut.LUT_INIT = 16'h3222;
    SB_LUT4 mult_17_i412_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n612));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i412_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i741_2_lut (.I0(\Kp[15] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n1102_adj_4889));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i741_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i457_2_lut (.I0(\Kp[9] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n679));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i457_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i367_2_lut (.I0(\Kp[7] ), .I1(n1[11]), .I2(GND_net), 
            .I3(GND_net), .O(n545));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i367_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_26_inv_0_i6_1_lut (.I0(PWMLimit[5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5401[5]));   // verilog/motorControl.v(55[22:31])
    defparam unary_minus_26_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_16_i506_2_lut (.I0(\Kp[10] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n752));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i506_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i302_2_lut (.I0(\Kp[6] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n448_adj_4890));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i302_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_14_i4_3_lut (.I0(n130[3]), .I1(n182[3]), .I2(n181), .I3(GND_net), 
            .O(n207[3]));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_14_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_15_i4_3_lut (.I0(n207[3]), .I1(IntegralLimit[3]), .I2(n155), 
            .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3996 [3]));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_15_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_26_inv_0_i7_1_lut (.I0(PWMLimit[6]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5401[6]));   // verilog/motorControl.v(55[22:31])
    defparam unary_minus_26_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_26_inv_0_i8_1_lut (.I0(PWMLimit[7]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5401[7]));   // verilog/motorControl.v(55[22:31])
    defparam unary_minus_26_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_17_i55_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n80));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i55_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i461_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n685));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i461_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i510_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n758));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i510_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_26_inv_0_i9_1_lut (.I0(PWMLimit[8]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5401[8]));   // verilog/motorControl.v(55[22:31])
    defparam unary_minus_26_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_26_inv_0_i10_1_lut (.I0(PWMLimit[9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5401[9]));   // verilog/motorControl.v(55[22:31])
    defparam unary_minus_26_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_17_i559_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n831));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i559_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i416_2_lut (.I0(\Kp[8] ), .I1(n1[11]), .I2(GND_net), 
            .I3(GND_net), .O(n618));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i416_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i747_2_lut (.I0(\Kp[15] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n1111));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i747_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i8_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n11));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i8_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i555_2_lut (.I0(\Kp[11] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n825));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i555_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i351_2_lut (.I0(\Kp[7] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n521_adj_4891));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i351_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i104_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n153));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i104_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i608_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n904));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i608_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_26_inv_0_i11_1_lut (.I0(PWMLimit[10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5401[10]));   // verilog/motorControl.v(55[22:31])
    defparam unary_minus_26_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_17_i153_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n226));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i153_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i465_2_lut (.I0(\Kp[9] ), .I1(n1[11]), .I2(GND_net), 
            .I3(GND_net), .O(n691));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i465_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5115_5_lut (.I0(GND_net), .I1(n13346[2]), .I2(n299), .I3(n44879), 
            .O(n12422[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5115_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_i657_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n977));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i657_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i706_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n1050));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i706_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_14_i10_3_lut (.I0(n130[9]), .I1(n182[9]), .I2(n181), .I3(GND_net), 
            .O(n207[9]));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_14_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_15_i10_3_lut (.I0(n207[9]), .I1(IntegralLimit[9]), .I2(n155), 
            .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3996 [9]));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_15_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_17_i67_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n98));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i67_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i20_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n29));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i20_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_26_inv_0_i12_1_lut (.I0(PWMLimit[11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5401[11]));   // verilog/motorControl.v(55[22:31])
    defparam unary_minus_26_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_16_i514_2_lut (.I0(\Kp[10] ), .I1(n1[11]), .I2(GND_net), 
            .I3(GND_net), .O(n764));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i514_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i202_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n299));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i202_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_26_inv_0_i13_1_lut (.I0(PWMLimit[12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5401[12]));   // verilog/motorControl.v(55[22:31])
    defparam unary_minus_26_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_17_i116_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n171));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i116_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i504_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n749));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i504_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i604_2_lut (.I0(\Kp[12] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n898));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i604_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i251_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n372));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i251_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i653_2_lut (.I0(\Kp[13] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n971));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i653_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i165_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n244));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i165_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i553_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n822));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i553_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i300_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n445));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i300_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i349_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n518));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i349_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i398_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n591));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i398_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i702_2_lut (.I0(\Kp[14] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n1044));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i702_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i214_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n317));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i214_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i563_2_lut (.I0(\Kp[11] ), .I1(n1[11]), .I2(GND_net), 
            .I3(GND_net), .O(n837));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i563_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i396_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n588));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i396_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_26_inv_0_i14_1_lut (.I0(PWMLimit[13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5401[13]));   // verilog/motorControl.v(55[22:31])
    defparam unary_minus_26_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_26_inv_0_i15_1_lut (.I0(PWMLimit[14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5401[14]));   // verilog/motorControl.v(55[22:31])
    defparam unary_minus_26_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_17_i263_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n390));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i263_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_26_inv_0_i16_1_lut (.I0(PWMLimit[15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5401[15]));   // verilog/motorControl.v(55[22:31])
    defparam unary_minus_26_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_26_inv_0_i17_1_lut (.I0(PWMLimit[16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5401[16]));   // verilog/motorControl.v(55[22:31])
    defparam unary_minus_26_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_17_i312_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n463));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i312_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i14847_3_lut (.I0(n356[23]), .I1(n436[23]), .I2(n10860), .I3(GND_net), 
            .O(n28918));   // verilog/motorControl.v(41[14] 61[8])
    defparam i14847_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14852_3_lut (.I0(n356[22]), .I1(n436[22]), .I2(n10860), .I3(GND_net), 
            .O(n28923));   // verilog/motorControl.v(41[14] 61[8])
    defparam i14852_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14857_3_lut (.I0(n356[21]), .I1(n436[21]), .I2(n10860), .I3(GND_net), 
            .O(n28928));   // verilog/motorControl.v(41[14] 61[8])
    defparam i14857_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_16_i612_2_lut (.I0(\Kp[12] ), .I1(n1[11]), .I2(GND_net), 
            .I3(GND_net), .O(n910));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i612_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_26_inv_0_i18_1_lut (.I0(PWMLimit[17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5401[17]));   // verilog/motorControl.v(55[22:31])
    defparam unary_minus_26_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i14862_3_lut (.I0(n356[20]), .I1(n436[20]), .I2(n10860), .I3(GND_net), 
            .O(n28933));   // verilog/motorControl.v(41[14] 61[8])
    defparam i14862_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14867_3_lut (.I0(n356[19]), .I1(n436[19]), .I2(n10860), .I3(GND_net), 
            .O(n28938));   // verilog/motorControl.v(41[14] 61[8])
    defparam i14867_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14872_3_lut (.I0(n356[18]), .I1(n436[18]), .I2(n10860), .I3(GND_net), 
            .O(n28943));   // verilog/motorControl.v(41[14] 61[8])
    defparam i14872_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14877_3_lut (.I0(n363), .I1(n436[17]), .I2(n10860), .I3(GND_net), 
            .O(n28948));   // verilog/motorControl.v(41[14] 61[8])
    defparam i14877_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14882_3_lut (.I0(n356[16]), .I1(n436[16]), .I2(n10860), .I3(GND_net), 
            .O(n28953));   // verilog/motorControl.v(41[14] 61[8])
    defparam i14882_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_5115_5 (.CI(n44879), .I0(n13346[2]), .I1(n299), .CO(n44880));
    SB_CARRY add_5316_13 (.CI(n45021), .I0(n17041[10]), .I1(n898), .CO(n45022));
    SB_LUT4 add_5115_4_lut (.I0(GND_net), .I1(n13346[1]), .I2(n226), .I3(n44878), 
            .O(n12422[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5115_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5115_4 (.CI(n44878), .I0(n13346[1]), .I1(n226), .CO(n44879));
    SB_LUT4 add_5115_3_lut (.I0(GND_net), .I1(n13346[0]), .I2(n153), .I3(n44877), 
            .O(n12422[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5115_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5115_3 (.CI(n44877), .I0(n13346[0]), .I1(n153), .CO(n44878));
    SB_LUT4 add_5176_8_lut (.I0(GND_net), .I1(n14585[5]), .I2(n521_adj_4891), 
            .I3(n45097), .O(n13786[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5176_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5316_12_lut (.I0(GND_net), .I1(n17041[9]), .I2(n825), 
            .I3(n45020), .O(n16530[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5316_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5115_2_lut (.I0(GND_net), .I1(n11), .I2(n80), .I3(GND_net), 
            .O(n12422[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5115_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5093_18 (.CI(n45146), .I0(n12905[15]), .I1(GND_net), 
            .CO(n45147));
    SB_CARRY add_5115_2 (.CI(GND_net), .I0(n11), .I1(n80), .CO(n44877));
    SB_CARRY add_5176_8 (.CI(n45097), .I0(n14585[5]), .I1(n521_adj_4891), 
            .CO(n45098));
    SB_LUT4 add_5156_21_lut (.I0(GND_net), .I1(n14186[18]), .I2(GND_net), 
            .I3(n44876), .O(n13346[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5156_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5156_20_lut (.I0(GND_net), .I1(n14186[17]), .I2(GND_net), 
            .I3(n44875), .O(n13346[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5156_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5316_12 (.CI(n45020), .I0(n17041[9]), .I1(n825), .CO(n45021));
    SB_CARRY add_5156_20 (.CI(n44875), .I0(n14186[17]), .I1(GND_net), 
            .CO(n44876));
    SB_LUT4 LessThan_10_i45_2_lut (.I0(IntegralLimit[22]), .I1(n130[22]), 
            .I2(GND_net), .I3(GND_net), .O(n45));   // verilog/motorControl.v(45[12:34])
    defparam LessThan_10_i45_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_5176_7_lut (.I0(GND_net), .I1(n14585[4]), .I2(n448_adj_4890), 
            .I3(n45096), .O(n13786[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5176_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5316_11_lut (.I0(GND_net), .I1(n17041[8]), .I2(n752), 
            .I3(n45019), .O(n16530[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5316_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_10_i41_2_lut (.I0(IntegralLimit[20]), .I1(n130[20]), 
            .I2(GND_net), .I3(GND_net), .O(n41));   // verilog/motorControl.v(45[12:34])
    defparam LessThan_10_i41_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_5316_11 (.CI(n45019), .I0(n17041[8]), .I1(n752), .CO(n45020));
    SB_LUT4 LessThan_10_i43_2_lut (.I0(IntegralLimit[21]), .I1(n130[21]), 
            .I2(GND_net), .I3(GND_net), .O(n43));   // verilog/motorControl.v(45[12:34])
    defparam LessThan_10_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_5156_19_lut (.I0(GND_net), .I1(n14186[16]), .I2(GND_net), 
            .I3(n44874), .O(n13346[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5156_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_10_i39_2_lut (.I0(IntegralLimit[19]), .I1(n130[19]), 
            .I2(GND_net), .I3(GND_net), .O(n39));   // verilog/motorControl.v(45[12:34])
    defparam LessThan_10_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_10_i35_2_lut (.I0(IntegralLimit[17]), .I1(n130[17]), 
            .I2(GND_net), .I3(GND_net), .O(n35));   // verilog/motorControl.v(45[12:34])
    defparam LessThan_10_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_10_i37_2_lut (.I0(IntegralLimit[18]), .I1(n130[18]), 
            .I2(GND_net), .I3(GND_net), .O(n37));   // verilog/motorControl.v(45[12:34])
    defparam LessThan_10_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_5316_10_lut (.I0(GND_net), .I1(n17041[7]), .I2(n679), 
            .I3(n45018), .O(n16530[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5316_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_10_i29_2_lut (.I0(IntegralLimit[14]), .I1(n130[14]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_4899));   // verilog/motorControl.v(45[12:34])
    defparam LessThan_10_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_10_i31_2_lut (.I0(IntegralLimit[15]), .I1(n130[15]), 
            .I2(GND_net), .I3(GND_net), .O(n31));   // verilog/motorControl.v(45[12:34])
    defparam LessThan_10_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_10_i33_2_lut (.I0(IntegralLimit[16]), .I1(n130[16]), 
            .I2(GND_net), .I3(GND_net), .O(n33));   // verilog/motorControl.v(45[12:34])
    defparam LessThan_10_i33_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_5156_19 (.CI(n44874), .I0(n14186[16]), .I1(GND_net), 
            .CO(n44875));
    SB_LUT4 add_5156_18_lut (.I0(GND_net), .I1(n14186[15]), .I2(GND_net), 
            .I3(n44873), .O(n13346[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5156_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5156_18 (.CI(n44873), .I0(n14186[15]), .I1(GND_net), 
            .CO(n44874));
    SB_DFF control_update_37 (.Q(control_update), .C(clk16MHz), .D(counter_31__N_3995));   // verilog/motorControl.v(23[10] 30[6])
    SB_CARRY add_5316_10 (.CI(n45018), .I0(n17041[7]), .I1(n679), .CO(n45019));
    SB_LUT4 add_5156_17_lut (.I0(GND_net), .I1(n14186[14]), .I2(GND_net), 
            .I3(n44872), .O(n13346[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5156_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i265_2_lut (.I0(\Kp[5] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n393));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i265_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i14887_3_lut (.I0(n356[15]), .I1(n436[15]), .I2(n10860), .I3(GND_net), 
            .O(n28958));   // verilog/motorControl.v(41[14] 61[8])
    defparam i14887_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14892_3_lut (.I0(n356[14]), .I1(n436[14]), .I2(n10860), .I3(GND_net), 
            .O(n28963));   // verilog/motorControl.v(41[14] 61[8])
    defparam i14892_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_5156_17 (.CI(n44872), .I0(n14186[14]), .I1(GND_net), 
            .CO(n44873));
    SB_LUT4 LessThan_10_i27_2_lut (.I0(IntegralLimit[13]), .I1(n130[13]), 
            .I2(GND_net), .I3(GND_net), .O(n27));   // verilog/motorControl.v(45[12:34])
    defparam LessThan_10_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i39095_4_lut (.I0(n21), .I1(n19_adj_4901), .I2(n17_adj_4902), 
            .I3(n9_adj_4903), .O(n54925));
    defparam i39095_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 add_5156_16_lut (.I0(GND_net), .I1(n14186[13]), .I2(n1105_adj_4885), 
            .I3(n44871), .O(n13346[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5156_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5156_16 (.CI(n44871), .I0(n14186[13]), .I1(n1105_adj_4885), 
            .CO(n44872));
    SB_LUT4 add_5093_17_lut (.I0(GND_net), .I1(n12905[14]), .I2(GND_net), 
            .I3(n45145), .O(n11935[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5093_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5176_7 (.CI(n45096), .I0(n14585[4]), .I1(n448_adj_4890), 
            .CO(n45097));
    SB_LUT4 add_5176_6_lut (.I0(GND_net), .I1(n14585[3]), .I2(n375_adj_4884), 
            .I3(n45095), .O(n13786[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5176_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5156_15_lut (.I0(GND_net), .I1(n14186[12]), .I2(n1032_adj_4883), 
            .I3(n44870), .O(n13346[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5156_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i39088_4_lut (.I0(n27), .I1(n15_adj_4904), .I2(n13_adj_4905), 
            .I3(n11_adj_4906), .O(n54918));
    defparam i39088_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i14897_3_lut (.I0(n356[13]), .I1(n436[13]), .I2(n10860), .I3(GND_net), 
            .O(n28968));   // verilog/motorControl.v(41[14] 61[8])
    defparam i14897_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_10_i12_3_lut (.I0(n130[7]), .I1(n130[16]), .I2(n33), 
            .I3(GND_net), .O(n12_adj_4907));   // verilog/motorControl.v(45[12:34])
    defparam LessThan_10_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14902_3_lut (.I0(n356[12]), .I1(n436[12]), .I2(n10860), .I3(GND_net), 
            .O(n28973));   // verilog/motorControl.v(41[14] 61[8])
    defparam i14902_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14907_3_lut (.I0(n356[11]), .I1(n436[11]), .I2(n10860), .I3(GND_net), 
            .O(n28978));   // verilog/motorControl.v(41[14] 61[8])
    defparam i14907_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_5316_9_lut (.I0(GND_net), .I1(n17041[6]), .I2(n606), .I3(n45017), 
            .O(n16530[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5316_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5156_15 (.CI(n44870), .I0(n14186[12]), .I1(n1032_adj_4883), 
            .CO(n44871));
    SB_CARRY add_5316_9 (.CI(n45017), .I0(n17041[6]), .I1(n606), .CO(n45018));
    SB_LUT4 add_5156_14_lut (.I0(GND_net), .I1(n14186[11]), .I2(n959_adj_4881), 
            .I3(n44869), .O(n13346[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5156_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5156_14 (.CI(n44869), .I0(n14186[11]), .I1(n959_adj_4881), 
            .CO(n44870));
    SB_LUT4 add_5156_13_lut (.I0(GND_net), .I1(n14186[10]), .I2(n886_adj_4880), 
            .I3(n44868), .O(n13346[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5156_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5156_13 (.CI(n44868), .I0(n14186[10]), .I1(n886_adj_4880), 
            .CO(n44869));
    SB_CARRY add_5176_6 (.CI(n45095), .I0(n14585[3]), .I1(n375_adj_4884), 
            .CO(n45096));
    SB_LUT4 add_5316_8_lut (.I0(GND_net), .I1(n17041[5]), .I2(n533), .I3(n45016), 
            .O(n16530[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5316_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14912_3_lut (.I0(n356[10]), .I1(n436[10]), .I2(n10860), .I3(GND_net), 
            .O(n28983));   // verilog/motorControl.v(41[14] 61[8])
    defparam i14912_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14917_3_lut (.I0(n356[9]), .I1(n436[9]), .I2(n10860), .I3(GND_net), 
            .O(n28988));   // verilog/motorControl.v(41[14] 61[8])
    defparam i14917_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_10_i10_3_lut (.I0(n130[5]), .I1(n130[6]), .I2(n13_adj_4905), 
            .I3(GND_net), .O(n10_adj_4910));   // verilog/motorControl.v(45[12:34])
    defparam LessThan_10_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_5316_8 (.CI(n45016), .I0(n17041[5]), .I1(n533), .CO(n45017));
    SB_LUT4 i14922_3_lut (.I0(n356[8]), .I1(n436[8]), .I2(n10860), .I3(GND_net), 
            .O(n28993));   // verilog/motorControl.v(41[14] 61[8])
    defparam i14922_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_10_i30_3_lut (.I0(n12_adj_4907), .I1(n130[17]), .I2(n35), 
            .I3(GND_net), .O(n30));   // verilog/motorControl.v(45[12:34])
    defparam LessThan_10_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i39480_4_lut (.I0(n13_adj_4905), .I1(n11_adj_4906), .I2(n9_adj_4903), 
            .I3(n54935), .O(n55311));
    defparam i39480_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i39476_4_lut (.I0(n19_adj_4901), .I1(n17_adj_4902), .I2(n15_adj_4904), 
            .I3(n55311), .O(n55307));
    defparam i39476_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i39927_4_lut (.I0(n25), .I1(n23_adj_4912), .I2(n21), .I3(n55307), 
            .O(n55758));
    defparam i39927_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i39681_4_lut (.I0(n31), .I1(n29_adj_4899), .I2(n27), .I3(n55758), 
            .O(n55512));
    defparam i39681_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 add_5156_12_lut (.I0(GND_net), .I1(n14186[9]), .I2(n813_adj_4879), 
            .I3(n44867), .O(n13346[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5156_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5316_7_lut (.I0(GND_net), .I1(n17041[4]), .I2(n460), .I3(n45015), 
            .O(n16530[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5316_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i39971_4_lut (.I0(n37), .I1(n35), .I2(n33), .I3(n55512), 
            .O(n55802));
    defparam i39971_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 LessThan_10_i16_3_lut (.I0(n130[9]), .I1(n130[21]), .I2(n43), 
            .I3(GND_net), .O(n16_adj_4913));   // verilog/motorControl.v(45[12:34])
    defparam LessThan_10_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_5316_7 (.CI(n45015), .I0(n17041[4]), .I1(n460), .CO(n45016));
    SB_CARRY add_5156_12 (.CI(n44867), .I0(n14186[9]), .I1(n813_adj_4879), 
            .CO(n44868));
    SB_LUT4 add_5156_11_lut (.I0(GND_net), .I1(n14186[8]), .I2(n740_adj_4878), 
            .I3(n44866), .O(n13346[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5156_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14927_3_lut (.I0(n356[7]), .I1(n436[7]), .I2(n10860), .I3(GND_net), 
            .O(n28998));   // verilog/motorControl.v(41[14] 61[8])
    defparam i14927_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14932_3_lut (.I0(n356[6]), .I1(n436[6]), .I2(n10860), .I3(GND_net), 
            .O(n29003));   // verilog/motorControl.v(41[14] 61[8])
    defparam i14932_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14937_3_lut (.I0(n356[5]), .I1(n436[5]), .I2(n10860), .I3(GND_net), 
            .O(n29008));   // verilog/motorControl.v(41[14] 61[8])
    defparam i14937_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14942_3_lut (.I0(n356[4]), .I1(n436[4]), .I2(n10860), .I3(GND_net), 
            .O(n29013));   // verilog/motorControl.v(41[14] 61[8])
    defparam i14942_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14947_3_lut (.I0(n356[3]), .I1(n436[3]), .I2(n10860), .I3(GND_net), 
            .O(n29018));   // verilog/motorControl.v(41[14] 61[8])
    defparam i14947_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i39755_3_lut (.I0(n6_adj_4915), .I1(n130[10]), .I2(n21), .I3(GND_net), 
            .O(n55586));   // verilog/motorControl.v(45[12:34])
    defparam i39755_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i39756_3_lut (.I0(n55586), .I1(n130[11]), .I2(n23_adj_4912), 
            .I3(GND_net), .O(n55587));   // verilog/motorControl.v(45[12:34])
    defparam i39756_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_5156_11 (.CI(n44866), .I0(n14186[8]), .I1(n740_adj_4878), 
            .CO(n44867));
    SB_LUT4 i14952_3_lut (.I0(n356[2]), .I1(n436[2]), .I2(n10860), .I3(GND_net), 
            .O(n29023));   // verilog/motorControl.v(41[14] 61[8])
    defparam i14952_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_10_i8_3_lut (.I0(n130[4]), .I1(n130[8]), .I2(n17_adj_4902), 
            .I3(GND_net), .O(n8_adj_4916));   // verilog/motorControl.v(45[12:34])
    defparam LessThan_10_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_5156_10_lut (.I0(GND_net), .I1(n14186[7]), .I2(n667_adj_4877), 
            .I3(n44865), .O(n13346[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5156_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_10_i24_3_lut (.I0(n16_adj_4913), .I1(n130[22]), .I2(n45), 
            .I3(GND_net), .O(n24));   // verilog/motorControl.v(45[12:34])
    defparam LessThan_10_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i39074_4_lut (.I0(n43), .I1(n25), .I2(n23_adj_4912), .I3(n54925), 
            .O(n54904));
    defparam i39074_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i39631_4_lut (.I0(n24), .I1(n8_adj_4916), .I2(n45), .I3(n54902), 
            .O(n55462));   // verilog/motorControl.v(45[12:34])
    defparam i39631_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i39352_3_lut (.I0(n55587), .I1(n130[12]), .I2(n25), .I3(GND_net), 
            .O(n55183));   // verilog/motorControl.v(45[12:34])
    defparam i39352_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_5156_10 (.CI(n44865), .I0(n14186[7]), .I1(n667_adj_4877), 
            .CO(n44866));
    SB_LUT4 add_5176_5_lut (.I0(GND_net), .I1(n14585[2]), .I2(n302_adj_4876), 
            .I3(n45094), .O(n13786[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5176_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5316_6_lut (.I0(GND_net), .I1(n17041[3]), .I2(n387), .I3(n45014), 
            .O(n16530[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5316_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i308_2_lut (.I0(\Kp[6] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n457_adj_4917));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i308_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5156_9_lut (.I0(GND_net), .I1(n14186[6]), .I2(n594_adj_4875), 
            .I3(n44864), .O(n13346[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5156_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5093_17 (.CI(n45145), .I0(n12905[14]), .I1(GND_net), 
            .CO(n45146));
    SB_CARRY add_5176_5 (.CI(n45094), .I0(n14585[2]), .I1(n302_adj_4876), 
            .CO(n45095));
    SB_CARRY add_5156_9 (.CI(n44864), .I0(n14186[6]), .I1(n594_adj_4875), 
            .CO(n44865));
    SB_CARRY add_5316_6 (.CI(n45014), .I0(n17041[3]), .I1(n387), .CO(n45015));
    SB_LUT4 add_5316_5_lut (.I0(GND_net), .I1(n17041[2]), .I2(n314), .I3(n45013), 
            .O(n16530[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5316_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_10_i4_4_lut (.I0(n130[0]), .I1(n130[1]), .I2(IntegralLimit[1]), 
            .I3(IntegralLimit[0]), .O(n4));   // verilog/motorControl.v(45[12:34])
    defparam LessThan_10_i4_4_lut.LUT_INIT = 16'h0c8e;
    SB_LUT4 add_5176_4_lut (.I0(GND_net), .I1(n14585[1]), .I2(n229_adj_4874), 
            .I3(n45093), .O(n13786[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5176_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5093_16_lut (.I0(GND_net), .I1(n12905[13]), .I2(n1099_adj_4873), 
            .I3(n45144), .O(n11935[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5093_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5176_4 (.CI(n45093), .I0(n14585[1]), .I1(n229_adj_4874), 
            .CO(n45094));
    SB_LUT4 add_5156_8_lut (.I0(GND_net), .I1(n14186[5]), .I2(n521), .I3(n44863), 
            .O(n13346[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5156_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5316_5 (.CI(n45013), .I0(n17041[2]), .I1(n314), .CO(n45014));
    SB_LUT4 LessThan_23_i41_2_lut (.I0(PWMLimit[20]), .I1(n356[20]), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4919));   // verilog/motorControl.v(52[14:29])
    defparam LessThan_23_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_23_i39_2_lut (.I0(PWMLimit[19]), .I1(n356[19]), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4920));   // verilog/motorControl.v(52[14:29])
    defparam LessThan_23_i39_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_5156_8 (.CI(n44863), .I0(n14186[5]), .I1(n521), .CO(n44864));
    SB_LUT4 LessThan_23_i45_2_lut (.I0(PWMLimit[22]), .I1(n356[22]), .I2(GND_net), 
            .I3(GND_net), .O(n45_adj_4921));   // verilog/motorControl.v(52[14:29])
    defparam LessThan_23_i45_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_5316_4_lut (.I0(GND_net), .I1(n17041[1]), .I2(n241), .I3(n45012), 
            .O(n16530[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5316_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i39753_3_lut (.I0(n4), .I1(n130[13]), .I2(n27), .I3(GND_net), 
            .O(n55584));   // verilog/motorControl.v(45[12:34])
    defparam i39753_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i39754_3_lut (.I0(n55584), .I1(n130[14]), .I2(n29_adj_4899), 
            .I3(GND_net), .O(n55585));   // verilog/motorControl.v(45[12:34])
    defparam i39754_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i39084_4_lut (.I0(n33), .I1(n31), .I2(n29_adj_4899), .I3(n54918), 
            .O(n54914));
    defparam i39084_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 add_5156_7_lut (.I0(GND_net), .I1(n14186[4]), .I2(n448), .I3(n44862), 
            .O(n13346[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5156_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_23_i43_2_lut (.I0(PWMLimit[21]), .I1(n356[21]), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_4922));   // verilog/motorControl.v(52[14:29])
    defparam LessThan_23_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_23_i29_2_lut (.I0(PWMLimit[14]), .I1(n356[14]), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4923));   // verilog/motorControl.v(52[14:29])
    defparam LessThan_23_i29_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_5156_7 (.CI(n44862), .I0(n14186[4]), .I1(n448), .CO(n44863));
    SB_LUT4 LessThan_23_i31_2_lut (.I0(PWMLimit[15]), .I1(n356[15]), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_4924));   // verilog/motorControl.v(52[14:29])
    defparam LessThan_23_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_23_i37_2_lut (.I0(PWMLimit[18]), .I1(n356[18]), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_4925));   // verilog/motorControl.v(52[14:29])
    defparam LessThan_23_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_5156_6_lut (.I0(GND_net), .I1(n14186[3]), .I2(n375), .I3(n44861), 
            .O(n13346[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5156_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_23_i23_2_lut (.I0(PWMLimit[11]), .I1(n356[11]), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_4926));   // verilog/motorControl.v(52[14:29])
    defparam LessThan_23_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_23_i25_2_lut (.I0(PWMLimit[12]), .I1(n356[12]), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_4927));   // verilog/motorControl.v(52[14:29])
    defparam LessThan_23_i25_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_5156_6 (.CI(n44861), .I0(n14186[3]), .I1(n375), .CO(n44862));
    SB_LUT4 i39945_4_lut (.I0(n30), .I1(n10_adj_4910), .I2(n35), .I3(n54912), 
            .O(n55776));   // verilog/motorControl.v(45[12:34])
    defparam i39945_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 add_5156_5_lut (.I0(GND_net), .I1(n14186[2]), .I2(n302), .I3(n44860), 
            .O(n13346[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5156_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5156_5 (.CI(n44860), .I0(n14186[2]), .I1(n302), .CO(n44861));
    SB_CARRY add_5316_4 (.CI(n45012), .I0(n17041[1]), .I1(n241), .CO(n45013));
    SB_LUT4 add_5156_4_lut (.I0(GND_net), .I1(n14186[1]), .I2(n229), .I3(n44859), 
            .O(n13346[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5156_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5093_16 (.CI(n45144), .I0(n12905[13]), .I1(n1099_adj_4873), 
            .CO(n45145));
    SB_CARRY add_5156_4 (.CI(n44859), .I0(n14186[1]), .I1(n229), .CO(n44860));
    SB_LUT4 i39354_3_lut (.I0(n55585), .I1(n130[15]), .I2(n31), .I3(GND_net), 
            .O(n55185));   // verilog/motorControl.v(45[12:34])
    defparam i39354_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_18_25_lut (.I0(GND_net), .I1(n11428[0]), .I2(n10897[0]), 
            .I3(n43771), .O(n356[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_18_24_lut (.I0(GND_net), .I1(n257[22]), .I2(n306[22]), 
            .I3(n43770), .O(n356[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_23_i11_2_lut (.I0(PWMLimit[5]), .I1(n356[5]), .I2(GND_net), 
            .I3(GND_net), .O(n11_adj_4929));   // verilog/motorControl.v(52[14:29])
    defparam LessThan_23_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i40029_4_lut (.I0(n55185), .I1(n55776), .I2(n35), .I3(n54914), 
            .O(n55860));   // verilog/motorControl.v(45[12:34])
    defparam i40029_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i40030_3_lut (.I0(n55860), .I1(n130[18]), .I2(n37), .I3(GND_net), 
            .O(n55861));   // verilog/motorControl.v(45[12:34])
    defparam i40030_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_23_i13_2_lut (.I0(PWMLimit[6]), .I1(n356[6]), .I2(GND_net), 
            .I3(GND_net), .O(n13_adj_4930));   // verilog/motorControl.v(52[14:29])
    defparam LessThan_23_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_23_i15_2_lut (.I0(PWMLimit[7]), .I1(n356[7]), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_4931));   // verilog/motorControl.v(52[14:29])
    defparam LessThan_23_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_23_i27_2_lut (.I0(PWMLimit[13]), .I1(n356[13]), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_4932));   // verilog/motorControl.v(52[14:29])
    defparam LessThan_23_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_23_i33_2_lut (.I0(PWMLimit[16]), .I1(n356[16]), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_4933));   // verilog/motorControl.v(52[14:29])
    defparam LessThan_23_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_23_i9_2_lut (.I0(PWMLimit[4]), .I1(n356[4]), .I2(GND_net), 
            .I3(GND_net), .O(n9_adj_4934));   // verilog/motorControl.v(52[14:29])
    defparam LessThan_23_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_23_i17_2_lut (.I0(PWMLimit[8]), .I1(n356[8]), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_4935));   // verilog/motorControl.v(52[14:29])
    defparam LessThan_23_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_23_i19_2_lut (.I0(PWMLimit[9]), .I1(n356[9]), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_4936));   // verilog/motorControl.v(52[14:29])
    defparam LessThan_23_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i40000_3_lut (.I0(n55861), .I1(n130[19]), .I2(n39), .I3(GND_net), 
            .O(n55831));   // verilog/motorControl.v(45[12:34])
    defparam i40000_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_5176_3_lut (.I0(GND_net), .I1(n14585[0]), .I2(n156_adj_4872), 
            .I3(n45092), .O(n13786[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5176_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5316_3_lut (.I0(GND_net), .I1(n17041[0]), .I2(n168), .I3(n45011), 
            .O(n16530[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5316_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5093_15_lut (.I0(GND_net), .I1(n12905[12]), .I2(n1026_adj_4871), 
            .I3(n45143), .O(n11935[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5093_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i39076_4_lut (.I0(n43), .I1(n41), .I2(n39), .I3(n55802), 
            .O(n54906));
    defparam i39076_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 LessThan_23_i21_2_lut (.I0(PWMLimit[10]), .I1(n356[10]), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_4937));   // verilog/motorControl.v(52[14:29])
    defparam LessThan_23_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_5156_3_lut (.I0(GND_net), .I1(n14186[0]), .I2(n156), .I3(n44858), 
            .O(n13346[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5156_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i38882_4_lut (.I0(n21_adj_4937), .I1(n19_adj_4936), .I2(n17_adj_4935), 
            .I3(n9_adj_4934), .O(n54712));
    defparam i38882_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i38874_4_lut (.I0(n27_adj_4932), .I1(n15_adj_4931), .I2(n13_adj_4930), 
            .I3(n11_adj_4929), .O(n54704));
    defparam i38874_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i39885_4_lut (.I0(n55183), .I1(n55462), .I2(n45), .I3(n54904), 
            .O(n55716));   // verilog/motorControl.v(45[12:34])
    defparam i39885_4_lut.LUT_INIT = 16'hccca;
    SB_CARRY add_5176_3 (.CI(n45092), .I0(n14585[0]), .I1(n156_adj_4872), 
            .CO(n45093));
    SB_LUT4 LessThan_23_i12_3_lut (.I0(n356[7]), .I1(n356[16]), .I2(n33_adj_4933), 
            .I3(GND_net), .O(n12_adj_4938));   // verilog/motorControl.v(52[14:29])
    defparam LessThan_23_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_5316_3 (.CI(n45011), .I0(n17041[0]), .I1(n168), .CO(n45012));
    SB_CARRY add_5156_3 (.CI(n44858), .I0(n14186[0]), .I1(n156), .CO(n44859));
    SB_LUT4 add_5176_2_lut (.I0(GND_net), .I1(n14_adj_4870), .I2(n83_adj_4869), 
            .I3(GND_net), .O(n13786[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5176_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i39360_3_lut (.I0(n55831), .I1(n130[20]), .I2(n41), .I3(GND_net), 
            .O(n55191));   // verilog/motorControl.v(45[12:34])
    defparam i39360_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_18_24 (.CI(n43770), .I0(n257[22]), .I1(n306[22]), .CO(n43771));
    SB_LUT4 i39963_4_lut (.I0(n55191), .I1(n55716), .I2(n45), .I3(n54906), 
            .O(n55794));   // verilog/motorControl.v(45[12:34])
    defparam i39963_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 add_18_23_lut (.I0(GND_net), .I1(n257[21]), .I2(n306[21]), 
            .I3(n43769), .O(n356[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5316_2_lut (.I0(GND_net), .I1(n26), .I2(n95), .I3(GND_net), 
            .O(n16530[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5316_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_23_i10_3_lut (.I0(n356[5]), .I1(n356[6]), .I2(n13_adj_4930), 
            .I3(GND_net), .O(n10_adj_4939));   // verilog/motorControl.v(52[14:29])
    defparam LessThan_23_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i39964_3_lut (.I0(n55794), .I1(IntegralLimit[23]), .I2(n130[23]), 
            .I3(GND_net), .O(n155));   // verilog/motorControl.v(45[12:34])
    defparam i39964_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 LessThan_23_i30_3_lut (.I0(n12_adj_4938), .I1(n363), .I2(n32464), 
            .I3(GND_net), .O(n30_adj_4940));   // verilog/motorControl.v(52[14:29])
    defparam LessThan_23_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_5156_2_lut (.I0(GND_net), .I1(n14), .I2(n83), .I3(GND_net), 
            .O(n13346[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5156_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5316_2 (.CI(GND_net), .I0(n26), .I1(n95), .CO(n45011));
    SB_LUT4 LessThan_12_i41_2_lut (.I0(n130[20]), .I1(n182[20]), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4942));   // verilog/motorControl.v(47[21:44])
    defparam LessThan_12_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i39273_4_lut (.I0(n13_adj_4930), .I1(n11_adj_4929), .I2(n9_adj_4934), 
            .I3(n54723), .O(n55103));
    defparam i39273_4_lut.LUT_INIT = 16'heeef;
    SB_CARRY add_5156_2 (.CI(GND_net), .I0(n14), .I1(n83), .CO(n44858));
    SB_LUT4 add_5466_11_lut (.I0(GND_net), .I1(n18945[8]), .I2(n770), 
            .I3(n44857), .O(n18746[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5466_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i298_2_lut (.I0(\Kp[6] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n442_adj_4943));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i298_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i39269_4_lut (.I0(n19_adj_4936), .I1(n17_adj_4935), .I2(n15_adj_4931), 
            .I3(n55103), .O(n55099));
    defparam i39269_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i39857_4_lut (.I0(n25_adj_4927), .I1(n23_adj_4926), .I2(n21_adj_4937), 
            .I3(n55099), .O(n55688));
    defparam i39857_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i39591_4_lut (.I0(n31_adj_4924), .I1(n29_adj_4923), .I2(n27_adj_4932), 
            .I3(n55688), .O(n55422));
    defparam i39591_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i39957_4_lut (.I0(n37_adj_4925), .I1(n32464), .I2(n33_adj_4933), 
            .I3(n55422), .O(n55788));
    defparam i39957_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 LessThan_23_i16_3_lut (.I0(n356[9]), .I1(n356[21]), .I2(n43_adj_4922), 
            .I3(GND_net), .O(n16_adj_4944));   // verilog/motorControl.v(52[14:29])
    defparam LessThan_23_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_12_i43_2_lut (.I0(n130[21]), .I1(n182[21]), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_4945));   // verilog/motorControl.v(47[21:44])
    defparam LessThan_12_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i39825_3_lut (.I0(n6_adj_4946), .I1(n356[10]), .I2(n21_adj_4937), 
            .I3(GND_net), .O(n55656));   // verilog/motorControl.v(52[14:29])
    defparam i39825_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_5466_10_lut (.I0(GND_net), .I1(n18945[7]), .I2(n697), 
            .I3(n44856), .O(n18746[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5466_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_12_i45_2_lut (.I0(n130[22]), .I1(n182[22]), .I2(GND_net), 
            .I3(GND_net), .O(n45_adj_4947));   // verilog/motorControl.v(47[21:44])
    defparam LessThan_12_i45_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i39826_3_lut (.I0(n55656), .I1(n356[11]), .I2(n23_adj_4926), 
            .I3(GND_net), .O(n55657));   // verilog/motorControl.v(52[14:29])
    defparam i39826_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_23_i8_3_lut (.I0(n356[4]), .I1(n356[8]), .I2(n17_adj_4935), 
            .I3(GND_net), .O(n8_adj_4948));   // verilog/motorControl.v(52[14:29])
    defparam LessThan_23_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_5346_16_lut (.I0(GND_net), .I1(n17490[13]), .I2(n1120), 
            .I3(n45010), .O(n17041[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5346_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5466_10 (.CI(n44856), .I0(n18945[7]), .I1(n697), .CO(n44857));
    SB_LUT4 LessThan_23_i24_3_lut (.I0(n16_adj_4944), .I1(n356[22]), .I2(n45_adj_4921), 
            .I3(GND_net), .O(n24_adj_4949));   // verilog/motorControl.v(52[14:29])
    defparam LessThan_23_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i38858_4_lut (.I0(n43_adj_4922), .I1(n25_adj_4927), .I2(n23_adj_4926), 
            .I3(n54712), .O(n54688));
    defparam i38858_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i39639_4_lut (.I0(n24_adj_4949), .I1(n8_adj_4948), .I2(n45_adj_4921), 
            .I3(n54686), .O(n55470));   // verilog/motorControl.v(52[14:29])
    defparam i39639_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 LessThan_12_i37_2_lut (.I0(n130[18]), .I1(n182[18]), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_4950));   // verilog/motorControl.v(47[21:44])
    defparam LessThan_12_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i39778_3_lut (.I0(n55657), .I1(n356[12]), .I2(n25_adj_4927), 
            .I3(GND_net), .O(n55609));   // verilog/motorControl.v(52[14:29])
    defparam i39778_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_23_i4_4_lut (.I0(PWMLimit[0]), .I1(n356[1]), .I2(PWMLimit[1]), 
            .I3(n356[0]), .O(n4_adj_4951));   // verilog/motorControl.v(52[14:29])
    defparam LessThan_23_i4_4_lut.LUT_INIT = 16'h4d0c;
    SB_LUT4 mult_16_i357_2_lut (.I0(\Kp[7] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n530_adj_4952));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i357_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_12_i39_2_lut (.I0(n130[19]), .I1(n182[19]), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4953));   // verilog/motorControl.v(47[21:44])
    defparam LessThan_12_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_12_i35_2_lut (.I0(n130[17]), .I1(n182[17]), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4954));   // verilog/motorControl.v(47[21:44])
    defparam LessThan_12_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i39837_3_lut (.I0(n4_adj_4951), .I1(n356[13]), .I2(n27_adj_4932), 
            .I3(GND_net), .O(n55668));   // verilog/motorControl.v(52[14:29])
    defparam i39837_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i39838_3_lut (.I0(n55668), .I1(n356[14]), .I2(n29_adj_4923), 
            .I3(GND_net), .O(n55669));   // verilog/motorControl.v(52[14:29])
    defparam i39838_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_5346_15_lut (.I0(GND_net), .I1(n17490[12]), .I2(n1047), 
            .I3(n45009), .O(n17041[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5346_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5466_9_lut (.I0(GND_net), .I1(n18945[6]), .I2(n624), .I3(n44855), 
            .O(n18746[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5466_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5466_9 (.CI(n44855), .I0(n18945[6]), .I1(n624), .CO(n44856));
    SB_CARRY add_5346_15 (.CI(n45009), .I0(n17490[12]), .I1(n1047), .CO(n45010));
    SB_LUT4 add_5466_8_lut (.I0(GND_net), .I1(n18945[5]), .I2(n551), .I3(n44854), 
            .O(n18746[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5466_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i38870_4_lut (.I0(n33_adj_4933), .I1(n31_adj_4924), .I2(n29_adj_4923), 
            .I3(n54704), .O(n54700));
    defparam i38870_4_lut.LUT_INIT = 16'haaab;
    SB_CARRY add_5466_8 (.CI(n44854), .I0(n18945[5]), .I1(n551), .CO(n44855));
    SB_LUT4 i39981_4_lut (.I0(n30_adj_4940), .I1(n10_adj_4939), .I2(n32464), 
            .I3(n54698), .O(n55812));   // verilog/motorControl.v(52[14:29])
    defparam i39981_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i39780_3_lut (.I0(n55669), .I1(n356[15]), .I2(n31_adj_4924), 
            .I3(GND_net), .O(n55611));   // verilog/motorControl.v(52[14:29])
    defparam i39780_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_18_23 (.CI(n43769), .I0(n257[21]), .I1(n306[21]), .CO(n43770));
    SB_LUT4 i40059_4_lut (.I0(n55611), .I1(n55812), .I2(n32464), .I3(n54700), 
            .O(n55890));   // verilog/motorControl.v(52[14:29])
    defparam i40059_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i40060_3_lut (.I0(n55890), .I1(n356[18]), .I2(n37_adj_4925), 
            .I3(GND_net), .O(n55891));   // verilog/motorControl.v(52[14:29])
    defparam i40060_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i40022_3_lut (.I0(n55891), .I1(n356[19]), .I2(n39_adj_4920), 
            .I3(GND_net), .O(n55853));   // verilog/motorControl.v(52[14:29])
    defparam i40022_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i38860_4_lut (.I0(n43_adj_4922), .I1(n41_adj_4919), .I2(n39_adj_4920), 
            .I3(n55788), .O(n54690));
    defparam i38860_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 LessThan_12_i29_2_lut (.I0(n130[14]), .I1(n182[14]), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4956));   // verilog/motorControl.v(47[21:44])
    defparam LessThan_12_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_5466_7_lut (.I0(GND_net), .I1(n18945[4]), .I2(n478), .I3(n44853), 
            .O(n18746[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5466_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14639_3_lut (.I0(n356[0]), .I1(n436[0]), .I2(n10860), .I3(GND_net), 
            .O(n28710));   // verilog/motorControl.v(41[14] 61[8])
    defparam i14639_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i39903_4_lut (.I0(n55609), .I1(n55470), .I2(n45_adj_4921), 
            .I3(n54688), .O(n55734));   // verilog/motorControl.v(52[14:29])
    defparam i39903_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 mult_16_i100_2_lut (.I0(\Kp[2] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n147_adj_4958));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i100_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i602_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n895));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i602_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i40008_3_lut (.I0(n55853), .I1(n356[20]), .I2(n41_adj_4919), 
            .I3(GND_net), .O(n40));   // verilog/motorControl.v(52[14:29])
    defparam i40008_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_12_i31_2_lut (.I0(n130[15]), .I1(n182[15]), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_4959));   // verilog/motorControl.v(47[21:44])
    defparam LessThan_12_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i39905_4_lut (.I0(n40), .I1(n55734), .I2(n45_adj_4921), .I3(n54690), 
            .O(n55736));   // verilog/motorControl.v(52[14:29])
    defparam i39905_4_lut.LUT_INIT = 16'hccca;
    SB_CARRY add_5466_7 (.CI(n44853), .I0(n18945[4]), .I1(n478), .CO(n44854));
    SB_LUT4 LessThan_12_i33_2_lut (.I0(n130[16]), .I1(n182[16]), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_4960));   // verilog/motorControl.v(47[21:44])
    defparam LessThan_12_i33_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_5176_2 (.CI(GND_net), .I0(n14_adj_4870), .I1(n83_adj_4869), 
            .CO(n45092));
    SB_LUT4 i39906_3_lut (.I0(n55736), .I1(PWMLimit[23]), .I2(n356[23]), 
            .I3(GND_net), .O(n409));   // verilog/motorControl.v(52[14:29])
    defparam i39906_3_lut.LUT_INIT = 16'h8e8e;
    SB_CARRY add_5093_15 (.CI(n45143), .I0(n12905[12]), .I1(n1026_adj_4871), 
            .CO(n45144));
    SB_LUT4 LessThan_12_i27_2_lut (.I0(n130[13]), .I1(n182[13]), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_4961));   // verilog/motorControl.v(47[21:44])
    defparam LessThan_12_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_5214_20_lut (.I0(GND_net), .I1(n15306[17]), .I2(GND_net), 
            .I3(n45091), .O(n14585[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5214_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5346_14_lut (.I0(GND_net), .I1(n17490[11]), .I2(n974), 
            .I3(n45008), .O(n17041[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5346_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_18_22_lut (.I0(GND_net), .I1(n257[20]), .I2(n306[20]), 
            .I3(n43768), .O(n356[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i314_2_lut (.I0(\Kp[6] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n466_adj_4962));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i314_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_18_22 (.CI(n43768), .I0(n257[20]), .I1(n306[20]), .CO(n43769));
    SB_LUT4 i39060_4_lut (.I0(n21_adj_4963), .I1(n19_adj_4964), .I2(n17_adj_4965), 
            .I3(n9_adj_4966), .O(n54890));
    defparam i39060_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 mult_16_i255_2_lut (.I0(\Kp[5] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n378_adj_4967));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i255_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_25_i39_2_lut (.I0(n356[19]), .I1(n436[19]), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4968));   // verilog/motorControl.v(54[23:39])
    defparam LessThan_25_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_25_i41_2_lut (.I0(n356[20]), .I1(n436[20]), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4969));   // verilog/motorControl.v(54[23:39])
    defparam LessThan_25_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_25_i45_2_lut (.I0(n356[22]), .I1(n436[22]), .I2(GND_net), 
            .I3(GND_net), .O(n45_adj_4970));   // verilog/motorControl.v(54[23:39])
    defparam LessThan_25_i45_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_17_i651_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n968));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i651_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i39053_4_lut (.I0(n27_adj_4961), .I1(n15_adj_4971), .I2(n13_adj_4972), 
            .I3(n11_adj_4973), .O(n54883));
    defparam i39053_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 LessThan_12_i12_3_lut (.I0(n182[7]), .I1(n182[16]), .I2(n33_adj_4960), 
            .I3(GND_net), .O(n12_adj_4974));   // verilog/motorControl.v(47[21:44])
    defparam LessThan_12_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_25_i43_2_lut (.I0(n356[21]), .I1(n436[21]), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_4975));   // verilog/motorControl.v(54[23:39])
    defparam LessThan_25_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_25_i37_2_lut (.I0(n356[18]), .I1(n436[18]), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_4976));   // verilog/motorControl.v(54[23:39])
    defparam LessThan_25_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_25_i29_2_lut (.I0(n356[14]), .I1(n436[14]), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4977));   // verilog/motorControl.v(54[23:39])
    defparam LessThan_25_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_25_i31_2_lut (.I0(n356[15]), .I1(n436[15]), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_4978));   // verilog/motorControl.v(54[23:39])
    defparam LessThan_25_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_12_i10_3_lut (.I0(n182[5]), .I1(n182[6]), .I2(n13_adj_4972), 
            .I3(GND_net), .O(n10_adj_4979));   // verilog/motorControl.v(47[21:44])
    defparam LessThan_12_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_25_i23_2_lut (.I0(n356[11]), .I1(n436[11]), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_4980));   // verilog/motorControl.v(54[23:39])
    defparam LessThan_25_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_25_i25_2_lut (.I0(n356[12]), .I1(n436[12]), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_4981));   // verilog/motorControl.v(54[23:39])
    defparam LessThan_25_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_16_i363_2_lut (.I0(\Kp[7] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n539_adj_4982));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i363_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_12_i30_3_lut (.I0(n12_adj_4974), .I1(n182[17]), .I2(n35_adj_4954), 
            .I3(GND_net), .O(n30_adj_4983));   // verilog/motorControl.v(47[21:44])
    defparam LessThan_12_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_16_i347_2_lut (.I0(\Kp[7] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n515_adj_4984));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i347_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_25_i35_2_lut (.I0(n363), .I1(n436[17]), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4985));   // verilog/motorControl.v(54[23:39])
    defparam LessThan_25_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_25_i33_2_lut (.I0(n356[16]), .I1(n436[16]), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_4986));   // verilog/motorControl.v(54[23:39])
    defparam LessThan_25_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_25_i11_2_lut (.I0(n356[5]), .I1(n436[5]), .I2(GND_net), 
            .I3(GND_net), .O(n11_adj_4987));   // verilog/motorControl.v(54[23:39])
    defparam LessThan_25_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 unary_minus_26_inv_0_i19_1_lut (.I0(PWMLimit[18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5401[18]));   // verilog/motorControl.v(55[22:31])
    defparam unary_minus_26_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 LessThan_25_i13_2_lut (.I0(n356[6]), .I1(n436[6]), .I2(GND_net), 
            .I3(GND_net), .O(n13_adj_4988));   // verilog/motorControl.v(54[23:39])
    defparam LessThan_25_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_17_i361_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n536));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i361_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_25_i15_2_lut (.I0(n356[7]), .I1(n436[7]), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_4989));   // verilog/motorControl.v(54[23:39])
    defparam LessThan_25_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_25_i27_2_lut (.I0(n356[13]), .I1(n436[13]), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_4990));   // verilog/motorControl.v(54[23:39])
    defparam LessThan_25_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i39436_4_lut (.I0(n13_adj_4972), .I1(n11_adj_4973), .I2(n9_adj_4966), 
            .I3(n54900), .O(n55267));
    defparam i39436_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i39432_4_lut (.I0(n19_adj_4964), .I1(n17_adj_4965), .I2(n15_adj_4971), 
            .I3(n55267), .O(n55263));
    defparam i39432_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i39921_4_lut (.I0(n25_adj_4991), .I1(n23_adj_4992), .I2(n21_adj_4963), 
            .I3(n55263), .O(n55752));
    defparam i39921_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 LessThan_25_i9_2_lut (.I0(n356[4]), .I1(n436[4]), .I2(GND_net), 
            .I3(GND_net), .O(n9_adj_4993));   // verilog/motorControl.v(54[23:39])
    defparam LessThan_25_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_25_i17_2_lut (.I0(n356[8]), .I1(n436[8]), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_4994));   // verilog/motorControl.v(54[23:39])
    defparam LessThan_25_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_25_i19_2_lut (.I0(n356[9]), .I1(n436[9]), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_4995));   // verilog/motorControl.v(54[23:39])
    defparam LessThan_25_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_25_i21_2_lut (.I0(n356[10]), .I1(n436[10]), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_4996));   // verilog/motorControl.v(54[23:39])
    defparam LessThan_25_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i38842_4_lut (.I0(n21_adj_4996), .I1(n19_adj_4995), .I2(n17_adj_4994), 
            .I3(n9_adj_4993), .O(n54672));
    defparam i38842_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i38836_4_lut (.I0(n27_adj_4990), .I1(n15_adj_4989), .I2(n13_adj_4988), 
            .I3(n11_adj_4987), .O(n54666));
    defparam i38836_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i39663_4_lut (.I0(n31_adj_4959), .I1(n29_adj_4956), .I2(n27_adj_4961), 
            .I3(n55752), .O(n55494));
    defparam i39663_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 LessThan_25_i12_3_lut (.I0(n436[7]), .I1(n436[16]), .I2(n33_adj_4986), 
            .I3(GND_net), .O(n12_adj_4997));   // verilog/motorControl.v(54[23:39])
    defparam LessThan_25_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i39969_4_lut (.I0(n37_adj_4950), .I1(n35_adj_4954), .I2(n33_adj_4960), 
            .I3(n55494), .O(n55800));
    defparam i39969_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 LessThan_12_i16_3_lut (.I0(n182[9]), .I1(n182[21]), .I2(n43_adj_4945), 
            .I3(GND_net), .O(n16_adj_4998));   // verilog/motorControl.v(47[21:44])
    defparam LessThan_12_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_25_i10_3_lut (.I0(n436[5]), .I1(n436[6]), .I2(n13_adj_4988), 
            .I3(GND_net), .O(n10_adj_4999));   // verilog/motorControl.v(54[23:39])
    defparam LessThan_25_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_25_i30_3_lut (.I0(n12_adj_4997), .I1(n436[17]), .I2(n35_adj_4985), 
            .I3(GND_net), .O(n30_adj_5000));   // verilog/motorControl.v(54[23:39])
    defparam LessThan_25_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i39241_4_lut (.I0(n13_adj_4988), .I1(n11_adj_4987), .I2(n9_adj_4993), 
            .I3(n54684), .O(n55071));
    defparam i39241_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i39237_4_lut (.I0(n19_adj_4995), .I1(n17_adj_4994), .I2(n15_adj_4989), 
            .I3(n55071), .O(n55067));
    defparam i39237_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i39851_4_lut (.I0(n25_adj_4981), .I1(n23_adj_4980), .I2(n21_adj_4996), 
            .I3(n55067), .O(n55682));
    defparam i39851_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i39575_4_lut (.I0(n31_adj_4978), .I1(n29_adj_4977), .I2(n27_adj_4990), 
            .I3(n55682), .O(n55406));
    defparam i39575_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i39955_4_lut (.I0(n37_adj_4976), .I1(n35_adj_4985), .I2(n33_adj_4986), 
            .I3(n55406), .O(n55786));
    defparam i39955_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i39833_3_lut (.I0(n6_adj_5001), .I1(n436[10]), .I2(n21_adj_4996), 
            .I3(GND_net), .O(n55664));   // verilog/motorControl.v(54[23:39])
    defparam i39833_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_25_i16_3_lut (.I0(n436[9]), .I1(n436[21]), .I2(n43_adj_4975), 
            .I3(GND_net), .O(n16_adj_5002));   // verilog/motorControl.v(54[23:39])
    defparam LessThan_25_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_25_i8_3_lut (.I0(n436[4]), .I1(n436[8]), .I2(n17_adj_4994), 
            .I3(GND_net), .O(n8_adj_5003));   // verilog/motorControl.v(54[23:39])
    defparam LessThan_25_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_25_i24_3_lut (.I0(n16_adj_5002), .I1(n436[22]), .I2(n45_adj_4970), 
            .I3(GND_net), .O(n24_adj_5004));   // verilog/motorControl.v(54[23:39])
    defparam LessThan_25_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i39834_3_lut (.I0(n55664), .I1(n436[11]), .I2(n23_adj_4980), 
            .I3(GND_net), .O(n55665));   // verilog/motorControl.v(54[23:39])
    defparam i39834_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i38816_4_lut (.I0(n43_adj_4975), .I1(n25_adj_4981), .I2(n23_adj_4980), 
            .I3(n54672), .O(n54646));
    defparam i38816_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i39749_3_lut (.I0(n6_adj_5005), .I1(n182[10]), .I2(n21_adj_4963), 
            .I3(GND_net), .O(n55580));   // verilog/motorControl.v(47[21:44])
    defparam i39749_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i39641_4_lut (.I0(n24_adj_5004), .I1(n8_adj_5003), .I2(n45_adj_4970), 
            .I3(n54644), .O(n55472));   // verilog/motorControl.v(54[23:39])
    defparam i39641_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i39750_3_lut (.I0(n55580), .I1(n182[11]), .I2(n23_adj_4992), 
            .I3(GND_net), .O(n55581));   // verilog/motorControl.v(47[21:44])
    defparam i39750_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_12_i8_3_lut (.I0(n182[4]), .I1(n182[8]), .I2(n17_adj_4965), 
            .I3(GND_net), .O(n8_adj_5006));   // verilog/motorControl.v(47[21:44])
    defparam LessThan_12_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_5346_14 (.CI(n45008), .I0(n17490[11]), .I1(n974), .CO(n45009));
    SB_LUT4 add_5466_6_lut (.I0(GND_net), .I1(n18945[3]), .I2(n405), .I3(n44852), 
            .O(n18746[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5466_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5466_6 (.CI(n44852), .I0(n18945[3]), .I1(n405), .CO(n44853));
    SB_LUT4 i39784_3_lut (.I0(n55665), .I1(n436[12]), .I2(n25_adj_4981), 
            .I3(GND_net), .O(n55615));   // verilog/motorControl.v(54[23:39])
    defparam i39784_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_25_i4_4_lut (.I0(n436[0]), .I1(n436[1]), .I2(n356[1]), 
            .I3(n356[0]), .O(n4_adj_5007));   // verilog/motorControl.v(54[23:39])
    defparam LessThan_25_i4_4_lut.LUT_INIT = 16'h0c8e;
    SB_LUT4 i39831_3_lut (.I0(n4_adj_5007), .I1(n436[13]), .I2(n27_adj_4990), 
            .I3(GND_net), .O(n55662));   // verilog/motorControl.v(54[23:39])
    defparam i39831_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i39832_3_lut (.I0(n55662), .I1(n436[14]), .I2(n29_adj_4977), 
            .I3(GND_net), .O(n55663));   // verilog/motorControl.v(54[23:39])
    defparam i39832_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i38828_4_lut (.I0(n33_adj_4986), .I1(n31_adj_4978), .I2(n29_adj_4977), 
            .I3(n54666), .O(n54658));
    defparam i38828_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i39983_4_lut (.I0(n30_adj_5000), .I1(n10_adj_4999), .I2(n35_adj_4985), 
            .I3(n54656), .O(n55814));   // verilog/motorControl.v(54[23:39])
    defparam i39983_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 add_5466_5_lut (.I0(GND_net), .I1(n18945[2]), .I2(n332), .I3(n44851), 
            .O(n18746[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5466_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_12_i24_3_lut (.I0(n16_adj_4998), .I1(n182[22]), .I2(n45_adj_4947), 
            .I3(GND_net), .O(n24_adj_5008));   // verilog/motorControl.v(47[21:44])
    defparam LessThan_12_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i39786_3_lut (.I0(n55663), .I1(n436[15]), .I2(n31_adj_4978), 
            .I3(GND_net), .O(n55617));   // verilog/motorControl.v(54[23:39])
    defparam i39786_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i40061_4_lut (.I0(n55617), .I1(n55814), .I2(n35_adj_4985), 
            .I3(n54658), .O(n55892));   // verilog/motorControl.v(54[23:39])
    defparam i40061_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i39038_4_lut (.I0(n43_adj_4945), .I1(n25_adj_4991), .I2(n23_adj_4992), 
            .I3(n54890), .O(n54868));
    defparam i39038_4_lut.LUT_INIT = 16'haaab;
    SB_CARRY add_5466_5 (.CI(n44851), .I0(n18945[2]), .I1(n332), .CO(n44852));
    SB_LUT4 i39633_4_lut (.I0(n24_adj_5008), .I1(n8_adj_5006), .I2(n45_adj_4947), 
            .I3(n54866), .O(n55464));   // verilog/motorControl.v(47[21:44])
    defparam i39633_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 add_5466_4_lut (.I0(GND_net), .I1(n18945[1]), .I2(n259), .I3(n44850), 
            .O(n18746[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5466_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_i700_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n1041));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i700_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i40062_3_lut (.I0(n55892), .I1(n436[18]), .I2(n37_adj_4976), 
            .I3(GND_net), .O(n55893));   // verilog/motorControl.v(54[23:39])
    defparam i40062_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i40020_3_lut (.I0(n55893), .I1(n436[19]), .I2(n39_adj_4968), 
            .I3(GND_net), .O(n55851));   // verilog/motorControl.v(54[23:39])
    defparam i40020_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i39362_3_lut (.I0(n55581), .I1(n182[12]), .I2(n25_adj_4991), 
            .I3(GND_net), .O(n55193));   // verilog/motorControl.v(47[21:44])
    defparam i39362_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i38818_4_lut (.I0(n43_adj_4975), .I1(n41_adj_4969), .I2(n39_adj_4968), 
            .I3(n55786), .O(n54648));
    defparam i38818_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i39909_4_lut (.I0(n55615), .I1(n55472), .I2(n45_adj_4970), 
            .I3(n54646), .O(n55740));   // verilog/motorControl.v(54[23:39])
    defparam i39909_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 add_5346_13_lut (.I0(GND_net), .I1(n17490[10]), .I2(n901), 
            .I3(n45007), .O(n17041[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5346_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5214_19_lut (.I0(GND_net), .I1(n15306[16]), .I2(GND_net), 
            .I3(n45090), .O(n14585[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5214_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_i749_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n1114));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i749_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5466_4 (.CI(n44850), .I0(n18945[1]), .I1(n259), .CO(n44851));
    SB_LUT4 i40010_3_lut (.I0(n55851), .I1(n436[20]), .I2(n41_adj_4969), 
            .I3(GND_net), .O(n40_adj_5009));   // verilog/motorControl.v(54[23:39])
    defparam i40010_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i39911_4_lut (.I0(n40_adj_5009), .I1(n55740), .I2(n45_adj_4970), 
            .I3(n54648), .O(n55742));   // verilog/motorControl.v(54[23:39])
    defparam i39911_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i39912_3_lut (.I0(n55742), .I1(n356[23]), .I2(n436[23]), .I3(GND_net), 
            .O(n55743));   // verilog/motorControl.v(54[23:39])
    defparam i39912_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i4991_3_lut (.I0(control_update), .I1(n409), .I2(n55743), 
            .I3(GND_net), .O(n10860));   // verilog/motorControl.v(20[7:21])
    defparam i4991_3_lut.LUT_INIT = 16'ha8a8;
    SB_LUT4 mult_17_i85_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [17]), 
            .I2(GND_net), .I3(GND_net), .O(n125_adj_5010));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i85_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i38_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [18]), 
            .I2(GND_net), .I3(GND_net), .O(n56));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i38_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i412_2_lut (.I0(\Kp[8] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n612_adj_5011));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i412_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_19_i41_2_lut (.I0(deadband[20]), .I1(n356[20]), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_5012));   // verilog/motorControl.v(51[12:29])
    defparam LessThan_19_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_19_i39_2_lut (.I0(deadband[19]), .I1(n356[19]), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_5013));   // verilog/motorControl.v(51[12:29])
    defparam LessThan_19_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_19_i45_2_lut (.I0(deadband[22]), .I1(n356[22]), .I2(GND_net), 
            .I3(GND_net), .O(n45_adj_5014));   // verilog/motorControl.v(51[12:29])
    defparam LessThan_19_i45_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_19_i43_2_lut (.I0(deadband[21]), .I1(n356[21]), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_5015));   // verilog/motorControl.v(51[12:29])
    defparam LessThan_19_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_19_i37_2_lut (.I0(deadband[18]), .I1(n356[18]), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_5016));   // verilog/motorControl.v(51[12:29])
    defparam LessThan_19_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_19_i21_2_lut (.I0(deadband[10]), .I1(n356[10]), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_5017));   // verilog/motorControl.v(51[12:29])
    defparam LessThan_19_i21_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_5346_13 (.CI(n45007), .I0(n17490[10]), .I1(n901), .CO(n45008));
    SB_LUT4 add_5346_12_lut (.I0(GND_net), .I1(n17490[9]), .I2(n828), 
            .I3(n45006), .O(n17041[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5346_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_19_i23_2_lut (.I0(deadband[11]), .I1(n356[11]), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_5018));   // verilog/motorControl.v(51[12:29])
    defparam LessThan_19_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_19_i25_2_lut (.I0(deadband[12]), .I1(n356[12]), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_5019));   // verilog/motorControl.v(51[12:29])
    defparam LessThan_19_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_19_i29_2_lut (.I0(deadband[14]), .I1(n356[14]), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_5020));   // verilog/motorControl.v(51[12:29])
    defparam LessThan_19_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_5466_3_lut (.I0(GND_net), .I1(n18945[0]), .I2(n186), .I3(n44849), 
            .O(n18746[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5466_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_19_i31_2_lut (.I0(deadband[15]), .I1(n356[15]), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_5021));   // verilog/motorControl.v(51[12:29])
    defparam LessThan_19_i31_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_5466_3 (.CI(n44849), .I0(n18945[0]), .I1(n186), .CO(n44850));
    SB_LUT4 LessThan_12_i4_4_lut (.I0(n130[0]), .I1(n182[1]), .I2(n130[1]), 
            .I3(n182[0]), .O(n4_adj_5022));   // verilog/motorControl.v(47[21:44])
    defparam LessThan_12_i4_4_lut.LUT_INIT = 16'h4d0c;
    SB_LUT4 i39747_3_lut (.I0(n4_adj_5022), .I1(n182[13]), .I2(n27_adj_4961), 
            .I3(GND_net), .O(n55578));   // verilog/motorControl.v(47[21:44])
    defparam i39747_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i39748_3_lut (.I0(n55578), .I1(n182[14]), .I2(n29_adj_4956), 
            .I3(GND_net), .O(n55579));   // verilog/motorControl.v(47[21:44])
    defparam i39748_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_5466_2_lut (.I0(GND_net), .I1(n44), .I2(n113), .I3(GND_net), 
            .O(n18746[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5466_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i39048_4_lut (.I0(n33_adj_4960), .I1(n31_adj_4959), .I2(n29_adj_4956), 
            .I3(n54883), .O(n54878));
    defparam i39048_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 mult_16_i149_2_lut (.I0(\Kp[3] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n220));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i149_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i39949_4_lut (.I0(n30_adj_4983), .I1(n10_adj_4979), .I2(n35_adj_4954), 
            .I3(n54876), .O(n55780));   // verilog/motorControl.v(47[21:44])
    defparam i39949_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i39364_3_lut (.I0(n55579), .I1(n182[15]), .I2(n31_adj_4959), 
            .I3(GND_net), .O(n55195));   // verilog/motorControl.v(47[21:44])
    defparam i39364_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i40035_4_lut (.I0(n55195), .I1(n55780), .I2(n35_adj_4954), 
            .I3(n54878), .O(n55866));   // verilog/motorControl.v(47[21:44])
    defparam i40035_4_lut.LUT_INIT = 16'hccca;
    SB_CARRY add_5466_2 (.CI(GND_net), .I0(n44), .I1(n113), .CO(n44849));
    SB_LUT4 add_5195_20_lut (.I0(GND_net), .I1(n14946[17]), .I2(GND_net), 
            .I3(n44848), .O(n14186[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5195_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5346_12 (.CI(n45006), .I0(n17490[9]), .I1(n828), .CO(n45007));
    SB_LUT4 LessThan_19_i17_2_lut (.I0(deadband[8]), .I1(n356[8]), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_5023));   // verilog/motorControl.v(51[12:29])
    defparam LessThan_19_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_18_21_lut (.I0(GND_net), .I1(n257[19]), .I2(n306[19]), 
            .I3(n43767), .O(n356[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i40036_3_lut (.I0(n55866), .I1(n182[18]), .I2(n37_adj_4950), 
            .I3(GND_net), .O(n55867));   // verilog/motorControl.v(47[21:44])
    defparam i40036_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_19_i19_2_lut (.I0(deadband[9]), .I1(n356[9]), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_5024));   // verilog/motorControl.v(51[12:29])
    defparam LessThan_19_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i39994_3_lut (.I0(n55867), .I1(n182[19]), .I2(n39_adj_4953), 
            .I3(GND_net), .O(n55825));   // verilog/motorControl.v(47[21:44])
    defparam i39994_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_19_i9_2_lut (.I0(deadband[4]), .I1(n356[4]), .I2(GND_net), 
            .I3(GND_net), .O(n9_adj_5025));   // verilog/motorControl.v(51[12:29])
    defparam LessThan_19_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_5195_19_lut (.I0(GND_net), .I1(n14946[16]), .I2(GND_net), 
            .I3(n44847), .O(n14186[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5195_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_19_i35_2_lut (.I0(deadband[17]), .I1(n363), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_5026));   // verilog/motorControl.v(51[12:29])
    defparam LessThan_19_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_5093_14_lut (.I0(GND_net), .I1(n12905[11]), .I2(n953_adj_5027), 
            .I3(n45142), .O(n11935[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5093_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_19_i33_2_lut (.I0(deadband[16]), .I1(n356[16]), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_5028));   // verilog/motorControl.v(51[12:29])
    defparam LessThan_19_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_19_i11_2_lut (.I0(deadband[5]), .I1(n356[5]), .I2(GND_net), 
            .I3(GND_net), .O(n11_adj_5029));   // verilog/motorControl.v(51[12:29])
    defparam LessThan_19_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_19_i13_2_lut (.I0(deadband[6]), .I1(n356[6]), .I2(GND_net), 
            .I3(GND_net), .O(n13_adj_5030));   // verilog/motorControl.v(51[12:29])
    defparam LessThan_19_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_19_i15_2_lut (.I0(deadband[7]), .I1(n356[7]), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_5031));   // verilog/motorControl.v(51[12:29])
    defparam LessThan_19_i15_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_18_21 (.CI(n43767), .I0(n257[19]), .I1(n306[19]), .CO(n43768));
    SB_LUT4 LessThan_19_i27_2_lut (.I0(deadband[13]), .I1(n356[13]), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_5032));   // verilog/motorControl.v(51[12:29])
    defparam LessThan_19_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_16_i304_2_lut (.I0(\Kp[6] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n451_adj_5033));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i304_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i38931_4_lut (.I0(n356[6]), .I1(n356[5]), .I2(n382[6]), .I3(n382[5]), 
            .O(n54761));
    defparam i38931_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 i39313_3_lut (.I0(n356[7]), .I1(n54761), .I2(n382[7]), .I3(GND_net), 
            .O(n55144));
    defparam i39313_3_lut.LUT_INIT = 16'hdede;
    SB_CARRY add_5195_19 (.CI(n44847), .I0(n14946[16]), .I1(GND_net), 
            .CO(n44848));
    SB_LUT4 i39040_4_lut (.I0(n43_adj_4945), .I1(n41_adj_4942), .I2(n39_adj_4953), 
            .I3(n55800), .O(n54870));
    defparam i39040_4_lut.LUT_INIT = 16'haaab;
    SB_CARRY add_5214_19 (.CI(n45090), .I0(n15306[16]), .I1(GND_net), 
            .CO(n45091));
    SB_LUT4 LessThan_21_i27_rep_175_2_lut (.I0(n356[13]), .I1(n382[13]), 
            .I2(GND_net), .I3(GND_net), .O(n57142));   // verilog/motorControl.v(51[33:53])
    defparam LessThan_21_i27_rep_175_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i39292_4_lut (.I0(n356[14]), .I1(n57142), .I2(n382[14]), .I3(n55144), 
            .O(n55123));
    defparam i39292_4_lut.LUT_INIT = 16'hdeff;
    SB_LUT4 add_18_20_lut (.I0(GND_net), .I1(n257[18]), .I2(n306[18]), 
            .I3(n43766), .O(n356[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5195_18_lut (.I0(GND_net), .I1(n14946[15]), .I2(GND_net), 
            .I3(n44846), .O(n14186[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5195_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_21_i31_rep_169_2_lut (.I0(n356[15]), .I1(n382[15]), 
            .I2(GND_net), .I3(GND_net), .O(n57136));   // verilog/motorControl.v(51[33:53])
    defparam LessThan_21_i31_rep_169_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_5093_14 (.CI(n45142), .I0(n12905[11]), .I1(n953_adj_5027), 
            .CO(n45143));
    SB_LUT4 add_5346_11_lut (.I0(GND_net), .I1(n17490[8]), .I2(n755), 
            .I3(n45005), .O(n17041[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5346_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5195_18 (.CI(n44846), .I0(n14946[15]), .I1(GND_net), 
            .CO(n44847));
    SB_LUT4 add_5214_18_lut (.I0(GND_net), .I1(n15306[15]), .I2(GND_net), 
            .I3(n45089), .O(n14585[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5214_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i39887_4_lut (.I0(n55193), .I1(n55464), .I2(n45_adj_4947), 
            .I3(n54868), .O(n55718));   // verilog/motorControl.v(47[21:44])
    defparam i39887_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i38927_4_lut (.I0(n356[8]), .I1(n356[4]), .I2(n382[8]), .I3(n382[4]), 
            .O(n54757));
    defparam i38927_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 i39307_3_lut (.I0(n356[9]), .I1(n54757), .I2(n382[9]), .I3(GND_net), 
            .O(n55138));
    defparam i39307_3_lut.LUT_INIT = 16'hdede;
    SB_LUT4 LessThan_21_i21_rep_190_2_lut (.I0(n356[10]), .I1(n382[10]), 
            .I2(GND_net), .I3(GND_net), .O(n57157));   // verilog/motorControl.v(51[33:53])
    defparam LessThan_21_i21_rep_190_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i39303_4_lut (.I0(n356[11]), .I1(n57157), .I2(n382[11]), .I3(n55138), 
            .O(n55134));
    defparam i39303_4_lut.LUT_INIT = 16'hdeff;
    SB_LUT4 i39370_3_lut (.I0(n55825), .I1(n182[20]), .I2(n41_adj_4942), 
            .I3(GND_net), .O(n55201));   // verilog/motorControl.v(47[21:44])
    defparam i39370_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i39965_4_lut (.I0(n55201), .I1(n55718), .I2(n45_adj_4947), 
            .I3(n54870), .O(n55796));   // verilog/motorControl.v(47[21:44])
    defparam i39965_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i39966_3_lut (.I0(n55796), .I1(n130[23]), .I2(n182[23]), .I3(GND_net), 
            .O(n181));   // verilog/motorControl.v(47[21:44])
    defparam i39966_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 LessThan_21_i25_rep_184_2_lut (.I0(n356[12]), .I1(n382[12]), 
            .I2(GND_net), .I3(GND_net), .O(n57151));   // verilog/motorControl.v(51[33:53])
    defparam LessThan_21_i25_rep_184_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_21_i16_3_lut (.I0(n382[9]), .I1(n382[21]), .I2(n356[21]), 
            .I3(GND_net), .O(n16_adj_5035));   // verilog/motorControl.v(51[33:53])
    defparam LessThan_21_i16_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i38895_4_lut (.I0(n356[21]), .I1(n356[9]), .I2(n382[21]), 
            .I3(n382[9]), .O(n54725));
    defparam i38895_4_lut.LUT_INIT = 16'h7bde;
    SB_CARRY add_18_20 (.CI(n43766), .I0(n257[18]), .I1(n306[18]), .CO(n43767));
    SB_LUT4 mux_14_i2_3_lut (.I0(n130[1]), .I1(n182[1]), .I2(n181), .I3(GND_net), 
            .O(n207[1]));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_14_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_15_i2_3_lut (.I0(n207[1]), .I1(IntegralLimit[1]), .I2(n155), 
            .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3996 [1]));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_15_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_5195_17_lut (.I0(GND_net), .I1(n14946[14]), .I2(GND_net), 
            .I3(n44845), .O(n14186[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5195_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i406_2_lut (.I0(\Kp[8] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n603_adj_5036));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i406_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i445_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n661));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i445_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_18_19_lut (.I0(GND_net), .I1(n257[17]), .I2(n306[17]), 
            .I3(n43765), .O(n363)) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_18_19 (.CI(n43765), .I0(n257[17]), .I1(n306[17]), .CO(n43766));
    SB_LUT4 LessThan_21_i8_3_lut (.I0(n382[4]), .I1(n382[8]), .I2(n356[8]), 
            .I3(GND_net), .O(n8_adj_5037));   // verilog/motorControl.v(51[33:53])
    defparam LessThan_21_i8_3_lut.LUT_INIT = 16'h8e8e;
    SB_CARRY add_5195_17 (.CI(n44845), .I0(n14946[14]), .I1(GND_net), 
            .CO(n44846));
    SB_CARRY add_5214_18 (.CI(n45089), .I0(n15306[15]), .I1(GND_net), 
            .CO(n45090));
    SB_LUT4 LessThan_21_i24_3_lut (.I0(n16_adj_5035), .I1(n382[22]), .I2(n356[22]), 
            .I3(GND_net), .O(n24_adj_5039));   // verilog/motorControl.v(51[33:53])
    defparam LessThan_21_i24_3_lut.LUT_INIT = 16'h8e8e;
    SB_CARRY add_5346_11 (.CI(n45005), .I0(n17490[8]), .I1(n755), .CO(n45006));
    SB_LUT4 add_5346_10_lut (.I0(GND_net), .I1(n17490[7]), .I2(n682), 
            .I3(n45004), .O(n17041[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5346_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i38935_4_lut (.I0(n356[3]), .I1(n356[2]), .I2(n382[3]), .I3(n382[2]), 
            .O(n54765));
    defparam i38935_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 add_5195_16_lut (.I0(GND_net), .I1(n14946[13]), .I2(n1108), 
            .I3(n44844), .O(n14186[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5195_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_21_i9_rep_183_2_lut (.I0(n356[4]), .I1(n382[4]), .I2(GND_net), 
            .I3(GND_net), .O(n57150));   // verilog/motorControl.v(51[33:53])
    defparam LessThan_21_i9_rep_183_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i38933_4_lut (.I0(n356[5]), .I1(n57150), .I2(n382[5]), .I3(n54765), 
            .O(n54763));
    defparam i38933_4_lut.LUT_INIT = 16'h5a7b;
    SB_LUT4 LessThan_21_i13_rep_211_2_lut (.I0(n356[6]), .I1(n382[6]), .I2(GND_net), 
            .I3(GND_net), .O(n57178));   // verilog/motorControl.v(51[33:53])
    defparam LessThan_21_i13_rep_211_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i39619_4_lut (.I0(n356[7]), .I1(n57178), .I2(n382[7]), .I3(n54763), 
            .O(n55450));
    defparam i39619_4_lut.LUT_INIT = 16'hffde;
    SB_CARRY add_5195_16 (.CI(n44844), .I0(n14946[13]), .I1(n1108), .CO(n44845));
    SB_LUT4 add_5195_15_lut (.I0(GND_net), .I1(n14946[12]), .I2(n1035), 
            .I3(n44843), .O(n14186[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5195_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5346_10 (.CI(n45004), .I0(n17490[7]), .I1(n682), .CO(n45005));
    SB_CARRY add_5195_15 (.CI(n44843), .I0(n14946[12]), .I1(n1035), .CO(n44844));
    SB_LUT4 add_18_18_lut (.I0(GND_net), .I1(n257[16]), .I2(n306[16]), 
            .I3(n43764), .O(n356[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_18_18 (.CI(n43764), .I0(n257[16]), .I1(n306[16]), .CO(n43765));
    SB_LUT4 add_5093_13_lut (.I0(GND_net), .I1(n12905[10]), .I2(n880_adj_5041), 
            .I3(n45141), .O(n11935[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5093_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5195_14_lut (.I0(GND_net), .I1(n14946[11]), .I2(n962), 
            .I3(n44842), .O(n14186[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5195_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 counter_2283_add_4_33_lut (.I0(GND_net), .I1(GND_net), .I2(counter[31]), 
            .I3(n44563), .O(n28[31])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2283_add_4_33_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 counter_2283_add_4_32_lut (.I0(GND_net), .I1(GND_net), .I2(counter[30]), 
            .I3(n44562), .O(n28[30])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2283_add_4_32_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_2283_add_4_32 (.CI(n44562), .I0(GND_net), .I1(counter[30]), 
            .CO(n44563));
    SB_LUT4 counter_2283_add_4_31_lut (.I0(GND_net), .I1(GND_net), .I2(counter[29]), 
            .I3(n44561), .O(n28[29])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2283_add_4_31_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_2283_add_4_31 (.CI(n44561), .I0(GND_net), .I1(counter[29]), 
            .CO(n44562));
    SB_LUT4 counter_2283_add_4_30_lut (.I0(GND_net), .I1(GND_net), .I2(counter[28]), 
            .I3(n44560), .O(n28[28])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2283_add_4_30_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5346_9_lut (.I0(GND_net), .I1(n17490[6]), .I2(n609), .I3(n45003), 
            .O(n17041[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5346_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_2283_add_4_30 (.CI(n44560), .I0(GND_net), .I1(counter[28]), 
            .CO(n44561));
    SB_CARRY add_5195_14 (.CI(n44842), .I0(n14946[11]), .I1(n962), .CO(n44843));
    SB_LUT4 counter_2283_add_4_29_lut (.I0(GND_net), .I1(GND_net), .I2(counter[27]), 
            .I3(n44559), .O(n28[27])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2283_add_4_29_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_21_i17_rep_208_2_lut (.I0(n356[8]), .I1(n382[8]), .I2(GND_net), 
            .I3(GND_net), .O(n57175));   // verilog/motorControl.v(51[33:53])
    defparam LessThan_21_i17_rep_208_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i39311_4_lut (.I0(n356[9]), .I1(n57175), .I2(n382[9]), .I3(n55450), 
            .O(n55142));
    defparam i39311_4_lut.LUT_INIT = 16'hdeff;
    SB_LUT4 add_5214_17_lut (.I0(GND_net), .I1(n15306[14]), .I2(GND_net), 
            .I3(n45088), .O(n14585[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5214_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i39739_4_lut (.I0(n356[11]), .I1(n57157), .I2(n382[11]), .I3(n55142), 
            .O(n55570));
    defparam i39739_4_lut.LUT_INIT = 16'hffde;
    SB_CARRY counter_2283_add_4_29 (.CI(n44559), .I0(GND_net), .I1(counter[27]), 
            .CO(n44560));
    SB_LUT4 counter_2283_add_4_28_lut (.I0(GND_net), .I1(GND_net), .I2(counter[26]), 
            .I3(n44558), .O(n28[26])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2283_add_4_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5214_17 (.CI(n45088), .I0(n15306[14]), .I1(GND_net), 
            .CO(n45089));
    SB_CARRY add_5346_9 (.CI(n45003), .I0(n17490[6]), .I1(n609), .CO(n45004));
    SB_LUT4 add_5195_13_lut (.I0(GND_net), .I1(n14946[10]), .I2(n889), 
            .I3(n44841), .O(n14186[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5195_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i38918_4_lut (.I0(n356[13]), .I1(n57151), .I2(n382[13]), .I3(n55570), 
            .O(n54748));
    defparam i38918_4_lut.LUT_INIT = 16'h5a7b;
    SB_LUT4 LessThan_21_i29_rep_173_2_lut (.I0(n356[14]), .I1(n382[14]), 
            .I2(GND_net), .I3(GND_net), .O(n57140));   // verilog/motorControl.v(51[33:53])
    defparam LessThan_21_i29_rep_173_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_5195_13 (.CI(n44841), .I0(n14946[10]), .I1(n889), .CO(n44842));
    SB_LUT4 i39609_4_lut (.I0(n356[15]), .I1(n57140), .I2(n382[15]), .I3(n54748), 
            .O(n55440));
    defparam i39609_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 add_18_17_lut (.I0(GND_net), .I1(n257[15]), .I2(n306[15]), 
            .I3(n43763), .O(n356[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_2283_add_4_28 (.CI(n44558), .I0(GND_net), .I1(counter[26]), 
            .CO(n44559));
    SB_LUT4 mult_16_i198_2_lut (.I0(\Kp[4] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n293));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i198_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 counter_2283_add_4_27_lut (.I0(GND_net), .I1(GND_net), .I2(counter[25]), 
            .I3(n44557), .O(n28[25])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2283_add_4_27_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5346_8_lut (.I0(GND_net), .I1(n17490[5]), .I2(n536_adj_5049), 
            .I3(n45002), .O(n17041[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5346_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5346_8 (.CI(n45002), .I0(n17490[5]), .I1(n536_adj_5049), 
            .CO(n45003));
    SB_CARRY add_18_17 (.CI(n43763), .I0(n257[15]), .I1(n306[15]), .CO(n43764));
    SB_LUT4 add_5214_16_lut (.I0(GND_net), .I1(n15306[13]), .I2(n1108_adj_5050), 
            .I3(n45087), .O(n14585[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5214_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_18_16_lut (.I0(GND_net), .I1(n257[14]), .I2(n306[14]), 
            .I3(n43762), .O(n356[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_2283_add_4_27 (.CI(n44557), .I0(GND_net), .I1(counter[25]), 
            .CO(n44558));
    SB_LUT4 add_5346_7_lut (.I0(GND_net), .I1(n17490[4]), .I2(n463_adj_5051), 
            .I3(n45001), .O(n17041[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5346_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5195_12_lut (.I0(GND_net), .I1(n14946[9]), .I2(n816), 
            .I3(n44840), .O(n14186[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5195_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5195_12 (.CI(n44840), .I0(n14946[9]), .I1(n816), .CO(n44841));
    SB_CARRY add_5093_13 (.CI(n45141), .I0(n12905[10]), .I1(n880_adj_5041), 
            .CO(n45142));
    SB_CARRY add_5214_16 (.CI(n45087), .I0(n15306[13]), .I1(n1108_adj_5050), 
            .CO(n45088));
    SB_LUT4 counter_2283_add_4_26_lut (.I0(GND_net), .I1(GND_net), .I2(counter[24]), 
            .I3(n44556), .O(n28[24])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2283_add_4_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5346_7 (.CI(n45001), .I0(n17490[4]), .I1(n463_adj_5051), 
            .CO(n45002));
    SB_CARRY counter_2283_add_4_26 (.CI(n44556), .I0(GND_net), .I1(counter[24]), 
            .CO(n44557));
    SB_LUT4 add_5195_11_lut (.I0(GND_net), .I1(n14946[8]), .I2(n743), 
            .I3(n44839), .O(n14186[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5195_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5195_11 (.CI(n44839), .I0(n14946[8]), .I1(n743), .CO(n44840));
    SB_LUT4 counter_2283_add_4_25_lut (.I0(GND_net), .I1(GND_net), .I2(counter[23]), 
            .I3(n44555), .O(n28[23])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2283_add_4_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_2283_add_4_25 (.CI(n44555), .I0(GND_net), .I1(counter[23]), 
            .CO(n44556));
    SB_LUT4 counter_2283_add_4_24_lut (.I0(GND_net), .I1(GND_net), .I2(counter[22]), 
            .I3(n44554), .O(n28[22])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2283_add_4_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_21_i33_rep_201_2_lut (.I0(n356[16]), .I1(n382[16]), 
            .I2(GND_net), .I3(GND_net), .O(n57168));   // verilog/motorControl.v(51[33:53])
    defparam LessThan_21_i33_rep_201_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i39861_4_lut (.I0(n363), .I1(n57168), .I2(n382[17]), .I3(n55440), 
            .O(n55692));
    defparam i39861_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 LessThan_21_i37_rep_164_2_lut (.I0(n356[18]), .I1(n382[18]), 
            .I2(GND_net), .I3(GND_net), .O(n57131));   // verilog/motorControl.v(51[33:53])
    defparam LessThan_21_i37_rep_164_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i39989_4_lut (.I0(n356[19]), .I1(n57131), .I2(n382[19]), .I3(n55692), 
            .O(n55820));
    defparam i39989_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 add_5195_10_lut (.I0(GND_net), .I1(n14946[7]), .I2(n670), 
            .I3(n44838), .O(n14186[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5195_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_2283_add_4_24 (.CI(n44554), .I0(GND_net), .I1(counter[22]), 
            .CO(n44555));
    SB_LUT4 counter_2283_add_4_23_lut (.I0(GND_net), .I1(GND_net), .I2(counter[21]), 
            .I3(n44553), .O(n28[21])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2283_add_4_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5346_6_lut (.I0(GND_net), .I1(n17490[3]), .I2(n390_adj_5058), 
            .I3(n45000), .O(n17041[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5346_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5214_15_lut (.I0(GND_net), .I1(n15306[12]), .I2(n1035_adj_5059), 
            .I3(n45086), .O(n14585[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5214_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_18_16 (.CI(n43762), .I0(n257[14]), .I1(n306[14]), .CO(n43763));
    SB_CARRY add_5195_10 (.CI(n44838), .I0(n14946[7]), .I1(n670), .CO(n44839));
    SB_CARRY counter_2283_add_4_23 (.CI(n44553), .I0(GND_net), .I1(counter[21]), 
            .CO(n44554));
    SB_CARRY add_5346_6 (.CI(n45000), .I0(n17490[3]), .I1(n390_adj_5058), 
            .CO(n45001));
    SB_LUT4 counter_2283_add_4_22_lut (.I0(GND_net), .I1(GND_net), .I2(counter[20]), 
            .I3(n44552), .O(n28[20])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2283_add_4_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5195_9_lut (.I0(GND_net), .I1(n14946[6]), .I2(n597), .I3(n44837), 
            .O(n14186[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5195_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_2283_add_4_22 (.CI(n44552), .I0(GND_net), .I1(counter[20]), 
            .CO(n44553));
    SB_CARRY add_5195_9 (.CI(n44837), .I0(n14946[6]), .I1(n597), .CO(n44838));
    SB_LUT4 counter_2283_add_4_21_lut (.I0(GND_net), .I1(GND_net), .I2(counter[19]), 
            .I3(n44551), .O(n28[19])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2283_add_4_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_2283_add_4_21 (.CI(n44551), .I0(GND_net), .I1(counter[19]), 
            .CO(n44552));
    SB_LUT4 add_5195_8_lut (.I0(GND_net), .I1(n14946[5]), .I2(n524), .I3(n44836), 
            .O(n14186[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5195_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_21_i41_rep_161_2_lut (.I0(n356[20]), .I1(n382[20]), 
            .I2(GND_net), .I3(GND_net), .O(n57128));   // verilog/motorControl.v(51[33:53])
    defparam LessThan_21_i41_rep_161_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i39005_4_lut (.I0(n27_adj_5032), .I1(n15_adj_5031), .I2(n13_adj_5030), 
            .I3(n11_adj_5029), .O(n54835));
    defparam i39005_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 counter_2283_add_4_20_lut (.I0(GND_net), .I1(GND_net), .I2(counter[18]), 
            .I3(n44550), .O(n28[18])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2283_add_4_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_2283_add_4_20 (.CI(n44550), .I0(GND_net), .I1(counter[18]), 
            .CO(n44551));
    SB_LUT4 counter_2283_add_4_19_lut (.I0(GND_net), .I1(GND_net), .I2(counter[17]), 
            .I3(n44549), .O(n28[17])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2283_add_4_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_19_i12_3_lut (.I0(n356[7]), .I1(n356[16]), .I2(n33_adj_5028), 
            .I3(GND_net), .O(n12_adj_5064));   // verilog/motorControl.v(51[12:29])
    defparam LessThan_19_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY counter_2283_add_4_19 (.CI(n44549), .I0(GND_net), .I1(counter[17]), 
            .CO(n44550));
    SB_LUT4 add_5346_5_lut (.I0(GND_net), .I1(n17490[2]), .I2(n317_adj_5065), 
            .I3(n44999), .O(n17041[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5346_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5195_8 (.CI(n44836), .I0(n14946[5]), .I1(n524), .CO(n44837));
    SB_LUT4 LessThan_19_i10_3_lut (.I0(n356[5]), .I1(n356[6]), .I2(n13_adj_5030), 
            .I3(GND_net), .O(n10_adj_5066));   // verilog/motorControl.v(51[12:29])
    defparam LessThan_19_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 counter_2283_add_4_18_lut (.I0(GND_net), .I1(GND_net), .I2(counter[16]), 
            .I3(n44548), .O(n28[16])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2283_add_4_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_2283_add_4_18 (.CI(n44548), .I0(GND_net), .I1(counter[16]), 
            .CO(n44549));
    SB_CARRY add_5346_5 (.CI(n44999), .I0(n17490[2]), .I1(n317_adj_5065), 
            .CO(n45000));
    SB_LUT4 add_5195_7_lut (.I0(GND_net), .I1(n14946[4]), .I2(n451_adj_5068), 
            .I3(n44835), .O(n14186[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5195_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 counter_2283_add_4_17_lut (.I0(GND_net), .I1(GND_net), .I2(counter[15]), 
            .I3(n44547), .O(n28[15])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2283_add_4_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5195_7 (.CI(n44835), .I0(n14946[4]), .I1(n451_adj_5068), 
            .CO(n44836));
    SB_LUT4 LessThan_19_i30_3_lut (.I0(n12_adj_5064), .I1(n363), .I2(n35_adj_5026), 
            .I3(GND_net), .O(n30_adj_5070));   // verilog/motorControl.v(51[12:29])
    defparam LessThan_19_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY counter_2283_add_4_17 (.CI(n44547), .I0(GND_net), .I1(counter[15]), 
            .CO(n44548));
    SB_LUT4 counter_2283_add_4_16_lut (.I0(GND_net), .I1(GND_net), .I2(counter[14]), 
            .I3(n44546), .O(n28[14])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2283_add_4_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5195_6_lut (.I0(GND_net), .I1(n14946[3]), .I2(n378_adj_5072), 
            .I3(n44834), .O(n14186[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5195_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_2283_add_4_16 (.CI(n44546), .I0(GND_net), .I1(counter[14]), 
            .CO(n44547));
    SB_LUT4 i39398_4_lut (.I0(n13_adj_5030), .I1(n11_adj_5029), .I2(n9_adj_5025), 
            .I3(n54864), .O(n55229));
    defparam i39398_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 counter_2283_add_4_15_lut (.I0(GND_net), .I1(GND_net), .I2(counter[13]), 
            .I3(n44545), .O(n28[13])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2283_add_4_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5195_6 (.CI(n44834), .I0(n14946[3]), .I1(n378_adj_5072), 
            .CO(n44835));
    SB_CARRY counter_2283_add_4_15 (.CI(n44545), .I0(GND_net), .I1(counter[13]), 
            .CO(n44546));
    SB_LUT4 counter_2283_add_4_14_lut (.I0(GND_net), .I1(GND_net), .I2(counter[12]), 
            .I3(n44544), .O(n28[12])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2283_add_4_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5214_15 (.CI(n45086), .I0(n15306[12]), .I1(n1035_adj_5059), 
            .CO(n45087));
    SB_LUT4 add_5195_5_lut (.I0(GND_net), .I1(n14946[2]), .I2(n305_adj_5074), 
            .I3(n44833), .O(n14186[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5195_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5093_12_lut (.I0(GND_net), .I1(n12905[9]), .I2(n807), 
            .I3(n45140), .O(n11935[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5093_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_2283_add_4_14 (.CI(n44544), .I0(GND_net), .I1(counter[12]), 
            .CO(n44545));
    SB_CARRY add_5195_5 (.CI(n44833), .I0(n14946[2]), .I1(n305_adj_5074), 
            .CO(n44834));
    SB_LUT4 counter_2283_add_4_13_lut (.I0(GND_net), .I1(GND_net), .I2(counter[11]), 
            .I3(n44543), .O(n28[11])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2283_add_4_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i39394_4_lut (.I0(n19_adj_5024), .I1(n17_adj_5023), .I2(n15_adj_5031), 
            .I3(n55229), .O(n55225));
    defparam i39394_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 add_18_15_lut (.I0(GND_net), .I1(n257[13]), .I2(n306[13]), 
            .I3(n43761), .O(n356[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i39915_4_lut (.I0(n25_adj_5019), .I1(n23_adj_5018), .I2(n21_adj_5017), 
            .I3(n55225), .O(n55746));
    defparam i39915_4_lut.LUT_INIT = 16'hfffe;
    SB_CARRY counter_2283_add_4_13 (.CI(n44543), .I0(GND_net), .I1(counter[11]), 
            .CO(n44544));
    SB_LUT4 add_5214_14_lut (.I0(GND_net), .I1(n15306[11]), .I2(n962_adj_5076), 
            .I3(n45085), .O(n14585[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5214_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 counter_2283_add_4_12_lut (.I0(GND_net), .I1(GND_net), .I2(counter[10]), 
            .I3(n44542), .O(n28[10])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2283_add_4_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5346_4_lut (.I0(GND_net), .I1(n17490[1]), .I2(n244_adj_5078), 
            .I3(n44998), .O(n17041[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5346_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5346_4 (.CI(n44998), .I0(n17490[1]), .I1(n244_adj_5078), 
            .CO(n44999));
    SB_CARRY add_18_15 (.CI(n43761), .I0(n257[13]), .I1(n306[13]), .CO(n43762));
    SB_LUT4 add_5346_3_lut (.I0(GND_net), .I1(n17490[0]), .I2(n171_adj_5079), 
            .I3(n44997), .O(n17041[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5346_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_2283_add_4_12 (.CI(n44542), .I0(GND_net), .I1(counter[10]), 
            .CO(n44543));
    SB_CARRY add_5346_3 (.CI(n44997), .I0(n17490[0]), .I1(n171_adj_5079), 
            .CO(n44998));
    SB_LUT4 counter_2283_add_4_11_lut (.I0(GND_net), .I1(GND_net), .I2(counter[9]), 
            .I3(n44541), .O(n28[9])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2283_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5195_4_lut (.I0(GND_net), .I1(n14946[1]), .I2(n232_adj_5081), 
            .I3(n44832), .O(n14186[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5195_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_2283_add_4_11 (.CI(n44541), .I0(GND_net), .I1(counter[9]), 
            .CO(n44542));
    SB_LUT4 counter_2283_add_4_10_lut (.I0(GND_net), .I1(GND_net), .I2(counter[8]), 
            .I3(n44540), .O(n28[8])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2283_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i39647_4_lut (.I0(n31_adj_5021), .I1(n29_adj_5020), .I2(n27_adj_5032), 
            .I3(n55746), .O(n55478));
    defparam i39647_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i39967_4_lut (.I0(n37_adj_5016), .I1(n35_adj_5026), .I2(n33_adj_5028), 
            .I3(n55478), .O(n55798));
    defparam i39967_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i39735_3_lut (.I0(n6_adj_5082), .I1(n356[10]), .I2(n21_adj_5017), 
            .I3(GND_net), .O(n55566));   // verilog/motorControl.v(51[12:29])
    defparam i39735_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_19_i16_3_lut (.I0(n356[9]), .I1(n356[21]), .I2(n43_adj_5015), 
            .I3(GND_net), .O(n16_adj_5083));   // verilog/motorControl.v(51[12:29])
    defparam LessThan_19_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY counter_2283_add_4_10 (.CI(n44540), .I0(GND_net), .I1(counter[8]), 
            .CO(n44541));
    SB_CARRY add_5195_4 (.CI(n44832), .I0(n14946[1]), .I1(n232_adj_5081), 
            .CO(n44833));
    SB_LUT4 add_18_14_lut (.I0(GND_net), .I1(n257[12]), .I2(n306[12]), 
            .I3(n43760), .O(n356[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5195_3_lut (.I0(GND_net), .I1(n14946[0]), .I2(n159_adj_5085), 
            .I3(n44831), .O(n14186[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5195_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5346_2_lut (.I0(GND_net), .I1(n29_adj_5086), .I2(n98_adj_5087), 
            .I3(GND_net), .O(n17041[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5346_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 counter_2283_add_4_9_lut (.I0(GND_net), .I1(GND_net), .I2(counter[7]), 
            .I3(n44539), .O(n28[7])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2283_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_18_14 (.CI(n43760), .I0(n257[12]), .I1(n306[12]), .CO(n43761));
    SB_LUT4 LessThan_19_i8_3_lut (.I0(n356[4]), .I1(n356[8]), .I2(n17_adj_5023), 
            .I3(GND_net), .O(n8_adj_5088));   // verilog/motorControl.v(51[12:29])
    defparam LessThan_19_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_19_i24_3_lut (.I0(n16_adj_5083), .I1(n356[22]), .I2(n45_adj_5014), 
            .I3(GND_net), .O(n24_adj_5089));   // verilog/motorControl.v(51[12:29])
    defparam LessThan_19_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i39018_4_lut (.I0(n21_adj_5017), .I1(n19_adj_5024), .I2(n17_adj_5023), 
            .I3(n9_adj_5025), .O(n54848));
    defparam i39018_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 mult_16_i79_2_lut (.I0(\Kp[1] ), .I1(n1[14]), .I2(GND_net), 
            .I3(GND_net), .O(n116));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i79_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i32_2_lut (.I0(\Kp[0] ), .I1(n1[15]), .I2(GND_net), 
            .I3(GND_net), .O(n47));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i32_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i39736_3_lut (.I0(n55566), .I1(n356[11]), .I2(n23_adj_5018), 
            .I3(GND_net), .O(n55567));   // verilog/motorControl.v(51[12:29])
    defparam i39736_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_18_13_lut (.I0(GND_net), .I1(n257[11]), .I2(n306[11]), 
            .I3(n43759), .O(n356[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i38950_4_lut (.I0(n43_adj_5015), .I1(n25_adj_5019), .I2(n23_adj_5018), 
            .I3(n54848), .O(n54780));
    defparam i38950_4_lut.LUT_INIT = 16'haaab;
    SB_CARRY add_5195_3 (.CI(n44831), .I0(n14946[0]), .I1(n159_adj_5085), 
            .CO(n44832));
    SB_LUT4 add_5195_2_lut (.I0(GND_net), .I1(n17_adj_5091), .I2(n86), 
            .I3(GND_net), .O(n14186[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5195_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_2283_add_4_9 (.CI(n44539), .I0(GND_net), .I1(counter[7]), 
            .CO(n44540));
    SB_LUT4 i39635_4_lut (.I0(n24_adj_5089), .I1(n8_adj_5088), .I2(n45_adj_5014), 
            .I3(n54777), .O(n55466));   // verilog/motorControl.v(51[12:29])
    defparam i39635_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i39372_3_lut (.I0(n55567), .I1(n356[12]), .I2(n25_adj_5019), 
            .I3(GND_net), .O(n55203));   // verilog/motorControl.v(51[12:29])
    defparam i39372_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_21_i12_3_lut (.I0(n382[7]), .I1(n382[16]), .I2(n356[16]), 
            .I3(GND_net), .O(n12_adj_5092));   // verilog/motorControl.v(51[33:53])
    defparam LessThan_21_i12_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 LessThan_21_i4_3_lut (.I0(n54560), .I1(n382[1]), .I2(n356[1]), 
            .I3(GND_net), .O(n4_adj_5094));   // verilog/motorControl.v(51[33:53])
    defparam LessThan_21_i4_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i39839_3_lut (.I0(n4_adj_5094), .I1(n382[13]), .I2(n356[13]), 
            .I3(GND_net), .O(n55670));   // verilog/motorControl.v(51[33:53])
    defparam i39839_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i39840_3_lut (.I0(n55670), .I1(n382[14]), .I2(n356[14]), .I3(GND_net), 
            .O(n55671));   // verilog/motorControl.v(51[33:53])
    defparam i39840_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 counter_2283_add_4_8_lut (.I0(GND_net), .I1(GND_net), .I2(counter[6]), 
            .I3(n44538), .O(n28[6])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2283_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_2283_add_4_8 (.CI(n44538), .I0(GND_net), .I1(counter[6]), 
            .CO(n44539));
    SB_LUT4 counter_2283_add_4_7_lut (.I0(GND_net), .I1(GND_net), .I2(counter[5]), 
            .I3(n44537), .O(n28[5])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2283_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i38905_4_lut (.I0(n356[16]), .I1(n356[7]), .I2(n382[16]), 
            .I3(n382[7]), .O(n54735));
    defparam i38905_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 LessThan_21_i35_rep_196_2_lut (.I0(n363), .I1(n382[17]), .I2(GND_net), 
            .I3(GND_net), .O(n57163));   // verilog/motorControl.v(51[33:53])
    defparam LessThan_21_i35_rep_196_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_21_i10_3_lut (.I0(n382[5]), .I1(n382[6]), .I2(n356[6]), 
            .I3(GND_net), .O(n10_adj_5096));   // verilog/motorControl.v(51[33:53])
    defparam LessThan_21_i10_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 LessThan_21_i30_3_lut (.I0(n12_adj_5092), .I1(n382[17]), .I2(n363), 
            .I3(GND_net), .O(n30_adj_5097));   // verilog/motorControl.v(51[33:53])
    defparam LessThan_21_i30_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i38908_4_lut (.I0(n356[16]), .I1(n57136), .I2(n382[16]), .I3(n55123), 
            .O(n54738));
    defparam i38908_4_lut.LUT_INIT = 16'h5a7b;
    SB_LUT4 mult_16_i461_2_lut (.I0(\Kp[9] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n685_adj_5098));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i461_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_14_i15_3_lut (.I0(n130[14]), .I1(n182[14]), .I2(n181), 
            .I3(GND_net), .O(n207[14]));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_14_i15_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_15_i15_3_lut (.I0(n207[14]), .I1(IntegralLimit[14]), .I2(n155), 
            .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3996 [14]));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_15_i15_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_17_i77_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [13]), 
            .I2(GND_net), .I3(GND_net), .O(n113_adj_5099));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i77_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i39979_4_lut (.I0(n30_adj_5097), .I1(n10_adj_5096), .I2(n57163), 
            .I3(n54735), .O(n55810));   // verilog/motorControl.v(51[33:53])
    defparam i39979_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i39774_3_lut (.I0(n55671), .I1(n382[15]), .I2(n356[15]), .I3(GND_net), 
            .O(n55605));   // verilog/motorControl.v(51[33:53])
    defparam i39774_3_lut.LUT_INIT = 16'h8e8e;
    SB_CARRY counter_2283_add_4_7 (.CI(n44537), .I0(GND_net), .I1(counter[5]), 
            .CO(n44538));
    SB_LUT4 i40057_4_lut (.I0(n55605), .I1(n55810), .I2(n57163), .I3(n54738), 
            .O(n55888));   // verilog/motorControl.v(51[33:53])
    defparam i40057_4_lut.LUT_INIT = 16'hccca;
    SB_CARRY add_5195_2 (.CI(GND_net), .I0(n17_adj_5091), .I1(n86), .CO(n44831));
    SB_LUT4 i40058_3_lut (.I0(n55888), .I1(n382[18]), .I2(n356[18]), .I3(GND_net), 
            .O(n55889));   // verilog/motorControl.v(51[33:53])
    defparam i40058_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 counter_2283_add_4_6_lut (.I0(GND_net), .I1(GND_net), .I2(counter[4]), 
            .I3(n44536), .O(n28[4])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2283_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_2283_add_4_6 (.CI(n44536), .I0(GND_net), .I1(counter[4]), 
            .CO(n44537));
    SB_LUT4 LessThan_21_i6_3_lut (.I0(n382[2]), .I1(n382[3]), .I2(n356[3]), 
            .I3(GND_net), .O(n6_adj_5100));   // verilog/motorControl.v(51[33:53])
    defparam LessThan_21_i6_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 mult_17_i30_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [14]), 
            .I2(GND_net), .I3(GND_net), .O(n44_adj_5101));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i30_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5346_2 (.CI(GND_net), .I0(n29_adj_5086), .I1(n98_adj_5087), 
            .CO(n44997));
    SB_LUT4 add_5232_19_lut (.I0(GND_net), .I1(n15630[16]), .I2(GND_net), 
            .I3(n44830), .O(n14946[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5232_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5232_18_lut (.I0(GND_net), .I1(n15630[15]), .I2(GND_net), 
            .I3(n44829), .O(n14946[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5232_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 counter_2283_add_4_5_lut (.I0(GND_net), .I1(GND_net), .I2(counter[3]), 
            .I3(n44535), .O(n28[3])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2283_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_2283_add_4_5 (.CI(n44535), .I0(GND_net), .I1(counter[3]), 
            .CO(n44536));
    SB_LUT4 mult_16_i353_2_lut (.I0(\Kp[7] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n524_adj_5102));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i353_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i126_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [13]), 
            .I2(GND_net), .I3(GND_net), .O(n186_adj_5103));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i126_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i175_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [13]), 
            .I2(GND_net), .I3(GND_net), .O(n259_adj_5104));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i175_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_18_13 (.CI(n43759), .I0(n257[11]), .I1(n306[11]), .CO(n43760));
    SB_LUT4 counter_2283_add_4_4_lut (.I0(GND_net), .I1(GND_net), .I2(counter[2]), 
            .I3(n44534), .O(n28[2])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2283_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5232_18 (.CI(n44829), .I0(n15630[15]), .I1(GND_net), 
            .CO(n44830));
    SB_LUT4 i39841_3_lut (.I0(n6_adj_5100), .I1(n382[10]), .I2(n356[10]), 
            .I3(GND_net), .O(n55672));   // verilog/motorControl.v(51[33:53])
    defparam i39841_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 add_5232_17_lut (.I0(GND_net), .I1(n15630[14]), .I2(GND_net), 
            .I3(n44828), .O(n14946[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5232_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_18_12_lut (.I0(GND_net), .I1(n257[10]), .I2(n306[10]), 
            .I3(n43758), .O(n356[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i39842_3_lut (.I0(n55672), .I1(n382[11]), .I2(n356[11]), .I3(GND_net), 
            .O(n55673));   // verilog/motorControl.v(51[33:53])
    defparam i39842_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i38897_4_lut (.I0(n356[21]), .I1(n57151), .I2(n382[21]), .I3(n55134), 
            .O(n54727));
    defparam i38897_4_lut.LUT_INIT = 16'h5a7b;
    SB_CARRY counter_2283_add_4_4 (.CI(n44534), .I0(GND_net), .I1(counter[2]), 
            .CO(n44535));
    SB_LUT4 mult_16_i128_2_lut (.I0(\Kp[2] ), .I1(n1[14]), .I2(GND_net), 
            .I3(GND_net), .O(n189_adj_5105));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i128_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i224_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [13]), 
            .I2(GND_net), .I3(GND_net), .O(n332_adj_5106));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i224_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 counter_2283_add_4_3_lut (.I0(GND_net), .I1(GND_net), .I2(counter[1]), 
            .I3(n44533), .O(n28[1])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2283_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_2283_add_4_3 (.CI(n44533), .I0(GND_net), .I1(counter[1]), 
            .CO(n44534));
    SB_LUT4 counter_2283_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(counter[0]), 
            .I3(VCC_net), .O(n28[0])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2283_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5507_8_lut (.I0(GND_net), .I1(n19282[5]), .I2(n560), .I3(n44996), 
            .O(n19170[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5507_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5232_17 (.CI(n44828), .I0(n15630[14]), .I1(GND_net), 
            .CO(n44829));
    SB_LUT4 mult_16_i510_2_lut (.I0(\Kp[10] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n758_adj_5108));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i510_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5232_16_lut (.I0(GND_net), .I1(n15630[13]), .I2(n1111_adj_5109), 
            .I3(n44827), .O(n14946[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5232_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i39637_4_lut (.I0(n24_adj_5039), .I1(n8_adj_5037), .I2(n57126), 
            .I3(n54725), .O(n55468));   // verilog/motorControl.v(51[33:53])
    defparam i39637_4_lut.LUT_INIT = 16'haaac;
    SB_CARRY counter_2283_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(counter[0]), 
            .CO(n44533));
    SB_CARRY add_18_12 (.CI(n43758), .I0(n257[10]), .I1(n306[10]), .CO(n43759));
    SB_LUT4 i39772_3_lut (.I0(n55673), .I1(n382[12]), .I2(n356[12]), .I3(GND_net), 
            .O(n55603));   // verilog/motorControl.v(51[33:53])
    defparam i39772_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 add_18_11_lut (.I0(GND_net), .I1(n257[9]), .I2(n306[9]), .I3(n43757), 
            .O(n356[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i40024_3_lut (.I0(n55889), .I1(n382[19]), .I2(n356[19]), .I3(GND_net), 
            .O(n55855));   // verilog/motorControl.v(51[33:53])
    defparam i40024_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i38899_4_lut (.I0(n356[21]), .I1(n57128), .I2(n382[21]), .I3(n55820), 
            .O(n54729));
    defparam i38899_4_lut.LUT_INIT = 16'h5a7b;
    SB_LUT4 mult_16_i247_2_lut (.I0(\Kp[5] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n366_adj_5111));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i247_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_21_i45_rep_159_2_lut (.I0(n356[22]), .I1(n382[22]), 
            .I2(GND_net), .I3(GND_net), .O(n57126));   // verilog/motorControl.v(51[33:53])
    defparam LessThan_21_i45_rep_159_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i39897_4_lut (.I0(n55603), .I1(n55468), .I2(n57126), .I3(n54727), 
            .O(n55728));   // verilog/motorControl.v(51[33:53])
    defparam i39897_4_lut.LUT_INIT = 16'hccca;
    SB_CARRY add_18_11 (.CI(n43757), .I0(n257[9]), .I1(n306[9]), .CO(n43758));
    SB_LUT4 mult_17_i273_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [13]), 
            .I2(GND_net), .I3(GND_net), .O(n405_adj_5112));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i273_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i322_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [13]), 
            .I2(GND_net), .I3(GND_net), .O(n478_adj_5113));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i322_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i371_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [13]), 
            .I2(GND_net), .I3(GND_net), .O(n551_adj_5114));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i371_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i40006_3_lut (.I0(n55855), .I1(n382[20]), .I2(n356[20]), .I3(GND_net), 
            .O(n40_adj_5115));   // verilog/motorControl.v(51[33:53])
    defparam i40006_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 LessThan_19_i4_4_lut (.I0(deadband[0]), .I1(n356[1]), .I2(deadband[1]), 
            .I3(n356[0]), .O(n4_adj_5116));   // verilog/motorControl.v(51[12:29])
    defparam LessThan_19_i4_4_lut.LUT_INIT = 16'h4d0c;
    SB_LUT4 i39731_3_lut (.I0(n4_adj_5116), .I1(n356[13]), .I2(n27_adj_5032), 
            .I3(GND_net), .O(n55562));   // verilog/motorControl.v(51[12:29])
    defparam i39731_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_16_i177_2_lut (.I0(\Kp[3] ), .I1(n1[14]), .I2(GND_net), 
            .I3(GND_net), .O(n262));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i177_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i39732_3_lut (.I0(n55562), .I1(n356[14]), .I2(n29_adj_5020), 
            .I3(GND_net), .O(n55563));   // verilog/motorControl.v(51[12:29])
    defparam i39732_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i38998_4_lut (.I0(n33_adj_5028), .I1(n31_adj_5021), .I2(n29_adj_5020), 
            .I3(n54835), .O(n54828));
    defparam i38998_4_lut.LUT_INIT = 16'haaab;
    SB_DFFSR counter_2283__i31 (.Q(counter[31]), .C(clk16MHz), .D(n28[31]), 
            .R(counter_31__N_3995));   // verilog/motorControl.v(24[16:25])
    SB_LUT4 i39977_4_lut (.I0(n30_adj_5070), .I1(n10_adj_5066), .I2(n35_adj_5026), 
            .I3(n54826), .O(n55808));   // verilog/motorControl.v(51[12:29])
    defparam i39977_4_lut.LUT_INIT = 16'haaac;
    SB_DFFSR counter_2283__i30 (.Q(counter[30]), .C(clk16MHz), .D(n28[30]), 
            .R(counter_31__N_3995));   // verilog/motorControl.v(24[16:25])
    SB_LUT4 mult_17_i410_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n609_adj_5117));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i410_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i134_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [17]), 
            .I2(GND_net), .I3(GND_net), .O(n198_adj_5118));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i134_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_26_inv_0_i20_1_lut (.I0(PWMLimit[19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5401[19]));   // verilog/motorControl.v(55[22:31])
    defparam unary_minus_26_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_DFFSR counter_2283__i29 (.Q(counter[29]), .C(clk16MHz), .D(n28[29]), 
            .R(counter_31__N_3995));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_2283__i28 (.Q(counter[28]), .C(clk16MHz), .D(n28[28]), 
            .R(counter_31__N_3995));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_2283__i27 (.Q(counter[27]), .C(clk16MHz), .D(n28[27]), 
            .R(counter_31__N_3995));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_2283__i26 (.Q(counter[26]), .C(clk16MHz), .D(n28[26]), 
            .R(counter_31__N_3995));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_2283__i25 (.Q(counter[25]), .C(clk16MHz), .D(n28[25]), 
            .R(counter_31__N_3995));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_2283__i24 (.Q(counter[24]), .C(clk16MHz), .D(n28[24]), 
            .R(counter_31__N_3995));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_2283__i23 (.Q(counter[23]), .C(clk16MHz), .D(n28[23]), 
            .R(counter_31__N_3995));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_2283__i22 (.Q(counter[22]), .C(clk16MHz), .D(n28[22]), 
            .R(counter_31__N_3995));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_2283__i21 (.Q(counter[21]), .C(clk16MHz), .D(n28[21]), 
            .R(counter_31__N_3995));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_2283__i20 (.Q(counter[20]), .C(clk16MHz), .D(n28[20]), 
            .R(counter_31__N_3995));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_2283__i19 (.Q(counter[19]), .C(clk16MHz), .D(n28[19]), 
            .R(counter_31__N_3995));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_2283__i18 (.Q(counter[18]), .C(clk16MHz), .D(n28[18]), 
            .R(counter_31__N_3995));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_2283__i17 (.Q(counter[17]), .C(clk16MHz), .D(n28[17]), 
            .R(counter_31__N_3995));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_2283__i16 (.Q(counter[16]), .C(clk16MHz), .D(n28[16]), 
            .R(counter_31__N_3995));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_2283__i15 (.Q(counter[15]), .C(clk16MHz), .D(n28[15]), 
            .R(counter_31__N_3995));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_2283__i14 (.Q(counter[14]), .C(clk16MHz), .D(n28[14]), 
            .R(counter_31__N_3995));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_2283__i13 (.Q(counter[13]), .C(clk16MHz), .D(n28[13]), 
            .R(counter_31__N_3995));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_2283__i12 (.Q(counter[12]), .C(clk16MHz), .D(n28[12]), 
            .R(counter_31__N_3995));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_2283__i11 (.Q(counter[11]), .C(clk16MHz), .D(n28[11]), 
            .R(counter_31__N_3995));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_2283__i10 (.Q(counter[10]), .C(clk16MHz), .D(n28[10]), 
            .R(counter_31__N_3995));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_2283__i9 (.Q(counter[9]), .C(clk16MHz), .D(n28[9]), 
            .R(counter_31__N_3995));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_2283__i8 (.Q(counter[8]), .C(clk16MHz), .D(n28[8]), 
            .R(counter_31__N_3995));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_2283__i7 (.Q(counter[7]), .C(clk16MHz), .D(n28[7]), 
            .R(counter_31__N_3995));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_2283__i6 (.Q(counter[6]), .C(clk16MHz), .D(n28[6]), 
            .R(counter_31__N_3995));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_2283__i5 (.Q(counter[5]), .C(clk16MHz), .D(n28[5]), 
            .R(counter_31__N_3995));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_2283__i4 (.Q(counter[4]), .C(clk16MHz), .D(n28[4]), 
            .R(counter_31__N_3995));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_2283__i3 (.Q(counter[3]), .C(clk16MHz), .D(n28[3]), 
            .R(counter_31__N_3995));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_2283__i2 (.Q(counter[2]), .C(clk16MHz), .D(n28[2]), 
            .R(counter_31__N_3995));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_2283__i1 (.Q(counter[1]), .C(clk16MHz), .D(n28[1]), 
            .R(counter_31__N_3995));   // verilog/motorControl.v(24[16:25])
    SB_LUT4 i39374_3_lut (.I0(n55563), .I1(n356[15]), .I2(n31_adj_5021), 
            .I3(GND_net), .O(n55205));   // verilog/motorControl.v(51[12:29])
    defparam i39374_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_26_inv_0_i21_1_lut (.I0(PWMLimit[20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5401[20]));   // verilog/motorControl.v(55[22:31])
    defparam unary_minus_26_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i40055_4_lut (.I0(n55205), .I1(n55808), .I2(n35_adj_5026), 
            .I3(n54828), .O(n55886));   // verilog/motorControl.v(51[12:29])
    defparam i40055_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i40056_3_lut (.I0(n55886), .I1(n356[18]), .I2(n37_adj_5016), 
            .I3(GND_net), .O(n55887));   // verilog/motorControl.v(51[12:29])
    defparam i40056_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i40026_3_lut (.I0(n55887), .I1(n356[19]), .I2(n39_adj_5013), 
            .I3(GND_net), .O(n55857));   // verilog/motorControl.v(51[12:29])
    defparam i40026_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i38952_4_lut (.I0(n43_adj_5015), .I1(n41_adj_5012), .I2(n39_adj_5013), 
            .I3(n55798), .O(n54782));
    defparam i38952_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i39891_4_lut (.I0(n55203), .I1(n55466), .I2(n45_adj_5014), 
            .I3(n54780), .O(n55722));   // verilog/motorControl.v(51[12:29])
    defparam i39891_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 mult_16_i226_2_lut (.I0(\Kp[4] ), .I1(n1[14]), .I2(GND_net), 
            .I3(GND_net), .O(n335_adj_5121));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i226_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i420_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [13]), 
            .I2(GND_net), .I3(GND_net), .O(n624_adj_5122));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i420_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i402_2_lut (.I0(\Kp[8] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n597_adj_5123));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i402_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i469_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [13]), 
            .I2(GND_net), .I3(GND_net), .O(n697_adj_5124));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i469_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i40004_3_lut (.I0(n55857), .I1(n356[20]), .I2(n41_adj_5012), 
            .I3(GND_net), .O(n40_adj_5125));   // verilog/motorControl.v(51[12:29])
    defparam i40004_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i39893_4_lut (.I0(n40_adj_5125), .I1(n55722), .I2(n45_adj_5014), 
            .I3(n54782), .O(n55724));   // verilog/motorControl.v(51[12:29])
    defparam i39893_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i39899_4_lut (.I0(n40_adj_5115), .I1(n55728), .I2(n57126), 
            .I3(n54729), .O(n55730));   // verilog/motorControl.v(51[33:53])
    defparam i39899_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 mult_16_i396_2_lut (.I0(\Kp[8] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n588_adj_5126));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i396_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5507_7_lut (.I0(GND_net), .I1(n19282[4]), .I2(n487), .I3(n44995), 
            .O(n19170[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5507_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5232_16 (.CI(n44827), .I0(n15630[13]), .I1(n1111_adj_5109), 
            .CO(n44828));
    SB_LUT4 mux_14_i14_3_lut (.I0(n130[13]), .I1(n182[13]), .I2(n181), 
            .I3(GND_net), .O(n207[13]));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_14_i14_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_15_i14_3_lut (.I0(n207[13]), .I1(IntegralLimit[13]), .I2(n155), 
            .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3996 [13]));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_15_i14_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_17_i518_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [13]), 
            .I2(GND_net), .I3(GND_net), .O(n770_adj_5127));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i518_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut_adj_1680 (.I0(n55724), .I1(control_update), .I2(deadband[23]), 
            .I3(n356[23]), .O(n52322));
    defparam i1_4_lut_adj_1680.LUT_INIT = 16'h4c04;
    SB_LUT4 i1_4_lut_adj_1681 (.I0(n52322), .I1(n55730), .I2(n356[23]), 
            .I3(n47_adj_5128), .O(n29330));
    defparam i1_4_lut_adj_1681.LUT_INIT = 16'h0a22;
    SB_LUT4 add_18_10_lut (.I0(GND_net), .I1(n257[8]), .I2(n306[8]), .I3(n43756), 
            .O(n356[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_18_10 (.CI(n43756), .I0(n257[8]), .I1(n306[8]), .CO(n43757));
    SB_LUT4 add_5232_15_lut (.I0(GND_net), .I1(n15630[12]), .I2(n1038_adj_5129), 
            .I3(n44826), .O(n14946[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5232_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5232_15 (.CI(n44826), .I0(n15630[12]), .I1(n1038_adj_5129), 
            .CO(n44827));
    SB_LUT4 add_5232_14_lut (.I0(GND_net), .I1(n15630[11]), .I2(n965), 
            .I3(n44825), .O(n14946[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5232_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5093_12 (.CI(n45140), .I0(n12905[9]), .I1(n807), .CO(n45141));
    SB_CARRY add_5214_14 (.CI(n45085), .I0(n15306[11]), .I1(n962_adj_5076), 
            .CO(n45086));
    SB_LUT4 add_5093_11_lut (.I0(GND_net), .I1(n12905[8]), .I2(n734), 
            .I3(n45139), .O(n11935[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5093_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i275_2_lut (.I0(\Kp[5] ), .I1(n1[14]), .I2(GND_net), 
            .I3(GND_net), .O(n408));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i275_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_18_9_lut (.I0(GND_net), .I1(n257[7]), .I2(n306[7]), .I3(n43755), 
            .O(n356[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5214_13_lut (.I0(GND_net), .I1(n15306[10]), .I2(n889_adj_5130), 
            .I3(n45084), .O(n14585[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5214_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i324_2_lut (.I0(\Kp[6] ), .I1(n1[14]), .I2(GND_net), 
            .I3(GND_net), .O(n481));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i324_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5232_14 (.CI(n44825), .I0(n15630[11]), .I1(n965), .CO(n44826));
    SB_CARRY add_18_9 (.CI(n43755), .I0(n257[7]), .I1(n306[7]), .CO(n43756));
    SB_CARRY add_5507_7 (.CI(n44995), .I0(n19282[4]), .I1(n487), .CO(n44996));
    SB_LUT4 add_5507_6_lut (.I0(GND_net), .I1(n19282[3]), .I2(n414), .I3(n44994), 
            .O(n19170[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5507_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_18_8_lut (.I0(GND_net), .I1(n257[6]), .I2(n306[6]), .I3(n43754), 
            .O(n356[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5232_13_lut (.I0(GND_net), .I1(n15630[10]), .I2(n892), 
            .I3(n44824), .O(n14946[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5232_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5093_11 (.CI(n45139), .I0(n12905[8]), .I1(n734), .CO(n45140));
    SB_CARRY add_5232_13 (.CI(n44824), .I0(n15630[10]), .I1(n892), .CO(n44825));
    SB_CARRY add_5214_13 (.CI(n45084), .I0(n15306[10]), .I1(n889_adj_5130), 
            .CO(n45085));
    SB_CARRY add_18_8 (.CI(n43754), .I0(n257[6]), .I1(n306[6]), .CO(n43755));
    SB_LUT4 add_18_7_lut (.I0(GND_net), .I1(n257[5]), .I2(n306[5]), .I3(n43753), 
            .O(n356[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_18_7 (.CI(n43753), .I0(n257[5]), .I1(n306[5]), .CO(n43754));
    SB_LUT4 add_18_6_lut (.I0(GND_net), .I1(n257[4]), .I2(n306[4]), .I3(n43752), 
            .O(n356[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5507_6 (.CI(n44994), .I0(n19282[3]), .I1(n414), .CO(n44995));
    SB_LUT4 add_5507_5_lut (.I0(GND_net), .I1(n19282[2]), .I2(n341_adj_5132), 
            .I3(n44993), .O(n19170[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5507_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5232_12_lut (.I0(GND_net), .I1(n15630[9]), .I2(n819), 
            .I3(n44823), .O(n14946[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5232_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5232_12 (.CI(n44823), .I0(n15630[9]), .I1(n819), .CO(n44824));
    SB_LUT4 add_5214_12_lut (.I0(GND_net), .I1(n15306[9]), .I2(n816_adj_5133), 
            .I3(n45083), .O(n14585[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5214_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5507_5 (.CI(n44993), .I0(n19282[2]), .I1(n341_adj_5132), 
            .CO(n44994));
    SB_LUT4 add_5232_11_lut (.I0(GND_net), .I1(n15630[8]), .I2(n746), 
            .I3(n44822), .O(n14946[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5232_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_18_6 (.CI(n43752), .I0(n257[4]), .I1(n306[4]), .CO(n43753));
    SB_CARRY add_5232_11 (.CI(n44822), .I0(n15630[8]), .I1(n746), .CO(n44823));
    SB_LUT4 add_5232_10_lut (.I0(GND_net), .I1(n15630[7]), .I2(n673), 
            .I3(n44821), .O(n14946[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5232_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_18_5_lut (.I0(GND_net), .I1(n257[3]), .I2(n306[3]), .I3(n43751), 
            .O(n356[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_18_5 (.CI(n43751), .I0(n257[3]), .I1(n306[3]), .CO(n43752));
    SB_CARRY add_5232_10 (.CI(n44821), .I0(n15630[7]), .I1(n673), .CO(n44822));
    SB_LUT4 add_18_4_lut (.I0(GND_net), .I1(n257[2]), .I2(n306[2]), .I3(n43750), 
            .O(n356[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5232_9_lut (.I0(GND_net), .I1(n15630[6]), .I2(n600), .I3(n44820), 
            .O(n14946[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5232_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_18_4 (.CI(n43750), .I0(n257[2]), .I1(n306[2]), .CO(n43751));
    SB_CARRY add_5214_12 (.CI(n45083), .I0(n15306[9]), .I1(n816_adj_5133), 
            .CO(n45084));
    SB_LUT4 add_5507_4_lut (.I0(GND_net), .I1(n19282[1]), .I2(n268), .I3(n44992), 
            .O(n19170[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5507_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_18_3_lut (.I0(GND_net), .I1(n257[1]), .I2(n306[1]), .I3(n43749), 
            .O(n356[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_18_3 (.CI(n43749), .I0(n257[1]), .I1(n306[1]), .CO(n43750));
    SB_LUT4 add_18_2_lut (.I0(GND_net), .I1(n257[0]), .I2(n306[0]), .I3(GND_net), 
            .O(n356[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5507_4 (.CI(n44992), .I0(n19282[1]), .I1(n268), .CO(n44993));
    SB_CARRY add_5232_9 (.CI(n44820), .I0(n15630[6]), .I1(n600), .CO(n44821));
    SB_LUT4 add_5232_8_lut (.I0(GND_net), .I1(n15630[5]), .I2(n527), .I3(n44819), 
            .O(n14946[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5232_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_18_2 (.CI(GND_net), .I0(n257[0]), .I1(n306[0]), .CO(n43749));
    SB_LUT4 add_9_25_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [23]), 
            .I2(n1[23]), .I3(n43748), .O(n130[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5232_8 (.CI(n44819), .I0(n15630[5]), .I1(n527), .CO(n44820));
    SB_LUT4 add_9_24_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [22]), 
            .I2(n1[22]), .I3(n43747), .O(n130[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5214_11_lut (.I0(GND_net), .I1(n15306[8]), .I2(n743_adj_5136), 
            .I3(n45082), .O(n14585[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5214_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5232_7_lut (.I0(GND_net), .I1(n15630[4]), .I2(n454_adj_5137), 
            .I3(n44818), .O(n14946[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5232_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_9_24 (.CI(n43747), .I0(\PID_CONTROLLER.integral [22]), 
            .I1(n1[22]), .CO(n43748));
    SB_CARRY add_5232_7 (.CI(n44818), .I0(n15630[4]), .I1(n454_adj_5137), 
            .CO(n44819));
    SB_LUT4 add_9_23_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [21]), 
            .I2(n1[21]), .I3(n43746), .O(n130[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_9_23 (.CI(n43746), .I0(\PID_CONTROLLER.integral [21]), 
            .I1(n1[21]), .CO(n43747));
    SB_LUT4 add_9_22_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [20]), 
            .I2(n1[20]), .I3(n43745), .O(n130[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5214_11 (.CI(n45082), .I0(n15306[8]), .I1(n743_adj_5136), 
            .CO(n45083));
    SB_CARRY add_9_22 (.CI(n43745), .I0(\PID_CONTROLLER.integral [20]), 
            .I1(n1[20]), .CO(n43746));
    SB_LUT4 add_5232_6_lut (.I0(GND_net), .I1(n15630[3]), .I2(n381), .I3(n44817), 
            .O(n14946[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5232_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5507_3_lut (.I0(GND_net), .I1(n19282[0]), .I2(n195_adj_5138), 
            .I3(n44991), .O(n19170[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5507_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5232_6 (.CI(n44817), .I0(n15630[3]), .I1(n381), .CO(n44818));
    SB_LUT4 add_9_21_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [19]), 
            .I2(n1[19]), .I3(n43744), .O(n130[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i373_2_lut (.I0(\Kp[7] ), .I1(n1[14]), .I2(GND_net), 
            .I3(GND_net), .O(n554));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i373_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5093_10_lut (.I0(GND_net), .I1(n12905[7]), .I2(n661_adj_5139), 
            .I3(n45138), .O(n11935[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5093_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5214_10_lut (.I0(GND_net), .I1(n15306[7]), .I2(n670_adj_5140), 
            .I3(n45081), .O(n14585[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5214_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_9_21 (.CI(n43744), .I0(\PID_CONTROLLER.integral [19]), 
            .I1(n1[19]), .CO(n43745));
    SB_CARRY add_5507_3 (.CI(n44991), .I0(n19282[0]), .I1(n195_adj_5138), 
            .CO(n44992));
    SB_LUT4 add_5507_2_lut (.I0(GND_net), .I1(n53), .I2(n122_adj_5141), 
            .I3(GND_net), .O(n19170[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5507_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_9_20_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [18]), 
            .I2(n1[18]), .I3(n43743), .O(n130[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_9_20 (.CI(n43743), .I0(\PID_CONTROLLER.integral [18]), 
            .I1(n1[18]), .CO(n43744));
    SB_LUT4 add_5232_5_lut (.I0(GND_net), .I1(n15630[2]), .I2(n308), .I3(n44816), 
            .O(n14946[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5232_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5232_5 (.CI(n44816), .I0(n15630[2]), .I1(n308), .CO(n44817));
    SB_LUT4 add_9_19_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [17]), 
            .I2(n1[17]), .I3(n43742), .O(n130[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_9_19 (.CI(n43742), .I0(\PID_CONTROLLER.integral [17]), 
            .I1(n1[17]), .CO(n43743));
    SB_LUT4 add_9_18_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [16]), 
            .I2(n1[16]), .I3(n43741), .O(n130[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5093_10 (.CI(n45138), .I0(n12905[7]), .I1(n661_adj_5139), 
            .CO(n45139));
    SB_CARRY add_9_18 (.CI(n43741), .I0(\PID_CONTROLLER.integral [16]), 
            .I1(n1[16]), .CO(n43742));
    SB_LUT4 add_9_17_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [15]), 
            .I2(n1[15]), .I3(n43740), .O(n130[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5214_10 (.CI(n45081), .I0(n15306[7]), .I1(n670_adj_5140), 
            .CO(n45082));
    SB_CARRY add_9_17 (.CI(n43740), .I0(\PID_CONTROLLER.integral [15]), 
            .I1(n1[15]), .CO(n43741));
    SB_LUT4 add_9_16_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [14]), 
            .I2(n1[14]), .I3(n43739), .O(n130[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_9_16 (.CI(n43739), .I0(\PID_CONTROLLER.integral [14]), 
            .I1(n1[14]), .CO(n43740));
    SB_LUT4 add_9_15_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [13]), 
            .I2(n1[13]), .I3(n43738), .O(n130[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_9_15 (.CI(n43738), .I0(\PID_CONTROLLER.integral [13]), 
            .I1(n1[13]), .CO(n43739));
    SB_CARRY add_5507_2 (.CI(GND_net), .I0(n53), .I1(n122_adj_5141), .CO(n44991));
    SB_LUT4 add_9_14_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [12]), 
            .I2(n1[12]), .I3(n43737), .O(n130[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5232_4_lut (.I0(GND_net), .I1(n15630[1]), .I2(n235), .I3(n44815), 
            .O(n14946[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5232_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5232_4 (.CI(n44815), .I0(n15630[1]), .I1(n235), .CO(n44816));
    SB_LUT4 add_5232_3_lut (.I0(GND_net), .I1(n15630[0]), .I2(n162_adj_5143), 
            .I3(n44814), .O(n14946[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5232_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i296_2_lut (.I0(\Kp[6] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n439_adj_5144));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i296_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_9_14 (.CI(n43737), .I0(\PID_CONTROLLER.integral [12]), 
            .I1(n1[12]), .CO(n43738));
    SB_LUT4 add_5374_15_lut (.I0(GND_net), .I1(n17881[12]), .I2(n1050_adj_5145), 
            .I3(n44990), .O(n17490[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5374_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_9_13_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [11]), 
            .I2(n1[11]), .I3(n43736), .O(n130[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_i51_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n74_adj_5146));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i51_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i4_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n5_adj_5147));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i4_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_9_13 (.CI(n43736), .I0(\PID_CONTROLLER.integral [11]), 
            .I1(n1[11]), .CO(n43737));
    SB_LUT4 add_9_12_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [10]), 
            .I2(n1[10]), .I3(n43735), .O(n130[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_9_12 (.CI(n43735), .I0(\PID_CONTROLLER.integral [10]), 
            .I1(n1[10]), .CO(n43736));
    SB_LUT4 mult_16_i345_2_lut (.I0(\Kp[7] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n512));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i345_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5374_14_lut (.I0(GND_net), .I1(n17881[11]), .I2(n977_adj_5148), 
            .I3(n44989), .O(n17490[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5374_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_9_11_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(n1[9]), .I3(n43734), .O(n130[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_9_11 (.CI(n43734), .I0(\PID_CONTROLLER.integral [9]), .I1(n1[9]), 
            .CO(n43735));
    SB_CARRY add_5232_3 (.CI(n44814), .I0(n15630[0]), .I1(n162_adj_5143), 
            .CO(n44815));
    SB_LUT4 add_9_10_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(n1[8]), .I3(n43733), .O(n130[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_9_10 (.CI(n43733), .I0(\PID_CONTROLLER.integral [8]), .I1(n1[8]), 
            .CO(n43734));
    SB_LUT4 mult_16_i455_2_lut (.I0(\Kp[9] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n676_adj_5149));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i455_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i100_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n147_adj_5150));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i100_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_9_9_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(n1[7]), .I3(n43732), .O(n130[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_9_9 (.CI(n43732), .I0(\PID_CONTROLLER.integral [7]), .I1(n1[7]), 
            .CO(n43733));
    SB_LUT4 add_5232_2_lut (.I0(GND_net), .I1(n20_adj_5151), .I2(n89), 
            .I3(GND_net), .O(n14946[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5232_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5232_2 (.CI(GND_net), .I0(n20_adj_5151), .I1(n89), .CO(n44814));
    SB_CARRY add_5374_14 (.CI(n44989), .I0(n17881[11]), .I1(n977_adj_5148), 
            .CO(n44990));
    SB_LUT4 add_9_8_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(n1[6]), .I3(n43731), .O(n130[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i559_2_lut (.I0(\Kp[11] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n831_adj_5152));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i559_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i422_2_lut (.I0(\Kp[8] ), .I1(n1[14]), .I2(GND_net), 
            .I3(GND_net), .O(n627));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i422_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i149_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n220_adj_5153));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i149_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i55_2_lut (.I0(\Kp[1] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n80_adj_5154));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i55_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_9_8 (.CI(n43731), .I0(\PID_CONTROLLER.integral [6]), .I1(n1[6]), 
            .CO(n43732));
    SB_LUT4 add_5484_10_lut (.I0(GND_net), .I1(n19106[7]), .I2(n700), 
            .I3(n44813), .O(n18945[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5484_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_9_7_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(n1[5]), .I3(n43730), .O(n130[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_9_7 (.CI(n43730), .I0(\PID_CONTROLLER.integral [5]), .I1(n1[5]), 
            .CO(n43731));
    SB_LUT4 add_9_6_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(n1[4]), .I3(n43729), .O(n130[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i8_2_lut (.I0(\Kp[0] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n11_adj_5155));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i8_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5374_13_lut (.I0(GND_net), .I1(n17881[10]), .I2(n904_adj_5156), 
            .I3(n44988), .O(n17490[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5374_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_9_6 (.CI(n43729), .I0(\PID_CONTROLLER.integral [4]), .I1(n1[4]), 
            .CO(n43730));
    SB_LUT4 add_9_5_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(n1[3]), .I3(n43728), .O(n130[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5484_9_lut (.I0(GND_net), .I1(n19106[6]), .I2(n627), .I3(n44812), 
            .O(n18945[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5484_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5374_13 (.CI(n44988), .I0(n17881[10]), .I1(n904_adj_5156), 
            .CO(n44989));
    SB_CARRY add_5484_9 (.CI(n44812), .I0(n19106[6]), .I1(n627), .CO(n44813));
    SB_LUT4 add_5374_12_lut (.I0(GND_net), .I1(n17881[9]), .I2(n831_adj_5152), 
            .I3(n44987), .O(n17490[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5374_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5484_8_lut (.I0(GND_net), .I1(n19106[5]), .I2(n554), .I3(n44811), 
            .O(n18945[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5484_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_9_5 (.CI(n43728), .I0(\PID_CONTROLLER.integral [3]), .I1(n1[3]), 
            .CO(n43729));
    SB_LUT4 add_9_4_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(n1[2]), .I3(n43727), .O(n130[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_9_4 (.CI(n43727), .I0(\PID_CONTROLLER.integral [2]), .I1(n1[2]), 
            .CO(n43728));
    SB_LUT4 add_9_3_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(n1[1]), .I3(n43726), .O(n130[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_i198_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n293_adj_5158));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i198_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i504_2_lut (.I0(\Kp[10] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n749_adj_5159));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i504_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i608_2_lut (.I0(\Kp[12] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n904_adj_5156));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i608_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5484_8 (.CI(n44811), .I0(n19106[5]), .I1(n554), .CO(n44812));
    SB_LUT4 mult_17_i247_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n366_adj_5160));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i247_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i394_2_lut (.I0(\Kp[8] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n585));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i394_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5484_7_lut (.I0(GND_net), .I1(n19106[4]), .I2(n481), .I3(n44810), 
            .O(n18945[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5484_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5484_7 (.CI(n44810), .I0(n19106[4]), .I1(n481), .CO(n44811));
    SB_CARRY add_9_3 (.CI(n43726), .I0(\PID_CONTROLLER.integral [1]), .I1(n1[1]), 
            .CO(n43727));
    SB_LUT4 add_9_2_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [0]), 
            .I2(n1[0]), .I3(GND_net), .O(n130[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5484_6_lut (.I0(GND_net), .I1(n19106[3]), .I2(n408), .I3(n44809), 
            .O(n18945[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5484_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5456_11_lut (.I0(GND_net), .I1(n18846[8]), .I2(n770_adj_5127), 
            .I3(n43931), .O(n18626[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5456_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5093_9_lut (.I0(GND_net), .I1(n12905[6]), .I2(n588_adj_5126), 
            .I3(n45137), .O(n11935[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5093_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5456_10_lut (.I0(GND_net), .I1(n18846[7]), .I2(n697_adj_5124), 
            .I3(n43930), .O(n18626[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5456_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5484_6 (.CI(n44809), .I0(n19106[3]), .I1(n408), .CO(n44810));
    SB_CARRY add_5456_10 (.CI(n43930), .I0(n18846[7]), .I1(n697_adj_5124), 
            .CO(n43931));
    SB_LUT4 add_5214_9_lut (.I0(GND_net), .I1(n15306[6]), .I2(n597_adj_5123), 
            .I3(n45080), .O(n14585[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5214_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5374_12 (.CI(n44987), .I0(n17881[9]), .I1(n831_adj_5152), 
            .CO(n44988));
    SB_LUT4 add_5456_9_lut (.I0(GND_net), .I1(n18846[6]), .I2(n624_adj_5122), 
            .I3(n43929), .O(n18626[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5456_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5484_5_lut (.I0(GND_net), .I1(n19106[2]), .I2(n335_adj_5121), 
            .I3(n44808), .O(n18945[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5484_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i471_2_lut (.I0(\Kp[9] ), .I1(n1[14]), .I2(GND_net), 
            .I3(GND_net), .O(n700));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i471_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_14_i7_3_lut (.I0(n130[6]), .I1(n182[6]), .I2(n181), .I3(GND_net), 
            .O(n207[6]));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_14_i7_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_9_2 (.CI(GND_net), .I0(\PID_CONTROLLER.integral [0]), .I1(n1[0]), 
            .CO(n43726));
    SB_LUT4 mult_17_i296_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n439_adj_5161));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i296_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5484_5 (.CI(n44808), .I0(n19106[2]), .I1(n335_adj_5121), 
            .CO(n44809));
    SB_LUT4 mux_15_i7_3_lut (.I0(n207[6]), .I1(IntegralLimit[6]), .I2(n155), 
            .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3996 [6]));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_15_i7_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_17_i61_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n89));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i61_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i14_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n20_adj_5151));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i14_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i553_2_lut (.I0(\Kp[11] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n822_adj_5162));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i553_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i345_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n512_adj_5163));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i345_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5484_4_lut (.I0(GND_net), .I1(n19106[1]), .I2(n262), .I3(n44807), 
            .O(n18945[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5484_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5456_9 (.CI(n43929), .I0(n18846[6]), .I1(n624_adj_5122), 
            .CO(n43930));
    SB_LUT4 mult_16_i104_2_lut (.I0(\Kp[2] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n153_adj_5164));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i104_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i602_2_lut (.I0(\Kp[12] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n895_adj_5165));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i602_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5456_8_lut (.I0(GND_net), .I1(n18846[5]), .I2(n551_adj_5114), 
            .I3(n43928), .O(n18626[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5456_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5456_8 (.CI(n43928), .I0(n18846[5]), .I1(n551_adj_5114), 
            .CO(n43929));
    SB_LUT4 add_5456_7_lut (.I0(GND_net), .I1(n18846[4]), .I2(n478_adj_5113), 
            .I3(n43927), .O(n18626[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5456_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_i394_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n585_adj_5166));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i394_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5456_7 (.CI(n43927), .I0(n18846[4]), .I1(n478_adj_5113), 
            .CO(n43928));
    SB_LUT4 mult_16_i657_2_lut (.I0(\Kp[13] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n977_adj_5148));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i657_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i153_2_lut (.I0(\Kp[3] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n226_adj_5167));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i153_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5484_4 (.CI(n44807), .I0(n19106[1]), .I1(n262), .CO(n44808));
    SB_LUT4 add_5456_6_lut (.I0(GND_net), .I1(n18846[3]), .I2(n405_adj_5112), 
            .I3(n43926), .O(n18626[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5456_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14957_3_lut (.I0(n356[1]), .I1(n436[1]), .I2(n10860), .I3(GND_net), 
            .O(n29028));   // verilog/motorControl.v(41[14] 61[8])
    defparam i14957_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_5374_11_lut (.I0(GND_net), .I1(n17881[8]), .I2(n758_adj_5108), 
            .I3(n44986), .O(n17490[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5374_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5093_9 (.CI(n45137), .I0(n12905[6]), .I1(n588_adj_5126), 
            .CO(n45138));
    SB_LUT4 mult_17_i443_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n658));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i443_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5456_6 (.CI(n43926), .I0(n18846[3]), .I1(n405_adj_5112), 
            .CO(n43927));
    SB_LUT4 mult_16_i443_2_lut (.I0(\Kp[9] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n658_adj_5168));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i443_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5456_5_lut (.I0(GND_net), .I1(n18846[2]), .I2(n332_adj_5106), 
            .I3(n43925), .O(n18626[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5456_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i651_2_lut (.I0(\Kp[13] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n968_adj_5169));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i651_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5484_3_lut (.I0(GND_net), .I1(n19106[0]), .I2(n189_adj_5105), 
            .I3(n44806), .O(n18945[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5484_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5456_5 (.CI(n43925), .I0(n18846[2]), .I1(n332_adj_5106), 
            .CO(n43926));
    SB_LUT4 add_5456_4_lut (.I0(GND_net), .I1(n18846[1]), .I2(n259_adj_5104), 
            .I3(n43924), .O(n18626[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5456_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5374_11 (.CI(n44986), .I0(n17881[8]), .I1(n758_adj_5108), 
            .CO(n44987));
    SB_CARRY add_5456_4 (.CI(n43924), .I0(n18846[1]), .I1(n259_adj_5104), 
            .CO(n43925));
    SB_LUT4 add_5456_3_lut (.I0(GND_net), .I1(n18846[0]), .I2(n186_adj_5103), 
            .I3(n43923), .O(n18626[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5456_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5214_9 (.CI(n45080), .I0(n15306[6]), .I1(n597_adj_5123), 
            .CO(n45081));
    SB_CARRY add_5456_3 (.CI(n43923), .I0(n18846[0]), .I1(n186_adj_5103), 
            .CO(n43924));
    SB_LUT4 add_5214_8_lut (.I0(GND_net), .I1(n15306[5]), .I2(n524_adj_5102), 
            .I3(n45079), .O(n14585[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5214_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i706_2_lut (.I0(\Kp[14] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n1050_adj_5145));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i706_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5456_2_lut (.I0(GND_net), .I1(n44_adj_5101), .I2(n113_adj_5099), 
            .I3(GND_net), .O(n18626[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5456_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5484_3 (.CI(n44806), .I0(n19106[0]), .I1(n189_adj_5105), 
            .CO(n44807));
    SB_LUT4 add_5374_10_lut (.I0(GND_net), .I1(n17881[7]), .I2(n685_adj_5098), 
            .I3(n44985), .O(n17490[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5374_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5484_2_lut (.I0(GND_net), .I1(n47), .I2(n116), .I3(GND_net), 
            .O(n18945[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5484_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5456_2 (.CI(GND_net), .I0(n44_adj_5101), .I1(n113_adj_5099), 
            .CO(n43923));
    SB_CARRY add_5484_2 (.CI(GND_net), .I0(n47), .I1(n116), .CO(n44806));
    SB_LUT4 unary_minus_13_inv_0_i1_1_lut (.I0(IntegralLimit[0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5402[0]));   // verilog/motorControl.v(48[22:36])
    defparam unary_minus_13_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_5214_8 (.CI(n45079), .I0(n15306[5]), .I1(n524_adj_5102), 
            .CO(n45080));
    SB_LUT4 unary_minus_13_inv_0_i2_1_lut (.I0(IntegralLimit[1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5402[1]));   // verilog/motorControl.v(48[22:36])
    defparam unary_minus_13_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_5374_10 (.CI(n44985), .I0(n17881[7]), .I1(n685_adj_5098), 
            .CO(n44986));
    SB_LUT4 add_5267_18_lut (.I0(GND_net), .I1(n16242[15]), .I2(GND_net), 
            .I3(n44805), .O(n15630[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5267_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5267_17_lut (.I0(GND_net), .I1(n16242[14]), .I2(GND_net), 
            .I3(n44804), .O(n15630[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5267_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_13_inv_0_i3_1_lut (.I0(IntegralLimit[2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5402[2]));   // verilog/motorControl.v(48[22:36])
    defparam unary_minus_13_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_17_i110_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n162_adj_5143));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i110_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5214_7_lut (.I0(GND_net), .I1(n15306[4]), .I2(n451_adj_5033), 
            .I3(n45078), .O(n14585[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5214_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5267_17 (.CI(n44804), .I0(n16242[14]), .I1(GND_net), 
            .CO(n44805));
    SB_LUT4 mult_16_i700_2_lut (.I0(\Kp[14] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n1041_adj_5173));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i700_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i159_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n235));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i159_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5374_9_lut (.I0(GND_net), .I1(n17881[6]), .I2(n612_adj_5011), 
            .I3(n44984), .O(n17490[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5374_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5374_9 (.CI(n44984), .I0(n17881[6]), .I1(n612_adj_5011), 
            .CO(n44985));
    SB_LUT4 unary_minus_13_inv_0_i4_1_lut (.I0(IntegralLimit[3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5402[3]));   // verilog/motorControl.v(48[22:36])
    defparam unary_minus_13_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_5267_16_lut (.I0(GND_net), .I1(n16242[13]), .I2(n1114), 
            .I3(n44803), .O(n15630[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5267_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_i492_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n731));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i492_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5267_16 (.CI(n44803), .I0(n16242[13]), .I1(n1114), .CO(n44804));
    SB_LUT4 add_5267_15_lut (.I0(GND_net), .I1(n16242[12]), .I2(n1041), 
            .I3(n44802), .O(n15630[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5267_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5093_8_lut (.I0(GND_net), .I1(n12905[5]), .I2(n515_adj_4984), 
            .I3(n45136), .O(n11935[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5093_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5214_7 (.CI(n45078), .I0(n15306[4]), .I1(n451_adj_5033), 
            .CO(n45079));
    SB_LUT4 add_5374_8_lut (.I0(GND_net), .I1(n17881[5]), .I2(n539_adj_4982), 
            .I3(n44983), .O(n17490[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5374_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5267_15 (.CI(n44802), .I0(n16242[12]), .I1(n1041), .CO(n44803));
    SB_CARRY add_5374_8 (.CI(n44983), .I0(n17881[5]), .I1(n539_adj_4982), 
            .CO(n44984));
    SB_CARRY add_5093_8 (.CI(n45136), .I0(n12905[5]), .I1(n515_adj_4984), 
            .CO(n45137));
    SB_LUT4 unary_minus_13_inv_0_i5_1_lut (.I0(IntegralLimit[4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5402[4]));   // verilog/motorControl.v(48[22:36])
    defparam unary_minus_13_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_13_inv_0_i6_1_lut (.I0(IntegralLimit[5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5402[5]));   // verilog/motorControl.v(48[22:36])
    defparam unary_minus_13_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_13_inv_0_i7_1_lut (.I0(IntegralLimit[6]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5402[6]));   // verilog/motorControl.v(48[22:36])
    defparam unary_minus_13_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_5267_14_lut (.I0(GND_net), .I1(n16242[11]), .I2(n968), 
            .I3(n44801), .O(n15630[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5267_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5214_6_lut (.I0(GND_net), .I1(n15306[3]), .I2(n378_adj_4967), 
            .I3(n45077), .O(n14585[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5214_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5374_7_lut (.I0(GND_net), .I1(n17881[4]), .I2(n466_adj_4962), 
            .I3(n44982), .O(n17490[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5374_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5267_14 (.CI(n44801), .I0(n16242[11]), .I1(n968), .CO(n44802));
    SB_CARRY add_5374_7 (.CI(n44982), .I0(n17881[4]), .I1(n466_adj_4962), 
            .CO(n44983));
    SB_LUT4 add_5267_13_lut (.I0(GND_net), .I1(n16242[10]), .I2(n895), 
            .I3(n44800), .O(n15630[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5267_13_lut.LUT_INIT = 16'hC33C;
    SB_DFFESR result__i0 (.Q(duty[0]), .C(clk16MHz), .E(control_update), 
            .D(n28711), .R(n29330));   // verilog/motorControl.v(41[14] 61[8])
    SB_LUT4 add_5093_7_lut (.I0(GND_net), .I1(n12905[4]), .I2(n442_adj_4943), 
            .I3(n45135), .O(n11935[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5093_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_i541_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n804));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i541_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5267_13 (.CI(n44800), .I0(n16242[10]), .I1(n895), .CO(n44801));
    SB_LUT4 add_5374_6_lut (.I0(GND_net), .I1(n17881[3]), .I2(n393), .I3(n44981), 
            .O(n17490[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5374_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_i459_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n682_adj_5177));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i459_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i208_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n308));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i208_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5267_12_lut (.I0(GND_net), .I1(n16242[9]), .I2(n822), 
            .I3(n44799), .O(n15630[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5267_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5267_12 (.CI(n44799), .I0(n16242[9]), .I1(n822), .CO(n44800));
    SB_CARRY add_5214_6 (.CI(n45077), .I0(n15306[3]), .I1(n378_adj_4967), 
            .CO(n45078));
    SB_CARRY add_5093_7 (.CI(n45135), .I0(n12905[4]), .I1(n442_adj_4943), 
            .CO(n45136));
    SB_CARRY add_5374_6 (.CI(n44981), .I0(n17881[3]), .I1(n393), .CO(n44982));
    SB_LUT4 add_5267_11_lut (.I0(GND_net), .I1(n16242[8]), .I2(n749), 
            .I3(n44798), .O(n15630[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5267_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_13_inv_0_i8_1_lut (.I0(IntegralLimit[7]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5402[7]));   // verilog/motorControl.v(48[22:36])
    defparam unary_minus_13_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_13_inv_0_i9_1_lut (.I0(IntegralLimit[8]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5402[8]));   // verilog/motorControl.v(48[22:36])
    defparam unary_minus_13_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_13_inv_0_i10_1_lut (.I0(IntegralLimit[9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5402[9]));   // verilog/motorControl.v(48[22:36])
    defparam unary_minus_13_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_DFFSR counter_2283__i0 (.Q(counter[0]), .C(clk16MHz), .D(n28[0]), 
            .R(counter_31__N_3995));   // verilog/motorControl.v(24[16:25])
    SB_LUT4 unary_minus_13_inv_0_i11_1_lut (.I0(IntegralLimit[10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5402[10]));   // verilog/motorControl.v(48[22:36])
    defparam unary_minus_13_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_5093_6_lut (.I0(GND_net), .I1(n12905[3]), .I2(n369_adj_4886), 
            .I3(n45134), .O(n11935[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5093_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5214_5_lut (.I0(GND_net), .I1(n15306[2]), .I2(n305), .I3(n45076), 
            .O(n14585[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5214_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_14_i18_3_lut (.I0(n130[17]), .I1(n182[17]), .I2(n181), 
            .I3(GND_net), .O(n207[17]));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_14_i18_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_15_i18_3_lut (.I0(n207[17]), .I1(IntegralLimit[17]), .I2(n155), 
            .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3996 [17]));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_15_i18_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_17_i83_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [16]), 
            .I2(GND_net), .I3(GND_net), .O(n122_adj_5141));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i83_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_13_inv_0_i12_1_lut (.I0(IntegralLimit[11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5402[11]));   // verilog/motorControl.v(48[22:36])
    defparam unary_minus_13_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_13_inv_0_i13_1_lut (.I0(IntegralLimit[12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5402[12]));   // verilog/motorControl.v(48[22:36])
    defparam unary_minus_13_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_13_inv_0_i14_1_lut (.I0(IntegralLimit[13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5402[13]));   // verilog/motorControl.v(48[22:36])
    defparam unary_minus_13_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_17_i75_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n110_adj_5185));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i75_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i28_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [13]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_5186));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i28_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i124_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n183_adj_5187));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i124_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i173_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n256));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i173_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i590_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n877));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i590_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5093_6 (.CI(n45134), .I0(n12905[3]), .I1(n369_adj_4886), 
            .CO(n45135));
    SB_LUT4 unary_minus_13_inv_0_i15_1_lut (.I0(IntegralLimit[14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5402[14]));   // verilog/motorControl.v(48[22:36])
    defparam unary_minus_13_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_17_i222_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n329));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i222_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5374_5_lut (.I0(GND_net), .I1(n17881[2]), .I2(n320), .I3(n44980), 
            .O(n17490[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5374_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_i36_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [17]), 
            .I2(GND_net), .I3(GND_net), .O(n53));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i36_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5214_5 (.CI(n45076), .I0(n15306[2]), .I1(n305), .CO(n45077));
    SB_LUT4 unary_minus_13_inv_0_i16_1_lut (.I0(IntegralLimit[15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5402[15]));   // verilog/motorControl.v(48[22:36])
    defparam unary_minus_13_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_5093_5_lut (.I0(GND_net), .I1(n12905[2]), .I2(n296_adj_4882), 
            .I3(n45133), .O(n11935[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5093_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i451_2_lut (.I0(\Kp[9] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n670_adj_5140));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i451_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5093_5 (.CI(n45133), .I0(n12905[2]), .I1(n296_adj_4882), 
            .CO(n45134));
    SB_LUT4 mult_16_i445_2_lut (.I0(\Kp[9] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n661_adj_5139));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i445_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5214_4_lut (.I0(GND_net), .I1(n15306[1]), .I2(n232), .I3(n45075), 
            .O(n14585[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5214_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_i132_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [16]), 
            .I2(GND_net), .I3(GND_net), .O(n195_adj_5138));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i132_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i749_2_lut (.I0(\Kp[15] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n1114_adj_5190));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i749_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i639_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n950));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i639_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_13_inv_0_i17_1_lut (.I0(IntegralLimit[16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5402[16]));   // verilog/motorControl.v(48[22:36])
    defparam unary_minus_13_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_17_i257_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n381));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i257_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i271_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n402_adj_5192));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i271_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i306_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n454_adj_5137));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i306_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i688_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n1023));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i688_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i500_2_lut (.I0(\Kp[10] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n743_adj_5136));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i500_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i355_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n527));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i355_2_lut.LUT_INIT = 16'h8888;
    SB_DFF \PID_CONTROLLER.integral_i0_i0  (.Q(\PID_CONTROLLER.integral [0]), 
           .C(clk16MHz), .D(n29381));   // verilog/motorControl.v(41[14] 61[8])
    SB_CARRY add_5267_11 (.CI(n44798), .I0(n16242[8]), .I1(n749), .CO(n44799));
    SB_LUT4 add_5267_10_lut (.I0(GND_net), .I1(n16242[7]), .I2(n676), 
            .I3(n44797), .O(n15630[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5267_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_14_i1_3_lut (.I0(n130[0]), .I1(n182[0]), .I2(n181), .I3(GND_net), 
            .O(n207[0]));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_14_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_5374_5 (.CI(n44980), .I0(n17881[2]), .I1(n320), .CO(n44981));
    SB_LUT4 mult_17_i320_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n475));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i320_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5267_10 (.CI(n44797), .I0(n16242[7]), .I1(n676), .CO(n44798));
    SB_LUT4 add_5267_9_lut (.I0(GND_net), .I1(n16242[6]), .I2(n603), .I3(n44796), 
            .O(n15630[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5267_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5093_4_lut (.I0(GND_net), .I1(n12905[1]), .I2(n223_adj_4867), 
            .I3(n45132), .O(n11935[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5093_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5214_4 (.CI(n45075), .I0(n15306[1]), .I1(n232), .CO(n45076));
    SB_LUT4 unary_minus_13_inv_0_i18_1_lut (.I0(IntegralLimit[17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5402[17]));   // verilog/motorControl.v(48[22:36])
    defparam unary_minus_13_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_5093_4 (.CI(n45132), .I0(n12905[1]), .I1(n223_adj_4867), 
            .CO(n45133));
    SB_CARRY add_5267_9 (.CI(n44796), .I0(n16242[6]), .I1(n603), .CO(n44797));
    SB_LUT4 add_5214_3_lut (.I0(GND_net), .I1(n15306[0]), .I2(n159), .I3(n45074), 
            .O(n14585[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5214_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_13_inv_0_i19_1_lut (.I0(IntegralLimit[18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5402[18]));   // verilog/motorControl.v(48[22:36])
    defparam unary_minus_13_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_5093_3_lut (.I0(GND_net), .I1(n12905[0]), .I2(n150_adj_4866), 
            .I3(n45131), .O(n11935[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5093_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_i737_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n1096));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i737_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i369_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n548));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i369_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_13_inv_0_i20_1_lut (.I0(IntegralLimit[19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5402[19]));   // verilog/motorControl.v(48[22:36])
    defparam unary_minus_13_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_16_i202_2_lut (.I0(\Kp[4] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n299_adj_5196));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i202_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_15_i1_3_lut (.I0(n207[0]), .I1(IntegralLimit[0]), .I2(n155), 
            .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3996 [0]));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_15_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_17_i2_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n306[0]));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i2_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_13_inv_0_i21_1_lut (.I0(IntegralLimit[20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5402[20]));   // verilog/motorControl.v(48[22:36])
    defparam unary_minus_13_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_16_i492_2_lut (.I0(\Kp[10] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n731_adj_5198));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i492_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i418_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n621));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i418_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i2_2_lut (.I0(\Kp[0] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n257[0]));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i2_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5267_8_lut (.I0(GND_net), .I1(n16242[5]), .I2(n530), .I3(n44795), 
            .O(n15630[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5267_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5214_3 (.CI(n45074), .I0(n15306[0]), .I1(n159), .CO(n45075));
    SB_LUT4 unary_minus_13_inv_0_i22_1_lut (.I0(IntegralLimit[21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5402[21]));   // verilog/motorControl.v(48[22:36])
    defparam unary_minus_13_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_17_i467_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n694));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i467_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_13_inv_0_i23_1_lut (.I0(IntegralLimit[22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5402[22]));   // verilog/motorControl.v(48[22:36])
    defparam unary_minus_13_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_13_inv_0_i24_1_lut (.I0(IntegralLimit[23]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5402[23]));   // verilog/motorControl.v(48[22:36])
    defparam unary_minus_13_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_17_i516_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n767));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i516_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i565_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n840));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i565_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i85_2_lut (.I0(\Kp[1] ), .I1(n1[17]), .I2(GND_net), 
            .I3(GND_net), .O(n125_adj_5200));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i85_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5374_4_lut (.I0(GND_net), .I1(n17881[1]), .I2(n247), .I3(n44979), 
            .O(n17490[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5374_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i38_2_lut (.I0(\Kp[0] ), .I1(n1[18]), .I2(GND_net), 
            .I3(GND_net), .O(n56_adj_5201));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i38_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5374_4 (.CI(n44979), .I0(n17881[1]), .I1(n247), .CO(n44980));
    SB_CARRY add_5267_8 (.CI(n44795), .I0(n16242[5]), .I1(n530), .CO(n44796));
    SB_LUT4 i23136_1_lut (.I0(n356[0]), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n37221));   // verilog/motorControl.v(50[18:38])
    defparam i23136_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_5267_7_lut (.I0(GND_net), .I1(n16242[4]), .I2(n457_adj_5202), 
            .I3(n44794), .O(n15630[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5267_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_20_inv_0_i1_1_lut (.I0(deadband[0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5403[0]));   // verilog/motorControl.v(51[43:52])
    defparam unary_minus_20_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_5267_7 (.CI(n44794), .I0(n16242[4]), .I1(n457_adj_5202), 
            .CO(n44795));
    SB_LUT4 unary_minus_26_inv_0_i22_1_lut (.I0(PWMLimit[21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5401[21]));   // verilog/motorControl.v(55[22:31])
    defparam unary_minus_26_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_26_inv_0_i23_1_lut (.I0(PWMLimit[22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5401[22]));   // verilog/motorControl.v(55[22:31])
    defparam unary_minus_26_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_16_i134_2_lut (.I0(\Kp[2] ), .I1(n1[17]), .I2(GND_net), 
            .I3(GND_net), .O(n198_adj_5206));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i134_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5267_6_lut (.I0(GND_net), .I1(n16242[3]), .I2(n384_adj_5207), 
            .I3(n44793), .O(n15630[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5267_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i251_2_lut (.I0(\Kp[5] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n372_adj_5208));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i251_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i183_2_lut (.I0(\Kp[3] ), .I1(n1[17]), .I2(GND_net), 
            .I3(GND_net), .O(n271));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i183_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_26_inv_0_i24_1_lut (.I0(PWMLimit[23]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5401[23]));   // verilog/motorControl.v(55[22:31])
    defparam unary_minus_26_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_5374_3_lut (.I0(GND_net), .I1(n17881[0]), .I2(n174), .I3(n44978), 
            .O(n17490[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5374_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i541_2_lut (.I0(\Kp[11] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n804_adj_5210));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i541_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5374_3 (.CI(n44978), .I0(n17881[0]), .I1(n174), .CO(n44979));
    SB_LUT4 unary_minus_20_inv_0_i2_1_lut (.I0(deadband[1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5403[1]));   // verilog/motorControl.v(51[43:52])
    defparam unary_minus_20_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_5093_3 (.CI(n45131), .I0(n12905[0]), .I1(n150_adj_4866), 
            .CO(n45132));
    SB_CARRY add_5267_6 (.CI(n44793), .I0(n16242[3]), .I1(n384_adj_5207), 
            .CO(n44794));
    SB_LUT4 add_5093_2_lut (.I0(GND_net), .I1(n8_adj_5212), .I2(n77_adj_5213), 
            .I3(GND_net), .O(n11935[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5093_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5374_2_lut (.I0(GND_net), .I1(n32), .I2(n101), .I3(GND_net), 
            .O(n17490[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5374_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i232_2_lut (.I0(\Kp[4] ), .I1(n1[17]), .I2(GND_net), 
            .I3(GND_net), .O(n344_adj_5214));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i232_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5214_2_lut (.I0(GND_net), .I1(n17_adj_5215), .I2(n86_adj_5216), 
            .I3(GND_net), .O(n14585[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5214_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5267_5_lut (.I0(GND_net), .I1(n16242[2]), .I2(n311_adj_5217), 
            .I3(n44792), .O(n15630[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5267_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5214_2 (.CI(GND_net), .I0(n17_adj_5215), .I1(n86_adj_5216), 
            .CO(n45074));
    SB_CARRY add_5267_5 (.CI(n44792), .I0(n16242[2]), .I1(n311_adj_5217), 
            .CO(n44793));
    SB_CARRY add_5374_2 (.CI(GND_net), .I0(n32), .I1(n101), .CO(n44978));
    SB_LUT4 add_5400_14_lut (.I0(GND_net), .I1(n18218[11]), .I2(n980), 
            .I3(n44977), .O(n17881[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5400_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5267_4_lut (.I0(GND_net), .I1(n16242[1]), .I2(n238), .I3(n44791), 
            .O(n15630[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5267_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5093_2 (.CI(GND_net), .I0(n8_adj_5212), .I1(n77_adj_5213), 
            .CO(n45131));
    SB_CARRY add_5267_4 (.CI(n44791), .I0(n16242[1]), .I1(n238), .CO(n44792));
    SB_LUT4 add_5267_3_lut (.I0(GND_net), .I1(n16242[0]), .I2(n165_adj_5218), 
            .I3(n44790), .O(n15630[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5267_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5136_22_lut (.I0(GND_net), .I1(n13786[19]), .I2(GND_net), 
            .I3(n45130), .O(n12905[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5136_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5475_10_lut (.I0(GND_net), .I1(n19026[7]), .I2(n700_adj_5219), 
            .I3(n45073), .O(n18846[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5475_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5400_13_lut (.I0(GND_net), .I1(n18218[10]), .I2(n907), 
            .I3(n44976), .O(n17881[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5400_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5267_3 (.CI(n44790), .I0(n16242[0]), .I1(n165_adj_5218), 
            .CO(n44791));
    SB_CARRY add_5400_13 (.CI(n44976), .I0(n18218[10]), .I1(n907), .CO(n44977));
    SB_LUT4 add_5400_12_lut (.I0(GND_net), .I1(n18218[9]), .I2(n834), 
            .I3(n44975), .O(n17881[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5400_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_20_inv_0_i3_1_lut (.I0(deadband[2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5403[2]));   // verilog/motorControl.v(51[43:52])
    defparam unary_minus_20_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_17_i508_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n755_adj_5221));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i508_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5267_2_lut (.I0(GND_net), .I1(n23_adj_5222), .I2(n92_adj_5223), 
            .I3(GND_net), .O(n15630[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5267_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5475_9_lut (.I0(GND_net), .I1(n19026[6]), .I2(n627_adj_5224), 
            .I3(n45072), .O(n18846[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5475_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_i183_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [17]), 
            .I2(GND_net), .I3(GND_net), .O(n271_adj_5225));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i183_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5267_2 (.CI(GND_net), .I0(n23_adj_5222), .I1(n92_adj_5223), 
            .CO(n44790));
    SB_LUT4 add_5300_17_lut (.I0(GND_net), .I1(n16786[14]), .I2(GND_net), 
            .I3(n44789), .O(n16242[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5300_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_i557_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n828_adj_5226));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i557_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5300_16_lut (.I0(GND_net), .I1(n16786[13]), .I2(n1117_adj_5227), 
            .I3(n44788), .O(n16242[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5300_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5136_21_lut (.I0(GND_net), .I1(n13786[18]), .I2(GND_net), 
            .I3(n45129), .O(n12905[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5136_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_add_1225_24_lut (.I0(n1[23]), .I1(n11935[21]), .I2(GND_net), 
            .I3(n45173), .O(n11428[0])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_16_add_1225_24_lut.LUT_INIT = 16'h6996;
    SB_CARRY add_5475_9 (.CI(n45072), .I0(n19026[6]), .I1(n627_adj_5224), 
            .CO(n45073));
    SB_CARRY add_5300_16 (.CI(n44788), .I0(n16786[13]), .I1(n1117_adj_5227), 
            .CO(n44789));
    SB_LUT4 unary_minus_20_inv_0_i4_1_lut (.I0(deadband[3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5403[3]));   // verilog/motorControl.v(51[43:52])
    defparam unary_minus_20_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_5300_15_lut (.I0(GND_net), .I1(n16786[12]), .I2(n1044_adj_5229), 
            .I3(n44787), .O(n16242[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5300_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5400_12 (.CI(n44975), .I0(n18218[9]), .I1(n834), .CO(n44976));
    SB_LUT4 unary_minus_20_inv_0_i5_1_lut (.I0(deadband[4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5403[4]));   // verilog/motorControl.v(51[43:52])
    defparam unary_minus_20_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_5300_15 (.CI(n44787), .I0(n16786[12]), .I1(n1044_adj_5229), 
            .CO(n44788));
    SB_CARRY add_5136_21 (.CI(n45129), .I0(n13786[18]), .I1(GND_net), 
            .CO(n45130));
    SB_LUT4 add_5400_11_lut (.I0(GND_net), .I1(n18218[8]), .I2(n761), 
            .I3(n44974), .O(n17881[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5400_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5300_14_lut (.I0(GND_net), .I1(n16786[11]), .I2(n971_adj_5231), 
            .I3(n44786), .O(n16242[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5300_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5300_14 (.CI(n44786), .I0(n16786[11]), .I1(n971_adj_5231), 
            .CO(n44787));
    SB_LUT4 add_5475_8_lut (.I0(GND_net), .I1(n19026[5]), .I2(n554_adj_5232), 
            .I3(n45071), .O(n18846[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5475_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5400_11 (.CI(n44974), .I0(n18218[8]), .I1(n761), .CO(n44975));
    SB_LUT4 add_5300_13_lut (.I0(GND_net), .I1(n16786[10]), .I2(n898_adj_5233), 
            .I3(n44785), .O(n16242[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5300_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_20_inv_0_i6_1_lut (.I0(deadband[5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5403[5]));   // verilog/motorControl.v(51[43:52])
    defparam unary_minus_20_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_5300_13 (.CI(n44785), .I0(n16786[10]), .I1(n898_adj_5233), 
            .CO(n44786));
    SB_LUT4 add_5400_10_lut (.I0(GND_net), .I1(n18218[7]), .I2(n688), 
            .I3(n44973), .O(n17881[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5400_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5400_10 (.CI(n44973), .I0(n18218[7]), .I1(n688), .CO(n44974));
    SB_LUT4 add_5300_12_lut (.I0(GND_net), .I1(n16786[9]), .I2(n825_adj_5235), 
            .I3(n44784), .O(n16242[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5300_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5300_12 (.CI(n44784), .I0(n16786[9]), .I1(n825_adj_5235), 
            .CO(n44785));
    SB_CARRY add_5475_8 (.CI(n45071), .I0(n19026[5]), .I1(n554_adj_5232), 
            .CO(n45072));
    SB_LUT4 add_5400_9_lut (.I0(GND_net), .I1(n18218[6]), .I2(n615), .I3(n44972), 
            .O(n17881[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5400_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5300_11_lut (.I0(GND_net), .I1(n16786[8]), .I2(n752_adj_5236), 
            .I3(n44783), .O(n16242[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5300_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5300_11 (.CI(n44783), .I0(n16786[8]), .I1(n752_adj_5236), 
            .CO(n44784));
    SB_LUT4 mult_16_i281_2_lut (.I0(\Kp[5] ), .I1(n1[17]), .I2(GND_net), 
            .I3(GND_net), .O(n417));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i281_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut_adj_1682 (.I0(n19450[2]), .I1(n6_adj_5237), .I2(\Kp[4] ), 
            .I3(n1[18]), .O(n19401[3]));   // verilog/motorControl.v(50[18:24])
    defparam i1_4_lut_adj_1682.LUT_INIT = 16'h9666;
    SB_LUT4 mult_16_i138_2_lut (.I0(\Kp[2] ), .I1(n1[19]), .I2(GND_net), 
            .I3(GND_net), .O(n204));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i138_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5300_10_lut (.I0(GND_net), .I1(n16786[7]), .I2(n679_adj_5238), 
            .I3(n44782), .O(n16242[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5300_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5300_10 (.CI(n44782), .I0(n16786[7]), .I1(n679_adj_5238), 
            .CO(n44783));
    SB_LUT4 add_5300_9_lut (.I0(GND_net), .I1(n16786[6]), .I2(n606_adj_5239), 
            .I3(n44781), .O(n16242[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5300_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i29216_4_lut (.I0(\Kp[0] ), .I1(\Kp[1] ), .I2(n1[22]), .I3(n1[21]), 
            .O(n19498[0]));   // verilog/motorControl.v(50[18:24])
    defparam i29216_4_lut.LUT_INIT = 16'h6ca0;
    SB_LUT4 add_5475_7_lut (.I0(GND_net), .I1(n19026[4]), .I2(n481_adj_5240), 
            .I3(n45070), .O(n18846[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5475_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5300_9 (.CI(n44781), .I0(n16786[6]), .I1(n606_adj_5239), 
            .CO(n44782));
    SB_CARRY add_5400_9 (.CI(n44972), .I0(n18218[6]), .I1(n615), .CO(n44973));
    SB_LUT4 add_5300_8_lut (.I0(GND_net), .I1(n16786[5]), .I2(n533_adj_5241), 
            .I3(n44780), .O(n16242[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5300_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5300_8 (.CI(n44780), .I0(n16786[5]), .I1(n533_adj_5241), 
            .CO(n44781));
    SB_LUT4 add_5400_8_lut (.I0(GND_net), .I1(n18218[5]), .I2(n542), .I3(n44971), 
            .O(n17881[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5400_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5300_7_lut (.I0(GND_net), .I1(n16786[4]), .I2(n460_adj_5242), 
            .I3(n44779), .O(n16242[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5300_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5136_20_lut (.I0(GND_net), .I1(n13786[17]), .I2(GND_net), 
            .I3(n45128), .O(n12905[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5136_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5300_7 (.CI(n44779), .I0(n16786[4]), .I1(n460_adj_5242), 
            .CO(n44780));
    SB_LUT4 add_5300_6_lut (.I0(GND_net), .I1(n16786[3]), .I2(n387_adj_5243), 
            .I3(n44778), .O(n16242[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5300_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5136_20 (.CI(n45128), .I0(n13786[17]), .I1(GND_net), 
            .CO(n45129));
    SB_CARRY add_5475_7 (.CI(n45070), .I0(n19026[4]), .I1(n481_adj_5240), 
            .CO(n45071));
    SB_CARRY add_5400_8 (.CI(n44971), .I0(n18218[5]), .I1(n542), .CO(n44972));
    SB_LUT4 add_5400_7_lut (.I0(GND_net), .I1(n18218[4]), .I2(n469), .I3(n44970), 
            .O(n17881[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5400_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5300_6 (.CI(n44778), .I0(n16786[3]), .I1(n387_adj_5243), 
            .CO(n44779));
    SB_LUT4 add_5300_5_lut (.I0(GND_net), .I1(n16786[2]), .I2(n314_adj_5244), 
            .I3(n44777), .O(n16242[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5300_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5300_5 (.CI(n44777), .I0(n16786[2]), .I1(n314_adj_5244), 
            .CO(n44778));
    SB_LUT4 mult_16_add_1225_23_lut (.I0(GND_net), .I1(n11935[20]), .I2(GND_net), 
            .I3(n45172), .O(n257[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_16_add_1225_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5400_7 (.CI(n44970), .I0(n18218[4]), .I1(n469), .CO(n44971));
    SB_CARRY mult_16_add_1225_23 (.CI(n45172), .I0(n11935[20]), .I1(GND_net), 
            .CO(n45173));
    SB_LUT4 add_5300_4_lut (.I0(GND_net), .I1(n16786[1]), .I2(n241_adj_5245), 
            .I3(n44776), .O(n16242[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5300_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i89_2_lut (.I0(\Kp[1] ), .I1(n1[19]), .I2(GND_net), 
            .I3(GND_net), .O(n131_adj_5246));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i89_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i42_2_lut (.I0(\Kp[0] ), .I1(n1[20]), .I2(GND_net), 
            .I3(GND_net), .O(n62));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i42_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5136_19_lut (.I0(GND_net), .I1(n13786[16]), .I2(GND_net), 
            .I3(n45127), .O(n12905[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5136_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5475_6_lut (.I0(GND_net), .I1(n19026[3]), .I2(n408_adj_5247), 
            .I3(n45069), .O(n18846[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5475_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5136_19 (.CI(n45127), .I0(n13786[16]), .I1(GND_net), 
            .CO(n45128));
    SB_CARRY add_5475_6 (.CI(n45069), .I0(n19026[3]), .I1(n408_adj_5247), 
            .CO(n45070));
    SB_LUT4 mult_16_add_1225_22_lut (.I0(GND_net), .I1(n11935[19]), .I2(GND_net), 
            .I3(n45171), .O(n257[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_16_add_1225_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5475_5_lut (.I0(GND_net), .I1(n19026[2]), .I2(n335_adj_5248), 
            .I3(n45068), .O(n18846[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5475_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5400_6_lut (.I0(GND_net), .I1(n18218[3]), .I2(n396_adj_5249), 
            .I3(n44969), .O(n17881[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5400_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5400_6 (.CI(n44969), .I0(n18218[3]), .I1(n396_adj_5249), 
            .CO(n44970));
    SB_CARRY add_5300_4 (.CI(n44776), .I0(n16786[1]), .I1(n241_adj_5245), 
            .CO(n44777));
    SB_LUT4 add_5300_3_lut (.I0(GND_net), .I1(n16786[0]), .I2(n168_adj_5250), 
            .I3(n44775), .O(n16242[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5300_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5300_3 (.CI(n44775), .I0(n16786[0]), .I1(n168_adj_5250), 
            .CO(n44776));
    SB_CARRY add_5475_5 (.CI(n45068), .I0(n19026[2]), .I1(n335_adj_5248), 
            .CO(n45069));
    SB_LUT4 add_5400_5_lut (.I0(GND_net), .I1(n18218[2]), .I2(n323), .I3(n44968), 
            .O(n17881[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5400_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5300_2_lut (.I0(GND_net), .I1(n26_adj_5251), .I2(n95_adj_5252), 
            .I3(GND_net), .O(n16242[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5300_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5400_5 (.CI(n44968), .I0(n18218[2]), .I1(n323), .CO(n44969));
    SB_CARRY add_5300_2 (.CI(GND_net), .I0(n26_adj_5251), .I1(n95_adj_5252), 
            .CO(n44775));
    SB_LUT4 add_5500_9_lut (.I0(GND_net), .I1(n19233[6]), .I2(n630_adj_5253), 
            .I3(n44774), .O(n19106[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5500_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5400_4_lut (.I0(GND_net), .I1(n18218[1]), .I2(n250), .I3(n44967), 
            .O(n17881[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5400_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5475_4_lut (.I0(GND_net), .I1(n19026[1]), .I2(n262_adj_5254), 
            .I3(n45067), .O(n18846[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5475_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5500_8_lut (.I0(GND_net), .I1(n19233[5]), .I2(n557_adj_5255), 
            .I3(n44773), .O(n19106[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5500_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5500_8 (.CI(n44773), .I0(n19233[5]), .I1(n557_adj_5255), 
            .CO(n44774));
    SB_LUT4 add_5500_7_lut (.I0(GND_net), .I1(n19233[4]), .I2(n484_adj_5256), 
            .I3(n44772), .O(n19106[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5500_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5500_7 (.CI(n44772), .I0(n19233[4]), .I1(n484_adj_5256), 
            .CO(n44773));
    SB_CARRY add_5400_4 (.CI(n44967), .I0(n18218[1]), .I1(n250), .CO(n44968));
    SB_CARRY mult_16_add_1225_22 (.CI(n45171), .I0(n11935[19]), .I1(GND_net), 
            .CO(n45172));
    SB_LUT4 add_5136_18_lut (.I0(GND_net), .I1(n13786[15]), .I2(GND_net), 
            .I3(n45126), .O(n12905[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5136_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5400_3_lut (.I0(GND_net), .I1(n18218[0]), .I2(n177), .I3(n44966), 
            .O(n17881[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5400_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5475_4 (.CI(n45067), .I0(n19026[1]), .I1(n262_adj_5254), 
            .CO(n45068));
    SB_LUT4 add_5500_6_lut (.I0(GND_net), .I1(n19233[3]), .I2(n411_adj_5257), 
            .I3(n44771), .O(n19106[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5500_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5400_3 (.CI(n44966), .I0(n18218[0]), .I1(n177), .CO(n44967));
    SB_CARRY add_5500_6 (.CI(n44771), .I0(n19233[3]), .I1(n411_adj_5257), 
            .CO(n44772));
    SB_LUT4 add_5500_5_lut (.I0(GND_net), .I1(n19233[2]), .I2(n338_adj_5258), 
            .I3(n44770), .O(n19106[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5500_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5500_5 (.CI(n44770), .I0(n19233[2]), .I1(n338_adj_5258), 
            .CO(n44771));
    SB_LUT4 add_5500_4_lut (.I0(GND_net), .I1(n19233[1]), .I2(n265_adj_5259), 
            .I3(n44769), .O(n19106[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5500_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5500_4 (.CI(n44769), .I0(n19233[1]), .I1(n265_adj_5259), 
            .CO(n44770));
    SB_LUT4 add_5400_2_lut (.I0(GND_net), .I1(n35_adj_5260), .I2(n104), 
            .I3(GND_net), .O(n17881[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5400_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i330_2_lut (.I0(\Kp[6] ), .I1(n1[17]), .I2(GND_net), 
            .I3(GND_net), .O(n490));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i330_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut_adj_1683 (.I0(\Kp[4] ), .I1(\Kp[5] ), .I2(n1[19]), 
            .I3(n1[18]), .O(n52332));   // verilog/motorControl.v(50[18:24])
    defparam i1_4_lut_adj_1683.LUT_INIT = 16'h6ca0;
    SB_LUT4 i1_3_lut (.I0(\Kp[3] ), .I1(n52332), .I2(n1[20]), .I3(GND_net), 
            .O(n52334));   // verilog/motorControl.v(50[18:24])
    defparam i1_3_lut.LUT_INIT = 16'h6c6c;
    SB_LUT4 add_5475_3_lut (.I0(GND_net), .I1(n19026[0]), .I2(n189_adj_5261), 
            .I3(n45066), .O(n18846[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5475_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5500_3_lut (.I0(GND_net), .I1(n19233[0]), .I2(n192_adj_5262), 
            .I3(n44768), .O(n19106[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5500_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5400_2 (.CI(GND_net), .I0(n35_adj_5260), .I1(n104), .CO(n44966));
    SB_CARRY add_5500_3 (.CI(n44768), .I0(n19233[0]), .I1(n192_adj_5262), 
            .CO(n44769));
    SB_LUT4 add_5500_2_lut (.I0(GND_net), .I1(n50_adj_5263), .I2(n119_adj_5264), 
            .I3(GND_net), .O(n19106[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5500_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5500_2 (.CI(GND_net), .I0(n50_adj_5263), .I1(n119_adj_5264), 
            .CO(n44768));
    SB_CARRY add_5475_3 (.CI(n45066), .I0(n19026[0]), .I1(n189_adj_5261), 
            .CO(n45067));
    SB_LUT4 mult_16_i142_2_lut (.I0(\Kp[2] ), .I1(n1[21]), .I2(GND_net), 
            .I3(GND_net), .O(n210));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i142_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5520_7_lut (.I0(GND_net), .I1(n51074), .I2(n490_adj_5265), 
            .I3(n44965), .O(n19282[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5520_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5331_16_lut (.I0(GND_net), .I1(n17266[13]), .I2(n1120_adj_5266), 
            .I3(n44767), .O(n16786[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5331_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5475_2_lut (.I0(GND_net), .I1(n47_adj_5267), .I2(n116_adj_5268), 
            .I3(GND_net), .O(n18846[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5475_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5520_6_lut (.I0(GND_net), .I1(n19366[3]), .I2(n417_adj_5269), 
            .I3(n44964), .O(n19282[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5520_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5331_15_lut (.I0(GND_net), .I1(n17266[12]), .I2(n1047_adj_5270), 
            .I3(n44766), .O(n16786[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5331_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5475_2 (.CI(GND_net), .I0(n47_adj_5267), .I1(n116_adj_5268), 
            .CO(n45066));
    SB_LUT4 i1_4_lut_adj_1684 (.I0(\Kp[1] ), .I1(n210), .I2(n1[22]), .I3(n52334), 
            .O(n52338));   // verilog/motorControl.v(50[18:24])
    defparam i1_4_lut_adj_1684.LUT_INIT = 16'h936c;
    SB_CARRY add_5331_15 (.CI(n44766), .I0(n17266[12]), .I1(n1047_adj_5270), 
            .CO(n44767));
    SB_CARRY add_5520_6 (.CI(n44964), .I0(n19366[3]), .I1(n417_adj_5269), 
            .CO(n44965));
    SB_LUT4 add_5331_14_lut (.I0(GND_net), .I1(n17266[11]), .I2(n974_adj_5271), 
            .I3(n44765), .O(n16786[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5331_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5331_14 (.CI(n44765), .I0(n17266[11]), .I1(n974_adj_5271), 
            .CO(n44766));
    SB_LUT4 add_5520_5_lut (.I0(GND_net), .I1(n19366[2]), .I2(n344_adj_5272), 
            .I3(n44963), .O(n19282[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5520_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5331_13_lut (.I0(GND_net), .I1(n17266[10]), .I2(n901_adj_5273), 
            .I3(n44764), .O(n16786[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5331_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5331_13 (.CI(n44764), .I0(n17266[10]), .I1(n901_adj_5273), 
            .CO(n44765));
    SB_LUT4 i29218_4_lut (.I0(\Kp[0] ), .I1(\Kp[1] ), .I2(n1[22]), .I3(n1[21]), 
            .O(n43305));   // verilog/motorControl.v(50[18:24])
    defparam i29218_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 add_5331_12_lut (.I0(GND_net), .I1(n17266[9]), .I2(n828_adj_5226), 
            .I3(n44763), .O(n16786[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5331_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5520_5 (.CI(n44963), .I0(n19366[2]), .I1(n344_adj_5272), 
            .CO(n44964));
    SB_CARRY add_5331_12 (.CI(n44763), .I0(n17266[9]), .I1(n828_adj_5226), 
            .CO(n44764));
    SB_LUT4 i1_4_lut_adj_1685 (.I0(n43305), .I1(\Kp[0] ), .I2(n52338), 
            .I3(n1[23]), .O(n52342));   // verilog/motorControl.v(50[18:24])
    defparam i1_4_lut_adj_1685.LUT_INIT = 16'h695a;
    SB_LUT4 mult_17_i606_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n901_adj_5273));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i606_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5520_4_lut (.I0(GND_net), .I1(n19366[1]), .I2(n271_adj_5225), 
            .I3(n44962), .O(n19282[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5520_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5331_11_lut (.I0(GND_net), .I1(n17266[8]), .I2(n755_adj_5221), 
            .I3(n44762), .O(n16786[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5331_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_26_add_3_25_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5401[23]), 
            .I3(n43878), .O(n436[23])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_26_add_3_24_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5401[22]), 
            .I3(n43877), .O(n436[22])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_26_add_3_24 (.CI(n43877), .I0(GND_net), .I1(n1_adj_5401[22]), 
            .CO(n43878));
    SB_LUT4 unary_minus_26_add_3_23_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5401[21]), 
            .I3(n43876), .O(n436[21])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5331_11 (.CI(n44762), .I0(n17266[8]), .I1(n755_adj_5221), 
            .CO(n44763));
    SB_CARRY unary_minus_26_add_3_23 (.CI(n43876), .I0(GND_net), .I1(n1_adj_5401[21]), 
            .CO(n43877));
    SB_LUT4 mult_17_i232_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [17]), 
            .I2(GND_net), .I3(GND_net), .O(n344_adj_5272));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i232_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5331_10_lut (.I0(GND_net), .I1(n17266[7]), .I2(n682_adj_5177), 
            .I3(n44761), .O(n16786[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5331_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i29420_4_lut (.I0(n19450[2]), .I1(\Kp[4] ), .I2(n6_adj_5237), 
            .I3(n1[18]), .O(n8_adj_5274));   // verilog/motorControl.v(50[18:24])
    defparam i29420_4_lut.LUT_INIT = 16'he8a0;
    SB_CARRY add_5136_18 (.CI(n45126), .I0(n13786[15]), .I1(GND_net), 
            .CO(n45127));
    SB_LUT4 add_5250_19_lut (.I0(GND_net), .I1(n15953[16]), .I2(GND_net), 
            .I3(n45065), .O(n15306[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5250_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_26_add_3_22_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5401[20]), 
            .I3(n43875), .O(n436[20])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5250_18_lut (.I0(GND_net), .I1(n15953[15]), .I2(GND_net), 
            .I3(n45064), .O(n15306[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5250_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_26_add_3_22 (.CI(n43875), .I0(GND_net), .I1(n1_adj_5401[20]), 
            .CO(n43876));
    SB_CARRY add_5520_4 (.CI(n44962), .I0(n19366[1]), .I1(n271_adj_5225), 
            .CO(n44963));
    SB_LUT4 unary_minus_26_add_3_21_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5401[19]), 
            .I3(n43874), .O(n436[19])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5331_10 (.CI(n44761), .I0(n17266[7]), .I1(n682_adj_5177), 
            .CO(n44762));
    SB_LUT4 add_5520_3_lut (.I0(GND_net), .I1(n19366[0]), .I2(n198_adj_5118), 
            .I3(n44961), .O(n19282[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5520_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5331_9_lut (.I0(GND_net), .I1(n17266[6]), .I2(n609_adj_5117), 
            .I3(n44760), .O(n16786[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5331_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5331_9 (.CI(n44760), .I0(n17266[6]), .I1(n609_adj_5117), 
            .CO(n44761));
    SB_LUT4 i1_4_lut_adj_1686 (.I0(n6_adj_5275), .I1(n8_adj_5274), .I2(n4_adj_5276), 
            .I3(n52342), .O(n50980));   // verilog/motorControl.v(50[18:24])
    defparam i1_4_lut_adj_1686.LUT_INIT = 16'h6996;
    SB_CARRY add_5520_3 (.CI(n44961), .I0(n19366[0]), .I1(n198_adj_5118), 
            .CO(n44962));
    SB_CARRY unary_minus_26_add_3_21 (.CI(n43874), .I0(GND_net), .I1(n1_adj_5401[19]), 
            .CO(n43875));
    SB_LUT4 add_5520_2_lut (.I0(GND_net), .I1(n56), .I2(n125_adj_5010), 
            .I3(GND_net), .O(n19282[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5520_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5520_2 (.CI(GND_net), .I0(n56), .I1(n125_adj_5010), .CO(n44961));
    SB_LUT4 add_5331_8_lut (.I0(GND_net), .I1(n17266[5]), .I2(n536), .I3(n44759), 
            .O(n16786[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5331_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_26_add_3_20_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5401[18]), 
            .I3(n43873), .O(n436[18])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5331_8 (.CI(n44759), .I0(n17266[5]), .I1(n536), .CO(n44760));
    SB_CARRY unary_minus_26_add_3_20 (.CI(n43873), .I0(GND_net), .I1(n1_adj_5401[18]), 
            .CO(n43874));
    SB_LUT4 mult_17_i655_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n974_adj_5271));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i655_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_26_add_3_19_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5401[17]), 
            .I3(n43872), .O(n436[17])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_26_add_3_19 (.CI(n43872), .I0(GND_net), .I1(n1_adj_5401[17]), 
            .CO(n43873));
    SB_LUT4 add_5424_13_lut (.I0(GND_net), .I1(n18505[10]), .I2(n910), 
            .I3(n44960), .O(n18218[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5424_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5331_7_lut (.I0(GND_net), .I1(n17266[4]), .I2(n463), .I3(n44758), 
            .O(n16786[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5331_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_26_add_3_18_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5401[16]), 
            .I3(n43871), .O(n436[16])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_26_add_3_18 (.CI(n43871), .I0(GND_net), .I1(n1_adj_5401[16]), 
            .CO(n43872));
    SB_LUT4 unary_minus_26_add_3_17_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5401[15]), 
            .I3(n43870), .O(n436[15])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5331_7 (.CI(n44758), .I0(n17266[4]), .I1(n463), .CO(n44759));
    SB_CARRY unary_minus_26_add_3_17 (.CI(n43870), .I0(GND_net), .I1(n1_adj_5401[15]), 
            .CO(n43871));
    SB_LUT4 add_5331_6_lut (.I0(GND_net), .I1(n17266[3]), .I2(n390), .I3(n44757), 
            .O(n16786[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5331_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5331_6 (.CI(n44757), .I0(n17266[3]), .I1(n390), .CO(n44758));
    SB_LUT4 unary_minus_26_add_3_16_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5401[14]), 
            .I3(n43869), .O(n436[14])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_26_add_3_16 (.CI(n43869), .I0(GND_net), .I1(n1_adj_5401[14]), 
            .CO(n43870));
    SB_LUT4 unary_minus_26_add_3_15_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5401[13]), 
            .I3(n43868), .O(n436[13])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5424_12_lut (.I0(GND_net), .I1(n18505[9]), .I2(n837), 
            .I3(n44959), .O(n18218[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5424_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5331_5_lut (.I0(GND_net), .I1(n17266[2]), .I2(n317), .I3(n44756), 
            .O(n16786[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5331_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5331_5 (.CI(n44756), .I0(n17266[2]), .I1(n317), .CO(n44757));
    SB_CARRY unary_minus_26_add_3_15 (.CI(n43868), .I0(GND_net), .I1(n1_adj_5401[13]), 
            .CO(n43869));
    SB_LUT4 add_5331_4_lut (.I0(GND_net), .I1(n17266[1]), .I2(n244), .I3(n44755), 
            .O(n16786[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5331_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5331_4 (.CI(n44755), .I0(n17266[1]), .I1(n244), .CO(n44756));
    SB_LUT4 add_5331_3_lut (.I0(GND_net), .I1(n17266[0]), .I2(n171), .I3(n44754), 
            .O(n16786[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5331_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_26_add_3_14_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5401[12]), 
            .I3(n43867), .O(n436[12])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5250_18 (.CI(n45064), .I0(n15953[15]), .I1(GND_net), 
            .CO(n45065));
    SB_CARRY add_5424_12 (.CI(n44959), .I0(n18505[9]), .I1(n837), .CO(n44960));
    SB_LUT4 mux_14_i13_3_lut (.I0(n130[12]), .I1(n182[12]), .I2(n181), 
            .I3(GND_net), .O(n207[12]));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_14_i13_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_5250_17_lut (.I0(GND_net), .I1(n15953[14]), .I2(GND_net), 
            .I3(n45063), .O(n15306[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5250_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5331_3 (.CI(n44754), .I0(n17266[0]), .I1(n171), .CO(n44755));
    SB_CARRY add_5250_17 (.CI(n45063), .I0(n15953[14]), .I1(GND_net), 
            .CO(n45064));
    SB_LUT4 add_5424_11_lut (.I0(GND_net), .I1(n18505[8]), .I2(n764), 
            .I3(n44958), .O(n18218[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5424_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_26_add_3_14 (.CI(n43867), .I0(GND_net), .I1(n1_adj_5401[12]), 
            .CO(n43868));
    SB_LUT4 unary_minus_26_add_3_13_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5401[11]), 
            .I3(n43866), .O(n436[11])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5424_11 (.CI(n44958), .I0(n18505[8]), .I1(n764), .CO(n44959));
    SB_LUT4 add_5331_2_lut (.I0(GND_net), .I1(n29), .I2(n98), .I3(GND_net), 
            .O(n16786[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5331_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_15_i13_3_lut (.I0(n207[12]), .I1(IntegralLimit[12]), .I2(n155), 
            .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3996 [12]));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_15_i13_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_5331_2 (.CI(GND_net), .I0(n29), .I1(n98), .CO(n44754));
    SB_LUT4 add_5360_15_lut (.I0(GND_net), .I1(n17686[12]), .I2(n1050), 
            .I3(n44753), .O(n17266[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5360_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5360_14_lut (.I0(GND_net), .I1(n17686[11]), .I2(n977), 
            .I3(n44752), .O(n17266[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5360_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5424_10_lut (.I0(GND_net), .I1(n18505[7]), .I2(n691), 
            .I3(n44957), .O(n18218[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5424_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_i73_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n107_adj_5277));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i73_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY unary_minus_26_add_3_13 (.CI(n43866), .I0(GND_net), .I1(n1_adj_5401[11]), 
            .CO(n43867));
    SB_LUT4 mult_16_add_1225_21_lut (.I0(GND_net), .I1(n11935[18]), .I2(GND_net), 
            .I3(n45170), .O(n257[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_16_add_1225_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5360_14 (.CI(n44752), .I0(n17686[11]), .I1(n977), .CO(n44753));
    SB_CARRY add_5424_10 (.CI(n44957), .I0(n18505[7]), .I1(n691), .CO(n44958));
    SB_CARRY mult_16_add_1225_21 (.CI(n45170), .I0(n11935[18]), .I1(GND_net), 
            .CO(n45171));
    SB_LUT4 mult_17_i26_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n38));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i26_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5136_17_lut (.I0(GND_net), .I1(n13786[14]), .I2(GND_net), 
            .I3(n45125), .O(n12905[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5136_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_26_add_3_12_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5401[10]), 
            .I3(n43865), .O(n436[10])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5360_13_lut (.I0(GND_net), .I1(n17686[10]), .I2(n904), 
            .I3(n44751), .O(n17266[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5360_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5250_16_lut (.I0(GND_net), .I1(n15953[13]), .I2(n1111), 
            .I3(n45062), .O(n15306[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5250_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5360_13 (.CI(n44751), .I0(n17686[10]), .I1(n904), .CO(n44752));
    SB_LUT4 add_5424_9_lut (.I0(GND_net), .I1(n18505[6]), .I2(n618), .I3(n44956), 
            .O(n18218[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5424_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5360_12_lut (.I0(GND_net), .I1(n17686[9]), .I2(n831), 
            .I3(n44750), .O(n17266[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5360_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_26_add_3_12 (.CI(n43865), .I0(GND_net), .I1(n1_adj_5401[10]), 
            .CO(n43866));
    SB_LUT4 unary_minus_26_add_3_11_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5401[9]), 
            .I3(n43864), .O(n436[9])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_26_add_3_11 (.CI(n43864), .I0(GND_net), .I1(n1_adj_5401[9]), 
            .CO(n43865));
    SB_LUT4 unary_minus_26_add_3_10_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5401[8]), 
            .I3(n43863), .O(n436[8])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_26_add_3_10 (.CI(n43863), .I0(GND_net), .I1(n1_adj_5401[8]), 
            .CO(n43864));
    SB_CARRY add_5136_17 (.CI(n45125), .I0(n13786[14]), .I1(GND_net), 
            .CO(n45126));
    SB_CARRY add_5360_12 (.CI(n44750), .I0(n17686[9]), .I1(n831), .CO(n44751));
    SB_LUT4 add_5360_11_lut (.I0(GND_net), .I1(n17686[8]), .I2(n758), 
            .I3(n44749), .O(n17266[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5360_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5250_16 (.CI(n45062), .I0(n15953[13]), .I1(n1111), .CO(n45063));
    SB_CARRY add_5360_11 (.CI(n44749), .I0(n17686[8]), .I1(n758), .CO(n44750));
    SB_LUT4 add_5360_10_lut (.I0(GND_net), .I1(n17686[7]), .I2(n685), 
            .I3(n44748), .O(n17266[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5360_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_26_add_3_9_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5401[7]), 
            .I3(n43862), .O(n436[7])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_26_add_3_9 (.CI(n43862), .I0(GND_net), .I1(n1_adj_5401[7]), 
            .CO(n43863));
    SB_CARRY add_5360_10 (.CI(n44748), .I0(n17686[7]), .I1(n685), .CO(n44749));
    SB_LUT4 unary_minus_26_add_3_8_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5401[6]), 
            .I3(n43861), .O(n436[6])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_i122_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n180));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i122_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_20_inv_0_i7_1_lut (.I0(deadband[6]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5403[6]));   // verilog/motorControl.v(51[43:52])
    defparam unary_minus_20_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_16_i61_2_lut (.I0(\Kp[1] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n89_adj_5279));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i61_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY unary_minus_26_add_3_8 (.CI(n43861), .I0(GND_net), .I1(n1_adj_5401[6]), 
            .CO(n43862));
    SB_LUT4 mult_16_i14_2_lut (.I0(\Kp[0] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n20_adj_5280));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i14_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5424_9 (.CI(n44956), .I0(n18505[6]), .I1(n618), .CO(n44957));
    SB_LUT4 unary_minus_26_add_3_7_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5401[5]), 
            .I3(n43860), .O(n436[5])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_20_inv_0_i8_1_lut (.I0(deadband[7]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5403[7]));   // verilog/motorControl.v(51[43:52])
    defparam unary_minus_20_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_5424_8_lut (.I0(GND_net), .I1(n18505[5]), .I2(n545), .I3(n44955), 
            .O(n18218[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5424_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_add_1225_20_lut (.I0(GND_net), .I1(n11935[17]), .I2(GND_net), 
            .I3(n45169), .O(n257[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_16_add_1225_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5136_16_lut (.I0(GND_net), .I1(n13786[13]), .I2(n1102_adj_4889), 
            .I3(n45124), .O(n12905[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5136_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_20_inv_0_i9_1_lut (.I0(deadband[8]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5403[8]));   // verilog/motorControl.v(51[43:52])
    defparam unary_minus_20_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_5424_8 (.CI(n44955), .I0(n18505[5]), .I1(n545), .CO(n44956));
    SB_LUT4 add_5360_9_lut (.I0(GND_net), .I1(n17686[6]), .I2(n612), .I3(n44747), 
            .O(n17266[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5360_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_26_add_3_7 (.CI(n43860), .I0(GND_net), .I1(n1_adj_5401[5]), 
            .CO(n43861));
    SB_LUT4 sub_8_add_2_25_lut (.I0(GND_net), .I1(setpoint[23]), .I2(motor_state[23]), 
            .I3(n43687), .O(n1[23])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_8_add_2_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i300_2_lut (.I0(\Kp[6] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n445_adj_5283));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i300_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mult_16_add_1225_20 (.CI(n45169), .I0(n11935[17]), .I1(GND_net), 
            .CO(n45170));
    SB_LUT4 mult_16_add_1225_19_lut (.I0(GND_net), .I1(n11935[16]), .I2(GND_net), 
            .I3(n45168), .O(n257[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_16_add_1225_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5136_16 (.CI(n45124), .I0(n13786[13]), .I1(n1102_adj_4889), 
            .CO(n45125));
    SB_CARRY mult_16_add_1225_19 (.CI(n45168), .I0(n11935[16]), .I1(GND_net), 
            .CO(n45169));
    SB_CARRY add_5360_9 (.CI(n44747), .I0(n17686[6]), .I1(n612), .CO(n44748));
    SB_LUT4 add_5360_8_lut (.I0(GND_net), .I1(n17686[5]), .I2(n539), .I3(n44746), 
            .O(n17266[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5360_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i110_2_lut (.I0(\Kp[2] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n162_adj_5284));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i110_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_20_inv_0_i10_1_lut (.I0(deadband[9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5403[9]));   // verilog/motorControl.v(51[43:52])
    defparam unary_minus_20_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_5360_8 (.CI(n44746), .I0(n17686[5]), .I1(n539), .CO(n44747));
    SB_LUT4 mult_17_i171_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n253));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i171_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i220_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n326));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i220_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i39070_3_lut_4_lut (.I0(n130[3]), .I1(n182[3]), .I2(n182[2]), 
            .I3(n130[2]), .O(n54900));   // verilog/motorControl.v(47[21:44])
    defparam i39070_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 add_5250_15_lut (.I0(GND_net), .I1(n15953[12]), .I2(n1038), 
            .I3(n45061), .O(n15306[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5250_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_12_i6_3_lut_3_lut (.I0(n130[3]), .I1(n182[3]), .I2(n182[2]), 
            .I3(GND_net), .O(n6_adj_5005));   // verilog/motorControl.v(47[21:44])
    defparam LessThan_12_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 add_5360_7_lut (.I0(GND_net), .I1(n17686[4]), .I2(n466), .I3(n44745), 
            .O(n17266[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5360_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i39105_3_lut_4_lut (.I0(IntegralLimit[3]), .I1(n130[3]), .I2(n130[2]), 
            .I3(IntegralLimit[2]), .O(n54935));   // verilog/motorControl.v(45[12:34])
    defparam i39105_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 sub_8_add_2_24_lut (.I0(GND_net), .I1(setpoint[22]), .I2(motor_state[22]), 
            .I3(n43686), .O(n1[22])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_8_add_2_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_10_i6_3_lut_3_lut (.I0(IntegralLimit[3]), .I1(n130[3]), 
            .I2(n130[2]), .I3(GND_net), .O(n6_adj_4915));   // verilog/motorControl.v(45[12:34])
    defparam LessThan_10_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_DFF \PID_CONTROLLER.integral_i0_i1  (.Q(\PID_CONTROLLER.integral [1]), 
           .C(clk16MHz), .D(n29915));   // verilog/motorControl.v(41[14] 61[8])
    SB_LUT4 add_5424_7_lut (.I0(GND_net), .I1(n18505[4]), .I2(n472), .I3(n44954), 
            .O(n18218[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5424_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5136_15_lut (.I0(GND_net), .I1(n13786[12]), .I2(n1029), 
            .I3(n45123), .O(n12905[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5136_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5424_7 (.CI(n44954), .I0(n18505[4]), .I1(n472), .CO(n44955));
    SB_CARRY add_5136_15 (.CI(n45123), .I0(n13786[12]), .I1(n1029), .CO(n45124));
    SB_LUT4 mult_16_add_1225_18_lut (.I0(GND_net), .I1(n11935[15]), .I2(GND_net), 
            .I3(n45167), .O(n257[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_16_add_1225_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i590_2_lut (.I0(\Kp[12] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n877_adj_5287));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i590_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5360_7 (.CI(n44745), .I0(n17686[4]), .I1(n466), .CO(n44746));
    SB_CARRY sub_8_add_2_24 (.CI(n43686), .I0(setpoint[22]), .I1(motor_state[22]), 
            .CO(n43687));
    SB_LUT4 add_5424_6_lut (.I0(GND_net), .I1(n18505[3]), .I2(n399_adj_5288), 
            .I3(n44953), .O(n18218[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5424_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5360_6_lut (.I0(GND_net), .I1(n17686[3]), .I2(n393_adj_5289), 
            .I3(n44744), .O(n17266[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5360_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_16_add_1225_18 (.CI(n45167), .I0(n11935[15]), .I1(GND_net), 
            .CO(n45168));
    SB_LUT4 mult_16_add_1225_17_lut (.I0(GND_net), .I1(n11935[14]), .I2(GND_net), 
            .I3(n45166), .O(n257[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_16_add_1225_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5424_6 (.CI(n44953), .I0(n18505[3]), .I1(n399_adj_5288), 
            .CO(n44954));
    SB_LUT4 add_5136_14_lut (.I0(GND_net), .I1(n13786[11]), .I2(n956_adj_5290), 
            .I3(n45122), .O(n12905[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5136_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5424_5_lut (.I0(GND_net), .I1(n18505[2]), .I2(n326_adj_5291), 
            .I3(n44952), .O(n18218[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5424_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5360_6 (.CI(n44744), .I0(n17686[3]), .I1(n393_adj_5289), 
            .CO(n44745));
    SB_LUT4 add_5360_5_lut (.I0(GND_net), .I1(n17686[2]), .I2(n320_adj_5292), 
            .I3(n44743), .O(n17266[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5360_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5360_5 (.CI(n44743), .I0(n17686[2]), .I1(n320_adj_5292), 
            .CO(n44744));
    SB_CARRY add_5424_5 (.CI(n44952), .I0(n18505[2]), .I1(n326_adj_5291), 
            .CO(n44953));
    SB_LUT4 add_5360_4_lut (.I0(GND_net), .I1(n17686[1]), .I2(n247_adj_5293), 
            .I3(n44742), .O(n17266[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5360_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5360_4 (.CI(n44742), .I0(n17686[1]), .I1(n247_adj_5293), 
            .CO(n44743));
    SB_CARRY add_5250_15 (.CI(n45061), .I0(n15953[12]), .I1(n1038), .CO(n45062));
    SB_LUT4 add_5360_3_lut (.I0(GND_net), .I1(n17686[0]), .I2(n174_adj_5294), 
            .I3(n44741), .O(n17266[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5360_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5424_4_lut (.I0(GND_net), .I1(n18505[1]), .I2(n253_adj_5295), 
            .I3(n44951), .O(n18218[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5424_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_26_add_3_6_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5401[4]), 
            .I3(n43859), .O(n436[4])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5360_3 (.CI(n44741), .I0(n17686[0]), .I1(n174_adj_5294), 
            .CO(n44742));
    SB_LUT4 add_5360_2_lut (.I0(GND_net), .I1(n32_adj_5297), .I2(n101_adj_5298), 
            .I3(GND_net), .O(n17266[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5360_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_8_add_2_23_lut (.I0(GND_net), .I1(setpoint[21]), .I2(motor_state[21]), 
            .I3(n43685), .O(n1[21])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_8_add_2_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5424_4 (.CI(n44951), .I0(n18505[1]), .I1(n253_adj_5295), 
            .CO(n44952));
    SB_CARRY sub_8_add_2_23 (.CI(n43685), .I0(setpoint[21]), .I1(motor_state[21]), 
            .CO(n43686));
    SB_CARRY unary_minus_26_add_3_6 (.CI(n43859), .I0(GND_net), .I1(n1_adj_5401[4]), 
            .CO(n43860));
    SB_LUT4 unary_minus_26_add_3_5_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5401[3]), 
            .I3(n43858), .O(n436[3])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5360_2 (.CI(GND_net), .I0(n32_adj_5297), .I1(n101_adj_5298), 
            .CO(n44741));
    SB_LUT4 sub_8_add_2_22_lut (.I0(GND_net), .I1(setpoint[20]), .I2(motor_state[20]), 
            .I3(n43684), .O(n1[20])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_8_add_2_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5514_8_lut (.I0(GND_net), .I1(n19330[5]), .I2(n560_adj_5300), 
            .I3(n44740), .O(n19233[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5514_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_i269_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n399_adj_5301));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i269_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5514_7_lut (.I0(GND_net), .I1(n19330[4]), .I2(n487_adj_5302), 
            .I3(n44739), .O(n19233[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5514_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_26_add_3_5 (.CI(n43858), .I0(GND_net), .I1(n1_adj_5401[3]), 
            .CO(n43859));
    SB_CARRY sub_8_add_2_22 (.CI(n43684), .I0(setpoint[20]), .I1(motor_state[20]), 
            .CO(n43685));
    SB_LUT4 unary_minus_26_add_3_4_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5401[2]), 
            .I3(n43857), .O(n436[2])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_8_add_2_21_lut (.I0(GND_net), .I1(setpoint[19]), .I2(motor_state[19]), 
            .I3(n43683), .O(n1[19])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_8_add_2_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5514_7 (.CI(n44739), .I0(n19330[4]), .I1(n487_adj_5302), 
            .CO(n44740));
    SB_CARRY sub_8_add_2_21 (.CI(n43683), .I0(setpoint[19]), .I1(motor_state[19]), 
            .CO(n43684));
    SB_LUT4 sub_8_add_2_20_lut (.I0(GND_net), .I1(setpoint[18]), .I2(motor_state[18]), 
            .I3(n43682), .O(n1[18])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_8_add_2_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_8_add_2_20 (.CI(n43682), .I0(setpoint[18]), .I1(motor_state[18]), 
            .CO(n43683));
    SB_CARRY mult_16_add_1225_17 (.CI(n45166), .I0(n11935[14]), .I1(GND_net), 
            .CO(n45167));
    SB_CARRY add_5136_14 (.CI(n45122), .I0(n13786[11]), .I1(n956_adj_5290), 
            .CO(n45123));
    SB_LUT4 add_5136_13_lut (.I0(GND_net), .I1(n13786[10]), .I2(n883_adj_5304), 
            .I3(n45121), .O(n12905[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5136_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_20_inv_0_i11_1_lut (.I0(deadband[10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5403[10]));   // verilog/motorControl.v(51[43:52])
    defparam unary_minus_20_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY unary_minus_26_add_3_4 (.CI(n43857), .I0(GND_net), .I1(n1_adj_5401[2]), 
            .CO(n43858));
    SB_LUT4 unary_minus_26_add_3_3_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5401[1]), 
            .I3(n43856), .O(n436[1])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5136_13 (.CI(n45121), .I0(n13786[10]), .I1(n883_adj_5304), 
            .CO(n45122));
    SB_LUT4 add_5514_6_lut (.I0(GND_net), .I1(n19330[3]), .I2(n414_adj_5307), 
            .I3(n44738), .O(n19233[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5514_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i159_2_lut (.I0(\Kp[3] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n235_adj_5308));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i159_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5424_3_lut (.I0(GND_net), .I1(n18505[0]), .I2(n180_adj_5309), 
            .I3(n44950), .O(n18218[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5424_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5250_14_lut (.I0(GND_net), .I1(n15953[11]), .I2(n965_adj_5310), 
            .I3(n45060), .O(n15306[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5250_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5250_14 (.CI(n45060), .I0(n15953[11]), .I1(n965_adj_5310), 
            .CO(n45061));
    SB_LUT4 sub_8_add_2_19_lut (.I0(GND_net), .I1(setpoint[17]), .I2(motor_state[17]), 
            .I3(n43681), .O(n1[17])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_8_add_2_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_8_add_2_19 (.CI(n43681), .I0(setpoint[17]), .I1(motor_state[17]), 
            .CO(n43682));
    SB_LUT4 sub_8_add_2_18_lut (.I0(GND_net), .I1(setpoint[16]), .I2(motor_state[16]), 
            .I3(n43680), .O(n1[16])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_8_add_2_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5514_6 (.CI(n44738), .I0(n19330[3]), .I1(n414_adj_5307), 
            .CO(n44739));
    SB_CARRY add_5424_3 (.CI(n44950), .I0(n18505[0]), .I1(n180_adj_5309), 
            .CO(n44951));
    SB_LUT4 add_5424_2_lut (.I0(GND_net), .I1(n38_adj_5311), .I2(n107_adj_5312), 
            .I3(GND_net), .O(n18218[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5424_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_26_add_3_3 (.CI(n43856), .I0(GND_net), .I1(n1_adj_5401[1]), 
            .CO(n43857));
    SB_LUT4 add_5514_5_lut (.I0(GND_net), .I1(n19330[2]), .I2(n341_adj_5313), 
            .I3(n44737), .O(n19233[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5514_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_add_1225_16_lut (.I0(GND_net), .I1(n11935[13]), .I2(n1096_adj_5314), 
            .I3(n45165), .O(n257[15])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_16_add_1225_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_8_add_2_18 (.CI(n43680), .I0(setpoint[16]), .I1(motor_state[16]), 
            .CO(n43681));
    SB_CARRY add_5514_5 (.CI(n44737), .I0(n19330[2]), .I1(n341_adj_5313), 
            .CO(n44738));
    SB_LUT4 unary_minus_26_add_3_2_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5401[0]), 
            .I3(VCC_net), .O(n436[0])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5514_4_lut (.I0(GND_net), .I1(n19330[1]), .I2(n268_adj_5316), 
            .I3(n44736), .O(n19233[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5514_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5514_4 (.CI(n44736), .I0(n19330[1]), .I1(n268_adj_5316), 
            .CO(n44737));
    SB_LUT4 add_5250_13_lut (.I0(GND_net), .I1(n15953[10]), .I2(n892_adj_5317), 
            .I3(n45059), .O(n15306[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5250_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5424_2 (.CI(GND_net), .I0(n38_adj_5311), .I1(n107_adj_5312), 
            .CO(n44950));
    SB_LUT4 add_5136_12_lut (.I0(GND_net), .I1(n13786[9]), .I2(n810_adj_5318), 
            .I3(n45120), .O(n12905[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5136_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_8_add_2_17_lut (.I0(GND_net), .I1(setpoint[15]), .I2(motor_state[15]), 
            .I3(n43679), .O(n1[15])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_8_add_2_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5514_3_lut (.I0(GND_net), .I1(n19330[0]), .I2(n195_adj_5319), 
            .I3(n44735), .O(n19233[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5514_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_8_add_2_17 (.CI(n43679), .I0(setpoint[15]), .I1(motor_state[15]), 
            .CO(n43680));
    SB_LUT4 sub_8_add_2_16_lut (.I0(GND_net), .I1(setpoint[14]), .I2(motor_state[14]), 
            .I3(n43678), .O(n1[14])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_8_add_2_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5136_12 (.CI(n45120), .I0(n13786[9]), .I1(n810_adj_5318), 
            .CO(n45121));
    SB_CARRY add_5250_13 (.CI(n45059), .I0(n15953[10]), .I1(n892_adj_5317), 
            .CO(n45060));
    SB_CARRY unary_minus_26_add_3_2 (.CI(VCC_net), .I0(GND_net), .I1(n1_adj_5401[0]), 
            .CO(n43856));
    SB_LUT4 add_5250_12_lut (.I0(GND_net), .I1(n15953[9]), .I2(n819_adj_5320), 
            .I3(n45058), .O(n15306[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5250_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5250_12 (.CI(n45058), .I0(n15953[9]), .I1(n819_adj_5320), 
            .CO(n45059));
    SB_LUT4 add_5446_12_lut (.I0(GND_net), .I1(n18746[9]), .I2(n840_adj_5321), 
            .I3(n44949), .O(n18505[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5446_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5446_11_lut (.I0(GND_net), .I1(n18746[8]), .I2(n767_adj_5322), 
            .I3(n44948), .O(n18505[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5446_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_20_add_3_25_lut (.I0(n356[23]), .I1(GND_net), .I2(n1_adj_5403[23]), 
            .I3(n43855), .O(n47_adj_5128)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_25_lut.LUT_INIT = 16'h6996;
    SB_CARRY sub_8_add_2_16 (.CI(n43678), .I0(setpoint[14]), .I1(motor_state[14]), 
            .CO(n43679));
    SB_CARRY add_5514_3 (.CI(n44735), .I0(n19330[0]), .I1(n195_adj_5319), 
            .CO(n44736));
    SB_LUT4 sub_8_add_2_15_lut (.I0(GND_net), .I1(setpoint[13]), .I2(motor_state[13]), 
            .I3(n43677), .O(n1[13])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_8_add_2_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5514_2_lut (.I0(GND_net), .I1(n53_adj_5324), .I2(n122_adj_5325), 
            .I3(GND_net), .O(n19233[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5514_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_8_add_2_15 (.CI(n43677), .I0(setpoint[13]), .I1(motor_state[13]), 
            .CO(n43678));
    SB_LUT4 unary_minus_20_add_3_24_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5403[22]), 
            .I3(n43854), .O(n382[22])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5446_11 (.CI(n44948), .I0(n18746[8]), .I1(n767_adj_5322), 
            .CO(n44949));
    SB_CARRY add_5514_2 (.CI(GND_net), .I0(n53_adj_5324), .I1(n122_adj_5325), 
            .CO(n44735));
    SB_CARRY mult_16_add_1225_16 (.CI(n45165), .I0(n11935[13]), .I1(n1096_adj_5314), 
            .CO(n45166));
    SB_LUT4 add_5387_14_lut (.I0(GND_net), .I1(n18050[11]), .I2(n980_adj_5327), 
            .I3(n44734), .O(n17686[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5387_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_8_add_2_14_lut (.I0(GND_net), .I1(setpoint[12]), .I2(motor_state[12]), 
            .I3(n43676), .O(n1[12])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_8_add_2_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5387_13_lut (.I0(GND_net), .I1(n18050[10]), .I2(n907_adj_5328), 
            .I3(n44733), .O(n17686[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5387_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_24 (.CI(n43854), .I0(GND_net), .I1(n1_adj_5403[22]), 
            .CO(n43855));
    SB_CARRY add_5387_13 (.CI(n44733), .I0(n18050[10]), .I1(n907_adj_5328), 
            .CO(n44734));
    SB_CARRY sub_8_add_2_14 (.CI(n43676), .I0(setpoint[12]), .I1(motor_state[12]), 
            .CO(n43677));
    SB_LUT4 add_5446_10_lut (.I0(GND_net), .I1(n18746[7]), .I2(n694_adj_5329), 
            .I3(n44947), .O(n18505[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5446_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5387_12_lut (.I0(GND_net), .I1(n18050[9]), .I2(n834_adj_5330), 
            .I3(n44732), .O(n17686[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5387_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5387_12 (.CI(n44732), .I0(n18050[9]), .I1(n834_adj_5330), 
            .CO(n44733));
    SB_LUT4 unary_minus_20_add_3_23_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5403[21]), 
            .I3(n43853), .O(n382[21])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_8_add_2_13_lut (.I0(GND_net), .I1(setpoint[11]), .I2(motor_state[11]), 
            .I3(n43675), .O(n1[11])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_8_add_2_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5387_11_lut (.I0(GND_net), .I1(n18050[8]), .I2(n761_adj_5332), 
            .I3(n44731), .O(n17686[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5387_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5387_11 (.CI(n44731), .I0(n18050[8]), .I1(n761_adj_5332), 
            .CO(n44732));
    SB_CARRY unary_minus_20_add_3_23 (.CI(n43853), .I0(GND_net), .I1(n1_adj_5403[21]), 
            .CO(n43854));
    SB_LUT4 unary_minus_20_add_3_22_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5403[20]), 
            .I3(n43852), .O(n382[20])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_22 (.CI(n43852), .I0(GND_net), .I1(n1_adj_5403[20]), 
            .CO(n43853));
    SB_CARRY sub_8_add_2_13 (.CI(n43675), .I0(setpoint[11]), .I1(motor_state[11]), 
            .CO(n43676));
    SB_LUT4 unary_minus_20_add_3_21_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5403[19]), 
            .I3(n43851), .O(n382[19])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_8_add_2_12_lut (.I0(GND_net), .I1(setpoint[10]), .I2(motor_state[10]), 
            .I3(n43674), .O(n1[10])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_8_add_2_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5250_11_lut (.I0(GND_net), .I1(n15953[8]), .I2(n746_adj_5335), 
            .I3(n45057), .O(n15306[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5250_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5446_10 (.CI(n44947), .I0(n18746[7]), .I1(n694_adj_5329), 
            .CO(n44948));
    SB_LUT4 add_5446_9_lut (.I0(GND_net), .I1(n18746[6]), .I2(n621_adj_5336), 
            .I3(n44946), .O(n18505[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5446_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5387_10_lut (.I0(GND_net), .I1(n18050[7]), .I2(n688_adj_5337), 
            .I3(n44730), .O(n17686[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5387_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5387_10 (.CI(n44730), .I0(n18050[7]), .I1(n688_adj_5337), 
            .CO(n44731));
    SB_LUT4 add_5387_9_lut (.I0(GND_net), .I1(n18050[6]), .I2(n615_adj_5338), 
            .I3(n44729), .O(n17686[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5387_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_8_add_2_12 (.CI(n43674), .I0(setpoint[10]), .I1(motor_state[10]), 
            .CO(n43675));
    SB_CARRY add_5387_9 (.CI(n44729), .I0(n18050[6]), .I1(n615_adj_5338), 
            .CO(n44730));
    SB_LUT4 sub_8_add_2_11_lut (.I0(GND_net), .I1(setpoint[9]), .I2(motor_state[9]), 
            .I3(n43673), .O(n1[9])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_8_add_2_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_21 (.CI(n43851), .I0(GND_net), .I1(n1_adj_5403[19]), 
            .CO(n43852));
    SB_CARRY add_5446_9 (.CI(n44946), .I0(n18746[6]), .I1(n621_adj_5336), 
            .CO(n44947));
    SB_LUT4 add_5446_8_lut (.I0(GND_net), .I1(n18746[5]), .I2(n548_adj_5339), 
            .I3(n44945), .O(n18505[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5446_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5387_8_lut (.I0(GND_net), .I1(n18050[5]), .I2(n542_adj_5340), 
            .I3(n44728), .O(n17686[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5387_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5387_8 (.CI(n44728), .I0(n18050[5]), .I1(n542_adj_5340), 
            .CO(n44729));
    SB_LUT4 unary_minus_20_add_3_20_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5403[18]), 
            .I3(n43850), .O(n382[18])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5446_8 (.CI(n44945), .I0(n18746[5]), .I1(n548_adj_5339), 
            .CO(n44946));
    SB_LUT4 add_5446_7_lut (.I0(GND_net), .I1(n18746[4]), .I2(n475_adj_5342), 
            .I3(n44944), .O(n18505[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5446_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5387_7_lut (.I0(GND_net), .I1(n18050[4]), .I2(n469_adj_5343), 
            .I3(n44727), .O(n17686[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5387_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_20 (.CI(n43850), .I0(GND_net), .I1(n1_adj_5403[18]), 
            .CO(n43851));
    SB_CARRY sub_8_add_2_11 (.CI(n43673), .I0(setpoint[9]), .I1(motor_state[9]), 
            .CO(n43674));
    SB_LUT4 unary_minus_20_add_3_19_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5403[17]), 
            .I3(n43849), .O(n382[17])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5387_7 (.CI(n44727), .I0(n18050[4]), .I1(n469_adj_5343), 
            .CO(n44728));
    SB_LUT4 sub_8_add_2_10_lut (.I0(GND_net), .I1(setpoint[8]), .I2(motor_state[8]), 
            .I3(n43672), .O(n1[8])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_8_add_2_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5387_6_lut (.I0(GND_net), .I1(n18050[3]), .I2(n396_adj_5345), 
            .I3(n44726), .O(n17686[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5387_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_20_inv_0_i12_1_lut (.I0(deadband[11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5403[11]));   // verilog/motorControl.v(51[43:52])
    defparam unary_minus_20_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_5136_11_lut (.I0(GND_net), .I1(n13786[8]), .I2(n737_adj_5347), 
            .I3(n45119), .O(n12905[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5136_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_19 (.CI(n43849), .I0(GND_net), .I1(n1_adj_5403[17]), 
            .CO(n43850));
    SB_CARRY add_5446_7 (.CI(n44944), .I0(n18746[4]), .I1(n475_adj_5342), 
            .CO(n44945));
    SB_CARRY sub_8_add_2_10 (.CI(n43672), .I0(setpoint[8]), .I1(motor_state[8]), 
            .CO(n43673));
    SB_CARRY add_5387_6 (.CI(n44726), .I0(n18050[3]), .I1(n396_adj_5345), 
            .CO(n44727));
    SB_LUT4 add_5387_5_lut (.I0(GND_net), .I1(n18050[2]), .I2(n323_adj_5348), 
            .I3(n44725), .O(n17686[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5387_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_20_add_3_18_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5403[16]), 
            .I3(n43848), .O(n382[16])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5250_11 (.CI(n45057), .I0(n15953[8]), .I1(n746_adj_5335), 
            .CO(n45058));
    SB_CARRY add_5387_5 (.CI(n44725), .I0(n18050[2]), .I1(n323_adj_5348), 
            .CO(n44726));
    SB_CARRY add_5136_11 (.CI(n45119), .I0(n13786[8]), .I1(n737_adj_5347), 
            .CO(n45120));
    SB_LUT4 mult_16_add_1225_15_lut (.I0(GND_net), .I1(n11935[12]), .I2(n1023_adj_5350), 
            .I3(n45164), .O(n257[14])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_16_add_1225_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5387_4_lut (.I0(GND_net), .I1(n18050[1]), .I2(n250_adj_5351), 
            .I3(n44724), .O(n17686[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5387_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5136_10_lut (.I0(GND_net), .I1(n13786[7]), .I2(n664_adj_5352), 
            .I3(n45118), .O(n12905[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5136_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_18 (.CI(n43848), .I0(GND_net), .I1(n1_adj_5403[16]), 
            .CO(n43849));
    SB_LUT4 add_5250_10_lut (.I0(GND_net), .I1(n15953[7]), .I2(n673_adj_5353), 
            .I3(n45056), .O(n15306[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5250_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5387_4 (.CI(n44724), .I0(n18050[1]), .I1(n250_adj_5351), 
            .CO(n44725));
    SB_CARRY add_5250_10 (.CI(n45056), .I0(n15953[7]), .I1(n673_adj_5353), 
            .CO(n45057));
    SB_LUT4 mult_17_i318_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n472_adj_5354));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i318_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5446_6_lut (.I0(GND_net), .I1(n18746[3]), .I2(n402_adj_5355), 
            .I3(n44943), .O(n18505[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5446_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5387_3_lut (.I0(GND_net), .I1(n18050[0]), .I2(n177_adj_5356), 
            .I3(n44723), .O(n17686[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5387_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i208_2_lut (.I0(\Kp[4] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n308_adj_5357));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i208_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5446_6 (.CI(n44943), .I0(n18746[3]), .I1(n402_adj_5355), 
            .CO(n44944));
    SB_LUT4 unary_minus_20_add_3_17_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5403[15]), 
            .I3(n43847), .O(n382[15])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5387_3 (.CI(n44723), .I0(n18050[0]), .I1(n177_adj_5356), 
            .CO(n44724));
    SB_LUT4 sub_8_add_2_9_lut (.I0(GND_net), .I1(setpoint[7]), .I2(motor_state[7]), 
            .I3(n43671), .O(n1[7])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_8_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_17 (.CI(n43847), .I0(GND_net), .I1(n1_adj_5403[15]), 
            .CO(n43848));
    SB_LUT4 add_5387_2_lut (.I0(GND_net), .I1(n35_adj_5359), .I2(n104_adj_5360), 
            .I3(GND_net), .O(n17686[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5387_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_i367_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n545_adj_5361));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i367_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5250_9_lut (.I0(GND_net), .I1(n15953[6]), .I2(n600_adj_5362), 
            .I3(n45055), .O(n15306[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5250_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5250_9 (.CI(n45055), .I0(n15953[6]), .I1(n600_adj_5362), 
            .CO(n45056));
    SB_LUT4 mult_17_i704_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n1047_adj_5270));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i704_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i75_2_lut (.I0(\Kp[1] ), .I1(n1[12]), .I2(GND_net), 
            .I3(GND_net), .O(n110_adj_5363));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i75_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5446_5_lut (.I0(GND_net), .I1(n18746[2]), .I2(n329_adj_5364), 
            .I3(n44942), .O(n18505[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5446_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5136_10 (.CI(n45118), .I0(n13786[7]), .I1(n664_adj_5352), 
            .CO(n45119));
    SB_CARRY add_5387_2 (.CI(GND_net), .I0(n35_adj_5359), .I1(n104_adj_5360), 
            .CO(n44723));
    SB_LUT4 add_5412_13_lut (.I0(GND_net), .I1(n18362[10]), .I2(n910_adj_5365), 
            .I3(n44722), .O(n18050[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5412_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5250_8_lut (.I0(GND_net), .I1(n15953[5]), .I2(n527_adj_5366), 
            .I3(n45054), .O(n15306[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5250_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i28_2_lut (.I0(\Kp[0] ), .I1(n1[13]), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_5367));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i28_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5446_5 (.CI(n44942), .I0(n18746[2]), .I1(n329_adj_5364), 
            .CO(n44943));
    SB_LUT4 add_5412_12_lut (.I0(GND_net), .I1(n18362[9]), .I2(n837_adj_5368), 
            .I3(n44721), .O(n18050[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5412_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_16_add_1225_15 (.CI(n45164), .I0(n11935[12]), .I1(n1023_adj_5350), 
            .CO(n45165));
    SB_LUT4 add_5446_4_lut (.I0(GND_net), .I1(n18746[1]), .I2(n256_adj_5369), 
            .I3(n44941), .O(n18505[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5446_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_add_1225_14_lut (.I0(GND_net), .I1(n11935[11]), .I2(n950_adj_5370), 
            .I3(n45163), .O(n257[13])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_16_add_1225_14_lut.LUT_INIT = 16'hC33C;
    SB_DFF \PID_CONTROLLER.integral_i0_i2  (.Q(\PID_CONTROLLER.integral [2]), 
           .C(clk16MHz), .D(n29914));   // verilog/motorControl.v(41[14] 61[8])
    SB_CARRY add_5412_12 (.CI(n44721), .I0(n18362[9]), .I1(n837_adj_5368), 
            .CO(n44722));
    SB_LUT4 add_5136_9_lut (.I0(GND_net), .I1(n13786[6]), .I2(n591_adj_5371), 
            .I3(n45117), .O(n12905[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5136_9_lut.LUT_INIT = 16'hC33C;
    SB_DFF \PID_CONTROLLER.integral_i0_i3  (.Q(\PID_CONTROLLER.integral [3]), 
           .C(clk16MHz), .D(n29913));   // verilog/motorControl.v(41[14] 61[8])
    SB_DFF \PID_CONTROLLER.integral_i0_i4  (.Q(\PID_CONTROLLER.integral [4]), 
           .C(clk16MHz), .D(n29912));   // verilog/motorControl.v(41[14] 61[8])
    SB_CARRY sub_8_add_2_9 (.CI(n43671), .I0(setpoint[7]), .I1(motor_state[7]), 
            .CO(n43672));
    SB_DFF \PID_CONTROLLER.integral_i0_i5  (.Q(\PID_CONTROLLER.integral [5]), 
           .C(clk16MHz), .D(n29911));   // verilog/motorControl.v(41[14] 61[8])
    SB_LUT4 unary_minus_20_add_3_16_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5403[14]), 
            .I3(n43846), .O(n382[14])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_16_lut.LUT_INIT = 16'hC33C;
    SB_DFF \PID_CONTROLLER.integral_i0_i6  (.Q(\PID_CONTROLLER.integral [6]), 
           .C(clk16MHz), .D(n29910));   // verilog/motorControl.v(41[14] 61[8])
    SB_CARRY add_5250_8 (.CI(n45054), .I0(n15953[5]), .I1(n527_adj_5366), 
            .CO(n45055));
    SB_LUT4 add_5412_11_lut (.I0(GND_net), .I1(n18362[8]), .I2(n764_adj_5373), 
            .I3(n44720), .O(n18050[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5412_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5412_11 (.CI(n44720), .I0(n18362[8]), .I1(n764_adj_5373), 
            .CO(n44721));
    SB_LUT4 add_5412_10_lut (.I0(GND_net), .I1(n18362[7]), .I2(n691_adj_5374), 
            .I3(n44719), .O(n18050[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5412_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5250_7_lut (.I0(GND_net), .I1(n15953[4]), .I2(n454_adj_5375), 
            .I3(n45053), .O(n15306[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5250_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5136_9 (.CI(n45117), .I0(n13786[6]), .I1(n591_adj_5371), 
            .CO(n45118));
    SB_CARRY unary_minus_20_add_3_16 (.CI(n43846), .I0(GND_net), .I1(n1_adj_5403[14]), 
            .CO(n43847));
    SB_CARRY add_5446_4 (.CI(n44941), .I0(n18746[1]), .I1(n256_adj_5369), 
            .CO(n44942));
    SB_LUT4 unary_minus_20_add_3_15_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5403[13]), 
            .I3(n43845), .O(n382[13])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5250_7 (.CI(n45053), .I0(n15953[4]), .I1(n454_adj_5375), 
            .CO(n45054));
    SB_LUT4 add_5136_8_lut (.I0(GND_net), .I1(n13786[5]), .I2(n518_adj_5377), 
            .I3(n45116), .O(n12905[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5136_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5412_10 (.CI(n44719), .I0(n18362[7]), .I1(n691_adj_5374), 
            .CO(n44720));
    SB_LUT4 sub_8_add_2_8_lut (.I0(GND_net), .I1(setpoint[6]), .I2(motor_state[6]), 
            .I3(n43670), .O(n1[6])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_8_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5250_6_lut (.I0(GND_net), .I1(n15953[3]), .I2(n381_adj_5378), 
            .I3(n45052), .O(n15306[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5250_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_15 (.CI(n43845), .I0(GND_net), .I1(n1_adj_5403[13]), 
            .CO(n43846));
    SB_LUT4 unary_minus_20_add_3_14_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5403[12]), 
            .I3(n43844), .O(n382[12])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5446_3_lut (.I0(GND_net), .I1(n18746[0]), .I2(n183_adj_5380), 
            .I3(n44940), .O(n18505[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5446_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5412_9_lut (.I0(GND_net), .I1(n18362[6]), .I2(n618_adj_5381), 
            .I3(n44718), .O(n18050[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5412_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5446_3 (.CI(n44940), .I0(n18746[0]), .I1(n183_adj_5380), 
            .CO(n44941));
    SB_CARRY add_5412_9 (.CI(n44718), .I0(n18362[6]), .I1(n618_adj_5381), 
            .CO(n44719));
    SB_CARRY mult_16_add_1225_14 (.CI(n45163), .I0(n11935[11]), .I1(n950_adj_5370), 
            .CO(n45164));
    SB_CARRY add_5250_6 (.CI(n45052), .I0(n15953[3]), .I1(n381_adj_5378), 
            .CO(n45053));
    SB_LUT4 add_5446_2_lut (.I0(GND_net), .I1(n41_adj_5367), .I2(n110_adj_5363), 
            .I3(GND_net), .O(n18505[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5446_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5446_2 (.CI(GND_net), .I0(n41_adj_5367), .I1(n110_adj_5363), 
            .CO(n44940));
    SB_LUT4 add_5412_8_lut (.I0(GND_net), .I1(n18362[5]), .I2(n545_adj_5361), 
            .I3(n44717), .O(n18050[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5412_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_add_1225_24_lut (.I0(\PID_CONTROLLER.integral_23__N_3996 [23]), 
            .I1(n11404[21]), .I2(GND_net), .I3(n44939), .O(n10897[0])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1225_24_lut.LUT_INIT = 16'h6996;
    SB_CARRY add_5412_8 (.CI(n44717), .I0(n18362[5]), .I1(n545_adj_5361), 
            .CO(n44718));
    SB_LUT4 mult_17_i281_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [17]), 
            .I2(GND_net), .I3(GND_net), .O(n417_adj_5269));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i281_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_add_1225_23_lut (.I0(GND_net), .I1(n11404[20]), .I2(GND_net), 
            .I3(n44938), .O(n306[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1225_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5250_5_lut (.I0(GND_net), .I1(n15953[2]), .I2(n308_adj_5357), 
            .I3(n45051), .O(n15306[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5250_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5412_7_lut (.I0(GND_net), .I1(n18362[4]), .I2(n472_adj_5354), 
            .I3(n44716), .O(n18050[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5412_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_8_add_2_8 (.CI(n43670), .I0(setpoint[6]), .I1(motor_state[6]), 
            .CO(n43671));
    SB_CARRY add_5250_5 (.CI(n45051), .I0(n15953[2]), .I1(n308_adj_5357), 
            .CO(n45052));
    SB_LUT4 mult_17_i416_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n618_adj_5381));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i416_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mult_17_add_1225_23 (.CI(n44938), .I0(n11404[20]), .I1(GND_net), 
            .CO(n44939));
    SB_LUT4 i1_4_lut_adj_1687 (.I0(n19426[2]), .I1(n6_adj_5382), .I2(\Ki[4] ), 
            .I3(\PID_CONTROLLER.integral_23__N_3996 [18]), .O(n19366[3]));   // verilog/motorControl.v(50[27:38])
    defparam i1_4_lut_adj_1687.LUT_INIT = 16'h9666;
    SB_CARRY unary_minus_20_add_3_14 (.CI(n43844), .I0(GND_net), .I1(n1_adj_5403[12]), 
            .CO(n43845));
    SB_LUT4 sub_8_add_2_7_lut (.I0(GND_net), .I1(setpoint[5]), .I2(motor_state[5]), 
            .I3(n43669), .O(n1[5])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_8_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i124_2_lut (.I0(\Kp[2] ), .I1(n1[12]), .I2(GND_net), 
            .I3(GND_net), .O(n183_adj_5380));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i124_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_add_1225_22_lut (.I0(GND_net), .I1(n11404[19]), .I2(GND_net), 
            .I3(n44937), .O(n306[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1225_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5412_7 (.CI(n44716), .I0(n18362[4]), .I1(n472_adj_5354), 
            .CO(n44717));
    SB_LUT4 unary_minus_20_inv_0_i13_1_lut (.I0(deadband[12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5403[12]));   // verilog/motorControl.v(51[43:52])
    defparam unary_minus_20_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_20_add_3_13_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5403[11]), 
            .I3(n43843), .O(n382[11])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i257_2_lut (.I0(\Kp[5] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n381_adj_5378));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i257_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY unary_minus_20_add_3_13 (.CI(n43843), .I0(GND_net), .I1(n1_adj_5403[11]), 
            .CO(n43844));
    SB_LUT4 add_5250_4_lut (.I0(GND_net), .I1(n15953[1]), .I2(n235_adj_5308), 
            .I3(n45050), .O(n15306[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5250_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_20_add_3_12_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5403[10]), 
            .I3(n43842), .O(n382[10])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5412_6_lut (.I0(GND_net), .I1(n18362[3]), .I2(n399_adj_5301), 
            .I3(n44715), .O(n18050[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5412_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_add_1225_13_lut (.I0(GND_net), .I1(n11935[10]), .I2(n877_adj_5287), 
            .I3(n45162), .O(n257[12])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_16_add_1225_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_8_add_2_7 (.CI(n43669), .I0(setpoint[5]), .I1(motor_state[5]), 
            .CO(n43670));
    SB_CARRY unary_minus_20_add_3_12 (.CI(n43842), .I0(GND_net), .I1(n1_adj_5403[10]), 
            .CO(n43843));
    SB_CARRY add_5412_6 (.CI(n44715), .I0(n18362[3]), .I1(n399_adj_5301), 
            .CO(n44716));
    SB_CARRY mult_16_add_1225_13 (.CI(n45162), .I0(n11935[10]), .I1(n877_adj_5287), 
            .CO(n45163));
    SB_LUT4 sub_8_add_2_6_lut (.I0(GND_net), .I1(setpoint[4]), .I2(motor_state[4]), 
            .I3(n43668), .O(n1[4])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_8_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5250_4 (.CI(n45050), .I0(n15953[1]), .I1(n235_adj_5308), 
            .CO(n45051));
    SB_LUT4 add_5412_5_lut (.I0(GND_net), .I1(n18362[2]), .I2(n326), .I3(n44714), 
            .O(n18050[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5412_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5412_5 (.CI(n44714), .I0(n18362[2]), .I1(n326), .CO(n44715));
    SB_LUT4 mult_17_i79_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [14]), 
            .I2(GND_net), .I3(GND_net), .O(n116_adj_5268));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i79_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5412_4_lut (.I0(GND_net), .I1(n18362[1]), .I2(n253), .I3(n44713), 
            .O(n18050[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5412_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_17_add_1225_22 (.CI(n44937), .I0(n11404[19]), .I1(GND_net), 
            .CO(n44938));
    SB_CARRY add_5136_8 (.CI(n45116), .I0(n13786[5]), .I1(n518_adj_5377), 
            .CO(n45117));
    SB_LUT4 unary_minus_20_add_3_11_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5403[9]), 
            .I3(n43841), .O(n382[9])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5250_3_lut (.I0(GND_net), .I1(n15953[0]), .I2(n162_adj_5284), 
            .I3(n45049), .O(n15306[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5250_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5136_7_lut (.I0(GND_net), .I1(n13786[4]), .I2(n445_adj_5283), 
            .I3(n45115), .O(n12905[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5136_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i349_2_lut (.I0(\Kp[7] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n518_adj_5377));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i349_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5250_3 (.CI(n45049), .I0(n15953[0]), .I1(n162_adj_5284), 
            .CO(n45050));
    SB_CARRY unary_minus_20_add_3_11 (.CI(n43841), .I0(GND_net), .I1(n1_adj_5403[9]), 
            .CO(n43842));
    SB_LUT4 unary_minus_20_add_3_10_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5403[8]), 
            .I3(n43840), .O(n382[8])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_8_add_2_6 (.CI(n43668), .I0(setpoint[4]), .I1(motor_state[4]), 
            .CO(n43669));
    SB_LUT4 unary_minus_20_inv_0_i14_1_lut (.I0(deadband[13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5403[13]));   // verilog/motorControl.v(51[43:52])
    defparam unary_minus_20_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_5136_7 (.CI(n45115), .I0(n13786[4]), .I1(n445_adj_5283), 
            .CO(n45116));
    SB_LUT4 mult_16_i306_2_lut (.I0(\Kp[6] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n454_adj_5375));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i306_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i465_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n691_adj_5374));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i465_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_add_1225_21_lut (.I0(GND_net), .I1(n11404[18]), .I2(GND_net), 
            .I3(n44936), .O(n306[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1225_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_10 (.CI(n43840), .I0(GND_net), .I1(n1_adj_5403[8]), 
            .CO(n43841));
    SB_LUT4 unary_minus_20_add_3_9_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5403[7]), 
            .I3(n43839), .O(n382[7])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5412_4 (.CI(n44713), .I0(n18362[1]), .I1(n253), .CO(n44714));
    SB_LUT4 add_5250_2_lut (.I0(GND_net), .I1(n20_adj_5280), .I2(n89_adj_5279), 
            .I3(GND_net), .O(n15306[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5250_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_9 (.CI(n43839), .I0(GND_net), .I1(n1_adj_5403[7]), 
            .CO(n43840));
    SB_CARRY mult_17_add_1225_21 (.CI(n44936), .I0(n11404[18]), .I1(GND_net), 
            .CO(n44937));
    SB_LUT4 unary_minus_20_add_3_8_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5403[6]), 
            .I3(n43838), .O(n382[6])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5412_3_lut (.I0(GND_net), .I1(n18362[0]), .I2(n180), .I3(n44712), 
            .O(n18050[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5412_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5412_3 (.CI(n44712), .I0(n18362[0]), .I1(n180), .CO(n44713));
    SB_LUT4 mult_17_add_1225_20_lut (.I0(GND_net), .I1(n11404[17]), .I2(GND_net), 
            .I3(n44935), .O(n306[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1225_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_17_add_1225_20 (.CI(n44935), .I0(n11404[17]), .I1(GND_net), 
            .CO(n44936));
    SB_LUT4 add_5412_2_lut (.I0(GND_net), .I1(n38), .I2(n107_adj_5277), 
            .I3(GND_net), .O(n18050[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5412_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_8 (.CI(n43838), .I0(GND_net), .I1(n1_adj_5403[6]), 
            .CO(n43839));
    SB_CARRY add_5412_2 (.CI(GND_net), .I0(n38), .I1(n107_adj_5277), .CO(n44712));
    SB_LUT4 add_5526_7_lut (.I0(GND_net), .I1(n50980), .I2(n490), .I3(n44711), 
            .O(n19330[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5526_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5526_6_lut (.I0(GND_net), .I1(n19401[3]), .I2(n417), .I3(n44710), 
            .O(n19330[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5526_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_20_add_3_7_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5403[5]), 
            .I3(n43837), .O(n382[5])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_7 (.CI(n43837), .I0(GND_net), .I1(n1_adj_5403[5]), 
            .CO(n43838));
    SB_LUT4 unary_minus_20_add_3_6_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5403[4]), 
            .I3(n43836), .O(n382[4])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_6 (.CI(n43836), .I0(GND_net), .I1(n1_adj_5403[4]), 
            .CO(n43837));
    SB_LUT4 unary_minus_20_add_3_5_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5403[3]), 
            .I3(n43835), .O(n382[3])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5526_6 (.CI(n44710), .I0(n19401[3]), .I1(n417), .CO(n44711));
    SB_LUT4 sub_8_add_2_5_lut (.I0(GND_net), .I1(setpoint[3]), .I2(motor_state[3]), 
            .I3(n43667), .O(n1[3])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_8_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_8_add_2_5 (.CI(n43667), .I0(setpoint[3]), .I1(motor_state[3]), 
            .CO(n43668));
    SB_CARRY unary_minus_20_add_3_5 (.CI(n43835), .I0(GND_net), .I1(n1_adj_5403[3]), 
            .CO(n43836));
    SB_LUT4 sub_8_add_2_4_lut (.I0(GND_net), .I1(setpoint[2]), .I2(motor_state[2]), 
            .I3(n43666), .O(n1[2])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_8_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_i514_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n764_adj_5373));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i514_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_20_inv_0_i15_1_lut (.I0(deadband[14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5403[14]));   // verilog/motorControl.v(51[43:52])
    defparam unary_minus_20_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_20_add_3_4_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5403[2]), 
            .I3(n43834), .O(n382[2])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5526_5_lut (.I0(GND_net), .I1(n19401[2]), .I2(n344_adj_5214), 
            .I3(n44709), .O(n19330[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5526_5_lut.LUT_INIT = 16'hC33C;
    SB_DFF \PID_CONTROLLER.integral_i0_i7  (.Q(\PID_CONTROLLER.integral [7]), 
           .C(clk16MHz), .D(n29909));   // verilog/motorControl.v(41[14] 61[8])
    SB_CARRY unary_minus_20_add_3_4 (.CI(n43834), .I0(GND_net), .I1(n1_adj_5403[2]), 
            .CO(n43835));
    SB_LUT4 unary_minus_20_add_3_3_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5403[1]), 
            .I3(n43833), .O(n382[1])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_add_1225_12_lut (.I0(GND_net), .I1(n11935[9]), .I2(n804_adj_5210), 
            .I3(n45161), .O(n257[11])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_16_add_1225_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5526_5 (.CI(n44709), .I0(n19401[2]), .I1(n344_adj_5214), 
            .CO(n44710));
    SB_LUT4 add_5526_4_lut (.I0(GND_net), .I1(n19401[1]), .I2(n271), .I3(n44708), 
            .O(n19330[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5526_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5136_6_lut (.I0(GND_net), .I1(n13786[3]), .I2(n372_adj_5208), 
            .I3(n45114), .O(n12905[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5136_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5526_4 (.CI(n44708), .I0(n19401[1]), .I1(n271), .CO(n44709));
    SB_LUT4 add_5526_3_lut (.I0(GND_net), .I1(n19401[0]), .I2(n198_adj_5206), 
            .I3(n44707), .O(n19330[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5526_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_8_add_2_4 (.CI(n43666), .I0(setpoint[2]), .I1(motor_state[2]), 
            .CO(n43667));
    SB_CARRY unary_minus_20_add_3_3 (.CI(n43833), .I0(GND_net), .I1(n1_adj_5403[1]), 
            .CO(n43834));
    SB_LUT4 unary_minus_20_add_3_2_lut (.I0(n37221), .I1(GND_net), .I2(n1_adj_5403[0]), 
            .I3(VCC_net), .O(n54560)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY unary_minus_20_add_3_2 (.CI(VCC_net), .I0(GND_net), .I1(n1_adj_5403[0]), 
            .CO(n43833));
    SB_CARRY add_5250_2 (.CI(GND_net), .I0(n20_adj_5280), .I1(n89_adj_5279), 
            .CO(n45049));
    SB_LUT4 mult_17_add_1225_19_lut (.I0(GND_net), .I1(n11404[16]), .I2(GND_net), 
            .I3(n44934), .O(n306[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1225_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_8_add_2_3_lut (.I0(GND_net), .I1(setpoint[1]), .I2(motor_state[1]), 
            .I3(n43665), .O(n1[1])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_8_add_2_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_17_add_1225_19 (.CI(n44934), .I0(n11404[16]), .I1(GND_net), 
            .CO(n44935));
    SB_CARRY add_5526_3 (.CI(n44707), .I0(n19401[0]), .I1(n198_adj_5206), 
            .CO(n44708));
    SB_LUT4 add_5526_2_lut (.I0(GND_net), .I1(n56_adj_5201), .I2(n125_adj_5200), 
            .I3(GND_net), .O(n19330[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5526_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5526_2 (.CI(GND_net), .I0(n56_adj_5201), .I1(n125_adj_5200), 
            .CO(n44707));
    SB_LUT4 add_5435_12_lut (.I0(GND_net), .I1(n18626[9]), .I2(n840), 
            .I3(n44706), .O(n18362[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5435_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_add_1225_18_lut (.I0(GND_net), .I1(n11404[15]), .I2(GND_net), 
            .I3(n44933), .O(n306[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1225_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5435_11_lut (.I0(GND_net), .I1(n18626[8]), .I2(n767), 
            .I3(n44705), .O(n18362[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5435_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_13_add_3_25_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5402[23]), 
            .I3(n43832), .O(n182[23])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_17_add_1225_18 (.CI(n44933), .I0(n11404[15]), .I1(GND_net), 
            .CO(n44934));
    SB_CARRY sub_8_add_2_3 (.CI(n43665), .I0(setpoint[1]), .I1(motor_state[1]), 
            .CO(n43666));
    SB_CARRY add_5435_11 (.CI(n44705), .I0(n18626[8]), .I1(n767), .CO(n44706));
    SB_CARRY mult_16_add_1225_12 (.CI(n45161), .I0(n11935[9]), .I1(n804_adj_5210), 
            .CO(n45162));
    SB_LUT4 unary_minus_13_add_3_24_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5402[22]), 
            .I3(n43831), .O(n182[22])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5136_6 (.CI(n45114), .I0(n13786[3]), .I1(n372_adj_5208), 
            .CO(n45115));
    SB_LUT4 add_5284_18_lut (.I0(GND_net), .I1(n16530[15]), .I2(GND_net), 
            .I3(n45048), .O(n15953[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5284_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_add_1225_17_lut (.I0(GND_net), .I1(n11404[14]), .I2(GND_net), 
            .I3(n44932), .O(n306[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1225_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5435_10_lut (.I0(GND_net), .I1(n18626[7]), .I2(n694), 
            .I3(n44704), .O(n18362[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5435_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_13_add_3_24 (.CI(n43831), .I0(GND_net), .I1(n1_adj_5402[22]), 
            .CO(n43832));
    SB_CARRY add_5435_10 (.CI(n44704), .I0(n18626[7]), .I1(n694), .CO(n44705));
    SB_CARRY mult_17_add_1225_17 (.CI(n44932), .I0(n11404[14]), .I1(GND_net), 
            .CO(n44933));
    SB_LUT4 unary_minus_13_add_3_23_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5402[21]), 
            .I3(n43830), .O(n182[21])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5435_9_lut (.I0(GND_net), .I1(n18626[6]), .I2(n621), .I3(n44703), 
            .O(n18362[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5435_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_add_1225_11_lut (.I0(GND_net), .I1(n11935[8]), .I2(n731_adj_5198), 
            .I3(n45160), .O(n257[10])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_16_add_1225_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5435_9 (.CI(n44703), .I0(n18626[6]), .I1(n621), .CO(n44704));
    SB_CARRY unary_minus_13_add_3_23 (.CI(n43830), .I0(GND_net), .I1(n1_adj_5402[21]), 
            .CO(n43831));
    SB_LUT4 unary_minus_13_add_3_22_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5402[20]), 
            .I3(n43829), .O(n182[20])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_13_add_3_22 (.CI(n43829), .I0(GND_net), .I1(n1_adj_5402[20]), 
            .CO(n43830));
    SB_LUT4 add_5136_5_lut (.I0(GND_net), .I1(n13786[2]), .I2(n299_adj_5196), 
            .I3(n45113), .O(n12905[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5136_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5284_17_lut (.I0(GND_net), .I1(n16530[14]), .I2(GND_net), 
            .I3(n45047), .O(n15953[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5284_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_13_add_3_21_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5402[19]), 
            .I3(n43828), .O(n182[19])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5435_8_lut (.I0(GND_net), .I1(n18626[5]), .I2(n548), .I3(n44702), 
            .O(n18362[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5435_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_13_add_3_21 (.CI(n43828), .I0(GND_net), .I1(n1_adj_5402[19]), 
            .CO(n43829));
    SB_CARRY add_5284_17 (.CI(n45047), .I0(n16530[14]), .I1(GND_net), 
            .CO(n45048));
    SB_LUT4 mult_17_add_1225_16_lut (.I0(GND_net), .I1(n11404[13]), .I2(n1096), 
            .I3(n44931), .O(n306[15])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1225_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_13_add_3_20_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5402[18]), 
            .I3(n43827), .O(n182[18])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_13_add_3_20 (.CI(n43827), .I0(GND_net), .I1(n1_adj_5402[18]), 
            .CO(n43828));
    SB_LUT4 unary_minus_13_add_3_19_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5402[17]), 
            .I3(n43826), .O(n182[17])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_17_add_1225_16 (.CI(n44931), .I0(n11404[13]), .I1(n1096), 
            .CO(n44932));
    SB_LUT4 sub_8_add_2_2_lut (.I0(GND_net), .I1(setpoint[0]), .I2(motor_state[0]), 
            .I3(VCC_net), .O(n1[0])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_8_add_2_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5435_8 (.CI(n44702), .I0(n18626[5]), .I1(n548), .CO(n44703));
    SB_LUT4 add_5435_7_lut (.I0(GND_net), .I1(n18626[4]), .I2(n475), .I3(n44701), 
            .O(n18362[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5435_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5435_7 (.CI(n44701), .I0(n18626[4]), .I1(n475), .CO(n44702));
    SB_LUT4 mult_17_add_1225_15_lut (.I0(GND_net), .I1(n11404[12]), .I2(n1023), 
            .I3(n44930), .O(n306[14])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1225_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5435_6_lut (.I0(GND_net), .I1(n18626[3]), .I2(n402_adj_5192), 
            .I3(n44700), .O(n18362[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5435_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i398_2_lut (.I0(\Kp[8] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n591_adj_5371));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i398_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY unary_minus_13_add_3_19 (.CI(n43826), .I0(GND_net), .I1(n1_adj_5402[17]), 
            .CO(n43827));
    SB_LUT4 unary_minus_13_add_3_18_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5402[16]), 
            .I3(n43825), .O(n182[16])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_8_add_2_2 (.CI(VCC_net), .I0(setpoint[0]), .I1(motor_state[0]), 
            .CO(n43665));
    SB_LUT4 mult_17_i32_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [15]), 
            .I2(GND_net), .I3(GND_net), .O(n47_adj_5267));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i32_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5435_6 (.CI(n44700), .I0(n18626[3]), .I1(n402_adj_5192), 
            .CO(n44701));
    SB_CARRY mult_17_add_1225_15 (.CI(n44930), .I0(n11404[12]), .I1(n1023), 
            .CO(n44931));
    SB_LUT4 mult_17_add_1225_14_lut (.I0(GND_net), .I1(n11404[11]), .I2(n950), 
            .I3(n44929), .O(n306[13])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1225_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5284_16_lut (.I0(GND_net), .I1(n16530[13]), .I2(n1114_adj_5190), 
            .I3(n45046), .O(n15953[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5284_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_17_add_1225_14 (.CI(n44929), .I0(n11404[11]), .I1(n950), 
            .CO(n44930));
    SB_CARRY unary_minus_13_add_3_18 (.CI(n43825), .I0(GND_net), .I1(n1_adj_5402[16]), 
            .CO(n43826));
    SB_LUT4 unary_minus_13_add_3_17_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5402[15]), 
            .I3(n43824), .O(n182[15])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_13_add_3_17 (.CI(n43824), .I0(GND_net), .I1(n1_adj_5402[15]), 
            .CO(n43825));
    SB_LUT4 add_5435_5_lut (.I0(GND_net), .I1(n18626[2]), .I2(n329), .I3(n44699), 
            .O(n18362[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5435_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_13_add_3_16_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5402[14]), 
            .I3(n43823), .O(n182[14])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_16_add_1225_11 (.CI(n45160), .I0(n11935[8]), .I1(n731_adj_5198), 
            .CO(n45161));
    SB_LUT4 mult_16_i639_2_lut (.I0(\Kp[13] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n950_adj_5370));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i639_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY unary_minus_13_add_3_16 (.CI(n43823), .I0(GND_net), .I1(n1_adj_5402[14]), 
            .CO(n43824));
    SB_CARRY add_5435_5 (.CI(n44699), .I0(n18626[2]), .I1(n329), .CO(n44700));
    SB_LUT4 mult_17_add_1225_13_lut (.I0(GND_net), .I1(n11404[10]), .I2(n877), 
            .I3(n44928), .O(n306[12])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1225_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5435_4_lut (.I0(GND_net), .I1(n18626[1]), .I2(n256), .I3(n44698), 
            .O(n18362[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5435_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5435_4 (.CI(n44698), .I0(n18626[1]), .I1(n256), .CO(n44699));
    SB_LUT4 add_5435_3_lut (.I0(GND_net), .I1(n18626[0]), .I2(n183_adj_5187), 
            .I3(n44697), .O(n18362[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5435_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5435_3 (.CI(n44697), .I0(n18626[0]), .I1(n183_adj_5187), 
            .CO(n44698));
    SB_LUT4 add_5435_2_lut (.I0(GND_net), .I1(n41_adj_5186), .I2(n110_adj_5185), 
            .I3(GND_net), .O(n18362[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5435_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5435_2 (.CI(GND_net), .I0(n41_adj_5186), .I1(n110_adj_5185), 
            .CO(n44697));
    SB_LUT4 unary_minus_13_add_3_15_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5402[13]), 
            .I3(n43822), .O(n182[13])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_13_add_3_15 (.CI(n43822), .I0(GND_net), .I1(n1_adj_5402[13]), 
            .CO(n43823));
    SB_LUT4 unary_minus_13_add_3_14_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5402[12]), 
            .I3(n43821), .O(n182[12])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_13_add_3_14 (.CI(n43821), .I0(GND_net), .I1(n1_adj_5402[12]), 
            .CO(n43822));
    SB_LUT4 unary_minus_13_add_3_13_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5402[11]), 
            .I3(n43820), .O(n182[11])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_13_add_3_13 (.CI(n43820), .I0(GND_net), .I1(n1_adj_5402[11]), 
            .CO(n43821));
    SB_LUT4 unary_minus_13_add_3_12_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5402[10]), 
            .I3(n43819), .O(n182[10])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_13_add_3_12 (.CI(n43819), .I0(GND_net), .I1(n1_adj_5402[10]), 
            .CO(n43820));
    SB_LUT4 unary_minus_13_add_3_11_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5402[9]), 
            .I3(n43818), .O(n182[9])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_13_add_3_11 (.CI(n43818), .I0(GND_net), .I1(n1_adj_5402[9]), 
            .CO(n43819));
    SB_LUT4 unary_minus_13_add_3_10_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5402[8]), 
            .I3(n43817), .O(n182[8])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_13_add_3_10 (.CI(n43817), .I0(GND_net), .I1(n1_adj_5402[8]), 
            .CO(n43818));
    SB_LUT4 unary_minus_13_add_3_9_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5402[7]), 
            .I3(n43816), .O(n182[7])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_9_lut.LUT_INIT = 16'hC33C;
    SB_DFF \PID_CONTROLLER.integral_i0_i8  (.Q(\PID_CONTROLLER.integral [8]), 
           .C(clk16MHz), .D(n29908));   // verilog/motorControl.v(41[14] 61[8])
    SB_CARRY mult_17_add_1225_13 (.CI(n44928), .I0(n11404[10]), .I1(n877), 
            .CO(n44929));
    SB_DFF \PID_CONTROLLER.integral_i0_i9  (.Q(\PID_CONTROLLER.integral [9]), 
           .C(clk16MHz), .D(n29907));   // verilog/motorControl.v(41[14] 61[8])
    SB_DFF \PID_CONTROLLER.integral_i0_i10  (.Q(\PID_CONTROLLER.integral [10]), 
           .C(clk16MHz), .D(n29906));   // verilog/motorControl.v(41[14] 61[8])
    SB_LUT4 mult_17_add_1225_12_lut (.I0(GND_net), .I1(n11404[9]), .I2(n804), 
            .I3(n44927), .O(n306[11])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1225_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_13_add_3_9 (.CI(n43816), .I0(GND_net), .I1(n1_adj_5402[7]), 
            .CO(n43817));
    SB_LUT4 unary_minus_13_add_3_8_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5402[6]), 
            .I3(n43815), .O(n182[6])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_13_add_3_8 (.CI(n43815), .I0(GND_net), .I1(n1_adj_5402[6]), 
            .CO(n43816));
    SB_LUT4 unary_minus_13_add_3_7_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5402[5]), 
            .I3(n43814), .O(n182[5])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_13_add_3_7 (.CI(n43814), .I0(GND_net), .I1(n1_adj_5402[5]), 
            .CO(n43815));
    SB_LUT4 unary_minus_13_add_3_6_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5402[4]), 
            .I3(n43813), .O(n182[4])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5284_16 (.CI(n45046), .I0(n16530[13]), .I1(n1114_adj_5190), 
            .CO(n45047));
    SB_DFF \PID_CONTROLLER.integral_i0_i11  (.Q(\PID_CONTROLLER.integral [11]), 
           .C(clk16MHz), .D(n29905));   // verilog/motorControl.v(41[14] 61[8])
    SB_DFF \PID_CONTROLLER.integral_i0_i12  (.Q(\PID_CONTROLLER.integral [12]), 
           .C(clk16MHz), .D(n29904));   // verilog/motorControl.v(41[14] 61[8])
    SB_CARRY mult_17_add_1225_12 (.CI(n44927), .I0(n11404[9]), .I1(n804), 
            .CO(n44928));
    SB_DFF \PID_CONTROLLER.integral_i0_i13  (.Q(\PID_CONTROLLER.integral [13]), 
           .C(clk16MHz), .D(n29903));   // verilog/motorControl.v(41[14] 61[8])
    SB_LUT4 mult_17_add_1225_11_lut (.I0(GND_net), .I1(n11404[8]), .I2(n731), 
            .I3(n44926), .O(n306[10])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1225_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i173_2_lut (.I0(\Kp[3] ), .I1(n1[12]), .I2(GND_net), 
            .I3(GND_net), .O(n256_adj_5369));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i173_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY unary_minus_13_add_3_6 (.CI(n43813), .I0(GND_net), .I1(n1_adj_5402[4]), 
            .CO(n43814));
    SB_LUT4 unary_minus_13_add_3_5_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5402[3]), 
            .I3(n43812), .O(n182[3])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_13_add_3_5 (.CI(n43812), .I0(GND_net), .I1(n1_adj_5402[3]), 
            .CO(n43813));
    SB_LUT4 add_5284_15_lut (.I0(GND_net), .I1(n16530[12]), .I2(n1041_adj_5173), 
            .I3(n45045), .O(n15953[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5284_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_13_add_3_4_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5402[2]), 
            .I3(n43811), .O(n182[2])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_13_add_3_4 (.CI(n43811), .I0(GND_net), .I1(n1_adj_5402[2]), 
            .CO(n43812));
    SB_LUT4 unary_minus_13_add_3_3_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5402[1]), 
            .I3(n43810), .O(n182[1])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_13_add_3_3 (.CI(n43810), .I0(GND_net), .I1(n1_adj_5402[1]), 
            .CO(n43811));
    SB_LUT4 unary_minus_13_add_3_2_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5402[0]), 
            .I3(VCC_net), .O(n182[0])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_2_lut.LUT_INIT = 16'hC33C;
    SB_DFF \PID_CONTROLLER.integral_i0_i14  (.Q(\PID_CONTROLLER.integral [14]), 
           .C(clk16MHz), .D(n29902));   // verilog/motorControl.v(41[14] 61[8])
    SB_DFF \PID_CONTROLLER.integral_i0_i15  (.Q(\PID_CONTROLLER.integral [15]), 
           .C(clk16MHz), .D(n29901));   // verilog/motorControl.v(41[14] 61[8])
    SB_CARRY unary_minus_13_add_3_2 (.CI(VCC_net), .I0(GND_net), .I1(n1_adj_5402[0]), 
            .CO(n43810));
    SB_DFF \PID_CONTROLLER.integral_i0_i16  (.Q(\PID_CONTROLLER.integral [16]), 
           .C(clk16MHz), .D(n29900));   // verilog/motorControl.v(41[14] 61[8])
    SB_LUT4 mult_17_i563_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n837_adj_5368));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i563_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mult_17_add_1225_11 (.CI(n44926), .I0(n11404[8]), .I1(n731), 
            .CO(n44927));
    SB_LUT4 mult_16_i355_2_lut (.I0(\Kp[7] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n527_adj_5366));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i355_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5284_15 (.CI(n45045), .I0(n16530[12]), .I1(n1041_adj_5173), 
            .CO(n45046));
    SB_LUT4 add_5284_14_lut (.I0(GND_net), .I1(n16530[11]), .I2(n968_adj_5169), 
            .I3(n45044), .O(n15953[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5284_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_i612_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n910_adj_5365));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i612_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_add_1225_10_lut (.I0(GND_net), .I1(n11935[7]), .I2(n658_adj_5168), 
            .I3(n45159), .O(n257[9])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_16_add_1225_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_add_1225_10_lut (.I0(GND_net), .I1(n11404[7]), .I2(n658), 
            .I3(n44925), .O(n306[9])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1225_10_lut.LUT_INIT = 16'hC33C;
    SB_DFF \PID_CONTROLLER.integral_i0_i17  (.Q(\PID_CONTROLLER.integral [17]), 
           .C(clk16MHz), .D(n29899));   // verilog/motorControl.v(41[14] 61[8])
    SB_DFF \PID_CONTROLLER.integral_i0_i18  (.Q(\PID_CONTROLLER.integral [18]), 
           .C(clk16MHz), .D(n29898));   // verilog/motorControl.v(41[14] 61[8])
    SB_DFF \PID_CONTROLLER.integral_i0_i19  (.Q(\PID_CONTROLLER.integral [19]), 
           .C(clk16MHz), .D(n29897));   // verilog/motorControl.v(41[14] 61[8])
    SB_LUT4 mult_16_i222_2_lut (.I0(\Kp[4] ), .I1(n1[12]), .I2(GND_net), 
            .I3(GND_net), .O(n329_adj_5364));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i222_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i29376_3_lut_4_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [22]), 
            .I2(\PID_CONTROLLER.integral_23__N_3996 [21]), .I3(\Ki[1] ), 
            .O(n19490[0]));   // verilog/motorControl.v(50[27:38])
    defparam i29376_3_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 i29378_3_lut_4_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [22]), 
            .I2(\PID_CONTROLLER.integral_23__N_3996 [21]), .I3(\Ki[1] ), 
            .O(n43478));   // verilog/motorControl.v(50[27:38])
    defparam i29378_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_CARRY mult_17_add_1225_10 (.CI(n44925), .I0(n11404[7]), .I1(n658), 
            .CO(n44926));
    SB_LUT4 mult_16_i404_2_lut (.I0(\Kp[8] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n600_adj_5362));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i404_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i29193_2_lut_3_lut_4_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [21]), 
            .I2(\PID_CONTROLLER.integral_23__N_3996 [20]), .I3(\Ki[1] ), 
            .O(n19466[0]));   // verilog/motorControl.v(50[27:38])
    defparam i29193_2_lut_3_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 mux_14_i12_3_lut (.I0(n130[11]), .I1(n182[11]), .I2(n181), 
            .I3(GND_net), .O(n207[11]));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_14_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29195_2_lut_3_lut_4_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [21]), 
            .I2(\PID_CONTROLLER.integral_23__N_3996 [20]), .I3(\Ki[1] ), 
            .O(n43280));   // verilog/motorControl.v(50[27:38])
    defparam i29195_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_CARRY mult_16_add_1225_10 (.CI(n45159), .I0(n11935[7]), .I1(n658_adj_5168), 
            .CO(n45160));
    SB_CARRY add_5136_5 (.CI(n45113), .I0(n13786[2]), .I1(n299_adj_5196), 
            .CO(n45114));
    SB_LUT4 mux_15_i12_3_lut (.I0(n207[11]), .I1(IntegralLimit[11]), .I2(n155), 
            .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3996 [11]));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_15_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF \PID_CONTROLLER.integral_i0_i20  (.Q(\PID_CONTROLLER.integral [20]), 
           .C(clk16MHz), .D(n29896));   // verilog/motorControl.v(41[14] 61[8])
    SB_DFF \PID_CONTROLLER.integral_i0_i21  (.Q(\PID_CONTROLLER.integral [21]), 
           .C(clk16MHz), .D(n29895));   // verilog/motorControl.v(41[14] 61[8])
    SB_DFF \PID_CONTROLLER.integral_i0_i22  (.Q(\PID_CONTROLLER.integral [22]), 
           .C(clk16MHz), .D(n29894));   // verilog/motorControl.v(41[14] 61[8])
    SB_LUT4 add_5136_4_lut (.I0(GND_net), .I1(n13786[1]), .I2(n226_adj_5167), 
            .I3(n45112), .O(n12905[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5136_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5136_4 (.CI(n45112), .I0(n13786[1]), .I1(n226_adj_5167), 
            .CO(n45113));
    SB_CARRY add_5284_14 (.CI(n45044), .I0(n16530[11]), .I1(n968_adj_5169), 
            .CO(n45045));
    SB_LUT4 mult_17_add_1225_9_lut (.I0(GND_net), .I1(n11404[6]), .I2(n585_adj_5166), 
            .I3(n44924), .O(n306[8])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1225_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5284_13_lut (.I0(GND_net), .I1(n16530[10]), .I2(n895_adj_5165), 
            .I3(n45043), .O(n15953[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5284_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5136_3_lut (.I0(GND_net), .I1(n13786[0]), .I2(n153_adj_5164), 
            .I3(n45111), .O(n12905[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5136_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_i71_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n104_adj_5360));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i71_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mult_17_add_1225_9 (.CI(n44924), .I0(n11404[6]), .I1(n585_adj_5166), 
            .CO(n44925));
    SB_LUT4 mult_17_i24_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_5359));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i24_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5284_13 (.CI(n45043), .I0(n16530[10]), .I1(n895_adj_5165), 
            .CO(n45044));
    SB_LUT4 mult_17_add_1225_8_lut (.I0(GND_net), .I1(n11404[5]), .I2(n512_adj_5163), 
            .I3(n44923), .O(n306[7])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1225_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5284_12_lut (.I0(GND_net), .I1(n16530[9]), .I2(n822_adj_5162), 
            .I3(n45042), .O(n15953[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5284_12_lut.LUT_INIT = 16'hC33C;
    SB_DFF \PID_CONTROLLER.integral_i0_i23  (.Q(\PID_CONTROLLER.integral [23]), 
           .C(clk16MHz), .D(n29893));   // verilog/motorControl.v(41[14] 61[8])
    SB_LUT4 i29290_3_lut_4_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [18]), 
            .I2(n4_adj_5384), .I3(n19426[1]), .O(n6_adj_5382));   // verilog/motorControl.v(50[27:38])
    defparam i29290_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_CARRY mult_17_add_1225_8 (.CI(n44923), .I0(n11404[5]), .I1(n512_adj_5163), 
            .CO(n44924));
    SB_LUT4 mult_17_add_1225_7_lut (.I0(GND_net), .I1(n11404[4]), .I2(n439_adj_5161), 
            .I3(n44922), .O(n306[6])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1225_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_3_lut_4_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [18]), 
            .I2(n4_adj_5384), .I3(n19426[1]), .O(n19366[2]));   // verilog/motorControl.v(50[27:38])
    defparam i1_3_lut_4_lut.LUT_INIT = 16'h8778;
    SB_CARRY mult_17_add_1225_7 (.CI(n44922), .I0(n11404[4]), .I1(n439_adj_5161), 
            .CO(n44923));
    SB_LUT4 i1_3_lut_4_lut_adj_1688 (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [18]), 
            .I2(n43362), .I3(n19426[0]), .O(n19366[1]));   // verilog/motorControl.v(50[27:38])
    defparam i1_3_lut_4_lut_adj_1688.LUT_INIT = 16'h8778;
    SB_LUT4 i29282_3_lut_4_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [18]), 
            .I2(n43362), .I3(n19426[0]), .O(n4_adj_5384));   // verilog/motorControl.v(50[27:38])
    defparam i29282_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 mult_16_add_1225_9_lut (.I0(GND_net), .I1(n11935[6]), .I2(n585), 
            .I3(n45158), .O(n257[8])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_16_add_1225_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5284_12 (.CI(n45042), .I0(n16530[9]), .I1(n822_adj_5162), 
            .CO(n45043));
    SB_LUT4 mult_17_add_1225_6_lut (.I0(GND_net), .I1(n11404[3]), .I2(n366_adj_5160), 
            .I3(n44921), .O(n306[5])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1225_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i29269_2_lut_3_lut_4_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [19]), 
            .I2(\PID_CONTROLLER.integral_23__N_3996 [18]), .I3(\Ki[1] ), 
            .O(n19366[0]));   // verilog/motorControl.v(50[27:38])
    defparam i29269_2_lut_3_lut_4_lut.LUT_INIT = 16'h7888;
    SB_CARRY mult_17_add_1225_6 (.CI(n44921), .I0(n11404[3]), .I1(n366_adj_5160), 
            .CO(n44922));
    SB_CARRY add_5136_3 (.CI(n45111), .I0(n13786[0]), .I1(n153_adj_5164), 
            .CO(n45112));
    SB_LUT4 i29271_2_lut_3_lut_4_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [19]), 
            .I2(\PID_CONTROLLER.integral_23__N_3996 [18]), .I3(\Ki[1] ), 
            .O(n43362));   // verilog/motorControl.v(50[27:38])
    defparam i29271_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 unary_minus_20_inv_0_i16_1_lut (.I0(deadband[15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5403[15]));   // verilog/motorControl.v(51[43:52])
    defparam unary_minus_20_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_5284_11_lut (.I0(GND_net), .I1(n16530[8]), .I2(n749_adj_5159), 
            .I3(n45041), .O(n15953[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5284_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_add_1225_5_lut (.I0(GND_net), .I1(n11404[2]), .I2(n293_adj_5158), 
            .I3(n44920), .O(n306[4])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1225_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_17_add_1225_5 (.CI(n44920), .I0(n11404[2]), .I1(n293_adj_5158), 
            .CO(n44921));
    SB_LUT4 mult_16_i751_2_lut (.I0(\Kp[15] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n1117));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i751_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i447_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n664));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i447_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5136_2_lut (.I0(GND_net), .I1(n11_adj_5155), .I2(n80_adj_5154), 
            .I3(GND_net), .O(n12905[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5136_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_add_1225_4_lut (.I0(GND_net), .I1(n11404[1]), .I2(n220_adj_5153), 
            .I3(n44919), .O(n306[3])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1225_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_16_add_1225_9 (.CI(n45158), .I0(n11935[6]), .I1(n585), 
            .CO(n45159));
    SB_CARRY add_5284_11 (.CI(n45041), .I0(n16530[8]), .I1(n749_adj_5159), 
            .CO(n45042));
    SB_CARRY mult_17_add_1225_4 (.CI(n44919), .I0(n11404[1]), .I1(n220_adj_5153), 
            .CO(n44920));
    SB_LUT4 mult_17_add_1225_3_lut (.I0(GND_net), .I1(n11404[0]), .I2(n147_adj_5150), 
            .I3(n44918), .O(n306[2])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1225_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5284_10_lut (.I0(GND_net), .I1(n16530[7]), .I2(n676_adj_5149), 
            .I3(n45040), .O(n15953[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5284_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_add_1225_8_lut (.I0(GND_net), .I1(n11935[5]), .I2(n512), 
            .I3(n45157), .O(n257[7])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_16_add_1225_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_17_add_1225_3 (.CI(n44918), .I0(n11404[0]), .I1(n147_adj_5150), 
            .CO(n44919));
    SB_CARRY add_5136_2 (.CI(GND_net), .I0(n11_adj_5155), .I1(n80_adj_5154), 
            .CO(n45111));
    SB_LUT4 add_5176_21_lut (.I0(GND_net), .I1(n14585[18]), .I2(GND_net), 
            .I3(n45110), .O(n13786[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5176_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_add_1225_2_lut (.I0(GND_net), .I1(n5_adj_5147), .I2(n74_adj_5146), 
            .I3(GND_net), .O(n306[1])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1225_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_16_add_1225_8 (.CI(n45157), .I0(n11935[5]), .I1(n512), 
            .CO(n45158));
    SB_LUT4 mult_16_add_1225_7_lut (.I0(GND_net), .I1(n11935[4]), .I2(n439_adj_5144), 
            .I3(n45156), .O(n257[6])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_16_add_1225_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_17_add_1225_2 (.CI(GND_net), .I0(n5_adj_5147), .I1(n74_adj_5146), 
            .CO(n44918));
    SB_CARRY mult_16_add_1225_7 (.CI(n45156), .I0(n11935[4]), .I1(n439_adj_5144), 
            .CO(n45157));
    SB_LUT4 mult_16_i400_2_lut (.I0(\Kp[8] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n594));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i400_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5070_23_lut (.I0(GND_net), .I1(n12422[20]), .I2(GND_net), 
            .I3(n44917), .O(n11404[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5070_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5070_22_lut (.I0(GND_net), .I1(n12422[19]), .I2(GND_net), 
            .I3(n44916), .O(n11404[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5070_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i29252_3_lut_4_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [19]), 
            .I2(n4_adj_5385), .I3(n19466[1]), .O(n6_adj_5386));   // verilog/motorControl.v(50[27:38])
    defparam i29252_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 mult_17_i120_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n177_adj_5356));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i120_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i271_2_lut (.I0(\Kp[5] ), .I1(n1[12]), .I2(GND_net), 
            .I3(GND_net), .O(n402_adj_5355));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i271_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_3_lut_4_lut_adj_1689 (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [19]), 
            .I2(n4_adj_5385), .I3(n19466[1]), .O(n19426[2]));   // verilog/motorControl.v(50[27:38])
    defparam i1_3_lut_4_lut_adj_1689.LUT_INIT = 16'h8778;
    SB_LUT4 add_5176_20_lut (.I0(GND_net), .I1(n14585[17]), .I2(GND_net), 
            .I3(n45109), .O(n13786[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5176_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_add_1225_6_lut (.I0(GND_net), .I1(n11935[3]), .I2(n366_adj_5111), 
            .I3(n45155), .O(n257[5])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_16_add_1225_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_16_add_1225_6 (.CI(n45155), .I0(n11935[3]), .I1(n366_adj_5111), 
            .CO(n45156));
    SB_LUT4 mult_16_i453_2_lut (.I0(\Kp[9] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n673_adj_5353));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i453_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i447_2_lut (.I0(\Kp[9] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n664_adj_5352));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i447_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i449_2_lut (.I0(\Kp[9] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n667));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i449_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i169_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n250_adj_5351));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i169_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i688_2_lut (.I0(\Kp[14] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n1023_adj_5350));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i688_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5070_22 (.CI(n44916), .I0(n12422[19]), .I1(GND_net), 
            .CO(n44917));
    SB_CARRY add_5284_10 (.CI(n45040), .I0(n16530[7]), .I1(n676_adj_5149), 
            .CO(n45041));
    SB_LUT4 unary_minus_20_inv_0_i17_1_lut (.I0(deadband[16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5403[16]));   // verilog/motorControl.v(51[43:52])
    defparam unary_minus_20_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_16_add_1225_5_lut (.I0(GND_net), .I1(n11935[2]), .I2(n293), 
            .I3(n45154), .O(n257[4])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_16_add_1225_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5176_20 (.CI(n45109), .I0(n14585[17]), .I1(GND_net), 
            .CO(n45110));
    SB_CARRY mult_16_add_1225_5 (.CI(n45154), .I0(n11935[2]), .I1(n293), 
            .CO(n45155));
    SB_LUT4 mult_17_i218_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n323_adj_5348));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i218_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5284_9_lut (.I0(GND_net), .I1(n16530[6]), .I2(n603_adj_5036), 
            .I3(n45039), .O(n15953[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5284_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_3_lut_4_lut_adj_1690 (.I0(n62_adj_5387), .I1(n131_adj_5388), 
            .I2(n204_adj_5389), .I3(n19466[0]), .O(n19426[1]));   // verilog/motorControl.v(50[27:38])
    defparam i1_3_lut_4_lut_adj_1690.LUT_INIT = 16'h8778;
    SB_LUT4 mult_17_i496_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n737));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i496_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5176_19_lut (.I0(GND_net), .I1(n14585[16]), .I2(GND_net), 
            .I3(n45108), .O(n13786[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5176_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_add_1225_4_lut (.I0(GND_net), .I1(n11935[1]), .I2(n220), 
            .I3(n45153), .O(n257[3])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_16_add_1225_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5070_21_lut (.I0(GND_net), .I1(n12422[18]), .I2(GND_net), 
            .I3(n44915), .O(n11404[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5070_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5070_21 (.CI(n44915), .I0(n12422[18]), .I1(GND_net), 
            .CO(n44916));
    SB_CARRY mult_16_add_1225_4 (.CI(n45153), .I0(n11935[1]), .I1(n220), 
            .CO(n45154));
    SB_LUT4 mult_17_i545_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n810));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i545_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i29244_3_lut_4_lut (.I0(n62_adj_5387), .I1(n131_adj_5388), .I2(n204_adj_5389), 
            .I3(n19466[0]), .O(n4_adj_5385));   // verilog/motorControl.v(50[27:38])
    defparam i29244_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 mult_16_i496_2_lut (.I0(\Kp[10] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n737_adj_5347));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i496_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i267_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n396_adj_5345));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i267_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_14_i17_3_lut (.I0(n130[16]), .I1(n182[16]), .I2(n181), 
            .I3(GND_net), .O(n207[16]));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_14_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_15_i17_3_lut (.I0(n207[16]), .I1(IntegralLimit[16]), .I2(n155), 
            .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3996 [16]));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_15_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_5284_9 (.CI(n45039), .I0(n16530[6]), .I1(n603_adj_5036), 
            .CO(n45040));
    SB_CARRY add_5176_19 (.CI(n45108), .I0(n14585[16]), .I1(GND_net), 
            .CO(n45109));
    SB_LUT4 add_5176_18_lut (.I0(GND_net), .I1(n14585[15]), .I2(GND_net), 
            .I3(n45107), .O(n13786[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5176_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_20_inv_0_i18_1_lut (.I0(deadband[17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5403[17]));   // verilog/motorControl.v(51[43:52])
    defparam unary_minus_20_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_5070_20_lut (.I0(GND_net), .I1(n12422[17]), .I2(GND_net), 
            .I3(n44914), .O(n11404[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5070_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_i753_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n1120_adj_5266));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i753_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_add_1225_3_lut (.I0(GND_net), .I1(n11935[0]), .I2(n147_adj_4958), 
            .I3(n45152), .O(n257[2])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_16_add_1225_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5176_18 (.CI(n45107), .I0(n14585[15]), .I1(GND_net), 
            .CO(n45108));
    SB_LUT4 add_5284_8_lut (.I0(GND_net), .I1(n16530[5]), .I2(n530_adj_4952), 
            .I3(n45038), .O(n15953[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5284_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5284_8 (.CI(n45038), .I0(n16530[5]), .I1(n530_adj_4952), 
            .CO(n45039));
    SB_CARRY add_5070_20 (.CI(n44914), .I0(n12422[17]), .I1(GND_net), 
            .CO(n44915));
    SB_LUT4 add_5070_19_lut (.I0(GND_net), .I1(n12422[16]), .I2(GND_net), 
            .I3(n44913), .O(n11404[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5070_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5284_7_lut (.I0(GND_net), .I1(n16530[4]), .I2(n457_adj_4917), 
            .I3(n45037), .O(n15953[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5284_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5070_19 (.CI(n44913), .I0(n12422[16]), .I1(GND_net), 
            .CO(n44914));
    SB_LUT4 mult_17_i81_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [15]), 
            .I2(GND_net), .I3(GND_net), .O(n119));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i81_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5070_18_lut (.I0(GND_net), .I1(n12422[15]), .I2(GND_net), 
            .I3(n44912), .O(n11404[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5070_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i29231_2_lut_4_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [20]), 
            .I2(\Ki[1] ), .I3(\PID_CONTROLLER.integral_23__N_3996 [19]), 
            .O(n19426[0]));   // verilog/motorControl.v(50[27:38])
    defparam i29231_2_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 add_5176_17_lut (.I0(GND_net), .I1(n14585[14]), .I2(GND_net), 
            .I3(n45106), .O(n13786[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5176_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_16_add_1225_3 (.CI(n45152), .I0(n11935[0]), .I1(n147_adj_4958), 
            .CO(n45153));
    SB_CARRY add_5070_18 (.CI(n44912), .I0(n12422[15]), .I1(GND_net), 
            .CO(n44913));
    SB_LUT4 mult_17_i34_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [16]), 
            .I2(GND_net), .I3(GND_net), .O(n50));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i34_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i594_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n883));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i594_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i316_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n469_adj_5343));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i316_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i320_2_lut (.I0(\Kp[6] ), .I1(n1[12]), .I2(GND_net), 
            .I3(GND_net), .O(n475_adj_5342));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i320_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_20_inv_0_i19_1_lut (.I0(deadband[18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5403[18]));   // verilog/motorControl.v(51[43:52])
    defparam unary_minus_20_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_16_add_1225_2_lut (.I0(GND_net), .I1(n5), .I2(n74), .I3(GND_net), 
            .O(n257[1])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_16_add_1225_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5176_17 (.CI(n45106), .I0(n14585[14]), .I1(GND_net), 
            .CO(n45107));
    SB_LUT4 add_5070_17_lut (.I0(GND_net), .I1(n12422[14]), .I2(GND_net), 
            .I3(n44911), .O(n11404[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5070_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_i643_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n956));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i643_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5284_7 (.CI(n45037), .I0(n16530[4]), .I1(n457_adj_4917), 
            .CO(n45038));
    SB_CARRY add_5070_17 (.CI(n44911), .I0(n12422[14]), .I1(GND_net), 
            .CO(n44912));
    SB_LUT4 add_5284_6_lut (.I0(GND_net), .I1(n16530[3]), .I2(n384), .I3(n45036), 
            .O(n15953[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5284_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_i365_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n542_adj_5340));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i365_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i369_2_lut (.I0(\Kp[7] ), .I1(n1[12]), .I2(GND_net), 
            .I3(GND_net), .O(n548_adj_5339));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i369_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5070_16_lut (.I0(GND_net), .I1(n12422[13]), .I2(n1099), 
            .I3(n44910), .O(n11404[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5070_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5284_6 (.CI(n45036), .I0(n16530[3]), .I1(n384), .CO(n45037));
    SB_CARRY mult_16_add_1225_2 (.CI(GND_net), .I0(n5), .I1(n74), .CO(n45152));
    SB_LUT4 add_5176_16_lut (.I0(GND_net), .I1(n14585[13]), .I2(n1105), 
            .I3(n45105), .O(n13786[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5176_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5284_5_lut (.I0(GND_net), .I1(n16530[2]), .I2(n311), .I3(n45035), 
            .O(n15953[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5284_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5070_16 (.CI(n44910), .I0(n12422[13]), .I1(n1099), .CO(n44911));
    SB_LUT4 add_5070_15_lut (.I0(GND_net), .I1(n12422[12]), .I2(n1026), 
            .I3(n44909), .O(n11404[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5070_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5070_15 (.CI(n44909), .I0(n12422[12]), .I1(n1026), .CO(n44910));
    SB_LUT4 add_5070_14_lut (.I0(GND_net), .I1(n12422[11]), .I2(n953), 
            .I3(n44908), .O(n11404[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5070_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_i414_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n615_adj_5338));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i414_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i463_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n688_adj_5337));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i463_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5176_16 (.CI(n45105), .I0(n14585[13]), .I1(n1105), .CO(n45106));
    SB_LUT4 mult_16_i418_2_lut (.I0(\Kp[8] ), .I1(n1[12]), .I2(GND_net), 
            .I3(GND_net), .O(n621_adj_5336));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i418_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5284_5 (.CI(n45035), .I0(n16530[2]), .I1(n311), .CO(n45036));
    SB_CARRY add_5070_14 (.CI(n44908), .I0(n12422[11]), .I1(n953), .CO(n44909));
    SB_LUT4 add_5070_13_lut (.I0(GND_net), .I1(n12422[10]), .I2(n880), 
            .I3(n44907), .O(n11404[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5070_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5070_13 (.CI(n44907), .I0(n12422[10]), .I1(n880), .CO(n44908));
    SB_LUT4 mult_17_i130_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [15]), 
            .I2(GND_net), .I3(GND_net), .O(n192));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i130_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i498_2_lut (.I0(\Kp[10] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n740));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i498_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i502_2_lut (.I0(\Kp[10] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n746_adj_5335));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i502_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5284_4_lut (.I0(GND_net), .I1(n16530[1]), .I2(n238_adj_5390), 
            .I3(n45034), .O(n15953[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5284_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5284_4 (.CI(n45034), .I0(n16530[1]), .I1(n238_adj_5390), 
            .CO(n45035));
    SB_LUT4 add_5176_15_lut (.I0(GND_net), .I1(n14585[12]), .I2(n1032), 
            .I3(n45104), .O(n13786[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5176_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5070_12_lut (.I0(GND_net), .I1(n12422[9]), .I2(n807_adj_5391), 
            .I3(n44906), .O(n11404[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5070_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5093_23_lut (.I0(GND_net), .I1(n12905[20]), .I2(GND_net), 
            .I3(n45151), .O(n11935[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5093_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5070_12 (.CI(n44906), .I0(n12422[9]), .I1(n807_adj_5391), 
            .CO(n44907));
    SB_LUT4 add_5284_3_lut (.I0(GND_net), .I1(n16530[0]), .I2(n165), .I3(n45033), 
            .O(n15953[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5284_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5070_11_lut (.I0(GND_net), .I1(n12422[8]), .I2(n734_adj_5392), 
            .I3(n44905), .O(n11404[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5070_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5070_11 (.CI(n44905), .I0(n12422[8]), .I1(n734_adj_5392), 
            .CO(n44906));
    SB_LUT4 add_5070_10_lut (.I0(GND_net), .I1(n12422[7]), .I2(n661), 
            .I3(n44904), .O(n11404[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5070_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_i692_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n1029_adj_4864));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i692_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_20_inv_0_i20_1_lut (.I0(deadband[19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5403[19]));   // verilog/motorControl.v(51[43:52])
    defparam unary_minus_20_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_20_inv_0_i21_1_lut (.I0(deadband[20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5403[20]));   // verilog/motorControl.v(51[43:52])
    defparam unary_minus_20_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_17_i138_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [19]), 
            .I2(GND_net), .I3(GND_net), .O(n204_adj_5389));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i138_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i741_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n1102));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i741_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i512_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n761_adj_5332));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i512_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i179_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [15]), 
            .I2(GND_net), .I3(GND_net), .O(n265));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i179_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_3_lut_4_lut_adj_1691 (.I0(\Kp[2] ), .I1(n1[20]), .I2(n19498[0]), 
            .I3(n43412), .O(n19481[1]));   // verilog/motorControl.v(50[18:24])
    defparam i1_3_lut_4_lut_adj_1691.LUT_INIT = 16'h8778;
    SB_LUT4 unary_minus_20_inv_0_i22_1_lut (.I0(deadband[21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5403[21]));   // verilog/motorControl.v(51[43:52])
    defparam unary_minus_20_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_17_i561_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n834_adj_5330));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i561_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i467_2_lut (.I0(\Kp[9] ), .I1(n1[12]), .I2(GND_net), 
            .I3(GND_net), .O(n694_adj_5329));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i467_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i610_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n907_adj_5328));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i610_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i29328_3_lut_4_lut (.I0(\Kp[2] ), .I1(n1[20]), .I2(n43412), 
            .I3(n19498[0]), .O(n4_adj_5276));   // verilog/motorControl.v(50[18:24])
    defparam i29328_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 mult_17_i181_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [16]), 
            .I2(GND_net), .I3(GND_net), .O(n268));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i181_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i404_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n600));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i404_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i228_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [15]), 
            .I2(GND_net), .I3(GND_net), .O(n338));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i228_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i29315_2_lut_3_lut_4_lut (.I0(\Kp[0] ), .I1(n1[21]), .I2(n1[20]), 
            .I3(\Kp[1] ), .O(n19481[0]));   // verilog/motorControl.v(50[18:24])
    defparam i29315_2_lut_3_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 mult_16_i547_2_lut (.I0(\Kp[11] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n813));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i547_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i659_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n980_adj_5327));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i659_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_20_inv_0_i23_1_lut (.I0(deadband[22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5403[22]));   // verilog/motorControl.v(51[43:52])
    defparam unary_minus_20_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_16_i83_2_lut (.I0(\Kp[1] ), .I1(n1[16]), .I2(GND_net), 
            .I3(GND_net), .O(n122_adj_5325));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i83_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i36_2_lut (.I0(\Kp[0] ), .I1(n1[17]), .I2(GND_net), 
            .I3(GND_net), .O(n53_adj_5324));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i36_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i29317_2_lut_3_lut_4_lut (.I0(\Kp[0] ), .I1(n1[21]), .I2(n1[20]), 
            .I3(\Kp[1] ), .O(n43412));   // verilog/motorControl.v(50[18:24])
    defparam i29317_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 mult_17_i277_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [15]), 
            .I2(GND_net), .I3(GND_net), .O(n411));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i277_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i596_2_lut (.I0(\Kp[12] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n886));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i596_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_20_inv_0_i24_1_lut (.I0(deadband[23]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5403[23]));   // verilog/motorControl.v(51[43:52])
    defparam unary_minus_20_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_14_i3_3_lut (.I0(n130[2]), .I1(n182[2]), .I2(n181), .I3(GND_net), 
            .O(n207[2]));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_14_i3_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_16_i516_2_lut (.I0(\Kp[10] ), .I1(n1[12]), .I2(GND_net), 
            .I3(GND_net), .O(n767_adj_5322));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i516_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i565_2_lut (.I0(\Kp[11] ), .I1(n1[12]), .I2(GND_net), 
            .I3(GND_net), .O(n840_adj_5321));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i565_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i551_2_lut (.I0(\Kp[11] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n819_adj_5320));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i551_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_15_i3_3_lut (.I0(n207[2]), .I1(IntegralLimit[2]), .I2(n155), 
            .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3996 [2]));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_15_i3_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_17_i53_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n77));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i53_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i6_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n8));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i6_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i326_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [15]), 
            .I2(GND_net), .I3(GND_net), .O(n484));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i326_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i102_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n150));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i102_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i132_2_lut (.I0(\Kp[2] ), .I1(n1[16]), .I2(GND_net), 
            .I3(GND_net), .O(n195_adj_5319));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i132_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i29412_3_lut_4_lut (.I0(\Kp[3] ), .I1(n1[18]), .I2(n4_adj_5394), 
            .I3(n19450[1]), .O(n6_adj_5237));   // verilog/motorControl.v(50[18:24])
    defparam i29412_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 mult_16_i645_2_lut (.I0(\Kp[13] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n959));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i645_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i151_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n223));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i151_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_3_lut_4_lut_adj_1692 (.I0(\Kp[3] ), .I1(n1[18]), .I2(n19450[1]), 
            .I3(n4_adj_5394), .O(n19401[2]));   // verilog/motorControl.v(50[18:24])
    defparam i1_3_lut_4_lut_adj_1692.LUT_INIT = 16'h8778;
    SB_LUT4 mult_17_i375_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [15]), 
            .I2(GND_net), .I3(GND_net), .O(n557));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i375_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_3_lut_4_lut_adj_1693 (.I0(\Kp[2] ), .I1(n1[18]), .I2(n19450[0]), 
            .I3(n43494), .O(n19401[1]));   // verilog/motorControl.v(50[18:24])
    defparam i1_3_lut_4_lut_adj_1693.LUT_INIT = 16'h8778;
    SB_LUT4 mult_16_i545_2_lut (.I0(\Kp[11] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n810_adj_5318));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i545_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i600_2_lut (.I0(\Kp[12] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n892_adj_5317));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i600_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i181_2_lut (.I0(\Kp[3] ), .I1(n1[16]), .I2(GND_net), 
            .I3(GND_net), .O(n268_adj_5316));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i181_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut_adj_1694 (.I0(n19490[0]), .I1(n43280), .I2(\Ki[2] ), 
            .I3(\PID_CONTROLLER.integral_23__N_3996 [20]), .O(n19466[1]));   // verilog/motorControl.v(50[27:38])
    defparam i1_4_lut_adj_1694.LUT_INIT = 16'h9666;
    SB_LUT4 unary_minus_26_inv_0_i1_1_lut (.I0(PWMLimit[0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5401[0]));   // verilog/motorControl.v(55[22:31])
    defparam unary_minus_26_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_17_i200_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n296));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i200_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i737_2_lut (.I0(\Kp[15] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n1096_adj_5314));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i737_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i230_2_lut (.I0(\Kp[4] ), .I1(n1[16]), .I2(GND_net), 
            .I3(GND_net), .O(n341_adj_5313));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i230_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i73_2_lut (.I0(\Kp[1] ), .I1(n1[11]), .I2(GND_net), 
            .I3(GND_net), .O(n107_adj_5312));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i73_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i26_2_lut (.I0(\Kp[0] ), .I1(n1[12]), .I2(GND_net), 
            .I3(GND_net), .O(n38_adj_5311));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i26_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i29404_3_lut_4_lut (.I0(\Kp[2] ), .I1(n1[18]), .I2(n43494), 
            .I3(n19450[0]), .O(n4_adj_5394));   // verilog/motorControl.v(50[18:24])
    defparam i29404_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 i29391_2_lut_3_lut_4_lut (.I0(\Kp[0] ), .I1(n1[19]), .I2(n1[18]), 
            .I3(\Kp[1] ), .O(n19401[0]));   // verilog/motorControl.v(50[18:24])
    defparam i29391_2_lut_3_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 i29393_2_lut_3_lut_4_lut (.I0(\Kp[0] ), .I1(n1[19]), .I2(n1[18]), 
            .I3(\Kp[1] ), .O(n43494));   // verilog/motorControl.v(50[18:24])
    defparam i29393_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 mult_17_i89_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [19]), 
            .I2(GND_net), .I3(GND_net), .O(n131_adj_5388));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i89_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i649_2_lut (.I0(\Kp[13] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n965_adj_5310));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i649_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i122_2_lut (.I0(\Kp[2] ), .I1(n1[11]), .I2(GND_net), 
            .I3(GND_net), .O(n180_adj_5309));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i122_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i29366_3_lut_4_lut (.I0(\Kp[3] ), .I1(n1[19]), .I2(n4_adj_5395), 
            .I3(n19481[1]), .O(n6_adj_5275));   // verilog/motorControl.v(50[18:24])
    defparam i29366_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 i1_3_lut_4_lut_adj_1695 (.I0(\Kp[3] ), .I1(n1[19]), .I2(n19481[1]), 
            .I3(n4_adj_5395), .O(n19450[2]));   // verilog/motorControl.v(50[18:24])
    defparam i1_3_lut_4_lut_adj_1695.LUT_INIT = 16'h8778;
    SB_LUT4 mult_16_i279_2_lut (.I0(\Kp[5] ), .I1(n1[16]), .I2(GND_net), 
            .I3(GND_net), .O(n414_adj_5307));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i279_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i42_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [20]), 
            .I2(GND_net), .I3(GND_net), .O(n62_adj_5387));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i42_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_26_inv_0_i2_1_lut (.I0(PWMLimit[1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5401[1]));   // verilog/motorControl.v(55[22:31])
    defparam unary_minus_26_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_16_i594_2_lut (.I0(\Kp[12] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n883_adj_5304));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i594_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_3_lut_4_lut_adj_1696 (.I0(n62), .I1(n131_adj_5246), .I2(n204), 
            .I3(n19481[0]), .O(n19450[1]));   // verilog/motorControl.v(50[18:24])
    defparam i1_3_lut_4_lut_adj_1696.LUT_INIT = 16'h8778;
    SB_LUT4 i29358_3_lut_4_lut (.I0(n62), .I1(n131_adj_5246), .I2(n204), 
            .I3(n19481[0]), .O(n4_adj_5395));   // verilog/motorControl.v(50[18:24])
    defparam i29358_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 unary_minus_26_inv_0_i3_1_lut (.I0(PWMLimit[2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5401[2]));   // verilog/motorControl.v(55[22:31])
    defparam unary_minus_26_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_16_i328_2_lut (.I0(\Kp[6] ), .I1(n1[16]), .I2(GND_net), 
            .I3(GND_net), .O(n487_adj_5302));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i328_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i377_2_lut (.I0(\Kp[7] ), .I1(n1[16]), .I2(GND_net), 
            .I3(GND_net), .O(n560_adj_5300));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i377_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_26_inv_0_i4_1_lut (.I0(PWMLimit[3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5401[3]));   // verilog/motorControl.v(55[22:31])
    defparam unary_minus_26_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_14_i11_3_lut (.I0(n130[10]), .I1(n182[10]), .I2(n181), 
            .I3(GND_net), .O(n207[10]));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_14_i11_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_15_i11_3_lut (.I0(n207[10]), .I1(IntegralLimit[10]), .I2(n155), 
            .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3996 [10]));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_15_i11_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_17_i69_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n101_adj_5298));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i69_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i22_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n32_adj_5297));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i22_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_26_inv_0_i5_1_lut (.I0(PWMLimit[4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5401[4]));   // verilog/motorControl.v(55[22:31])
    defparam unary_minus_26_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_16_i171_2_lut (.I0(\Kp[3] ), .I1(n1[11]), .I2(GND_net), 
            .I3(GND_net), .O(n253_adj_5295));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i171_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i118_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n174_adj_5294));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i118_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i167_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n247_adj_5293));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i167_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i216_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n320_adj_5292));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i216_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i220_2_lut (.I0(\Kp[4] ), .I1(n1[11]), .I2(GND_net), 
            .I3(GND_net), .O(n326_adj_5291));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i220_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i29345_2_lut_4_lut (.I0(\Kp[0] ), .I1(n1[20]), .I2(\Kp[1] ), 
            .I3(n1[19]), .O(n19450[0]));   // verilog/motorControl.v(50[18:24])
    defparam i29345_2_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 mult_16_i643_2_lut (.I0(\Kp[13] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n956_adj_5290));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i643_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i265_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n393_adj_5289));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i265_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_14_i21_3_lut (.I0(n130[20]), .I1(n182[20]), .I2(n181), 
            .I3(GND_net), .O(n207[20]));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_14_i21_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_15_i21_3_lut (.I0(n207[20]), .I1(IntegralLimit[20]), .I2(n155), 
            .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3996 [20]));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_15_i21_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_17_i453_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n673));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i453_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_14_i20_3_lut (.I0(n130[19]), .I1(n182[19]), .I2(n181), 
            .I3(GND_net), .O(n207[19]));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_14_i20_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_17_i502_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n746));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i502_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_15_i20_3_lut (.I0(n207[19]), .I1(IntegralLimit[19]), .I2(n155), 
            .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3996 [19]));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_15_i20_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_16_i549_2_lut (.I0(\Kp[11] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n816_adj_5133));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i549_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i551_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n819));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i551_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i230_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [16]), 
            .I2(GND_net), .I3(GND_net), .O(n341_adj_5132));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i230_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_14_i19_3_lut (.I0(n130[18]), .I1(n182[18]), .I2(n181), 
            .I3(GND_net), .O(n207[18]));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_14_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_15_i19_3_lut (.I0(n207[18]), .I1(IntegralLimit[18]), .I2(n155), 
            .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3996 [18]));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_15_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_14_i22_3_lut (.I0(n130[21]), .I1(n182[21]), .I2(n181), 
            .I3(GND_net), .O(n207[21]));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_14_i22_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_17_i600_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n892));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i600_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i279_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [16]), 
            .I2(GND_net), .I3(GND_net), .O(n414));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i279_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_15_i22_3_lut (.I0(n207[21]), .I1(IntegralLimit[21]), .I2(n155), 
            .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3996 [21]));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_15_i22_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_16_i598_2_lut (.I0(\Kp[12] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n889_adj_5130));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i598_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i494_2_lut (.I0(\Kp[10] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n734));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i494_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i649_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n965));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i649_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_14_i24_3_lut (.I0(n130[23]), .I1(n182[23]), .I2(n181), 
            .I3(GND_net), .O(n207[23]));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_14_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_15_i24_3_lut (.I0(n207[23]), .I1(IntegralLimit[23]), .I2(n155), 
            .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3996 [23]));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_15_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_14_i23_3_lut (.I0(n130[22]), .I1(n182[22]), .I2(n181), 
            .I3(GND_net), .O(n207[22]));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_14_i23_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_15_i23_3_lut (.I0(n207[22]), .I1(IntegralLimit[22]), .I2(n155), 
            .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3996 [22]));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_15_i23_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_17_i330_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [17]), 
            .I2(GND_net), .I3(GND_net), .O(n490_adj_5265));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i330_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut_adj_1697 (.I0(\Ki[1] ), .I1(\Ki[0] ), .I2(\PID_CONTROLLER.integral_23__N_3996 [22]), 
            .I3(\PID_CONTROLLER.integral_23__N_3996 [23]), .O(n52300));   // verilog/motorControl.v(50[27:38])
    defparam i1_4_lut_adj_1697.LUT_INIT = 16'h93a0;
    SB_LUT4 i1_4_lut_adj_1698 (.I0(\Ki[5] ), .I1(\Ki[4] ), .I2(\PID_CONTROLLER.integral_23__N_3996 [18]), 
            .I3(\PID_CONTROLLER.integral_23__N_3996 [19]), .O(n52304));   // verilog/motorControl.v(50[27:38])
    defparam i1_4_lut_adj_1698.LUT_INIT = 16'h6ca0;
    SB_LUT4 i1_4_lut_adj_1699 (.I0(\Ki[3] ), .I1(\Ki[2] ), .I2(\PID_CONTROLLER.integral_23__N_3996 [20]), 
            .I3(\PID_CONTROLLER.integral_23__N_3996 [21]), .O(n52302));   // verilog/motorControl.v(50[27:38])
    defparam i1_4_lut_adj_1699.LUT_INIT = 16'h6ca0;
    SB_LUT4 i1_4_lut_adj_1700 (.I0(n52302), .I1(n43478), .I2(n52304), 
            .I3(n52300), .O(n52310));   // verilog/motorControl.v(50[27:38])
    defparam i1_4_lut_adj_1700.LUT_INIT = 16'h6996;
    SB_LUT4 i29206_4_lut (.I0(n19490[0]), .I1(\Ki[2] ), .I2(n43280), .I3(\PID_CONTROLLER.integral_23__N_3996 [20]), 
            .O(n4_adj_5397));   // verilog/motorControl.v(50[27:38])
    defparam i29206_4_lut.LUT_INIT = 16'he8a0;
    SB_LUT4 i29298_4_lut (.I0(n19426[2]), .I1(\Ki[4] ), .I2(n6_adj_5382), 
            .I3(\PID_CONTROLLER.integral_23__N_3996 [18]), .O(n8_adj_5398));   // verilog/motorControl.v(50[27:38])
    defparam i29298_4_lut.LUT_INIT = 16'he8a0;
    SB_LUT4 i1_4_lut_adj_1701 (.I0(n6_adj_5386), .I1(n8_adj_5398), .I2(n4_adj_5397), 
            .I3(n52310), .O(n51074));   // verilog/motorControl.v(50[27:38])
    defparam i1_4_lut_adj_1701.LUT_INIT = 16'h6996;
    SB_LUT4 mux_14_i16_3_lut (.I0(n130[15]), .I1(n182[15]), .I2(n181), 
            .I3(GND_net), .O(n207[15]));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_14_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_16_i81_2_lut (.I0(\Kp[1] ), .I1(n1[15]), .I2(GND_net), 
            .I3(GND_net), .O(n119_adj_5264));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i81_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_15_i16_3_lut (.I0(n207[15]), .I1(IntegralLimit[15]), .I2(n155), 
            .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3996 [15]));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_15_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_17_i424_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [15]), 
            .I2(GND_net), .I3(GND_net), .O(n630));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i424_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i249_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n369));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i249_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i34_2_lut (.I0(\Kp[0] ), .I1(n1[16]), .I2(GND_net), 
            .I3(GND_net), .O(n50_adj_5263));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i34_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i298_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n442));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i298_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i347_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n515));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i347_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i63_2_lut (.I0(\Kp[1] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n92));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i63_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i130_2_lut (.I0(\Kp[2] ), .I1(n1[15]), .I2(GND_net), 
            .I3(GND_net), .O(n192_adj_5262));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i130_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i16_2_lut (.I0(\Kp[0] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n23));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i16_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i39034_3_lut_4_lut (.I0(deadband[3]), .I1(n356[3]), .I2(n356[2]), 
            .I3(deadband[2]), .O(n54864));   // verilog/motorControl.v(51[12:29])
    defparam i39034_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 LessThan_19_i6_3_lut_3_lut (.I0(deadband[3]), .I1(n356[3]), 
            .I2(n356[2]), .I3(GND_net), .O(n6_adj_5082));   // verilog/motorControl.v(51[12:29])
    defparam LessThan_19_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 mult_16_i694_2_lut (.I0(\Kp[14] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n1032));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i694_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i112_2_lut (.I0(\Kp[2] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n165));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i112_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i128_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [14]), 
            .I2(GND_net), .I3(GND_net), .O(n189_adj_5261));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i128_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i71_2_lut (.I0(\Kp[1] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n104));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i71_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i24_2_lut (.I0(\Kp[0] ), .I1(n1[11]), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_5260));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i24_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i38947_2_lut_4_lut (.I0(deadband[21]), .I1(n356[21]), .I2(deadband[9]), 
            .I3(n356[9]), .O(n54777));
    defparam i38947_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 mult_16_i179_2_lut (.I0(\Kp[3] ), .I1(n1[15]), .I2(GND_net), 
            .I3(GND_net), .O(n265_adj_5259));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i179_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i38854_3_lut_4_lut (.I0(n356[3]), .I1(n436[3]), .I2(n436[2]), 
            .I3(n356[2]), .O(n54684));   // verilog/motorControl.v(54[23:39])
    defparam i38854_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 LessThan_25_i6_3_lut_3_lut (.I0(n356[3]), .I1(n436[3]), .I2(n436[2]), 
            .I3(GND_net), .O(n6_adj_5001));   // verilog/motorControl.v(54[23:39])
    defparam LessThan_25_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 mult_16_i228_2_lut (.I0(\Kp[4] ), .I1(n1[15]), .I2(GND_net), 
            .I3(GND_net), .O(n338_adj_5258));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i228_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i277_2_lut (.I0(\Kp[5] ), .I1(n1[15]), .I2(GND_net), 
            .I3(GND_net), .O(n411_adj_5257));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i277_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i120_2_lut (.I0(\Kp[2] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n177));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i120_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i38996_2_lut_4_lut (.I0(deadband[16]), .I1(n356[16]), .I2(deadband[7]), 
            .I3(n356[7]), .O(n54826));
    defparam i38996_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i38893_3_lut_4_lut (.I0(PWMLimit[3]), .I1(n356[3]), .I2(n356[2]), 
            .I3(PWMLimit[2]), .O(n54723));   // verilog/motorControl.v(52[14:29])
    defparam i38893_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 LessThan_23_i6_3_lut_3_lut (.I0(PWMLimit[3]), .I1(n356[3]), 
            .I2(n356[2]), .I3(GND_net), .O(n6_adj_4946));   // verilog/motorControl.v(52[14:29])
    defparam LessThan_23_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 mult_16_i326_2_lut (.I0(\Kp[6] ), .I1(n1[15]), .I2(GND_net), 
            .I3(GND_net), .O(n484_adj_5256));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i326_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i375_2_lut (.I0(\Kp[7] ), .I1(n1[15]), .I2(GND_net), 
            .I3(GND_net), .O(n557_adj_5255));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i375_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i177_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [14]), 
            .I2(GND_net), .I3(GND_net), .O(n262_adj_5254));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i177_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i169_2_lut (.I0(\Kp[3] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n250));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i169_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i14640_3_lut_4_lut (.I0(control_update), .I1(n409), .I2(n28710), 
            .I3(PWMLimit[0]), .O(n28711));
    defparam i14640_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i14958_3_lut_4_lut (.I0(control_update), .I1(n409), .I2(n29028), 
            .I3(PWMLimit[1]), .O(n29029));
    defparam i14958_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 mult_16_i424_2_lut (.I0(\Kp[8] ), .I1(n1[15]), .I2(GND_net), 
            .I3(GND_net), .O(n630_adj_5253));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i424_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i14848_3_lut_4_lut (.I0(control_update), .I1(n409), .I2(n28918), 
            .I3(PWMLimit[23]), .O(n28919));
    defparam i14848_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i14853_3_lut_4_lut (.I0(control_update), .I1(n409), .I2(n28923), 
            .I3(PWMLimit[22]), .O(n28924));
    defparam i14853_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i14858_3_lut_4_lut (.I0(control_update), .I1(n409), .I2(n28928), 
            .I3(PWMLimit[21]), .O(n28929));
    defparam i14858_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i14863_3_lut_4_lut (.I0(control_update), .I1(n409), .I2(n28933), 
            .I3(PWMLimit[20]), .O(n28934));
    defparam i14863_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i14868_3_lut_4_lut (.I0(control_update), .I1(n409), .I2(n28938), 
            .I3(PWMLimit[19]), .O(n28939));
    defparam i14868_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i14873_3_lut_4_lut (.I0(control_update), .I1(n409), .I2(n28943), 
            .I3(PWMLimit[18]), .O(n28944));
    defparam i14873_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i14878_3_lut_4_lut (.I0(control_update), .I1(n409), .I2(n28948), 
            .I3(PWMLimit[17]), .O(n28949));
    defparam i14878_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i14883_3_lut_4_lut (.I0(control_update), .I1(n409), .I2(n28953), 
            .I3(PWMLimit[16]), .O(n28954));
    defparam i14883_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 mux_14_i9_3_lut (.I0(n130[8]), .I1(n182[8]), .I2(n181), .I3(GND_net), 
            .O(n207[8]));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_14_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14888_3_lut_4_lut (.I0(control_update), .I1(n409), .I2(n28958), 
            .I3(PWMLimit[15]), .O(n28959));
    defparam i14888_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i14893_3_lut_4_lut (.I0(control_update), .I1(n409), .I2(n28963), 
            .I3(PWMLimit[14]), .O(n28964));
    defparam i14893_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i14898_3_lut_4_lut (.I0(control_update), .I1(n409), .I2(n28968), 
            .I3(PWMLimit[13]), .O(n28969));
    defparam i14898_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i14903_3_lut_4_lut (.I0(control_update), .I1(n409), .I2(n28973), 
            .I3(PWMLimit[12]), .O(n28974));
    defparam i14903_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 mux_15_i9_3_lut (.I0(n207[8]), .I1(IntegralLimit[8]), .I2(n155), 
            .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3996 [8]));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_15_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14908_3_lut_4_lut (.I0(control_update), .I1(n409), .I2(n28978), 
            .I3(PWMLimit[11]), .O(n28979));
    defparam i14908_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 mult_17_i65_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n95_adj_5252));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i65_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i18_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n26_adj_5251));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i18_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i14913_3_lut_4_lut (.I0(control_update), .I1(n409), .I2(n28983), 
            .I3(PWMLimit[10]), .O(n28984));
    defparam i14913_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 mult_16_i218_2_lut (.I0(\Kp[4] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n323));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i218_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i114_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n168_adj_5250));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i114_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i267_2_lut (.I0(\Kp[5] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n396_adj_5249));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i267_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i14918_3_lut_4_lut (.I0(control_update), .I1(n409), .I2(n28988), 
            .I3(PWMLimit[9]), .O(n28989));
    defparam i14918_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 mult_17_i226_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [14]), 
            .I2(GND_net), .I3(GND_net), .O(n335_adj_5248));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i226_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i14923_3_lut_4_lut (.I0(control_update), .I1(n409), .I2(n28993), 
            .I3(PWMLimit[8]), .O(n28994));
    defparam i14923_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i14928_3_lut_4_lut (.I0(control_update), .I1(n409), .I2(n28998), 
            .I3(PWMLimit[7]), .O(n28999));
    defparam i14928_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i14933_3_lut_4_lut (.I0(control_update), .I1(n409), .I2(n29003), 
            .I3(PWMLimit[6]), .O(n29004));
    defparam i14933_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i14938_3_lut_4_lut (.I0(control_update), .I1(n409), .I2(n29008), 
            .I3(PWMLimit[5]), .O(n29009));
    defparam i14938_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i14943_3_lut_4_lut (.I0(control_update), .I1(n409), .I2(n29013), 
            .I3(PWMLimit[4]), .O(n29014));
    defparam i14943_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 mult_17_i275_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [14]), 
            .I2(GND_net), .I3(GND_net), .O(n408_adj_5247));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i275_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i14948_3_lut_4_lut (.I0(control_update), .I1(n409), .I2(n29018), 
            .I3(PWMLimit[3]), .O(n29019));
    defparam i14948_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i14953_3_lut_4_lut (.I0(control_update), .I1(n409), .I2(n29023), 
            .I3(PWMLimit[2]), .O(n29024));
    defparam i14953_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 mult_17_i163_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n241_adj_5245));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i163_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i698_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n1038_adj_5129));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i698_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i328_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [16]), 
            .I2(GND_net), .I3(GND_net), .O(n487));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i328_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i212_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n314_adj_5244));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i212_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i316_2_lut (.I0(\Kp[6] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n469));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i316_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i261_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n387_adj_5243));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i261_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i310_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n460_adj_5242));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i310_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i365_2_lut (.I0(\Kp[7] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n542));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i365_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i359_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n533_adj_5241));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i359_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i39036_2_lut_4_lut (.I0(n130[21]), .I1(n182[21]), .I2(n130[9]), 
            .I3(n182[9]), .O(n54866));
    defparam i39036_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 mult_17_i324_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [14]), 
            .I2(GND_net), .I3(GND_net), .O(n481_adj_5240));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i324_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i38814_2_lut_4_lut (.I0(n356[21]), .I1(n436[21]), .I2(n356[9]), 
            .I3(n436[9]), .O(n54644));
    defparam i38814_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 mult_17_i408_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n606_adj_5239));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i408_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i457_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n679_adj_5238));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i457_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i506_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n752_adj_5236));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i506_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i414_2_lut (.I0(\Kp[8] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n615));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i414_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i555_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n825_adj_5235));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i555_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i463_2_lut (.I0(\Kp[9] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n688));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i463_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i38826_2_lut_4_lut (.I0(n356[16]), .I1(n436[16]), .I2(n356[7]), 
            .I3(n436[7]), .O(n54656));
    defparam i38826_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i39046_2_lut_4_lut (.I0(n130[16]), .I1(n182[16]), .I2(n130[7]), 
            .I3(n182[7]), .O(n54876));
    defparam i39046_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 mult_17_i747_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n1111_adj_5109));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i747_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i604_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n898_adj_5233));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i604_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i377_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [16]), 
            .I2(GND_net), .I3(GND_net), .O(n560));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i377_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i373_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [14]), 
            .I2(GND_net), .I3(GND_net), .O(n554_adj_5232));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i373_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i653_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n971_adj_5231));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i653_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i38856_2_lut_4_lut (.I0(PWMLimit[21]), .I1(n356[21]), .I2(PWMLimit[9]), 
            .I3(n356[9]), .O(n54686));
    defparam i38856_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 mult_16_i512_2_lut (.I0(\Kp[10] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n761));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i512_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i38868_2_lut_4_lut (.I0(PWMLimit[16]), .I1(n356[16]), .I2(PWMLimit[7]), 
            .I3(n356[7]), .O(n54698));
    defparam i38868_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 mult_17_i702_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n1044_adj_5229));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i702_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i751_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n1117_adj_5227));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i751_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i422_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [14]), 
            .I2(GND_net), .I3(GND_net), .O(n627_adj_5224));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i422_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_14_i8_3_lut (.I0(n130[7]), .I1(n182[7]), .I2(n181), .I3(GND_net), 
            .O(n207[7]));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_14_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_15_i8_3_lut (.I0(n207[7]), .I1(IntegralLimit[7]), .I2(n155), 
            .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3996 [7]));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_15_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_17_i63_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n92_adj_5223));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i63_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i16_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_5222));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i16_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i561_2_lut (.I0(\Kp[11] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n834));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i561_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i39072_2_lut_4_lut (.I0(IntegralLimit[21]), .I1(n130[21]), .I2(IntegralLimit[9]), 
            .I3(n130[9]), .O(n54902));
    defparam i39072_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 mult_16_i610_2_lut (.I0(\Kp[12] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n907));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i610_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i471_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [14]), 
            .I2(GND_net), .I3(GND_net), .O(n700_adj_5219));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i471_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i39082_2_lut_4_lut (.I0(IntegralLimit[16]), .I1(n130[16]), .I2(IntegralLimit[7]), 
            .I3(n130[7]), .O(n54912));
    defparam i39082_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 mult_17_i112_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n165_adj_5218));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i112_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_14_i6_3_lut (.I0(n130[5]), .I1(n182[5]), .I2(n181), .I3(GND_net), 
            .O(n207[5]));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_14_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_15_i6_3_lut (.I0(n207[5]), .I1(IntegralLimit[5]), .I2(n155), 
            .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3996 [5]));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_15_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_17_i161_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n238));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i161_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i59_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n86));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i59_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i12_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_5091));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i12_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i659_2_lut (.I0(\Kp[13] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n980));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i659_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i67_2_lut (.I0(\Kp[1] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n98_adj_5087));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i67_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i20_2_lut (.I0(\Kp[0] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_5086));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i20_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i210_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n311_adj_5217));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i210_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i108_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n159_adj_5085));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i108_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i59_2_lut (.I0(\Kp[1] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n86_adj_5216));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i59_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_10_i9_2_lut (.I0(IntegralLimit[4]), .I1(n130[4]), .I2(GND_net), 
            .I3(GND_net), .O(n9_adj_4903));   // verilog/motorControl.v(45[12:34])
    defparam LessThan_10_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_16_i12_2_lut (.I0(\Kp[0] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_5215));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i12_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i69_2_lut (.I0(\Kp[1] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n101));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i69_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_10_i11_2_lut (.I0(IntegralLimit[5]), .I1(n130[5]), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_4906));   // verilog/motorControl.v(45[12:34])
    defparam LessThan_10_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_10_i13_2_lut (.I0(IntegralLimit[6]), .I1(n130[6]), 
            .I2(GND_net), .I3(GND_net), .O(n13_adj_4905));   // verilog/motorControl.v(45[12:34])
    defparam LessThan_10_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_17_i157_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n232_adj_5081));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i157_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i22_2_lut (.I0(\Kp[0] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n32));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i22_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_10_i15_2_lut (.I0(IntegralLimit[7]), .I1(n130[7]), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_4904));   // verilog/motorControl.v(45[12:34])
    defparam LessThan_10_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_16_i116_2_lut (.I0(\Kp[2] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n171_adj_5079));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i116_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_10_i21_2_lut (.I0(IntegralLimit[10]), .I1(n130[10]), 
            .I2(GND_net), .I3(GND_net), .O(n21));   // verilog/motorControl.v(45[12:34])
    defparam LessThan_10_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_16_i53_2_lut (.I0(\Kp[1] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n77_adj_5213));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i53_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_10_i19_2_lut (.I0(IntegralLimit[9]), .I1(n130[9]), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_4901));   // verilog/motorControl.v(45[12:34])
    defparam LessThan_10_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_16_i165_2_lut (.I0(\Kp[3] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n244_adj_5078));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i165_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_10_i17_2_lut (.I0(IntegralLimit[8]), .I1(n130[8]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_4902));   // verilog/motorControl.v(45[12:34])
    defparam LessThan_10_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_16_i647_2_lut (.I0(\Kp[13] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n962_adj_5076));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i647_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i543_2_lut (.I0(\Kp[11] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n807));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i543_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_10_i23_2_lut (.I0(IntegralLimit[11]), .I1(n130[11]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_4912));   // verilog/motorControl.v(45[12:34])
    defparam LessThan_10_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_10_i25_2_lut (.I0(IntegralLimit[12]), .I1(n130[12]), 
            .I2(GND_net), .I3(GND_net), .O(n25));   // verilog/motorControl.v(45[12:34])
    defparam LessThan_10_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_12_i9_2_lut (.I0(n130[4]), .I1(n182[4]), .I2(GND_net), 
            .I3(GND_net), .O(n9_adj_4966));   // verilog/motorControl.v(47[21:44])
    defparam LessThan_12_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_12_i11_2_lut (.I0(n130[5]), .I1(n182[5]), .I2(GND_net), 
            .I3(GND_net), .O(n11_adj_4973));   // verilog/motorControl.v(47[21:44])
    defparam LessThan_12_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_12_i13_2_lut (.I0(n130[6]), .I1(n182[6]), .I2(GND_net), 
            .I3(GND_net), .O(n13_adj_4972));   // verilog/motorControl.v(47[21:44])
    defparam LessThan_12_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_12_i15_2_lut (.I0(n130[7]), .I1(n182[7]), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_4971));   // verilog/motorControl.v(47[21:44])
    defparam LessThan_12_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_12_i21_2_lut (.I0(n130[10]), .I1(n182[10]), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_4963));   // verilog/motorControl.v(47[21:44])
    defparam LessThan_12_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_12_i19_2_lut (.I0(n130[9]), .I1(n182[9]), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_4964));   // verilog/motorControl.v(47[21:44])
    defparam LessThan_12_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_12_i17_2_lut (.I0(n130[8]), .I1(n182[8]), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_4965));   // verilog/motorControl.v(47[21:44])
    defparam LessThan_12_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_12_i23_2_lut (.I0(n130[11]), .I1(n182[11]), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_4992));   // verilog/motorControl.v(47[21:44])
    defparam LessThan_12_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_12_i25_2_lut (.I0(n130[12]), .I1(n182[12]), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_4991));   // verilog/motorControl.v(47[21:44])
    defparam LessThan_12_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_16_i6_2_lut (.I0(\Kp[0] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n8_adj_5212));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i6_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i118_2_lut (.I0(\Kp[2] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n174));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i118_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i206_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n305_adj_5074));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i206_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i255_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n378_adj_5072));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i255_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i259_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n384_adj_5207));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i259_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i304_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n451_adj_5068));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i304_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i214_2_lut (.I0(\Kp[4] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n317_adj_5065));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i214_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i353_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n524));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i353_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i308_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n457_adj_5202));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i308_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i402_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n597));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i402_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i696_2_lut (.I0(\Kp[14] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n1035_adj_5059));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i696_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i263_2_lut (.I0(\Kp[5] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n390_adj_5058));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i263_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i451_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n670));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i451_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i500_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n743));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i500_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i549_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n816));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i549_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i312_2_lut (.I0(\Kp[6] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n463_adj_5051));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i312_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i745_2_lut (.I0(\Kp[15] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n1108_adj_5050));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i745_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i361_2_lut (.I0(\Kp[7] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n536_adj_5049));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i361_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i598_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n889));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i598_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i410_2_lut (.I0(\Kp[8] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n609));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i410_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i647_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n962));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i647_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i592_2_lut (.I0(\Kp[12] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n880_adj_5041));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i592_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i696_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n1035));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i696_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i745_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n1108));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i745_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i459_2_lut (.I0(\Kp[9] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n682));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i459_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i508_2_lut (.I0(\Kp[10] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n755));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i508_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i641_2_lut (.I0(\Kp[13] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n953_adj_5027));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i641_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i494_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n734_adj_5392));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i494_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i543_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n807_adj_5391));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i543_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i161_2_lut (.I0(\Kp[3] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n238_adj_5390));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i161_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i269_2_lut (.I0(\Kp[5] ), .I1(n1[11]), .I2(GND_net), 
            .I3(GND_net), .O(n399_adj_5288));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i269_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i77_2_lut (.I0(\Kp[1] ), .I1(n1[13]), .I2(GND_net), 
            .I3(GND_net), .O(n113));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i77_2_lut.LUT_INIT = 16'h8888;
    
endmodule
//
// Verilog Description of module EEPROM
//

module EEPROM (\state[3] , n6, GND_net, clk16MHz, read, \state[0] , 
            enable_slow_N_4393, n6271, \state[1] , n48526, VCC_net, 
            n48558, n29393, rw, n48670, data_ready, n36659, n49838, 
            n49919, \state_7__N_4290[0] , n4, n4_adj_18, n36542, n7354, 
            \state[2] , n26, \state_7__N_4306[3] , n7936, scl_enable, 
            \saved_addr[0] , \state[0]_adj_19 , n29452, sda_enable, 
            n29364, data, n29363, n29362, n29361, n29360, n29359, 
            n29358, n10, n10_adj_20, n8, n29835, n54609, n27243, 
            n27238, scl, sda_out) /* synthesis syn_noprune=1, syn_module_defined=1 */ ;
    output \state[3] ;
    output n6;
    input GND_net;
    input clk16MHz;
    input read;
    output \state[0] ;
    output enable_slow_N_4393;
    output [0:0]n6271;
    output \state[1] ;
    input n48526;
    input VCC_net;
    input n48558;
    input n29393;
    output rw;
    input n48670;
    output data_ready;
    output n36659;
    input n49838;
    output n49919;
    output \state_7__N_4290[0] ;
    output n4;
    output n4_adj_18;
    output n36542;
    output n7354;
    output \state[2] ;
    output n26;
    input \state_7__N_4306[3] ;
    input n7936;
    output scl_enable;
    output \saved_addr[0] ;
    output \state[0]_adj_19 ;
    input n29452;
    output sda_enable;
    input n29364;
    output [7:0]data;
    input n29363;
    input n29362;
    input n29361;
    input n29360;
    input n29359;
    input n29358;
    output n10;
    output n10_adj_20;
    input n8;
    input n29835;
    output n54609;
    output n27243;
    output n27238;
    output scl;
    output sda_out;
    
    wire clk16MHz /* synthesis SET_AS_NETWORK=clk16MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    
    wire n27106;
    wire [15:0]delay_counter_15__N_4192;
    
    wire n28916;
    wire [15:0]delay_counter;   // verilog/eeprom.v(24[12:25])
    
    wire n29315, n28, n26_c, n27, n25, enable;
    wire [15:0]n4876;
    
    wire n43809, n43808, n43807, n43806, n43805, n43804, n43803, 
        n43802, n43801, n43800, n43799, n43798, n43797, n43796, 
        n43795;
    
    SB_LUT4 i2_2_lut (.I0(\state[3] ), .I1(n27106), .I2(GND_net), .I3(GND_net), 
            .O(n6));   // verilog/eeprom.v(42[12:28])
    defparam i2_2_lut.LUT_INIT = 16'heeee;
    SB_DFFESR delay_counter_i0_i1 (.Q(delay_counter[1]), .C(clk16MHz), .E(n28916), 
            .D(delay_counter_15__N_4192[1]), .R(n29315));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFFESR delay_counter_i0_i2 (.Q(delay_counter[2]), .C(clk16MHz), .E(n28916), 
            .D(delay_counter_15__N_4192[2]), .R(n29315));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFFESR delay_counter_i0_i3 (.Q(delay_counter[3]), .C(clk16MHz), .E(n28916), 
            .D(delay_counter_15__N_4192[3]), .R(n29315));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFFESS delay_counter_i0_i4 (.Q(delay_counter[4]), .C(clk16MHz), .E(n28916), 
            .D(delay_counter_15__N_4192[4]), .S(n29315));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFFESR delay_counter_i0_i5 (.Q(delay_counter[5]), .C(clk16MHz), .E(n28916), 
            .D(delay_counter_15__N_4192[5]), .R(n29315));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFFESS delay_counter_i0_i6 (.Q(delay_counter[6]), .C(clk16MHz), .E(n28916), 
            .D(delay_counter_15__N_4192[6]), .S(n29315));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFFESS delay_counter_i0_i7 (.Q(delay_counter[7]), .C(clk16MHz), .E(n28916), 
            .D(delay_counter_15__N_4192[7]), .S(n29315));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFFESS delay_counter_i0_i8 (.Q(delay_counter[8]), .C(clk16MHz), .E(n28916), 
            .D(delay_counter_15__N_4192[8]), .S(n29315));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFFESS delay_counter_i0_i9 (.Q(delay_counter[9]), .C(clk16MHz), .E(n28916), 
            .D(delay_counter_15__N_4192[9]), .S(n29315));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFFESS delay_counter_i0_i10 (.Q(delay_counter[10]), .C(clk16MHz), 
            .E(n28916), .D(delay_counter_15__N_4192[10]), .S(n29315));   // verilog/eeprom.v(26[8] 58[4])
    SB_LUT4 i12_4_lut (.I0(delay_counter[6]), .I1(delay_counter[10]), .I2(delay_counter[12]), 
            .I3(delay_counter[8]), .O(n28));   // verilog/eeprom.v(42[12:28])
    defparam i12_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i10_4_lut (.I0(delay_counter[11]), .I1(delay_counter[2]), .I2(delay_counter[7]), 
            .I3(delay_counter[5]), .O(n26_c));   // verilog/eeprom.v(42[12:28])
    defparam i10_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i11_4_lut (.I0(delay_counter[15]), .I1(delay_counter[3]), .I2(delay_counter[14]), 
            .I3(delay_counter[1]), .O(n27));   // verilog/eeprom.v(42[12:28])
    defparam i11_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i9_4_lut (.I0(delay_counter[4]), .I1(delay_counter[9]), .I2(delay_counter[13]), 
            .I3(delay_counter[0]), .O(n25));   // verilog/eeprom.v(42[12:28])
    defparam i9_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut (.I0(n25), .I1(n27), .I2(n26_c), .I3(n28), .O(n27106));   // verilog/eeprom.v(42[12:28])
    defparam i15_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 mux_1487_Mux_0_i1_4_lut (.I0(read), .I1(n27106), .I2(\state[0] ), 
            .I3(enable_slow_N_4393), .O(n6271[0]));   // verilog/eeprom.v(29[3] 57[10])
    defparam mux_1487_Mux_0_i1_4_lut.LUT_INIT = 16'h0a3a;
    SB_DFFESR delay_counter_i0_i11 (.Q(delay_counter[11]), .C(clk16MHz), 
            .E(n28916), .D(delay_counter_15__N_4192[11]), .R(n29315));   // verilog/eeprom.v(26[8] 58[4])
    SB_LUT4 i15248_2_lut (.I0(n28916), .I1(\state[0] ), .I2(GND_net), 
            .I3(GND_net), .O(n29315));   // verilog/eeprom.v(26[8] 58[4])
    defparam i15248_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1_3_lut (.I0(read), .I1(\state[1] ), .I2(\state[0] ), .I3(GND_net), 
            .O(n28916));
    defparam i1_3_lut.LUT_INIT = 16'h3232;
    SB_DFFESR delay_counter_i0_i12 (.Q(delay_counter[12]), .C(clk16MHz), 
            .E(n28916), .D(delay_counter_15__N_4192[12]), .R(n29315));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFFSR enable_39 (.Q(enable), .C(clk16MHz), .D(n6271[0]), .R(\state[1] ));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFFESR delay_counter_i0_i13 (.Q(delay_counter[13]), .C(clk16MHz), 
            .E(n28916), .D(delay_counter_15__N_4192[13]), .R(n29315));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFFESR delay_counter_i0_i14 (.Q(delay_counter[14]), .C(clk16MHz), 
            .E(n28916), .D(delay_counter_15__N_4192[14]), .R(n29315));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFFESR delay_counter_i0_i15 (.Q(delay_counter[15]), .C(clk16MHz), 
            .E(n28916), .D(delay_counter_15__N_4192[15]), .R(n29315));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFFE state__i1 (.Q(\state[1] ), .C(clk16MHz), .E(VCC_net), .D(n48526));   // verilog/eeprom.v(26[8] 58[4])
    SB_LUT4 i40080_2_lut (.I0(n27106), .I1(enable_slow_N_4393), .I2(GND_net), 
            .I3(GND_net), .O(n4876[4]));   // verilog/eeprom.v(46[18] 48[12])
    defparam i40080_2_lut.LUT_INIT = 16'h2222;
    SB_DFF state__i0 (.Q(\state[0] ), .C(clk16MHz), .D(n48558));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFFESR delay_counter_i0_i0 (.Q(delay_counter[0]), .C(clk16MHz), .E(n28916), 
            .D(delay_counter_15__N_4192[0]), .R(n29315));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFF rw_43 (.Q(rw), .C(clk16MHz), .D(n29393));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFF data_ready_42 (.Q(data_ready), .C(clk16MHz), .D(n48670));   // verilog/eeprom.v(26[8] 58[4])
    SB_LUT4 i22595_2_lut_3_lut (.I0(\state[0] ), .I1(\state[1] ), .I2(enable_slow_N_4393), 
            .I3(GND_net), .O(n36659));   // verilog/eeprom.v(51[5:9])
    defparam i22595_2_lut_3_lut.LUT_INIT = 16'hfbfb;
    SB_LUT4 i34160_4_lut_4_lut (.I0(\state[0] ), .I1(\state[1] ), .I2(n49838), 
            .I3(enable_slow_N_4393), .O(n49919));   // verilog/eeprom.v(51[5:9])
    defparam i34160_4_lut_4_lut.LUT_INIT = 16'hfcf8;
    SB_LUT4 add_1035_17_lut (.I0(GND_net), .I1(delay_counter[15]), .I2(n4876[4]), 
            .I3(n43809), .O(delay_counter_15__N_4192[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1035_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_1035_16_lut (.I0(GND_net), .I1(delay_counter[14]), .I2(n4876[4]), 
            .I3(n43808), .O(delay_counter_15__N_4192[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1035_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1035_16 (.CI(n43808), .I0(delay_counter[14]), .I1(n4876[4]), 
            .CO(n43809));
    SB_LUT4 add_1035_15_lut (.I0(GND_net), .I1(delay_counter[13]), .I2(n4876[4]), 
            .I3(n43807), .O(delay_counter_15__N_4192[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1035_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1035_15 (.CI(n43807), .I0(delay_counter[13]), .I1(n4876[4]), 
            .CO(n43808));
    SB_LUT4 add_1035_14_lut (.I0(GND_net), .I1(delay_counter[12]), .I2(n4876[4]), 
            .I3(n43806), .O(delay_counter_15__N_4192[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1035_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1035_14 (.CI(n43806), .I0(delay_counter[12]), .I1(n4876[4]), 
            .CO(n43807));
    SB_LUT4 add_1035_13_lut (.I0(GND_net), .I1(delay_counter[11]), .I2(n4876[4]), 
            .I3(n43805), .O(delay_counter_15__N_4192[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1035_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1035_13 (.CI(n43805), .I0(delay_counter[11]), .I1(n4876[4]), 
            .CO(n43806));
    SB_LUT4 add_1035_12_lut (.I0(GND_net), .I1(delay_counter[10]), .I2(n4876[4]), 
            .I3(n43804), .O(delay_counter_15__N_4192[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1035_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1035_12 (.CI(n43804), .I0(delay_counter[10]), .I1(n4876[4]), 
            .CO(n43805));
    SB_LUT4 add_1035_11_lut (.I0(GND_net), .I1(delay_counter[9]), .I2(n4876[4]), 
            .I3(n43803), .O(delay_counter_15__N_4192[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1035_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1035_11 (.CI(n43803), .I0(delay_counter[9]), .I1(n4876[4]), 
            .CO(n43804));
    SB_LUT4 add_1035_10_lut (.I0(GND_net), .I1(delay_counter[8]), .I2(n4876[4]), 
            .I3(n43802), .O(delay_counter_15__N_4192[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1035_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1035_10 (.CI(n43802), .I0(delay_counter[8]), .I1(n4876[4]), 
            .CO(n43803));
    SB_LUT4 add_1035_9_lut (.I0(GND_net), .I1(delay_counter[7]), .I2(n4876[4]), 
            .I3(n43801), .O(delay_counter_15__N_4192[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1035_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1035_9 (.CI(n43801), .I0(delay_counter[7]), .I1(n4876[4]), 
            .CO(n43802));
    SB_LUT4 add_1035_8_lut (.I0(GND_net), .I1(delay_counter[6]), .I2(n4876[4]), 
            .I3(n43800), .O(delay_counter_15__N_4192[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1035_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1035_8 (.CI(n43800), .I0(delay_counter[6]), .I1(n4876[4]), 
            .CO(n43801));
    SB_LUT4 add_1035_7_lut (.I0(GND_net), .I1(delay_counter[5]), .I2(n4876[4]), 
            .I3(n43799), .O(delay_counter_15__N_4192[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1035_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1035_7 (.CI(n43799), .I0(delay_counter[5]), .I1(n4876[4]), 
            .CO(n43800));
    SB_LUT4 add_1035_6_lut (.I0(GND_net), .I1(delay_counter[4]), .I2(n4876[4]), 
            .I3(n43798), .O(delay_counter_15__N_4192[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1035_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1035_6 (.CI(n43798), .I0(delay_counter[4]), .I1(n4876[4]), 
            .CO(n43799));
    SB_LUT4 add_1035_5_lut (.I0(GND_net), .I1(delay_counter[3]), .I2(n4876[4]), 
            .I3(n43797), .O(delay_counter_15__N_4192[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1035_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1035_5 (.CI(n43797), .I0(delay_counter[3]), .I1(n4876[4]), 
            .CO(n43798));
    SB_LUT4 add_1035_4_lut (.I0(GND_net), .I1(delay_counter[2]), .I2(n4876[4]), 
            .I3(n43796), .O(delay_counter_15__N_4192[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1035_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1035_4 (.CI(n43796), .I0(delay_counter[2]), .I1(n4876[4]), 
            .CO(n43797));
    SB_LUT4 add_1035_3_lut (.I0(GND_net), .I1(delay_counter[1]), .I2(n4876[4]), 
            .I3(n43795), .O(delay_counter_15__N_4192[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1035_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1035_3 (.CI(n43795), .I0(delay_counter[1]), .I1(n4876[4]), 
            .CO(n43796));
    SB_LUT4 add_1035_2_lut (.I0(GND_net), .I1(delay_counter[0]), .I2(n4876[4]), 
            .I3(GND_net), .O(delay_counter_15__N_4192[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1035_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1035_2 (.CI(GND_net), .I0(delay_counter[0]), .I1(n4876[4]), 
            .CO(n43795));
    i2c_controller i2c (.\state_7__N_4290[0] (\state_7__N_4290[0] ), .enable_slow_N_4393(enable_slow_N_4393), 
            .GND_net(GND_net), .n4(n4), .n4_adj_16(n4_adj_18), .n36542(n36542), 
            .n7354(n7354), .\state[2] (\state[2] ), .\state[3] (\state[3] ), 
            .n26(n26), .\state_7__N_4306[3] (\state_7__N_4306[3] ), .n7936(n7936), 
            .clk16MHz(clk16MHz), .scl_enable(scl_enable), .\saved_addr[0] (\saved_addr[0] ), 
            .\state[0] (\state[0]_adj_19 ), .n29452(n29452), .VCC_net(VCC_net), 
            .sda_enable(sda_enable), .n29364(n29364), .data({data}), .n29363(n29363), 
            .n29362(n29362), .n29361(n29361), .n29360(n29360), .n29359(n29359), 
            .n29358(n29358), .n10(n10), .enable(enable), .n10_adj_17(n10_adj_20), 
            .n8(n8), .n29835(n29835), .n54609(n54609), .n27243(n27243), 
            .n27238(n27238), .scl(scl), .sda_out(sda_out)) /* synthesis syn_noprune=1, syn_module_defined=1 */ ;   // verilog/eeprom.v(60[16] 74[4])
    
endmodule
//
// Verilog Description of module i2c_controller
//

module i2c_controller (\state_7__N_4290[0] , enable_slow_N_4393, GND_net, 
            n4, n4_adj_16, n36542, n7354, \state[2] , \state[3] , 
            n26, \state_7__N_4306[3] , n7936, clk16MHz, scl_enable, 
            \saved_addr[0] , \state[0] , n29452, VCC_net, sda_enable, 
            n29364, data, n29363, n29362, n29361, n29360, n29359, 
            n29358, n10, enable, n10_adj_17, n8, n29835, n54609, 
            n27243, n27238, scl, sda_out) /* synthesis syn_noprune=1, syn_module_defined=1 */ ;
    output \state_7__N_4290[0] ;
    output enable_slow_N_4393;
    input GND_net;
    output n4;
    output n4_adj_16;
    output n36542;
    output n7354;
    output \state[2] ;
    output \state[3] ;
    output n26;
    input \state_7__N_4306[3] ;
    input n7936;
    input clk16MHz;
    output scl_enable;
    output \saved_addr[0] ;
    output \state[0] ;
    input n29452;
    input VCC_net;
    output sda_enable;
    input n29364;
    output [7:0]data;
    input n29363;
    input n29362;
    input n29361;
    input n29360;
    input n29359;
    input n29358;
    output n10;
    input enable;
    output n10_adj_17;
    input n8;
    input n29835;
    output n54609;
    output n27243;
    output n27238;
    output scl;
    output sda_out;
    
    wire i2c_clk /* synthesis is_clock=1, SET_AS_NETWORK=\eeprom/i2c/i2c_clk */ ;   // verilog/i2c_controller.v(41[6:13])
    wire clk16MHz /* synthesis SET_AS_NETWORK=clk16MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    
    wire enable_slow_N_4392;
    wire [7:0]counter;   // verilog/i2c_controller.v(36[12:19])
    
    wire n5;
    wire [7:0]state;   // verilog/i2c_controller.v(33[12:17])
    
    wire n37252, n36727, n36761, n48720, n51358;
    wire [7:0]counter2;   // verilog/i2c_controller.v(37[12:20])
    
    wire n10_c, n29177, i2c_clk_N_4379;
    wire [7:0]n119;
    
    wire n28838, n29228, n15, n49846, n7347, n37, scl_enable_N_4380, 
        n54555, n54527, n11, n54697, n28780;
    wire [5:0]n29;
    
    wire n4_adj_4849, n33_adj_4850, n29171, n7050, n34_adj_4851, n7849, 
        n43961, n43960, n43959, n43958, n43957, n43956, n43955, 
        n19508, n29168, sda_out_adj_4852, n7, n10_adj_4853, n54614, 
        n11_adj_4855, n12, n9, state_7__N_4289, n11_adj_4857, n36445, 
        n11_adj_4858, n11_adj_4859, n44658, n44657, n44656, n44655, 
        n44654;
    
    SB_LUT4 i40104_2_lut (.I0(\state_7__N_4290[0] ), .I1(enable_slow_N_4393), 
            .I2(GND_net), .I3(GND_net), .O(enable_slow_N_4392));   // verilog/i2c_controller.v(62[6:32])
    defparam i40104_2_lut.LUT_INIT = 16'h7777;
    SB_LUT4 equal_385_i4_2_lut (.I0(counter[1]), .I1(counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n4));   // verilog/i2c_controller.v(153[6:23])
    defparam equal_385_i4_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 equal_383_i4_2_lut (.I0(counter[1]), .I1(counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n4_adj_16));   // verilog/i2c_controller.v(153[6:23])
    defparam equal_383_i4_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 i22478_2_lut (.I0(counter[1]), .I1(counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n36542));
    defparam i22478_2_lut.LUT_INIT = 16'h8888;
    SB_DFFESS state_i0_i1 (.Q(state[1]), .C(i2c_clk), .E(n7354), .D(n5), 
            .S(n37252));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESS state_i0_i2 (.Q(\state[2] ), .C(i2c_clk), .E(n7354), .D(n36727), 
            .S(n36761));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESS state_i0_i3 (.Q(\state[3] ), .C(i2c_clk), .E(n7354), .D(n48720), 
            .S(n51358));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_LUT4 i4_4_lut (.I0(counter2[3]), .I1(counter2[5]), .I2(counter2[2]), 
            .I3(counter2[4]), .O(n10_c));
    defparam i4_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i5_3_lut (.I0(counter2[1]), .I1(n10_c), .I2(counter2[0]), 
            .I3(GND_net), .O(n29177));
    defparam i5_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i1_2_lut (.I0(i2c_clk), .I1(n29177), .I2(GND_net), .I3(GND_net), 
            .O(i2c_clk_N_4379));
    defparam i1_2_lut.LUT_INIT = 16'h6666;
    SB_DFFESS counter_i1 (.Q(counter[1]), .C(i2c_clk), .E(n28838), .D(n119[1]), 
            .S(n29228));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESS counter_i2 (.Q(counter[2]), .C(i2c_clk), .E(n28838), .D(n119[2]), 
            .S(n29228));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESR counter_i3 (.Q(counter[3]), .C(i2c_clk), .E(n28838), .D(n119[3]), 
            .R(n29228));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESR counter_i4 (.Q(counter[4]), .C(i2c_clk), .E(n28838), .D(n119[4]), 
            .R(n29228));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESR counter_i5 (.Q(counter[5]), .C(i2c_clk), .E(n28838), .D(n119[5]), 
            .R(n29228));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESR counter_i6 (.Q(counter[6]), .C(i2c_clk), .E(n28838), .D(n119[6]), 
            .R(n29228));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESR counter_i7 (.Q(counter[7]), .C(i2c_clk), .E(n28838), .D(n119[7]), 
            .R(n29228));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_LUT4 i1_2_lut_adj_1670 (.I0(\state[2] ), .I1(state[1]), .I2(GND_net), 
            .I3(GND_net), .O(n26));
    defparam i1_2_lut_adj_1670.LUT_INIT = 16'heeee;
    SB_LUT4 i34094_2_lut (.I0(\state_7__N_4306[3] ), .I1(n15), .I2(GND_net), 
            .I3(GND_net), .O(n49846));
    defparam i34094_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i17_4_lut (.I0(n7347), .I1(n49846), .I2(n7936), .I3(n37), 
            .O(n28838));
    defparam i17_4_lut.LUT_INIT = 16'h3a30;
    SB_DFF i2c_clk_121 (.Q(i2c_clk), .C(clk16MHz), .D(i2c_clk_N_4379));   // verilog/i2c_controller.v(58[9] 71[5])
    SB_DFFN i2c_scl_enable_123 (.Q(scl_enable), .C(i2c_clk), .D(scl_enable_N_4380));   // verilog/i2c_controller.v(76[12] 82[6])
    SB_LUT4 i38853_2_lut (.I0(counter[1]), .I1(\saved_addr[0] ), .I2(GND_net), 
            .I3(GND_net), .O(n54555));   // verilog/i2c_controller.v(198[28:35])
    defparam i38853_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i38926_4_lut (.I0(n54555), .I1(state[1]), .I2(counter[0]), 
            .I3(counter[2]), .O(n54527));   // verilog/i2c_controller.v(181[4] 214[11])
    defparam i38926_4_lut.LUT_INIT = 16'hc008;
    SB_LUT4 i39150_4_lut (.I0(n54527), .I1(\state[2] ), .I2(\state[0] ), 
            .I3(n11), .O(n54697));   // verilog/i2c_controller.v(181[4] 214[11])
    defparam i39150_4_lut.LUT_INIT = 16'h0322;
    SB_DFFE enable_slow_120 (.Q(\state_7__N_4290[0] ), .C(clk16MHz), .E(n28780), 
            .D(enable_slow_N_4392));   // verilog/i2c_controller.v(58[9] 71[5])
    SB_LUT4 i22_3_lut_3_lut (.I0(\state[0] ), .I1(state[1]), .I2(\state[3] ), 
            .I3(GND_net), .O(n11));   // verilog/i2c_controller.v(77[47:62])
    defparam i22_3_lut_3_lut.LUT_INIT = 16'h1a1a;
    SB_LUT4 i23188_3_lut_4_lut (.I0(\state[0] ), .I1(state[1]), .I2(\state[2] ), 
            .I3(n15), .O(scl_enable_N_4380));   // verilog/i2c_controller.v(77[47:62])
    defparam i23188_3_lut_4_lut.LUT_INIT = 16'hfe00;
    SB_DFFSR counter2_2294_2295__i6 (.Q(counter2[5]), .C(clk16MHz), .D(n29[5]), 
            .R(n29177));   // verilog/i2c_controller.v(69[20:35])
    SB_DFFSR counter2_2294_2295__i5 (.Q(counter2[4]), .C(clk16MHz), .D(n29[4]), 
            .R(n29177));   // verilog/i2c_controller.v(69[20:35])
    SB_DFFSR counter2_2294_2295__i4 (.Q(counter2[3]), .C(clk16MHz), .D(n29[3]), 
            .R(n29177));   // verilog/i2c_controller.v(69[20:35])
    SB_DFFSR counter2_2294_2295__i3 (.Q(counter2[2]), .C(clk16MHz), .D(n29[2]), 
            .R(n29177));   // verilog/i2c_controller.v(69[20:35])
    SB_DFFSR counter2_2294_2295__i2 (.Q(counter2[1]), .C(clk16MHz), .D(n29[1]), 
            .R(n29177));   // verilog/i2c_controller.v(69[20:35])
    SB_LUT4 i1_2_lut_adj_1671 (.I0(\state[2] ), .I1(state[1]), .I2(GND_net), 
            .I3(GND_net), .O(n4_adj_4849));   // verilog/i2c_controller.v(181[4] 214[11])
    defparam i1_2_lut_adj_1671.LUT_INIT = 16'h4444;
    SB_DFF saved_addr__i1 (.Q(\saved_addr[0] ), .C(i2c_clk), .D(n29452));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_LUT4 i1_3_lut (.I0(state[1]), .I1(n33_adj_4850), .I2(n37), .I3(GND_net), 
            .O(n29171));
    defparam i1_3_lut.LUT_INIT = 16'h5454;
    SB_LUT4 i40108_4_lut (.I0(n7050), .I1(n34_adj_4851), .I2(n4_adj_4849), 
            .I3(n37), .O(n7849));
    defparam i40108_4_lut.LUT_INIT = 16'haf8c;
    SB_LUT4 sub_39_add_2_9_lut (.I0(GND_net), .I1(counter[7]), .I2(VCC_net), 
            .I3(n43961), .O(n119[7])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_39_add_2_8_lut (.I0(GND_net), .I1(counter[6]), .I2(VCC_net), 
            .I3(n43960), .O(n119[6])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_39_add_2_8 (.CI(n43960), .I0(counter[6]), .I1(VCC_net), 
            .CO(n43961));
    SB_LUT4 sub_39_add_2_7_lut (.I0(GND_net), .I1(counter[5]), .I2(VCC_net), 
            .I3(n43959), .O(n119[5])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_39_add_2_7 (.CI(n43959), .I0(counter[5]), .I1(VCC_net), 
            .CO(n43960));
    SB_LUT4 sub_39_add_2_6_lut (.I0(GND_net), .I1(counter[4]), .I2(VCC_net), 
            .I3(n43958), .O(n119[4])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_39_add_2_6 (.CI(n43958), .I0(counter[4]), .I1(VCC_net), 
            .CO(n43959));
    SB_LUT4 sub_39_add_2_5_lut (.I0(GND_net), .I1(counter[3]), .I2(VCC_net), 
            .I3(n43957), .O(n119[3])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_39_add_2_5 (.CI(n43957), .I0(counter[3]), .I1(VCC_net), 
            .CO(n43958));
    SB_LUT4 sub_39_add_2_4_lut (.I0(GND_net), .I1(counter[2]), .I2(VCC_net), 
            .I3(n43956), .O(n119[2])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_39_add_2_4 (.CI(n43956), .I0(counter[2]), .I1(VCC_net), 
            .CO(n43957));
    SB_LUT4 sub_39_add_2_3_lut (.I0(GND_net), .I1(counter[1]), .I2(VCC_net), 
            .I3(n43955), .O(n119[1])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_39_add_2_3 (.CI(n43955), .I0(counter[1]), .I1(VCC_net), 
            .CO(n43956));
    SB_LUT4 sub_39_add_2_2_lut (.I0(GND_net), .I1(counter[0]), .I2(GND_net), 
            .I3(VCC_net), .O(n119[0])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_39_add_2_2 (.CI(VCC_net), .I0(counter[0]), .I1(GND_net), 
            .CO(n43955));
    SB_DFFNESS write_enable_131 (.Q(sda_enable), .C(i2c_clk), .E(n7849), 
            .D(n19508), .S(n29171));   // verilog/i2c_controller.v(180[12] 215[6])
    SB_DFFNE sda_out_132 (.Q(sda_out_adj_4852), .C(i2c_clk), .E(n29168), 
            .D(n54697));   // verilog/i2c_controller.v(180[12] 215[6])
    SB_DFFESS counter_i0 (.Q(counter[0]), .C(i2c_clk), .E(n28838), .D(n119[0]), 
            .S(n29228));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFSR counter2_2294_2295__i1 (.Q(counter2[0]), .C(clk16MHz), .D(n29[0]), 
            .R(n29177));   // verilog/i2c_controller.v(69[20:35])
    SB_DFF data_out_i0_i7 (.Q(data[7]), .C(i2c_clk), .D(n29364));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFF data_out_i0_i6 (.Q(data[6]), .C(i2c_clk), .D(n29363));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFF data_out_i0_i5 (.Q(data[5]), .C(i2c_clk), .D(n29362));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFF data_out_i0_i4 (.Q(data[4]), .C(i2c_clk), .D(n29361));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFF data_out_i0_i3 (.Q(data[3]), .C(i2c_clk), .D(n29360));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFF data_out_i0_i2 (.Q(data[2]), .C(i2c_clk), .D(n29359));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFF data_out_i0_i1 (.Q(data[1]), .C(i2c_clk), .D(n29358));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_LUT4 i1_2_lut_adj_1672 (.I0(\state[3] ), .I1(\state[2] ), .I2(GND_net), 
            .I3(GND_net), .O(n7));
    defparam i1_2_lut_adj_1672.LUT_INIT = 16'h2222;
    SB_LUT4 i39090_4_lut (.I0(n10_adj_4853), .I1(n10), .I2(\state_7__N_4306[3] ), 
            .I3(enable), .O(n54614));   // verilog/i2c_controller.v(92[4] 172[11])
    defparam i39090_4_lut.LUT_INIT = 16'h7073;
    SB_LUT4 i1_4_lut (.I0(state[1]), .I1(n7), .I2(n54614), .I3(\state[0] ), 
            .O(n48720));   // verilog/i2c_controller.v(92[4] 172[11])
    defparam i1_4_lut.LUT_INIT = 16'ha088;
    SB_LUT4 i40640_2_lut (.I0(\state_7__N_4306[3] ), .I1(n11_adj_4855), 
            .I2(GND_net), .I3(GND_net), .O(n36727));
    defparam i40640_2_lut.LUT_INIT = 16'h1111;
    SB_LUT4 i2_2_lut (.I0(counter[2]), .I1(counter[1]), .I2(GND_net), 
            .I3(GND_net), .O(n10_adj_17));   // verilog/i2c_controller.v(110[10:22])
    defparam i2_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 state_7__I_0_143_i10_2_lut (.I0(\state[2] ), .I1(\state[3] ), 
            .I2(GND_net), .I3(GND_net), .O(n10));   // verilog/i2c_controller.v(151[5:14])
    defparam state_7__I_0_143_i10_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 i5_4_lut (.I0(counter[3]), .I1(counter[5]), .I2(counter[0]), 
            .I3(counter[4]), .O(n12));   // verilog/i2c_controller.v(110[10:22])
    defparam i5_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i6_4_lut (.I0(counter[6]), .I1(n12), .I2(counter[7]), .I3(n10_adj_17), 
            .O(n7347));   // verilog/i2c_controller.v(110[10:22])
    defparam i6_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 equal_309_i10_2_lut (.I0(\state[2] ), .I1(\state[3] ), .I2(GND_net), 
            .I3(GND_net), .O(n10_adj_4853));   // verilog/i2c_controller.v(77[27:43])
    defparam equal_309_i10_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 state_7__I_0_143_i9_2_lut (.I0(\state[0] ), .I1(state[1]), .I2(GND_net), 
            .I3(GND_net), .O(n9));   // verilog/i2c_controller.v(151[5:14])
    defparam state_7__I_0_143_i9_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 i40086_4_lut (.I0(state_7__N_4289), .I1(n7347), .I2(n11_adj_4857), 
            .I3(n36445), .O(n7354));
    defparam i40086_4_lut.LUT_INIT = 16'h5111;
    SB_LUT4 i1_4_lut_adj_1673 (.I0(n11_adj_4858), .I1(n11_adj_4855), .I2(\state_7__N_4306[3] ), 
            .I3(\saved_addr[0] ), .O(n5));   // verilog/i2c_controller.v(92[4] 172[11])
    defparam i1_4_lut_adj_1673.LUT_INIT = 16'h5755;
    SB_DFFE state_i0_i0 (.Q(\state[0] ), .C(i2c_clk), .E(VCC_net), .D(n8));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFF data_out_i0_i0 (.Q(data[0]), .C(i2c_clk), .D(n29835));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_LUT4 i38983_3_lut_4_lut (.I0(n11_adj_4857), .I1(n11_adj_4859), .I2(enable_slow_N_4393), 
            .I3(\state_7__N_4290[0] ), .O(n54609));
    defparam i38983_3_lut_4_lut.LUT_INIT = 16'h8088;
    SB_LUT4 counter2_2294_2295_add_4_7_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter2[5]), .I3(n44658), .O(n29[5])) /* synthesis syn_instantiated=1 */ ;
    defparam counter2_2294_2295_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 counter2_2294_2295_add_4_6_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter2[4]), .I3(n44657), .O(n29[4])) /* synthesis syn_instantiated=1 */ ;
    defparam counter2_2294_2295_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter2_2294_2295_add_4_6 (.CI(n44657), .I0(GND_net), .I1(counter2[4]), 
            .CO(n44658));
    SB_LUT4 counter2_2294_2295_add_4_5_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter2[3]), .I3(n44656), .O(n29[3])) /* synthesis syn_instantiated=1 */ ;
    defparam counter2_2294_2295_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i40648_3_lut_4_lut (.I0(n11_adj_4857), .I1(n11_adj_4859), .I2(n15), 
            .I3(n7354), .O(n37252));
    defparam i40648_3_lut_4_lut.LUT_INIT = 16'h7f00;
    SB_CARRY counter2_2294_2295_add_4_5 (.CI(n44656), .I0(GND_net), .I1(counter2[3]), 
            .CO(n44657));
    SB_LUT4 i2_3_lut_4_lut (.I0(\state[0] ), .I1(state[1]), .I2(\state[2] ), 
            .I3(\state[3] ), .O(n11_adj_4859));   // verilog/i2c_controller.v(77[27:43])
    defparam i2_3_lut_4_lut.LUT_INIT = 16'hfdff;
    SB_LUT4 counter2_2294_2295_add_4_4_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter2[2]), .I3(n44655), .O(n29[2])) /* synthesis syn_instantiated=1 */ ;
    defparam counter2_2294_2295_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter2_2294_2295_add_4_4 (.CI(n44655), .I0(GND_net), .I1(counter2[2]), 
            .CO(n44656));
    SB_LUT4 counter2_2294_2295_add_4_3_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter2[1]), .I3(n44654), .O(n29[1])) /* synthesis syn_instantiated=1 */ ;
    defparam counter2_2294_2295_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter2_2294_2295_add_4_3 (.CI(n44654), .I0(GND_net), .I1(counter2[1]), 
            .CO(n44655));
    SB_LUT4 counter2_2294_2295_add_4_2_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter2[0]), .I3(VCC_net), .O(n29[0])) /* synthesis syn_instantiated=1 */ ;
    defparam counter2_2294_2295_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter2_2294_2295_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(counter2[0]), 
            .CO(n44654));
    SB_LUT4 i23039_3_lut_4_lut (.I0(\state[0] ), .I1(state[1]), .I2(\state[2] ), 
            .I3(\state[3] ), .O(state_7__N_4289));
    defparam i23039_3_lut_4_lut.LUT_INIT = 16'hf800;
    SB_LUT4 i1_2_lut_3_lut (.I0(n9), .I1(n10), .I2(counter[0]), .I3(GND_net), 
            .O(n27243));   // verilog/i2c_controller.v(151[5:14])
    defparam i1_2_lut_3_lut.LUT_INIT = 16'hefef;
    SB_LUT4 i1_2_lut_3_lut_adj_1674 (.I0(n9), .I1(n10), .I2(counter[0]), 
            .I3(GND_net), .O(n27238));   // verilog/i2c_controller.v(151[5:14])
    defparam i1_2_lut_3_lut_adj_1674.LUT_INIT = 16'hfefe;
    SB_LUT4 i40646_3_lut_4_lut (.I0(n9), .I1(n10), .I2(n11_adj_4859), 
            .I3(n7354), .O(n36761));   // verilog/i2c_controller.v(151[5:14])
    defparam i40646_3_lut_4_lut.LUT_INIT = 16'h1f00;
    SB_LUT4 state_7__I_0_139_i11_2_lut_3_lut_4_lut (.I0(\state[0] ), .I1(state[1]), 
            .I2(\state[2] ), .I3(\state[3] ), .O(n11_adj_4855));
    defparam state_7__I_0_139_i11_2_lut_3_lut_4_lut.LUT_INIT = 16'hfff7;
    SB_LUT4 state_7__I_0_144_i11_2_lut_3_lut_4_lut (.I0(\state[0] ), .I1(state[1]), 
            .I2(\state[2] ), .I3(\state[3] ), .O(n11_adj_4858));   // verilog/i2c_controller.v(77[27:43])
    defparam state_7__I_0_144_i11_2_lut_3_lut_4_lut.LUT_INIT = 16'hffdf;
    SB_LUT4 equal_309_i11_2_lut_3_lut_4_lut (.I0(\state[0] ), .I1(state[1]), 
            .I2(\state[2] ), .I3(\state[3] ), .O(n15));   // verilog/i2c_controller.v(77[27:43])
    defparam equal_309_i11_2_lut_3_lut_4_lut.LUT_INIT = 16'hfffd;
    SB_LUT4 state_7__I_0_138_i11_2_lut_4_lut (.I0(\state[0] ), .I1(state[1]), 
            .I2(\state[2] ), .I3(\state[3] ), .O(n11_adj_4857));   // verilog/i2c_controller.v(109[5:12])
    defparam state_7__I_0_138_i11_2_lut_4_lut.LUT_INIT = 16'hfffb;
    SB_LUT4 i23009_2_lut_3_lut (.I0(\state[2] ), .I1(\state[3] ), .I2(\state[0] ), 
            .I3(GND_net), .O(n36445));
    defparam i23009_2_lut_3_lut.LUT_INIT = 16'hfdfd;
    SB_LUT4 i40644_3_lut_4_lut (.I0(\state[2] ), .I1(\state[3] ), .I2(state[1]), 
            .I3(n7354), .O(n51358));
    defparam i40644_3_lut_4_lut.LUT_INIT = 16'h0200;
    SB_LUT4 i22476_2_lut (.I0(i2c_clk), .I1(scl_enable), .I2(GND_net), 
            .I3(GND_net), .O(scl));   // verilog/i2c_controller.v(45[19:61])
    defparam i22476_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 i40637_2_lut_4_lut (.I0(\state[0] ), .I1(\state[2] ), .I2(state[1]), 
            .I3(\state[3] ), .O(n19508));   // verilog/i2c_controller.v(181[4] 214[11])
    defparam i40637_2_lut_4_lut.LUT_INIT = 16'h0100;
    SB_LUT4 i2708_2_lut (.I0(sda_out_adj_4852), .I1(sda_enable), .I2(GND_net), 
            .I3(GND_net), .O(sda_out));   // verilog/i2c_controller.v(46[9:20])
    defparam i2708_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_4_lut (.I0(state[1]), .I1(\state[3] ), .I2(\state[2] ), 
            .I3(\state[0] ), .O(n34_adj_4851));
    defparam i1_2_lut_4_lut.LUT_INIT = 16'h1104;
    SB_LUT4 i56_3_lut_3_lut (.I0(\state[3] ), .I1(\state[2] ), .I2(\state[0] ), 
            .I3(GND_net), .O(n33_adj_4850));
    defparam i56_3_lut_3_lut.LUT_INIT = 16'h5252;
    SB_LUT4 i3_2_lut_4_lut (.I0(\state[2] ), .I1(\state[0] ), .I2(state[1]), 
            .I3(\state[3] ), .O(n7050));
    defparam i3_2_lut_4_lut.LUT_INIT = 16'h0144;
    SB_LUT4 equal_2273_i19_2_lut_3_lut_4_lut (.I0(\state[0] ), .I1(state[1]), 
            .I2(\state[2] ), .I3(\state[3] ), .O(enable_slow_N_4393));   // verilog/i2c_controller.v(77[47:62])
    defparam equal_2273_i19_2_lut_3_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_4_lut (.I0(\state[0] ), .I1(\state[3] ), .I2(state[1]), 
            .I3(\state[2] ), .O(n29168));
    defparam i1_4_lut_4_lut.LUT_INIT = 16'h0316;
    SB_LUT4 i34043_2_lut_4_lut (.I0(\state[0] ), .I1(\state[2] ), .I2(\state[3] ), 
            .I3(n49846), .O(n29228));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i34043_2_lut_4_lut.LUT_INIT = 16'h0002;
    SB_LUT4 i1_4_lut_4_lut_adj_1675 (.I0(\state[3] ), .I1(\state[2] ), .I2(state[1]), 
            .I3(\state[0] ), .O(n37));
    defparam i1_4_lut_4_lut_adj_1675.LUT_INIT = 16'h1154;
    SB_LUT4 i1_2_lut_3_lut_adj_1676 (.I0(enable), .I1(\state_7__N_4290[0] ), 
            .I2(enable_slow_N_4393), .I3(GND_net), .O(n28780));
    defparam i1_2_lut_3_lut_adj_1676.LUT_INIT = 16'heaea;
    
endmodule
//
// Verilog Description of module \quadrature_decoder(1) 
//

module \quadrature_decoder(1)  (encoder1_position, GND_net, b_prev, a_new, 
            position_31__N_4108, VCC_net, ENCODER1_B_N_keep, n2269, 
            ENCODER1_A_N_keep, n29500, n2274) /* synthesis lattice_noprune=1 */ ;
    output [31:0]encoder1_position;
    input GND_net;
    output b_prev;
    output [1:0]a_new;
    output position_31__N_4108;
    input VCC_net;
    input ENCODER1_B_N_keep;
    input n2269;
    input ENCODER1_A_N_keep;
    input n29500;
    output n2274;
    
    wire [31:0]n133;
    
    wire direction_N_4113, n44653, n44652, n44651, n44650, n44649, 
        n44648, n44647, n44646, n44645, n44644, n44643, n44642, 
        n44641, n44640, n44639, n44638, n44637, n44636, n44635, 
        n44634, n44633, n44632, n44631, n44630, n44629, n44628;
    wire [1:0]b_new;   // vhdl/quadrature_decoder.vhd(40[9:14])
    
    wire position_31__N_4111, debounce_cnt, a_prev;
    wire [1:0]a_new_c;   // vhdl/quadrature_decoder.vhd(39[9:14])
    
    wire a_prev_N_4116, n44627, n44626, n44625, n44624, n44623, 
        n29548, n29547;
    
    SB_LUT4 position_2293_add_4_33_lut (.I0(GND_net), .I1(direction_N_4113), 
            .I2(encoder1_position[31]), .I3(n44653), .O(n133[31])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2293_add_4_33_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 position_2293_add_4_32_lut (.I0(GND_net), .I1(direction_N_4113), 
            .I2(encoder1_position[30]), .I3(n44652), .O(n133[30])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2293_add_4_32_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2293_add_4_32 (.CI(n44652), .I0(direction_N_4113), 
            .I1(encoder1_position[30]), .CO(n44653));
    SB_LUT4 position_2293_add_4_31_lut (.I0(GND_net), .I1(direction_N_4113), 
            .I2(encoder1_position[29]), .I3(n44651), .O(n133[29])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2293_add_4_31_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2293_add_4_31 (.CI(n44651), .I0(direction_N_4113), 
            .I1(encoder1_position[29]), .CO(n44652));
    SB_LUT4 position_2293_add_4_30_lut (.I0(GND_net), .I1(direction_N_4113), 
            .I2(encoder1_position[28]), .I3(n44650), .O(n133[28])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2293_add_4_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2293_add_4_30 (.CI(n44650), .I0(direction_N_4113), 
            .I1(encoder1_position[28]), .CO(n44651));
    SB_LUT4 position_2293_add_4_29_lut (.I0(GND_net), .I1(direction_N_4113), 
            .I2(encoder1_position[27]), .I3(n44649), .O(n133[27])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2293_add_4_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2293_add_4_29 (.CI(n44649), .I0(direction_N_4113), 
            .I1(encoder1_position[27]), .CO(n44650));
    SB_LUT4 position_2293_add_4_28_lut (.I0(GND_net), .I1(direction_N_4113), 
            .I2(encoder1_position[26]), .I3(n44648), .O(n133[26])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2293_add_4_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2293_add_4_28 (.CI(n44648), .I0(direction_N_4113), 
            .I1(encoder1_position[26]), .CO(n44649));
    SB_LUT4 position_2293_add_4_27_lut (.I0(GND_net), .I1(direction_N_4113), 
            .I2(encoder1_position[25]), .I3(n44647), .O(n133[25])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2293_add_4_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2293_add_4_27 (.CI(n44647), .I0(direction_N_4113), 
            .I1(encoder1_position[25]), .CO(n44648));
    SB_LUT4 position_2293_add_4_26_lut (.I0(GND_net), .I1(direction_N_4113), 
            .I2(encoder1_position[24]), .I3(n44646), .O(n133[24])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2293_add_4_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2293_add_4_26 (.CI(n44646), .I0(direction_N_4113), 
            .I1(encoder1_position[24]), .CO(n44647));
    SB_LUT4 position_2293_add_4_25_lut (.I0(GND_net), .I1(direction_N_4113), 
            .I2(encoder1_position[23]), .I3(n44645), .O(n133[23])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2293_add_4_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2293_add_4_25 (.CI(n44645), .I0(direction_N_4113), 
            .I1(encoder1_position[23]), .CO(n44646));
    SB_LUT4 position_2293_add_4_24_lut (.I0(GND_net), .I1(direction_N_4113), 
            .I2(encoder1_position[22]), .I3(n44644), .O(n133[22])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2293_add_4_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2293_add_4_24 (.CI(n44644), .I0(direction_N_4113), 
            .I1(encoder1_position[22]), .CO(n44645));
    SB_LUT4 position_2293_add_4_23_lut (.I0(GND_net), .I1(direction_N_4113), 
            .I2(encoder1_position[21]), .I3(n44643), .O(n133[21])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2293_add_4_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2293_add_4_23 (.CI(n44643), .I0(direction_N_4113), 
            .I1(encoder1_position[21]), .CO(n44644));
    SB_LUT4 position_2293_add_4_22_lut (.I0(GND_net), .I1(direction_N_4113), 
            .I2(encoder1_position[20]), .I3(n44642), .O(n133[20])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2293_add_4_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2293_add_4_22 (.CI(n44642), .I0(direction_N_4113), 
            .I1(encoder1_position[20]), .CO(n44643));
    SB_LUT4 position_2293_add_4_21_lut (.I0(GND_net), .I1(direction_N_4113), 
            .I2(encoder1_position[19]), .I3(n44641), .O(n133[19])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2293_add_4_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2293_add_4_21 (.CI(n44641), .I0(direction_N_4113), 
            .I1(encoder1_position[19]), .CO(n44642));
    SB_LUT4 position_2293_add_4_20_lut (.I0(GND_net), .I1(direction_N_4113), 
            .I2(encoder1_position[18]), .I3(n44640), .O(n133[18])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2293_add_4_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2293_add_4_20 (.CI(n44640), .I0(direction_N_4113), 
            .I1(encoder1_position[18]), .CO(n44641));
    SB_LUT4 position_2293_add_4_19_lut (.I0(GND_net), .I1(direction_N_4113), 
            .I2(encoder1_position[17]), .I3(n44639), .O(n133[17])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2293_add_4_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2293_add_4_19 (.CI(n44639), .I0(direction_N_4113), 
            .I1(encoder1_position[17]), .CO(n44640));
    SB_LUT4 position_2293_add_4_18_lut (.I0(GND_net), .I1(direction_N_4113), 
            .I2(encoder1_position[16]), .I3(n44638), .O(n133[16])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2293_add_4_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2293_add_4_18 (.CI(n44638), .I0(direction_N_4113), 
            .I1(encoder1_position[16]), .CO(n44639));
    SB_LUT4 position_2293_add_4_17_lut (.I0(GND_net), .I1(direction_N_4113), 
            .I2(encoder1_position[15]), .I3(n44637), .O(n133[15])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2293_add_4_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2293_add_4_17 (.CI(n44637), .I0(direction_N_4113), 
            .I1(encoder1_position[15]), .CO(n44638));
    SB_LUT4 position_2293_add_4_16_lut (.I0(GND_net), .I1(direction_N_4113), 
            .I2(encoder1_position[14]), .I3(n44636), .O(n133[14])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2293_add_4_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2293_add_4_16 (.CI(n44636), .I0(direction_N_4113), 
            .I1(encoder1_position[14]), .CO(n44637));
    SB_LUT4 position_2293_add_4_15_lut (.I0(GND_net), .I1(direction_N_4113), 
            .I2(encoder1_position[13]), .I3(n44635), .O(n133[13])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2293_add_4_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2293_add_4_15 (.CI(n44635), .I0(direction_N_4113), 
            .I1(encoder1_position[13]), .CO(n44636));
    SB_LUT4 position_2293_add_4_14_lut (.I0(GND_net), .I1(direction_N_4113), 
            .I2(encoder1_position[12]), .I3(n44634), .O(n133[12])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2293_add_4_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2293_add_4_14 (.CI(n44634), .I0(direction_N_4113), 
            .I1(encoder1_position[12]), .CO(n44635));
    SB_LUT4 position_2293_add_4_13_lut (.I0(GND_net), .I1(direction_N_4113), 
            .I2(encoder1_position[11]), .I3(n44633), .O(n133[11])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2293_add_4_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2293_add_4_13 (.CI(n44633), .I0(direction_N_4113), 
            .I1(encoder1_position[11]), .CO(n44634));
    SB_LUT4 position_2293_add_4_12_lut (.I0(GND_net), .I1(direction_N_4113), 
            .I2(encoder1_position[10]), .I3(n44632), .O(n133[10])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2293_add_4_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2293_add_4_12 (.CI(n44632), .I0(direction_N_4113), 
            .I1(encoder1_position[10]), .CO(n44633));
    SB_LUT4 position_2293_add_4_11_lut (.I0(GND_net), .I1(direction_N_4113), 
            .I2(encoder1_position[9]), .I3(n44631), .O(n133[9])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2293_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2293_add_4_11 (.CI(n44631), .I0(direction_N_4113), 
            .I1(encoder1_position[9]), .CO(n44632));
    SB_LUT4 position_2293_add_4_10_lut (.I0(GND_net), .I1(direction_N_4113), 
            .I2(encoder1_position[8]), .I3(n44630), .O(n133[8])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2293_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2293_add_4_10 (.CI(n44630), .I0(direction_N_4113), 
            .I1(encoder1_position[8]), .CO(n44631));
    SB_LUT4 position_2293_add_4_9_lut (.I0(GND_net), .I1(direction_N_4113), 
            .I2(encoder1_position[7]), .I3(n44629), .O(n133[7])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2293_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2293_add_4_9 (.CI(n44629), .I0(direction_N_4113), 
            .I1(encoder1_position[7]), .CO(n44630));
    SB_LUT4 position_2293_add_4_8_lut (.I0(GND_net), .I1(direction_N_4113), 
            .I2(encoder1_position[6]), .I3(n44628), .O(n133[6])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2293_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2293_add_4_8 (.CI(n44628), .I0(direction_N_4113), 
            .I1(encoder1_position[6]), .CO(n44629));
    SB_LUT4 b_prev_I_0_43_2_lut (.I0(b_prev), .I1(b_new[1]), .I2(GND_net), 
            .I3(GND_net), .O(position_31__N_4111));   // vhdl/quadrature_decoder.vhd(63[37:56])
    defparam b_prev_I_0_43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 debounce_cnt_I_0_4_lut (.I0(debounce_cnt), .I1(a_prev), .I2(position_31__N_4111), 
            .I3(a_new[1]), .O(position_31__N_4108));   // vhdl/quadrature_decoder.vhd(62[7] 63[64])
    defparam debounce_cnt_I_0_4_lut.LUT_INIT = 16'ha2a8;
    SB_LUT4 i40095_4_lut (.I0(a_new_c[0]), .I1(b_new[0]), .I2(a_new[1]), 
            .I3(b_new[1]), .O(a_prev_N_4116));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    defparam i40095_4_lut.LUT_INIT = 16'h8421;
    SB_LUT4 position_2293_add_4_7_lut (.I0(GND_net), .I1(direction_N_4113), 
            .I2(encoder1_position[5]), .I3(n44627), .O(n133[5])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2293_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2293_add_4_7 (.CI(n44627), .I0(direction_N_4113), 
            .I1(encoder1_position[5]), .CO(n44628));
    SB_LUT4 position_2293_add_4_6_lut (.I0(GND_net), .I1(direction_N_4113), 
            .I2(encoder1_position[4]), .I3(n44626), .O(n133[4])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2293_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2293_add_4_6 (.CI(n44626), .I0(direction_N_4113), 
            .I1(encoder1_position[4]), .CO(n44627));
    SB_LUT4 position_2293_add_4_5_lut (.I0(GND_net), .I1(direction_N_4113), 
            .I2(encoder1_position[3]), .I3(n44625), .O(n133[3])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2293_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2293_add_4_5 (.CI(n44625), .I0(direction_N_4113), 
            .I1(encoder1_position[3]), .CO(n44626));
    SB_LUT4 position_2293_add_4_4_lut (.I0(GND_net), .I1(direction_N_4113), 
            .I2(encoder1_position[2]), .I3(n44624), .O(n133[2])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2293_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2293_add_4_4 (.CI(n44624), .I0(direction_N_4113), 
            .I1(encoder1_position[2]), .CO(n44625));
    SB_LUT4 position_2293_add_4_3_lut (.I0(GND_net), .I1(direction_N_4113), 
            .I2(encoder1_position[1]), .I3(n44623), .O(n133[1])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2293_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2293_add_4_3 (.CI(n44623), .I0(direction_N_4113), 
            .I1(encoder1_position[1]), .CO(n44624));
    SB_LUT4 position_2293_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(encoder1_position[0]), 
            .I3(VCC_net), .O(n133[0])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2293_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2293_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(encoder1_position[0]), 
            .CO(n44623));
    SB_LUT4 b_prev_I_0_45_2_lut (.I0(b_prev), .I1(a_new[1]), .I2(GND_net), 
            .I3(GND_net), .O(direction_N_4113));   // vhdl/quadrature_decoder.vhd(64[18:37])
    defparam b_prev_I_0_45_2_lut.LUT_INIT = 16'h9999;
    SB_DFF b_new_i0 (.Q(b_new[0]), .C(n2269), .D(ENCODER1_B_N_keep));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_DFF a_new_i0 (.Q(a_new_c[0]), .C(n2269), .D(ENCODER1_A_N_keep));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_DFF debounce_cnt_37 (.Q(debounce_cnt), .C(n2269), .D(a_prev_N_4116));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_DFF direction_40 (.Q(n2274), .C(n2269), .D(n29500));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_DFFE position_2293__i31 (.Q(encoder1_position[31]), .C(n2269), .E(position_31__N_4108), 
            .D(n133[31]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2293__i30 (.Q(encoder1_position[30]), .C(n2269), .E(position_31__N_4108), 
            .D(n133[30]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2293__i29 (.Q(encoder1_position[29]), .C(n2269), .E(position_31__N_4108), 
            .D(n133[29]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2293__i28 (.Q(encoder1_position[28]), .C(n2269), .E(position_31__N_4108), 
            .D(n133[28]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2293__i27 (.Q(encoder1_position[27]), .C(n2269), .E(position_31__N_4108), 
            .D(n133[27]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2293__i26 (.Q(encoder1_position[26]), .C(n2269), .E(position_31__N_4108), 
            .D(n133[26]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2293__i25 (.Q(encoder1_position[25]), .C(n2269), .E(position_31__N_4108), 
            .D(n133[25]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2293__i24 (.Q(encoder1_position[24]), .C(n2269), .E(position_31__N_4108), 
            .D(n133[24]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2293__i23 (.Q(encoder1_position[23]), .C(n2269), .E(position_31__N_4108), 
            .D(n133[23]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2293__i22 (.Q(encoder1_position[22]), .C(n2269), .E(position_31__N_4108), 
            .D(n133[22]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2293__i21 (.Q(encoder1_position[21]), .C(n2269), .E(position_31__N_4108), 
            .D(n133[21]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2293__i20 (.Q(encoder1_position[20]), .C(n2269), .E(position_31__N_4108), 
            .D(n133[20]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2293__i19 (.Q(encoder1_position[19]), .C(n2269), .E(position_31__N_4108), 
            .D(n133[19]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2293__i18 (.Q(encoder1_position[18]), .C(n2269), .E(position_31__N_4108), 
            .D(n133[18]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2293__i17 (.Q(encoder1_position[17]), .C(n2269), .E(position_31__N_4108), 
            .D(n133[17]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2293__i16 (.Q(encoder1_position[16]), .C(n2269), .E(position_31__N_4108), 
            .D(n133[16]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2293__i15 (.Q(encoder1_position[15]), .C(n2269), .E(position_31__N_4108), 
            .D(n133[15]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2293__i14 (.Q(encoder1_position[14]), .C(n2269), .E(position_31__N_4108), 
            .D(n133[14]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2293__i13 (.Q(encoder1_position[13]), .C(n2269), .E(position_31__N_4108), 
            .D(n133[13]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2293__i12 (.Q(encoder1_position[12]), .C(n2269), .E(position_31__N_4108), 
            .D(n133[12]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2293__i11 (.Q(encoder1_position[11]), .C(n2269), .E(position_31__N_4108), 
            .D(n133[11]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2293__i10 (.Q(encoder1_position[10]), .C(n2269), .E(position_31__N_4108), 
            .D(n133[10]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2293__i9 (.Q(encoder1_position[9]), .C(n2269), .E(position_31__N_4108), 
            .D(n133[9]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2293__i8 (.Q(encoder1_position[8]), .C(n2269), .E(position_31__N_4108), 
            .D(n133[8]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2293__i7 (.Q(encoder1_position[7]), .C(n2269), .E(position_31__N_4108), 
            .D(n133[7]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2293__i6 (.Q(encoder1_position[6]), .C(n2269), .E(position_31__N_4108), 
            .D(n133[6]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2293__i5 (.Q(encoder1_position[5]), .C(n2269), .E(position_31__N_4108), 
            .D(n133[5]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2293__i4 (.Q(encoder1_position[4]), .C(n2269), .E(position_31__N_4108), 
            .D(n133[4]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2293__i3 (.Q(encoder1_position[3]), .C(n2269), .E(position_31__N_4108), 
            .D(n133[3]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2293__i2 (.Q(encoder1_position[2]), .C(n2269), .E(position_31__N_4108), 
            .D(n133[2]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2293__i1 (.Q(encoder1_position[1]), .C(n2269), .E(position_31__N_4108), 
            .D(n133[1]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2293__i0 (.Q(encoder1_position[0]), .C(n2269), .E(position_31__N_4108), 
            .D(n133[0]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFF a_new_i1 (.Q(a_new[1]), .C(n2269), .D(a_new_c[0]));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_DFF b_new_i1 (.Q(b_new[1]), .C(n2269), .D(b_new[0]));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_LUT4 i15468_3_lut_4_lut (.I0(debounce_cnt), .I1(a_prev_N_4116), .I2(a_new[1]), 
            .I3(a_prev), .O(n29548));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    defparam i15468_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i15467_3_lut_4_lut (.I0(debounce_cnt), .I1(a_prev_N_4116), .I2(b_new[1]), 
            .I3(b_prev), .O(n29547));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    defparam i15467_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF a_prev_38 (.Q(a_prev), .C(n2269), .D(n29548));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_DFF b_prev_39 (.Q(b_prev), .C(n2269), .D(n29547));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    
endmodule
//
// Verilog Description of module coms
//

module coms (n29523, deadband, clk16MHz, n29522, n29521, \Kp[1] , 
            n29520, \Kp[2] , n29519, \Kp[3] , n29518, \Kp[4] , GND_net, 
            \data_in_frame[3] , n63, n3303, n27219, n48947, n48957, 
            \data_out_frame[16] , \data_out_frame[17] , \data_out_frame[18] , 
            \data_out_frame[19] , n27218, \FRAME_MATCHER.state[3] , \data_out_frame[22] , 
            \data_out_frame[23] , \data_out_frame[20] , \data_out_frame[21] , 
            \data_in_frame[2] , rx_data_ready, n22875, \data_out_frame[6] , 
            \data_out_frame[7] , \data_out_frame[4] , \data_out_frame[5] , 
            n29516, \Kp[5] , \data_in_frame[4] , \data_in_frame[5] , 
            PWMLimit, n50654, \data_in[0] , \data_in[1] , \data_in[2] , 
            \data_in[3] , n29515, \Kp[6] , n63_adj_6, n29514, \Kp[7] , 
            rx_data, n122, n8, n7, \data_in_frame[1] , \data_in_frame[8] , 
            ID, \data_out_frame[8] , \data_out_frame[9] , \data_out_frame[10] , 
            \data_out_frame[11] , \data_out_frame[14] , \data_out_frame[15] , 
            \data_out_frame[12] , \data_out_frame[13] , tx_active, \data_in_frame[13] , 
            \data_in_frame[15] , \FRAME_MATCHER.state[0] , n29513, \Kp[8] , 
            n29512, \Kp[9] , setpoint, n19602, \data_in_frame[8][2] , 
            n29511, \Kp[10] , \data_in_frame[9] , n29510, \Kp[11] , 
            n29509, \Kp[12] , \data_in_frame[10][2] , n29508, \Kp[13] , 
            n29507, \Kp[14] , n363, n32464, \data_in_frame[12] , \data_in_frame[10][1] , 
            n29506, \Kp[15] , \data_in_frame[16] , n29505, \Ki[1] , 
            n29504, \Ki[2] , n29503, \Ki[3] , n29502, \Ki[4] , n29499, 
            \Ki[5] , n29498, \Ki[6] , n29497, \Ki[7] , n29496, \Ki[8] , 
            n29495, \Ki[9] , n29494, \Ki[10] , n29493, \Ki[11] , 
            n29492, \Ki[12] , n29491, \Ki[13] , n29490, \Ki[14] , 
            n29486, \Ki[15] , n29485, n29484, n29483, n29482, n29481, 
            n29480, n29479, n29478, n29477, n29476, \data_in_frame[14] , 
            n29472, n4, n29471, \data_in_frame[8][6] , \data_in_frame[11] , 
            n29470, n29469, DE_c, n29468, n29467, n29466, n29465, 
            n29464, n29463, n29462, n29461, n29460, n29456, n29455, 
            n29454, n29453, n29451, \data_out_frame[25] , n29450, 
            \data_in_frame[21] , \data_in_frame[20] , n29449, n29448, 
            n29447, n29446, n29445, n29444, n29443, n29442, n29441, 
            n29440, n29439, n29438, n29437, n29436, n29435, n29434, 
            n29433, n29432, n29431, n29430, n29429, n29428, n29427, 
            n29426, n29425, n29424, n29423, n29422, n29421, n29420, 
            n29419, \data_out_frame[24] , \data_in_frame[8][4] , \data_in_frame[8][5] , 
            n29418, n30058, n30057, n30056, n30055, n30054, n30053, 
            n30052, n30051, n30050, n30049, n30048, n30047, n30046, 
            n30045, n30044, n30043, n30042, n30041, n30040, n30039, 
            n30038, n30037, n30036, n30035, n30034, n30033, n30032, 
            n30031, n30030, n30029, n30028, n30027, n30026, n30025, 
            n30024, n30023, n30022, n30021, n30020, n30019, n30018, 
            n30017, n30016, n30015, n30014, n30013, n30012, n30011, 
            n30010, n30009, n30008, n30007, n30006, n30005, n30004, 
            n30003, n30002, n30001, n30000, n29999, n29998, n29997, 
            n29996, n29995, n29994, n29993, n29992, n29991, n29990, 
            n29989, n29988, n29987, n29986, n29985, n29984, n29983, 
            n29982, n29981, n29980, n29979, n29978, n29977, n29976, 
            n29417, n29416, n29415, n29414, n29412, n29411, n29410, 
            n29408, n29406, n29405, n29404, n29403, n29402, n29401, 
            n29400, n29397, n29396, n29395, n29394, LED_c, n29975, 
            n29974, n29973, n29972, n29971, n29970, n29969, n29968, 
            n29967, n29962, control_mode, n29961, n29960, n29959, 
            n29958, n29957, n29956, n29955, current_limit, n29954, 
            n29953, n29952, n29951, n29950, n29949, n29948, n29947, 
            n29946, n29945, n29944, n29943, n29942, n29941, n29940, 
            n29939, n29390, n29938, n29389, n29937, n29936, n29935, 
            n29934, n29388, n29387, n29386, n29385, n29384, n29383, 
            n29382, n29380, n29379, n29378, n50741, n29375, n29374, 
            neopxl_color, n29371, n29370, \Ki[0] , n29369, \Kp[0] , 
            n29368, IntegralLimit, n29933, n29932, n29931, n29930, 
            n29929, n29928, n29927, n29926, n6, n29925, n29923, 
            n29922, n29356, n29355, n29921, n29920, n29919, n29918, 
            n57033, n29353, n29874, n29873, n29872, n29870, n29868, 
            n29867, n29866, n29865, n29864, n29863, n29862, n29861, 
            n29834, n29833, n29832, n29831, n29830, n29827, n29826, 
            n29825, n29824, \data_in_frame[10][3] , \data_in_frame[10][4] , 
            \data_in_frame[10][5] , \data_in_frame[10][6] , \data_in_frame[10][7] , 
            n29571, n29570, n29569, n29568, n29567, n29566, n29565, 
            n29564, n29563, n29562, n29561, n29560, n29559, n29558, 
            n29557, n29556, n29555, n29554, n29553, n29552, n29551, 
            n29550, n29549, n29546, n29545, n29544, n29543, n29542, 
            n29541, n29540, n29539, n29538, n29537, n29536, n29534, 
            n29533, n29532, n29531, n29530, n29529, n29527, n29526, 
            n29525, n29524, n24210, \state[0] , \state[2] , \state[3] , 
            n7936, \FRAME_MATCHER.state_31__N_3007[2] , n28848, n29280, 
            r_SM_Main, \r_SM_Main_2__N_3848[1] , \r_Bit_Index[0] , VCC_net, 
            tx_o, n19728, n29842, n29413, n57032, n4_adj_7, tx_enable, 
            r_SM_Main_adj_15, \r_SM_Main_2__N_3777[2] , r_Rx_Data, n28852, 
            n29282, RX_N_10, \r_Bit_Index[0]_adj_11 , n4_adj_12, n36556, 
            n4_adj_13, n4_adj_14, n29845, n48522, n48878, n29880, 
            n29878, n29877, n29871, n29860, n29849, n29759, n29528, 
            n27208, n27203) /* synthesis syn_module_defined=1 */ ;
    input n29523;
    output [23:0]deadband;
    input clk16MHz;
    input n29522;
    input n29521;
    output \Kp[1] ;
    input n29520;
    output \Kp[2] ;
    input n29519;
    output \Kp[3] ;
    input n29518;
    output \Kp[4] ;
    input GND_net;
    output [7:0]\data_in_frame[3] ;
    output n63;
    output n3303;
    output n27219;
    output n48947;
    output n48957;
    output [7:0]\data_out_frame[16] ;
    output [7:0]\data_out_frame[17] ;
    output [7:0]\data_out_frame[18] ;
    output [7:0]\data_out_frame[19] ;
    output n27218;
    output \FRAME_MATCHER.state[3] ;
    output [7:0]\data_out_frame[22] ;
    output [7:0]\data_out_frame[23] ;
    output [7:0]\data_out_frame[20] ;
    output [7:0]\data_out_frame[21] ;
    output [7:0]\data_in_frame[2] ;
    output rx_data_ready;
    output n22875;
    output [7:0]\data_out_frame[6] ;
    output [7:0]\data_out_frame[7] ;
    output [7:0]\data_out_frame[4] ;
    output [7:0]\data_out_frame[5] ;
    input n29516;
    output \Kp[5] ;
    output [7:0]\data_in_frame[4] ;
    output [7:0]\data_in_frame[5] ;
    output [23:0]PWMLimit;
    output n50654;
    output [7:0]\data_in[0] ;
    output [7:0]\data_in[1] ;
    output [7:0]\data_in[2] ;
    output [7:0]\data_in[3] ;
    input n29515;
    output \Kp[6] ;
    output n63_adj_6;
    input n29514;
    output \Kp[7] ;
    output [7:0]rx_data;
    output n122;
    output n8;
    output n7;
    output [7:0]\data_in_frame[1] ;
    output [7:0]\data_in_frame[8] ;
    input [7:0]ID;
    output [7:0]\data_out_frame[8] ;
    output [7:0]\data_out_frame[9] ;
    output [7:0]\data_out_frame[10] ;
    output [7:0]\data_out_frame[11] ;
    output [7:0]\data_out_frame[14] ;
    output [7:0]\data_out_frame[15] ;
    output [7:0]\data_out_frame[12] ;
    output [7:0]\data_out_frame[13] ;
    output tx_active;
    output [7:0]\data_in_frame[13] ;
    output [7:0]\data_in_frame[15] ;
    output \FRAME_MATCHER.state[0] ;
    input n29513;
    output \Kp[8] ;
    input n29512;
    output \Kp[9] ;
    output [23:0]setpoint;
    output n19602;
    output \data_in_frame[8][2] ;
    input n29511;
    output \Kp[10] ;
    output [7:0]\data_in_frame[9] ;
    input n29510;
    output \Kp[11] ;
    input n29509;
    output \Kp[12] ;
    output \data_in_frame[10][2] ;
    input n29508;
    output \Kp[13] ;
    input n29507;
    output \Kp[14] ;
    input n363;
    output n32464;
    output [7:0]\data_in_frame[12] ;
    output \data_in_frame[10][1] ;
    input n29506;
    output \Kp[15] ;
    output [7:0]\data_in_frame[16] ;
    input n29505;
    output \Ki[1] ;
    input n29504;
    output \Ki[2] ;
    input n29503;
    output \Ki[3] ;
    input n29502;
    output \Ki[4] ;
    input n29499;
    output \Ki[5] ;
    input n29498;
    output \Ki[6] ;
    input n29497;
    output \Ki[7] ;
    input n29496;
    output \Ki[8] ;
    input n29495;
    output \Ki[9] ;
    input n29494;
    output \Ki[10] ;
    input n29493;
    output \Ki[11] ;
    input n29492;
    output \Ki[12] ;
    input n29491;
    output \Ki[13] ;
    input n29490;
    output \Ki[14] ;
    input n29486;
    output \Ki[15] ;
    input n29485;
    input n29484;
    input n29483;
    input n29482;
    input n29481;
    input n29480;
    input n29479;
    input n29478;
    input n29477;
    input n29476;
    output [7:0]\data_in_frame[14] ;
    input n29472;
    output n4;
    input n29471;
    output \data_in_frame[8][6] ;
    output [7:0]\data_in_frame[11] ;
    input n29470;
    input n29469;
    output DE_c;
    input n29468;
    input n29467;
    input n29466;
    input n29465;
    input n29464;
    input n29463;
    input n29462;
    input n29461;
    input n29460;
    input n29456;
    input n29455;
    input n29454;
    input n29453;
    input n29451;
    output [7:0]\data_out_frame[25] ;
    input n29450;
    output [7:0]\data_in_frame[21] ;
    output [7:0]\data_in_frame[20] ;
    input n29449;
    input n29448;
    input n29447;
    input n29446;
    input n29445;
    input n29444;
    input n29443;
    input n29442;
    input n29441;
    input n29440;
    input n29439;
    input n29438;
    input n29437;
    input n29436;
    input n29435;
    input n29434;
    input n29433;
    input n29432;
    input n29431;
    input n29430;
    input n29429;
    input n29428;
    input n29427;
    input n29426;
    input n29425;
    input n29424;
    input n29423;
    input n29422;
    input n29421;
    input n29420;
    input n29419;
    output [7:0]\data_out_frame[24] ;
    output \data_in_frame[8][4] ;
    output \data_in_frame[8][5] ;
    input n29418;
    input n30058;
    input n30057;
    input n30056;
    input n30055;
    input n30054;
    input n30053;
    input n30052;
    input n30051;
    input n30050;
    input n30049;
    input n30048;
    input n30047;
    input n30046;
    input n30045;
    input n30044;
    input n30043;
    input n30042;
    input n30041;
    input n30040;
    input n30039;
    input n30038;
    input n30037;
    input n30036;
    input n30035;
    input n30034;
    input n30033;
    input n30032;
    input n30031;
    input n30030;
    input n30029;
    input n30028;
    input n30027;
    input n30026;
    input n30025;
    input n30024;
    input n30023;
    input n30022;
    input n30021;
    input n30020;
    input n30019;
    input n30018;
    input n30017;
    input n30016;
    input n30015;
    input n30014;
    input n30013;
    input n30012;
    input n30011;
    input n30010;
    input n30009;
    input n30008;
    input n30007;
    input n30006;
    input n30005;
    input n30004;
    input n30003;
    input n30002;
    input n30001;
    input n30000;
    input n29999;
    input n29998;
    input n29997;
    input n29996;
    input n29995;
    input n29994;
    input n29993;
    input n29992;
    input n29991;
    input n29990;
    input n29989;
    input n29988;
    input n29987;
    input n29986;
    input n29985;
    input n29984;
    input n29983;
    input n29982;
    input n29981;
    input n29980;
    input n29979;
    input n29978;
    input n29977;
    input n29976;
    input n29417;
    input n29416;
    input n29415;
    input n29414;
    input n29412;
    input n29411;
    input n29410;
    input n29408;
    input n29406;
    input n29405;
    input n29404;
    input n29403;
    input n29402;
    input n29401;
    input n29400;
    input n29397;
    input n29396;
    input n29395;
    input n29394;
    output LED_c;
    input n29975;
    input n29974;
    input n29973;
    input n29972;
    input n29971;
    input n29970;
    input n29969;
    input n29968;
    input n29967;
    input n29962;
    output [7:0]control_mode;
    input n29961;
    input n29960;
    input n29959;
    input n29958;
    input n29957;
    input n29956;
    input n29955;
    output [15:0]current_limit;
    input n29954;
    input n29953;
    input n29952;
    input n29951;
    input n29950;
    input n29949;
    input n29948;
    input n29947;
    input n29946;
    input n29945;
    input n29944;
    input n29943;
    input n29942;
    input n29941;
    input n29940;
    input n29939;
    input n29390;
    input n29938;
    input n29389;
    input n29937;
    input n29936;
    input n29935;
    input n29934;
    input n29388;
    input n29387;
    input n29386;
    input n29385;
    input n29384;
    input n29383;
    input n29382;
    input n29380;
    input n29379;
    input n29378;
    input n50741;
    input n29375;
    input n29374;
    output [23:0]neopxl_color;
    input n29371;
    input n29370;
    output \Ki[0] ;
    input n29369;
    output \Kp[0] ;
    input n29368;
    output [23:0]IntegralLimit;
    input n29933;
    input n29932;
    input n29931;
    input n29930;
    input n29929;
    input n29928;
    input n29927;
    input n29926;
    output n6;
    input n29925;
    input n29923;
    input n29922;
    input n29356;
    input n29355;
    input n29921;
    input n29920;
    input n29919;
    input n29918;
    input n57033;
    input n29353;
    input n29874;
    input n29873;
    input n29872;
    input n29870;
    input n29868;
    input n29867;
    input n29866;
    input n29865;
    input n29864;
    input n29863;
    input n29862;
    input n29861;
    input n29834;
    input n29833;
    input n29832;
    input n29831;
    input n29830;
    input n29827;
    input n29826;
    input n29825;
    input n29824;
    output \data_in_frame[10][3] ;
    output \data_in_frame[10][4] ;
    output \data_in_frame[10][5] ;
    output \data_in_frame[10][6] ;
    output \data_in_frame[10][7] ;
    input n29571;
    input n29570;
    input n29569;
    input n29568;
    input n29567;
    input n29566;
    input n29565;
    input n29564;
    input n29563;
    input n29562;
    input n29561;
    input n29560;
    input n29559;
    input n29558;
    input n29557;
    input n29556;
    input n29555;
    input n29554;
    input n29553;
    input n29552;
    input n29551;
    input n29550;
    input n29549;
    input n29546;
    input n29545;
    input n29544;
    input n29543;
    input n29542;
    input n29541;
    input n29540;
    input n29539;
    input n29538;
    input n29537;
    input n29536;
    input n29534;
    input n29533;
    input n29532;
    input n29531;
    input n29530;
    input n29529;
    input n29527;
    input n29526;
    input n29525;
    input n29524;
    output n24210;
    input \state[0] ;
    input \state[2] ;
    input \state[3] ;
    output n7936;
    output \FRAME_MATCHER.state_31__N_3007[2] ;
    output n28848;
    output n29280;
    output [2:0]r_SM_Main;
    output \r_SM_Main_2__N_3848[1] ;
    output \r_Bit_Index[0] ;
    input VCC_net;
    output tx_o;
    output n19728;
    input n29842;
    input n29413;
    input n57032;
    output n4_adj_7;
    output tx_enable;
    output [2:0]r_SM_Main_adj_15;
    output \r_SM_Main_2__N_3777[2] ;
    output r_Rx_Data;
    output n28852;
    output n29282;
    input RX_N_10;
    output \r_Bit_Index[0]_adj_11 ;
    output n4_adj_12;
    output n36556;
    output n4_adj_13;
    output n4_adj_14;
    input n29845;
    input n48522;
    input n48878;
    input n29880;
    input n29878;
    input n29877;
    input n29871;
    input n29860;
    input n29849;
    input n29759;
    input n29528;
    output n27208;
    output n27203;
    
    wire clk16MHz /* synthesis SET_AS_NETWORK=clk16MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    
    wire n56910, n56859, n7_c;
    wire [7:0]byte_transmit_counter;   // verilog/coms.v(103[12:33])
    wire [7:0]tx_data;   // verilog/coms.v(106[13:20])
    
    wire n56703, n54602, n56904, n2;
    wire [31:0]\FRAME_MATCHER.i ;   // verilog/coms.v(116[11:12])
    
    wire n3, n2_adj_4620, n3_adj_4621, n56751, n7_adj_4622;
    wire [7:0]\data_in_frame[19] ;   // verilog/coms.v(97[12:25])
    
    wire n49097, n46832, n25607, n4623, n3_adj_4623, n2_adj_4624, 
        n3_adj_4625;
    wire [31:0]\FRAME_MATCHER.state ;   // verilog/coms.v(113[11:16])
    
    wire n36483, n7678, n7679;
    wire [31:0]\FRAME_MATCHER.state_31__N_2879 ;
    
    wire n5, n1, n57034, n36546, n6_c, n48306, n53225, n53226, 
        n5_adj_4626, n110, n24251, n50640;
    wire [31:0]\FRAME_MATCHER.state_31__N_2943 ;
    
    wire n60, n48404, n53259, n53258, n53195, n7680, n4_c, n49, 
        n48308, n11, n48310, n53196, n53274, n53273, n53318;
    wire [7:0]\data_in_frame[18] ;   // verilog/coms.v(97[12:25])
    
    wire n7681, n53319, n48368, \FRAME_MATCHER.rx_data_ready_prev , 
        n161, n53181, n53180, n53201, n36451, n48984, n53202, 
        n53280, n53279, n12, n48222, n48366, n45364, n27110, n49948, 
        n7682, n27217, n48314, n38, n3_adj_4627, n3_adj_4628, n48224, 
        n53307, n53306, n3_adj_4629, n49094, n160, n48470, n48478, 
        n3_adj_4630, n3_adj_4631, \FRAME_MATCHER.i_31__N_2845 , n39, 
        n27180, n4452, n12_adj_4632, n48220, n7_adj_4633, n3_adj_4634, 
        Kp_23__N_1098, n27862;
    wire [7:0]\data_in_frame[0] ;   // verilog/coms.v(97[12:25])
    
    wire n27863, n48216;
    wire [7:0]\data_in_frame[10] ;   // verilog/coms.v(97[12:25])
    
    wire n29376, n7683, n48214, n27304, n3_adj_4635, n4_adj_4636, 
        n24280, n48250, n7684, n14, n27268, n15, n27088, n3_adj_4637, 
        n3_adj_4638, n3_adj_4639, n48212, n16, n17, n27226, n10, 
        n3_adj_4640, n10_adj_4641, n14_adj_4642, n27255, n18, n20, 
        n15_adj_4643, n63_adj_4644, n20_adj_4645, n19, n6_adj_4646, 
        n53065, n16_adj_4648, n17_adj_4649, n63_adj_4650, n44, n42, 
        n3_adj_4651, n3_adj_4652, n3_adj_4653, n3_adj_4654, n48218, 
        n43, n41, n40, n39_adj_4655, n50, n45, n27108, n3_adj_4656, 
        n3_adj_4657, n3_adj_4658, n4599, n6_adj_4659, n3_adj_4660, 
        n2_adj_4661, n63_adj_4662, n6_adj_4663, n37171;
    wire [7:0]\data_in_frame[23] ;   // verilog/coms.v(97[12:25])
    
    wire n29487, n7685, n7686, n3_adj_4665, n31, n31_adj_4666, n23548, 
        n49218, n49221, n49399, n49608, n7687, n7688, Kp_23__N_1324, 
        n7_adj_4667, n49258;
    wire [7:0]\data_in_frame[7] ;   // verilog/coms.v(97[12:25])
    
    wire n49226, n28263, n52864, n27659, n12_adj_4668, n10_adj_4669, 
        n11_adj_4670, n9, n24549, n49064, n49021, n45758, n49206, 
        n10_adj_4671, Kp_23__N_1296, n4_adj_4672, n49038;
    wire [7:0]\data_in_frame[8]_c ;   // verilog/coms.v(97[12:25])
    
    wire n51412, n7_adj_4673, n27669, n49120, n28, n27962, n3_adj_4674, 
        n27954, n27604, n26, n27928, n46188, n27;
    wire [7:0]\data_in_frame[17] ;   // verilog/coms.v(97[12:25])
    
    wire n7689, n45804, n49688, n28082, n25, n52680, n48979, n48871, 
        n28716, n56895, n54596;
    wire [0:0]n6223;
    wire [2:0]r_SM_Main_2__N_3851;
    
    wire n49887, n7690, n7691, n53264, n53265, n53172, n7692, 
        n53171, n7693, n4_adj_4675, n4_adj_4676, tx_transmit_N_3748, 
        n36465, n7694, n49824, n7828, n8_adj_4677, n7695, n7696, 
        n49111, n49246, Kp_23__N_1602, n28406, n7673, n48993, n29631, 
        n29632, n49911, n27235, n50359, n51106, n29633, n8_adj_4678, 
        n46800, n49288, n49432, n52608, n52614, n45766, n51108, 
        Kp_23__N_1895, n51124, n52474, n48905, n50995, n52418, n49122, 
        n52422, n49699, n29634, n56715, n56898;
    wire [7:0]\data_in_frame[6] ;   // verilog/coms.v(97[12:25])
    
    wire n52916, n2_adj_4679, n49229, n28268, n49646, n52690, n52696, 
        n46727, n29635, n2_adj_4680, n29636, n49637, n29637, n19836, 
        n2_adj_4681, n2_adj_4682, n28527, n29638, n25500, n49060, 
        n2_adj_4683, n52934, n49495, n27307, n27223, n2_adj_4684, 
        n2_adj_4685, n2_adj_4686, n2_adj_4687, n49492, n51163, n4_adj_4688, 
        n27461, n52728, n28132, n49376, n27706, n2_adj_4689, n2_adj_4690, 
        n49543, n2_adj_4691, n2_adj_4692, n56955, n28138, n49373, 
        n2_adj_4693, n49667, n12_adj_4694, n49203, n2_adj_4695, n2_adj_4696, 
        n8_adj_4697, n29623, n29624, n2_adj_4698, n2_adj_4699, n53183, 
        n29625, n49466, n53184, n56799, n7_adj_4700, n53292, n53291, 
        n53207, n53208, n29626, n2_adj_4701, n53214, n53213, n29627, 
        n29628, n29629, n49652, n49328, n52836, n29630;
    wire [7:0]n9046;
    
    wire n28738, n29306, n26844, n27400, n46749, n49249, n49085, 
        n49117, n49032, Kp_23__N_1079, n28037, n49165, n28066, n49074, 
        n50429, n52566, n49664, n49517, n52574, n52588, n49522, 
        n52572, n52580, n49042, n52592, n49540, n52552, n49705, 
        n28303, n49702;
    wire [7:0]\data_out_frame[26] ;   // verilog/coms.v(98[12:26])
    wire [7:0]\data_out_frame[27] ;   // verilog/coms.v(98[12:26])
    
    wire n56892, n56928, n56835, n7_adj_4703, n56922, n56829, n7_adj_4704, 
        n49475, n56637, n54592, n56940, n15_adj_4705, n55901, n49525, 
        n28017, Kp_23__N_1209, n2_adj_4706, n3_adj_4707, n8_adj_4708, 
        n29615, n56916, n56823, n7_adj_4709, n27248, n48390, n56685, 
        n54598, n29616, n28030, n28050, n49162, n52708, n52710, 
        n27680, n14_adj_4710, n49569, n27577, n52716, n46699, n46413, 
        n52722, n50767, n46793, n29617, n52524, n49612, n52528, 
        n45864, n46708, n49234, n52530, n52536, n53228, n53229, 
        n49335, n28403, n52542, n29618, n49446, n49582, n48, n56847, 
        n7_adj_4711, n37153, n12_adj_4712, n49633, n27692, n49696, 
        n46673, n49331, n49599, n49451, n49578, n10_adj_4713, n48866, 
        n46738, n50764, n46718, n45830, n51314, n25418, n12_adj_4714, 
        n14_adj_4715, n45802, n52394, n46827, n49412, n46420, n51417, 
        n15_adj_4716, n48864, n10_adj_4717, n52740, n49590, n52670, 
        n4_adj_4718, n29619, n45939, n45874, n50279, n27557, Kp_23__N_1203, 
        n45811, n46666, n51092, n56886, n56889, Kp_23__N_1305, n56880, 
        n56883, n29620, n51209, n51166, n28807, n49352, n6_adj_4719, 
        n28069, n27599, n49457, n49138, n29621, n28020, n28539, 
        Kp_23__N_985, n45762, n4_adj_4720, n52650, n52900, n49252, 
        Kp_23__N_1206, n49237, n53192, n53193, n56856, n53190, n53189, 
        n53135, n53136, n56844, n53262, n53261, n53177, n53178, 
        n56838, n53244, n53243, n56841, n52948, n53198, n53199, 
        n56832, n53235, n53234, n53238, n53237, n45897, n52656, 
        n49395, n49605, n10_adj_4721, n49301, n28368, n28272, n27811, 
        n52658, n52664, n49384, n51154, n46852, n50744, n29622, 
        n28124, n55899, n46686, n45834, n49482, n52486, n52488, 
        n52490, n49682, n52494, n46682, n45512, n52500, n46917, 
        n46823, n52506, n49640, n52512, n46031, n52362, n52368, 
        n49596, n50545, n49180, n49370, n49340, n2_adj_4722, n3_adj_4723, 
        n50639, n50933, n2_adj_4724, n3_adj_4725, n49440, n45782, 
        n49035, n12_adj_4726, n50929, n49685, n50579, n27720, n46744, 
        n10_adj_4727, n49379, n46865, n51110, n2_adj_4728, n3_adj_4729, 
        Kp_23__N_1720, n49175, n49071, Kp_23__N_1103, n26302, n2_adj_4730, 
        n3_adj_4731, n2_adj_4732, n3_adj_4733, n49456, n49567, n51440, 
        n7_adj_4734, n46905, n27352, n49711, n49144, n27478, n49265, 
        n49418, n49615, n49443, n49444, n27554, n7_adj_4735, n49324, 
        n28079, n52382, n7_adj_4736, n7_adj_4737, n49581, n52762, 
        n50862, n56826, n36478, n49172, n49404, n53174, n43725, 
        n53175, n43724, n45884, n49460, n49010, n46834, n49415, 
        n6_adj_4738, n43723, n53322, n53321, n43722, n43721, n43720, 
        n43719, n8_adj_4739, n29607, n56820, n49046, n29608, n52632, 
        n56796, n29136, n29609, n46868, n49272, n29966, n29965, 
        n29964, n29963, n56748, n28_adj_4740, n32, n49670, n30, 
        n52640, n49478, n31_adj_4741, n50867, n52426, n52430, n29373, 
        n29372, n49690, n52436, n29, n49188, n45770, n49364, n10_adj_4742, 
        n56712, n56700, n50453, n49367, n56694, n56697, n27378, 
        n14_adj_4743, n56682, n10_adj_4744, n46458, n46753, n7677, 
        n7676, n7675, n7674, n48446, n48316, n29610, n29611, n28496, 
        n43718, n3746, n27455, n6_adj_4745, n49016, n43717, n43716, 
        n49618, n49693, n15_adj_4746, n43715, n49426, n14_adj_4747, 
        n27701, n43714, n49631, n46697, n29612, n49355, n46172, 
        n28322, n43713, n2_adj_4748, n43712, n49555, n28448, n12_adj_4749, 
        n49332, n1995, n27214, n29613, n46033, n49708, n36, n28151, 
        n46913, n14_adj_4751, n28176, n49321, n15_adj_4752, n50725, 
        n51346, n49673, n34, n29614, n26_adj_4753, n40_adj_4754, 
        n8_adj_4755, n29599, n24278, n27569, n38_adj_4756, n39_adj_4757, 
        n49593, n49304, n37, n29924, n2_adj_4758, n43711, n52970, 
        n29600, n6_adj_4759, n49275, n46808, n49255, n46403, n27715, 
        n49552, n49339, n6_adj_4760, n46729, n50817, n50449, n6_adj_4761, 
        n14_adj_4762, n48370, n10_adj_4763, n48364, n2_adj_4764, n43710, 
        n48362, n43709, n48360, n45838, n50641, n48358, n43708, 
        n46710, n10_adj_4765, n43707, n26774, n49559, n10_adj_4766, 
        n43706, n49624, n49621, n46821, n43705, n43704, n48356, 
        n48354, n48350, n43703, n46804, n27359, n48348, n43702, 
        n43701, n43700, n43699, n48346, n29601, n48456, n2_adj_4767, 
        n43698, n48458, n43697, n48460, n43696, n49534, n48462, 
        n29602, n43695, n48480, n43694, n43693, n36472, n49454, 
        n50240, n36474, n7_adj_4768, n43692, n36476, n48482, n1945, 
        n46695, n49284, n36480, n48484, n43691, n49655, n49318, 
        n48408, n48486, n27612, n52442, n43690, n43689, n43688, 
        n29603, n12_adj_4769, n28346, n46897, n46842, n46677, n49347, 
        n49268, n49240, n52448, n49295, n49223, n50375, n49350, 
        n49630, n49052, n27319, n49181, n6_adj_4770, n52454, n37148, 
        n37146, n37142, n37140, n37136, n7_adj_4771, n48454, n48452, 
        n7_adj_4772, n48450, n48448, n45750, n28180, n49472, n3_adj_4773, 
        n45914, n52460, n54597, n28196, n3_adj_4774, n46802, n3_adj_4775, 
        n3_adj_4776, n53222, n53223, n56670, n49197, n49184, n27424, 
        n49679, n49537, n16_adj_4777, n8_adj_4778, n49514, n53232, 
        n53231, n56673, n1168, n49649, n10_adj_4779, n27584, n53186, 
        n53187, n56664, n49392, n17_adj_4780, n26802, n49429, n28170, 
        n53241, n53240, n56667, n49546, n49280, n53401, n53399, 
        n7_adj_4781, n53317, n53315, n46848, n53155, n53153, n53149, 
        n53147, n53143, n53141, n49358, n52466, n49528, n49572, 
        n49178, n53164, n53162, n53159, n53160, n56646, n53252, 
        n53170, n53168, n53253, n56649, n53308, n52556, n51147, 
        n49261, n49409, n29604, n49498, n28573, n49661, n6_adj_4782, 
        n6_adj_4783, n46816, n27894, n49091, n46370, n28296, n49147, 
        n1191, n49200, n49135, n28318, n27915, n38_adj_4784, n28_adj_4785, 
        n29605, n13, n11_adj_4786, n51468, n49107, n49502, n51399, 
        n49658, n6_adj_4787, n27335, n50291, n28_adj_4788, n26_adj_4789, 
        n29606, n1169, n10_adj_4790, n56634, n49298, n49562, n49531, 
        n27_adj_4791, n6_adj_4792, n25_adj_4793, n27747, n12_adj_4794, 
        n46894, n27785, n26777, n27890, n49168, n10_adj_4795, n29787, 
        n29786, n29781, n46693, n29780, n29779, n29778, n29777, 
        n29776, n29775, n29774, n29773, n29772, n29771, n29770, 
        n29769, n29768, n29767, n29766, n29765, n29764, n29763, 
        n29762, n29761, n29760, n29757, n29756, n29755, n29754, 
        n29753, n29752, n29751, n29750, n29749, n29748, n29747, 
        n29746, n29745, n29744, n29743, n29742, n29741, n29740, 
        n29739, n29738, n29737, n29736, n29735, n29734, n29733, 
        n29732, n29731, n29730, n29729, n29728, n29727, n29726, 
        n29725, n29724, n29723, n29722, n29721, n29720, n29719, 
        n29718, n29717, n29716, n29715, n29714, n29713, n49566, 
        n29712, n29711, n29710, n29709, n29708, n29707, n29706, 
        n29705, n29704, n29703, n29702, n29701, n29700, n29699, 
        n29698, n29697, n29695, n6_adj_4796, n29694, n29693, n29692, 
        n29691, n29690, n29689, n29688, n29687, n29686, n29685, 
        n29684, n29683, n29682, n29681, n29680, n29679, n29678, 
        n29677, n29676, n29675, n29674, n29673, n29672, n29671, 
        n29670, n29669, n29668, n29667, n29666, n56976, n29665, 
        n29664, n29663, n29662, n29661, n29660, n29659, n29658, 
        n29657, n29656, n29655, n29654, n29653, n29652, n29651, 
        n29650, n29649, n29648, n29647, n29646, n29645, n29644, 
        n29643, n29642, n29641, n29640, n29639, n8_adj_4797, n29591, 
        n29598, n29597, n29596, n29595, n29594, n29593, n29592, 
        n29590, n29589, n29588, n29587, n29586, n29585, n29584, 
        n29583, n29582;
    wire [7:0]\data_in_frame[22] ;   // verilog/coms.v(97[12:25])
    
    wire n29581, n29580, n29579, n29578, n29577, n29576, n29575, 
        n29574, n29573, n29572, n56979, n49082, n75, n10_adj_4798, 
        n56961, n49151, n48970, n49342, n57052, n50_adj_4799, n46844, 
        n49549, n49132, n46915, n45836, n12_adj_4800, n49602, n49126, 
        n27535, n27922, n1563, n49024, n49505, n49114, n10_adj_4801, 
        n49511, n49129, n10_adj_4802, n14_adj_4803, n49307, n6_adj_4804, 
        n49067, n12_adj_4805, n6_adj_4806, n49489, n49508, n50853, 
        n27323, n27906, n4_adj_4807, n54603, n56934, n45980, n12_adj_4808, 
        n45752, n50716, n35, n49469, n34_adj_4809, n51236, n8_adj_4810, 
        n40_adj_4811, n38_adj_4812, n52400, n42_adj_4813, n37_adj_4814, 
        n49013, n10_adj_4815, n53163, n16_adj_4816, n15_adj_4817, 
        n17_adj_4818, n33, n52402, n41_adj_4819, n27347, n49191, 
        n51469, n43_adj_4820, n49243, n40_adj_4821, n46, n8_adj_4822, 
        n49212, n39_adj_4823, n47, n8_adj_4824, n50913, n52404, 
        n7_adj_4825, n49643, n54601, n52856, n1519, n1516, n46186, 
        n52408, n27339, n54599, n51299, n49057, n52862, n1193, 
        n27959, n14_adj_4826, n15_adj_4827, n12_adj_4828, n49101, 
        n56970, n52412, n49028, n12_adj_4829, n27938, n12_adj_4830, 
        n52750, n10_adj_4831, n14_adj_4832, n51304, n45844, n12_adj_4833, 
        n56973, n52414, n56964, n56967, n26_adj_4834, n52972, n23, 
        n22, n4_adj_4835, n52974, n32_adj_4836, n27_adj_4837, n48882, 
        n52744, n53040, n24055, n53142, n56958, n53154, n53148, 
        n28382, n52774, n46100, n12_adj_4838, n56952;
    
    SB_LUT4 n56910_bdd_4_lut (.I0(n56910), .I1(n56859), .I2(n7_c), .I3(byte_transmit_counter[4]), 
            .O(tx_data[2]));
    defparam n56910_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_41027 (.I0(byte_transmit_counter[3]), 
            .I1(n56703), .I2(n54602), .I3(byte_transmit_counter[4]), .O(n56904));
    defparam byte_transmit_counter_3__bdd_4_lut_41027.LUT_INIT = 16'he4aa;
    SB_DFF deadband_i0_i22 (.Q(deadband[22]), .C(clk16MHz), .D(n29523));   // verilog/coms.v(128[12] 303[6])
    SB_DFF deadband_i0_i23 (.Q(deadband[23]), .C(clk16MHz), .D(n29522));   // verilog/coms.v(128[12] 303[6])
    SB_DFF Kp_i1 (.Q(\Kp[1] ), .C(clk16MHz), .D(n29521));   // verilog/coms.v(128[12] 303[6])
    SB_DFF Kp_i2 (.Q(\Kp[2] ), .C(clk16MHz), .D(n29520));   // verilog/coms.v(128[12] 303[6])
    SB_DFF Kp_i3 (.Q(\Kp[3] ), .C(clk16MHz), .D(n29519));   // verilog/coms.v(128[12] 303[6])
    SB_DFFSS \FRAME_MATCHER.i_i22  (.Q(\FRAME_MATCHER.i [22]), .C(clk16MHz), 
            .D(n2), .S(n3));   // verilog/coms.v(128[12] 303[6])
    SB_DFFSS \FRAME_MATCHER.i_i21  (.Q(\FRAME_MATCHER.i [21]), .C(clk16MHz), 
            .D(n2_adj_4620), .S(n3_adj_4621));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 n56904_bdd_4_lut (.I0(n56904), .I1(n56751), .I2(n7_adj_4622), 
            .I3(byte_transmit_counter[4]), .O(tx_data[1]));
    defparam n56904_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF Kp_i4 (.Q(\Kp[4] ), .C(clk16MHz), .D(n29518));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i3_4_lut (.I0(\data_in_frame[19] [3]), .I1(n49097), .I2(n46832), 
            .I3(\data_in_frame[19] [2]), .O(n25607));
    defparam i3_4_lut.LUT_INIT = 16'h9669;
    SB_LUT4 select_713_Select_13_i3_2_lut (.I0(\FRAME_MATCHER.i [13]), .I1(n4623), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4623));
    defparam select_713_Select_13_i3_2_lut.LUT_INIT = 16'h8888;
    SB_DFFSS \FRAME_MATCHER.i_i0  (.Q(\FRAME_MATCHER.i [0]), .C(clk16MHz), 
            .D(n2_adj_4624), .S(n3_adj_4625));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 mux_2112_i6_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n36483), 
            .I2(\data_in_frame[3] [5]), .I3(\data_in_frame[19] [5]), .O(n7678));
    defparam mux_2112_i6_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 mux_2112_i7_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n36483), 
            .I2(\data_in_frame[3] [6]), .I3(\data_in_frame[19] [6]), .O(n7679));
    defparam mux_2112_i7_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_4_lut (.I0(n63), .I1(n3303), .I2(n27219), .I3(\FRAME_MATCHER.state_31__N_2879 [1]), 
            .O(n5));
    defparam i1_4_lut.LUT_INIT = 16'h5f5d;
    SB_LUT4 i3_4_lut_adj_955 (.I0(n5), .I1(\FRAME_MATCHER.state_31__N_2879 [1]), 
            .I2(n1), .I3(n48947), .O(n57034));
    defparam i3_4_lut_adj_955.LUT_INIT = 16'hfefa;
    SB_LUT4 i1_4_lut_adj_956 (.I0(\FRAME_MATCHER.state_31__N_2879 [1]), .I1(n36546), 
            .I2(n48957), .I3(n6_c), .O(n48306));
    defparam i1_4_lut_adj_956.LUT_INIT = 16'ha8a0;
    SB_LUT4 i37395_3_lut (.I0(\data_out_frame[16] [3]), .I1(\data_out_frame[17] [3]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n53225));
    defparam i37395_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i37396_3_lut (.I0(\data_out_frame[18] [3]), .I1(\data_out_frame[19] [3]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n53226));
    defparam i37396_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2_4_lut (.I0(n5_adj_4626), .I1(n27218), .I2(n110), .I3(n24251), 
            .O(n50640));
    defparam i2_4_lut.LUT_INIT = 16'hfbfa;
    SB_LUT4 i1_4_lut_adj_957 (.I0(\FRAME_MATCHER.state_31__N_2943 [3]), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(n60), .I3(n50640), .O(n48404));
    defparam i1_4_lut_adj_957.LUT_INIT = 16'hce0a;
    SB_LUT4 i37429_3_lut (.I0(\data_out_frame[22] [3]), .I1(\data_out_frame[23] [3]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n53259));
    defparam i37429_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i37428_3_lut (.I0(\data_out_frame[20] [3]), .I1(\data_out_frame[21] [3]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n53258));
    defparam i37428_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i37365_3_lut (.I0(\data_out_frame[16] [2]), .I1(\data_out_frame[17] [2]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n53195));
    defparam i37365_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_2112_i8_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n36483), 
            .I2(\data_in_frame[3] [7]), .I3(\data_in_frame[19] [7]), .O(n7680));
    defparam mux_2112_i8_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_3_lut (.I0(\FRAME_MATCHER.state[3] ), .I1(n4_c), .I2(n49), 
            .I3(GND_net), .O(n48308));
    defparam i1_3_lut.LUT_INIT = 16'ha8a8;
    SB_LUT4 i1_2_lut (.I0(\FRAME_MATCHER.state [4]), .I1(n11), .I2(GND_net), 
            .I3(GND_net), .O(n48310));
    defparam i1_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i37366_3_lut (.I0(\data_out_frame[18] [2]), .I1(\data_out_frame[19] [2]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n53196));
    defparam i37366_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i37444_3_lut (.I0(\data_out_frame[22] [2]), .I1(\data_out_frame[23] [2]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n53274));
    defparam i37444_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i37443_3_lut (.I0(\data_out_frame[20] [2]), .I1(\data_out_frame[21] [2]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n53273));
    defparam i37443_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i37488_3_lut (.I0(\data_out_frame[16] [1]), .I1(\data_out_frame[17] [1]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n53318));
    defparam i37488_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_2112_i9_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n36483), 
            .I2(\data_in_frame[2] [0]), .I3(\data_in_frame[18] [0]), .O(n7681));
    defparam mux_2112_i9_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i37489_3_lut (.I0(\data_out_frame[18] [1]), .I1(\data_out_frame[19] [1]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n53319));
    defparam i37489_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_958 (.I0(\FRAME_MATCHER.state [5]), .I1(n11), .I2(GND_net), 
            .I3(GND_net), .O(n48368));
    defparam i1_2_lut_adj_958.LUT_INIT = 16'h8888;
    SB_LUT4 i14_2_lut (.I0(rx_data_ready), .I1(\FRAME_MATCHER.rx_data_ready_prev ), 
            .I2(GND_net), .I3(GND_net), .O(n161));   // verilog/coms.v(154[9:50])
    defparam i14_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i37351_3_lut (.I0(\data_out_frame[22] [1]), .I1(\data_out_frame[23] [1]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n53181));
    defparam i37351_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i37350_3_lut (.I0(\data_out_frame[20] [1]), .I1(\data_out_frame[21] [1]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n53180));
    defparam i37350_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i37371_3_lut (.I0(\data_out_frame[16] [0]), .I1(\data_out_frame[17] [0]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n53201));
    defparam i37371_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3_4_lut_adj_959 (.I0(n36451), .I1(\FRAME_MATCHER.i [5]), .I2(\FRAME_MATCHER.i [4]), 
            .I3(\FRAME_MATCHER.i [3]), .O(n48984));   // verilog/coms.v(155[7:23])
    defparam i3_4_lut_adj_959.LUT_INIT = 16'hffdf;
    SB_LUT4 i37372_3_lut (.I0(\data_out_frame[18] [0]), .I1(\data_out_frame[19] [0]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n53202));
    defparam i37372_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i37450_3_lut (.I0(\data_out_frame[22] [0]), .I1(\data_out_frame[23] [0]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n53280));
    defparam i37450_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i37449_3_lut (.I0(\data_out_frame[20] [0]), .I1(\data_out_frame[21] [0]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n53279));
    defparam i37449_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_960 (.I0(\FRAME_MATCHER.state [6]), .I1(n12), .I2(GND_net), 
            .I3(GND_net), .O(n48222));
    defparam i1_2_lut_adj_960.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_961 (.I0(\FRAME_MATCHER.state [7]), .I1(n11), .I2(GND_net), 
            .I3(GND_net), .O(n48366));
    defparam i1_2_lut_adj_961.LUT_INIT = 16'h8888;
    SB_LUT4 i34187_4_lut (.I0(\FRAME_MATCHER.i [31]), .I1(n45364), .I2(n27110), 
            .I3(\FRAME_MATCHER.state [2]), .O(n49948));
    defparam i34187_4_lut.LUT_INIT = 16'h5044;
    SB_LUT4 mux_2112_i10_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n36483), 
            .I2(\data_in_frame[2] [1]), .I3(\data_in_frame[18] [1]), .O(n7682));
    defparam mux_2112_i10_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_4_lut_adj_962 (.I0(n4_c), .I1(n49948), .I2(n27217), .I3(n22875), 
            .O(n11));
    defparam i1_4_lut_adj_962.LUT_INIT = 16'habaa;
    SB_LUT4 i1_2_lut_adj_963 (.I0(\FRAME_MATCHER.state [8]), .I1(n11), .I2(GND_net), 
            .I3(GND_net), .O(n48314));
    defparam i1_2_lut_adj_963.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut_adj_964 (.I0(n38), .I1(n27217), .I2(n3_adj_4627), 
            .I3(n3_adj_4628), .O(n12));
    defparam i1_4_lut_adj_964.LUT_INIT = 16'hbbba;
    SB_LUT4 i1_2_lut_adj_965 (.I0(\FRAME_MATCHER.state [9]), .I1(n12), .I2(GND_net), 
            .I3(GND_net), .O(n48224));
    defparam i1_2_lut_adj_965.LUT_INIT = 16'h8888;
    SB_LUT4 i37477_3_lut (.I0(\data_out_frame[6] [0]), .I1(\data_out_frame[7] [0]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n53307));
    defparam i37477_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i37476_3_lut (.I0(\data_out_frame[4] [0]), .I1(\data_out_frame[5] [0]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n53306));
    defparam i37476_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF Kp_i5 (.Q(\Kp[5] ), .C(clk16MHz), .D(n29516));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 select_713_Select_14_i3_2_lut (.I0(\FRAME_MATCHER.i [14]), .I1(n4623), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4629));
    defparam select_713_Select_14_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut_adj_966 (.I0(\data_in_frame[4] [7]), .I1(\data_in_frame[3] [1]), 
            .I2(\data_in_frame[5] [2]), .I3(\data_in_frame[5] [1]), .O(n49094));   // verilog/coms.v(86[17:70])
    defparam i1_4_lut_adj_966.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_967 (.I0(\FRAME_MATCHER.state [14]), .I1(n160), 
            .I2(GND_net), .I3(GND_net), .O(n48470));
    defparam i1_2_lut_adj_967.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_968 (.I0(\FRAME_MATCHER.state [15]), .I1(n160), 
            .I2(GND_net), .I3(GND_net), .O(n48478));
    defparam i1_2_lut_adj_968.LUT_INIT = 16'h8888;
    SB_LUT4 select_713_Select_12_i3_2_lut (.I0(\FRAME_MATCHER.i [12]), .I1(n4623), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4630));
    defparam select_713_Select_12_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_713_Select_10_i3_2_lut (.I0(\FRAME_MATCHER.i [10]), .I1(n4623), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4631));
    defparam select_713_Select_10_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i163_4_lut (.I0(\FRAME_MATCHER.i_31__N_2845 ), .I1(n39), .I2(n27180), 
            .I3(n4452), .O(n160));   // verilog/coms.v(116[11:12])
    defparam i163_4_lut.LUT_INIT = 16'hccec;
    SB_LUT4 i1_2_lut_adj_969 (.I0(\FRAME_MATCHER.state [16]), .I1(n12_adj_4632), 
            .I2(GND_net), .I3(GND_net), .O(n48220));
    defparam i1_2_lut_adj_969.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_970 (.I0(\FRAME_MATCHER.state [16]), .I1(n160), 
            .I2(GND_net), .I3(GND_net), .O(n7_adj_4633));   // verilog/coms.v(213[5:16])
    defparam i1_2_lut_adj_970.LUT_INIT = 16'h8888;
    SB_LUT4 select_713_Select_9_i3_2_lut (.I0(\FRAME_MATCHER.i [9]), .I1(n4623), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4634));
    defparam select_713_Select_9_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_3_lut_adj_971 (.I0(Kp_23__N_1098), .I1(n27862), .I2(\data_in_frame[0] [7]), 
            .I3(GND_net), .O(n27863));   // verilog/coms.v(72[16:69])
    defparam i1_3_lut_adj_971.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_972 (.I0(\FRAME_MATCHER.state [18]), .I1(n12_adj_4632), 
            .I2(GND_net), .I3(GND_net), .O(n48216));   // verilog/coms.v(116[11:12])
    defparam i1_2_lut_adj_972.LUT_INIT = 16'h8888;
    SB_LUT4 i18377_3_lut (.I0(PWMLimit[0]), .I1(\data_in_frame[10] [0]), 
            .I2(n50654), .I3(GND_net), .O(n29376));
    defparam i18377_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_2112_i11_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n36483), 
            .I2(\data_in_frame[2] [2]), .I3(\data_in_frame[18] [2]), .O(n7683));
    defparam mux_2112_i11_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_adj_973 (.I0(\FRAME_MATCHER.state [20]), .I1(n12_adj_4632), 
            .I2(GND_net), .I3(GND_net), .O(n48214));   // verilog/coms.v(116[11:12])
    defparam i1_2_lut_adj_973.LUT_INIT = 16'h8888;
    SB_LUT4 i22594_4_lut (.I0(\FRAME_MATCHER.i [3]), .I1(\FRAME_MATCHER.i [31]), 
            .I2(n27304), .I3(\FRAME_MATCHER.i [4]), .O(n4452));   // verilog/coms.v(260[9:58])
    defparam i22594_4_lut.LUT_INIT = 16'h3230;
    SB_LUT4 select_713_Select_8_i3_2_lut (.I0(\FRAME_MATCHER.i [8]), .I1(n4623), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4635));
    defparam select_713_Select_8_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i22593_2_lut (.I0(n27110), .I1(\FRAME_MATCHER.i [31]), .I2(GND_net), 
            .I3(GND_net), .O(n3303));   // verilog/coms.v(228[9:54])
    defparam i22593_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1_2_lut_adj_974 (.I0(n5_adj_4626), .I1(n38), .I2(GND_net), 
            .I3(GND_net), .O(n4_adj_4636));
    defparam i1_2_lut_adj_974.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_975 (.I0(\FRAME_MATCHER.i_31__N_2845 ), .I1(n4452), 
            .I2(GND_net), .I3(GND_net), .O(n48947));
    defparam i1_2_lut_adj_975.LUT_INIT = 16'h2222;
    SB_LUT4 i1_4_lut_adj_976 (.I0(\FRAME_MATCHER.state [22]), .I1(n24280), 
            .I2(n4_adj_4636), .I3(n27218), .O(n48250));
    defparam i1_4_lut_adj_976.LUT_INIT = 16'ha0a8;
    SB_LUT4 i1_2_lut_adj_977 (.I0(\FRAME_MATCHER.state [2]), .I1(n27217), 
            .I2(GND_net), .I3(GND_net), .O(n27219));   // verilog/coms.v(223[5:21])
    defparam i1_2_lut_adj_977.LUT_INIT = 16'hdddd;
    SB_LUT4 mux_2112_i12_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n36483), 
            .I2(\data_in_frame[2] [3]), .I3(\data_in_frame[18] [3]), .O(n7684));
    defparam mux_2112_i12_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5_3_lut (.I0(\data_in[0] [3]), .I1(\data_in[1] [4]), .I2(\data_in[1] [5]), 
            .I3(GND_net), .O(n14));
    defparam i5_3_lut.LUT_INIT = 16'hdfdf;
    SB_LUT4 i6_4_lut (.I0(\data_in[0] [6]), .I1(n27268), .I2(\data_in[2] [4]), 
            .I3(\data_in[1] [0]), .O(n15));
    defparam i6_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i8_4_lut (.I0(n15), .I1(\data_in[3] [0]), .I2(n14), .I3(\data_in[2] [2]), 
            .O(n27088));
    defparam i8_4_lut.LUT_INIT = 16'hfbff;
    SB_LUT4 select_713_Select_7_i3_2_lut (.I0(\FRAME_MATCHER.i [7]), .I1(n4623), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4637));
    defparam select_713_Select_7_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_713_Select_6_i3_2_lut (.I0(\FRAME_MATCHER.i [6]), .I1(n4623), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4638));
    defparam select_713_Select_6_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_713_Select_15_i3_2_lut (.I0(\FRAME_MATCHER.i [15]), .I1(n4623), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4639));
    defparam select_713_Select_15_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_978 (.I0(\FRAME_MATCHER.state [24]), .I1(n12_adj_4632), 
            .I2(GND_net), .I3(GND_net), .O(n48212));   // verilog/coms.v(116[11:12])
    defparam i1_2_lut_adj_978.LUT_INIT = 16'h8888;
    SB_LUT4 i6_4_lut_adj_979 (.I0(\data_in[1] [3]), .I1(\data_in[0] [1]), 
            .I2(\data_in[3] [2]), .I3(\data_in[0] [5]), .O(n16));
    defparam i6_4_lut_adj_979.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_4_lut (.I0(\data_in[2] [6]), .I1(\data_in[2] [5]), .I2(\data_in[2] [0]), 
            .I3(\data_in[1] [2]), .O(n17));
    defparam i7_4_lut.LUT_INIT = 16'hfffd;
    SB_LUT4 i9_4_lut (.I0(n17), .I1(\data_in[1] [6]), .I2(n16), .I3(\data_in[3] [7]), 
            .O(n27226));
    defparam i9_4_lut.LUT_INIT = 16'hfbff;
    SB_LUT4 i4_4_lut (.I0(\data_in[1] [7]), .I1(\data_in[0] [0]), .I2(\data_in[1] [1]), 
            .I3(\data_in[0] [4]), .O(n10));
    defparam i4_4_lut.LUT_INIT = 16'hfdff;
    SB_LUT4 i5_3_lut_adj_980 (.I0(\data_in[3] [4]), .I1(n10), .I2(\data_in[2] [7]), 
            .I3(GND_net), .O(n27268));
    defparam i5_3_lut_adj_980.LUT_INIT = 16'hdfdf;
    SB_LUT4 select_713_Select_16_i3_2_lut (.I0(\FRAME_MATCHER.i [16]), .I1(n4623), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4640));
    defparam select_713_Select_16_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_2_lut (.I0(\data_in[2] [3]), .I1(\data_in[3] [5]), .I2(GND_net), 
            .I3(GND_net), .O(n10_adj_4641));
    defparam i2_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i6_4_lut_adj_981 (.I0(\data_in[0] [2]), .I1(\data_in[3] [3]), 
            .I2(\data_in[3] [1]), .I3(\data_in[0] [7]), .O(n14_adj_4642));
    defparam i6_4_lut_adj_981.LUT_INIT = 16'hfeff;
    SB_LUT4 i7_4_lut_adj_982 (.I0(\data_in[3] [6]), .I1(n14_adj_4642), .I2(n10_adj_4641), 
            .I3(\data_in[2] [1]), .O(n27255));
    defparam i7_4_lut_adj_982.LUT_INIT = 16'hfffd;
    SB_LUT4 i7_4_lut_adj_983 (.I0(\data_in[2] [4]), .I1(n27255), .I2(\data_in[1] [5]), 
            .I3(n27268), .O(n18));
    defparam i7_4_lut_adj_983.LUT_INIT = 16'hfffd;
    SB_LUT4 i9_4_lut_adj_984 (.I0(\data_in[0] [6]), .I1(n18), .I2(\data_in[3] [0]), 
            .I3(n27226), .O(n20));
    defparam i9_4_lut_adj_984.LUT_INIT = 16'hfffd;
    SB_LUT4 i4_2_lut (.I0(\data_in[1] [0]), .I1(\data_in[0] [3]), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_4643));
    defparam i4_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i10_4_lut (.I0(n15_adj_4643), .I1(n20), .I2(\data_in[2] [2]), 
            .I3(\data_in[1] [4]), .O(n63_adj_4644));
    defparam i10_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i8_4_lut_adj_985 (.I0(n27255), .I1(\data_in[1] [3]), .I2(n27088), 
            .I3(\data_in[1] [2]), .O(n20_adj_4645));
    defparam i8_4_lut_adj_985.LUT_INIT = 16'hfbff;
    SB_LUT4 i7_4_lut_adj_986 (.I0(\data_in[2] [6]), .I1(\data_in[1] [6]), 
            .I2(\data_in[3] [7]), .I3(\data_in[0] [1]), .O(n19));
    defparam i7_4_lut_adj_986.LUT_INIT = 16'hfeff;
    SB_LUT4 i1_2_lut_adj_987 (.I0(n24280), .I1(\FRAME_MATCHER.state [2]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_4646));   // verilog/coms.v(116[11:12])
    defparam i1_2_lut_adj_987.LUT_INIT = 16'h2222;
    SB_LUT4 i1_4_lut_adj_988 (.I0(n38), .I1(n27217), .I2(n3_adj_4628), 
            .I3(n6_adj_4646), .O(n12_adj_4632));   // verilog/coms.v(116[11:12])
    defparam i1_4_lut_adj_988.LUT_INIT = 16'hbbba;
    SB_LUT4 i37299_4_lut (.I0(\data_in[2] [5]), .I1(\data_in[2] [0]), .I2(\data_in[3] [2]), 
            .I3(\data_in[0] [5]), .O(n53065));
    defparam i37299_4_lut.LUT_INIT = 16'h8000;
    SB_DFF Kp_i6 (.Q(\Kp[6] ), .C(clk16MHz), .D(n29515));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i11_3_lut (.I0(n53065), .I1(n19), .I2(n20_adj_4645), .I3(GND_net), 
            .O(n63_adj_6));
    defparam i11_3_lut.LUT_INIT = 16'hfdfd;
    SB_LUT4 i6_4_lut_adj_989 (.I0(\data_in[3] [6]), .I1(\data_in[0] [7]), 
            .I2(\data_in[2] [1]), .I3(n27088), .O(n16_adj_4648));
    defparam i6_4_lut_adj_989.LUT_INIT = 16'hffef;
    SB_LUT4 i7_4_lut_adj_990 (.I0(n27226), .I1(\data_in[2] [3]), .I2(\data_in[0] [2]), 
            .I3(\data_in[3] [1]), .O(n17_adj_4649));
    defparam i7_4_lut_adj_990.LUT_INIT = 16'hbfff;
    SB_LUT4 i9_4_lut_adj_991 (.I0(n17_adj_4649), .I1(\data_in[3] [5]), .I2(n16_adj_4648), 
            .I3(\data_in[3] [3]), .O(n63_adj_4650));
    defparam i9_4_lut_adj_991.LUT_INIT = 16'hfbff;
    SB_LUT4 i2_3_lut (.I0(n63_adj_4650), .I1(n63_adj_6), .I2(n63_adj_4644), 
            .I3(GND_net), .O(n22875));   // verilog/coms.v(158[6] 160[9])
    defparam i2_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i18_4_lut (.I0(\FRAME_MATCHER.i [30]), .I1(\FRAME_MATCHER.i [21]), 
            .I2(\FRAME_MATCHER.i [24]), .I3(\FRAME_MATCHER.i [17]), .O(n44));
    defparam i18_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut (.I0(\FRAME_MATCHER.i [29]), .I1(\FRAME_MATCHER.i [6]), 
            .I2(\FRAME_MATCHER.i [18]), .I3(\FRAME_MATCHER.i [23]), .O(n42));
    defparam i16_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 select_713_Select_5_i3_2_lut (.I0(\FRAME_MATCHER.i [5]), .I1(n4623), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4651));
    defparam select_713_Select_5_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_713_Select_17_i3_2_lut (.I0(\FRAME_MATCHER.i [17]), .I1(n4623), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4652));
    defparam select_713_Select_17_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_713_Select_18_i3_2_lut (.I0(\FRAME_MATCHER.i [18]), .I1(n4623), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4653));
    defparam select_713_Select_18_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_713_Select_4_i3_2_lut (.I0(\FRAME_MATCHER.i [4]), .I1(n4623), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4654));
    defparam select_713_Select_4_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_992 (.I0(\FRAME_MATCHER.state [26]), .I1(n12_adj_4632), 
            .I2(GND_net), .I3(GND_net), .O(n48218));
    defparam i1_2_lut_adj_992.LUT_INIT = 16'h8888;
    SB_LUT4 i17_4_lut (.I0(\FRAME_MATCHER.i [7]), .I1(\FRAME_MATCHER.i [20]), 
            .I2(\FRAME_MATCHER.i [12]), .I3(\FRAME_MATCHER.i [14]), .O(n43));
    defparam i17_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut (.I0(\FRAME_MATCHER.i [22]), .I1(\FRAME_MATCHER.i [11]), 
            .I2(\FRAME_MATCHER.i [26]), .I3(\FRAME_MATCHER.i [16]), .O(n41));
    defparam i15_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i14_4_lut (.I0(\FRAME_MATCHER.i [13]), .I1(\FRAME_MATCHER.i [15]), 
            .I2(\FRAME_MATCHER.i [10]), .I3(\FRAME_MATCHER.i [28]), .O(n40));
    defparam i14_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_2_lut (.I0(\FRAME_MATCHER.i [9]), .I1(\FRAME_MATCHER.i [27]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_4655));
    defparam i13_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i24_4_lut (.I0(n41), .I1(n43), .I2(n42), .I3(n44), .O(n50));
    defparam i24_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i19_4_lut (.I0(\FRAME_MATCHER.i [8]), .I1(\FRAME_MATCHER.i [25]), 
            .I2(\FRAME_MATCHER.i [5]), .I3(\FRAME_MATCHER.i [19]), .O(n45));
    defparam i19_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i25_4_lut (.I0(n45), .I1(n50), .I2(n39_adj_4655), .I3(n40), 
            .O(n27304));
    defparam i25_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_adj_993 (.I0(\FRAME_MATCHER.i [4]), .I1(n27304), .I2(GND_net), 
            .I3(GND_net), .O(n27108));   // verilog/coms.v(155[7:23])
    defparam i1_2_lut_adj_993.LUT_INIT = 16'heeee;
    SB_LUT4 select_713_Select_19_i3_2_lut (.I0(\FRAME_MATCHER.i [19]), .I1(n4623), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4656));
    defparam select_713_Select_19_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_713_Select_3_i3_2_lut (.I0(\FRAME_MATCHER.i [3]), .I1(n4623), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4657));
    defparam select_713_Select_3_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_713_Select_2_i3_2_lut (.I0(\FRAME_MATCHER.i [2]), .I1(n4623), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4658));
    defparam select_713_Select_2_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i111_2_lut (.I0(n4599), .I1(n22875), .I2(GND_net), .I3(GND_net), 
            .O(n38));
    defparam i111_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_2_lut_adj_994 (.I0(\FRAME_MATCHER.i [2]), .I1(\FRAME_MATCHER.i [3]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_4659));
    defparam i2_2_lut_adj_994.LUT_INIT = 16'heeee;
    SB_LUT4 i3_4_lut_adj_995 (.I0(\FRAME_MATCHER.i [0]), .I1(n6_adj_4659), 
            .I2(n27108), .I3(\FRAME_MATCHER.i [1]), .O(n45364));
    defparam i3_4_lut_adj_995.LUT_INIT = 16'hfefc;
    SB_LUT4 select_713_Select_1_i3_2_lut (.I0(\FRAME_MATCHER.i [1]), .I1(n4623), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4660));
    defparam select_713_Select_1_i3_2_lut.LUT_INIT = 16'h8888;
    SB_DFF Kp_i7 (.Q(\Kp[7] ), .C(clk16MHz), .D(n29514));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i4_4_lut_adj_996 (.I0(n60), .I1(n2_adj_4661), .I2(n63_adj_4662), 
            .I3(n6_adj_4663), .O(n4599));
    defparam i4_4_lut_adj_996.LUT_INIT = 16'h8000;
    SB_LUT4 i1_2_lut_adj_997 (.I0(\FRAME_MATCHER.state [2]), .I1(n27217), 
            .I2(GND_net), .I3(GND_net), .O(n27218));   // verilog/coms.v(152[5:27])
    defparam i1_2_lut_adj_997.LUT_INIT = 16'heeee;
    SB_LUT4 i15407_3_lut_4_lut (.I0(n37171), .I1(n48984), .I2(rx_data[3]), 
            .I3(\data_in_frame[23] [3]), .O(n29487));
    defparam i15407_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 mux_2112_i13_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n36483), 
            .I2(\data_in_frame[2] [4]), .I3(\data_in_frame[18] [4]), .O(n7685));
    defparam mux_2112_i13_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i22455_3_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n63_adj_4644), 
            .I2(n63_adj_4650), .I3(GND_net), .O(n122));   // verilog/coms.v(140[4] 142[7])
    defparam i22455_3_lut.LUT_INIT = 16'hb3b3;
    SB_LUT4 select_751_Select_2_i8_3_lut (.I0(n122), .I1(n4599), .I2(n63_adj_6), 
            .I3(GND_net), .O(n8));
    defparam select_751_Select_2_i8_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 select_751_Select_2_i7_4_lut (.I0(n122), .I1(\FRAME_MATCHER.i_31__N_2845 ), 
            .I2(n4452), .I3(n63_adj_6), .O(n7));
    defparam select_751_Select_2_i7_4_lut.LUT_INIT = 16'hc8c0;
    SB_LUT4 mux_2112_i14_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n36483), 
            .I2(\data_in_frame[2] [5]), .I3(\data_in_frame[18] [5]), .O(n7686));
    defparam mux_2112_i14_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 select_713_Select_20_i3_2_lut (.I0(\FRAME_MATCHER.i [20]), .I1(n4623), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4665));
    defparam select_713_Select_20_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i4694_3_lut (.I0(n31), .I1(n31_adj_4666), .I2(\FRAME_MATCHER.state [1]), 
            .I3(GND_net), .O(n23548));
    defparam i4694_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_998 (.I0(n49218), .I1(n49221), .I2(\data_in_frame[1] [4]), 
            .I3(\data_in_frame[5] [6]), .O(n49399));
    defparam i1_4_lut_adj_998.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_999 (.I0(\data_in_frame[8] [0]), .I1(n49399), .I2(GND_net), 
            .I3(GND_net), .O(n49608));
    defparam i1_2_lut_adj_999.LUT_INIT = 16'h6666;
    SB_LUT4 mux_2112_i15_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n36483), 
            .I2(\data_in_frame[2] [6]), .I3(\data_in_frame[18] [6]), .O(n7687));
    defparam mux_2112_i15_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 mux_2112_i16_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n36483), 
            .I2(\data_in_frame[2] [7]), .I3(\data_in_frame[18] [7]), .O(n7688));
    defparam mux_2112_i16_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2_2_lut_adj_1000 (.I0(\data_in_frame[8] [7]), .I1(Kp_23__N_1324), 
            .I2(GND_net), .I3(GND_net), .O(n7_adj_4667));
    defparam i2_2_lut_adj_1000.LUT_INIT = 16'h6666;
    SB_LUT4 i1_3_lut_adj_1001 (.I0(\data_in_frame[5] [2]), .I1(n49258), 
            .I2(\data_in_frame[7] [4]), .I3(GND_net), .O(n49226));
    defparam i1_3_lut_adj_1001.LUT_INIT = 16'h9696;
    SB_LUT4 i1_4_lut_adj_1002 (.I0(n28263), .I1(n27862), .I2(n49226), 
            .I3(n52864), .O(n27659));
    defparam i1_4_lut_adj_1002.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1003 (.I0(\data_in_frame[0] [4]), .I1(\data_in_frame[0] [6]), 
            .I2(ID[4]), .I3(ID[6]), .O(n12_adj_4668));   // verilog/coms.v(239[12:32])
    defparam i4_4_lut_adj_1003.LUT_INIT = 16'h7bde;
    SB_LUT4 i2_4_lut_adj_1004 (.I0(\data_in_frame[0] [1]), .I1(\data_in_frame[0] [2]), 
            .I2(ID[1]), .I3(ID[2]), .O(n10_adj_4669));   // verilog/coms.v(239[12:32])
    defparam i2_4_lut_adj_1004.LUT_INIT = 16'h7bde;
    SB_LUT4 i3_4_lut_adj_1005 (.I0(\data_in_frame[0] [7]), .I1(\data_in_frame[0] [5]), 
            .I2(ID[7]), .I3(ID[5]), .O(n11_adj_4670));   // verilog/coms.v(239[12:32])
    defparam i3_4_lut_adj_1005.LUT_INIT = 16'h7bde;
    SB_LUT4 i1_4_lut_adj_1006 (.I0(\data_in_frame[0] [0]), .I1(\data_in_frame[0] [3]), 
            .I2(ID[0]), .I3(ID[3]), .O(n9));   // verilog/coms.v(239[12:32])
    defparam i1_4_lut_adj_1006.LUT_INIT = 16'h7bde;
    SB_LUT4 i7_4_lut_adj_1007 (.I0(n9), .I1(n11_adj_4670), .I2(n10_adj_4669), 
            .I3(n12_adj_4668), .O(n24549));   // verilog/coms.v(239[12:32])
    defparam i7_4_lut_adj_1007.LUT_INIT = 16'hfffe;
    SB_LUT4 i4_4_lut_adj_1008 (.I0(n49064), .I1(n49021), .I2(n45758), 
            .I3(n49206), .O(n10_adj_4671));   // verilog/coms.v(79[16:27])
    defparam i4_4_lut_adj_1008.LUT_INIT = 16'h6996;
    SB_LUT4 equal_2277_i4_2_lut (.I0(Kp_23__N_1296), .I1(\data_in_frame[8] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_4672));   // verilog/coms.v(237[9:81])
    defparam equal_2277_i4_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i5_3_lut_adj_1009 (.I0(n49038), .I1(n10_adj_4671), .I2(\data_in_frame[8]_c [1]), 
            .I3(GND_net), .O(n51412));   // verilog/coms.v(79[16:27])
    defparam i5_3_lut_adj_1009.LUT_INIT = 16'h9696;
    SB_LUT4 i12_4_lut (.I0(n7_adj_4673), .I1(n27669), .I2(n49120), .I3(n27659), 
            .O(n28));
    defparam i12_4_lut.LUT_INIT = 16'hbfff;
    SB_LUT4 i10_4_lut_adj_1010 (.I0(n27962), .I1(n3_adj_4674), .I2(n27954), 
            .I3(n27604), .O(n26));
    defparam i10_4_lut_adj_1010.LUT_INIT = 16'hfffe;
    SB_LUT4 i11_4_lut (.I0(n27928), .I1(n51412), .I2(n46188), .I3(n4_adj_4672), 
            .O(n27));
    defparam i11_4_lut.LUT_INIT = 16'hffef;
    SB_LUT4 mux_2112_i17_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n36483), 
            .I2(\data_in_frame[1] [0]), .I3(\data_in_frame[17] [0]), .O(n7689));
    defparam mux_2112_i17_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i9_4_lut_adj_1011 (.I0(n45804), .I1(n49688), .I2(n7_adj_4667), 
            .I3(n28082), .O(n25));
    defparam i9_4_lut_adj_1011.LUT_INIT = 16'hfffb;
    SB_LUT4 i15_4_lut_adj_1012 (.I0(n25), .I1(n27), .I2(n26), .I3(n28), 
            .O(n31_adj_4666));
    defparam i15_4_lut_adj_1012.LUT_INIT = 16'hfffe;
    SB_LUT4 i22419_2_lut (.I0(n31_adj_4666), .I1(n24549), .I2(GND_net), 
            .I3(GND_net), .O(n36483));
    defparam i22419_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_1013 (.I0(\FRAME_MATCHER.state [2]), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(GND_net), .I3(GND_net), .O(n52680));
    defparam i1_2_lut_adj_1013.LUT_INIT = 16'hdddd;
    SB_LUT4 i40091_4_lut (.I0(n48979), .I1(n23548), .I2(n48871), .I3(n52680), 
            .O(n28716));
    defparam i40091_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i39050_2_lut (.I0(n56895), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n54596));
    defparam i39050_2_lut.LUT_INIT = 16'h2222;
    SB_DFFSR tx_transmit_4011 (.Q(r_SM_Main_2__N_3851[0]), .C(clk16MHz), 
            .D(n6223[0]), .R(n49887));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 mux_2112_i18_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n36483), 
            .I2(\data_in_frame[1] [1]), .I3(\data_in_frame[17] [1]), .O(n7690));
    defparam mux_2112_i18_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 mux_2112_i19_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n36483), 
            .I2(\data_in_frame[1] [2]), .I3(\data_in_frame[17] [2]), .O(n7691));
    defparam mux_2112_i19_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i37434_3_lut (.I0(\data_out_frame[8] [1]), .I1(\data_out_frame[9] [1]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n53264));
    defparam i37434_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i37435_3_lut (.I0(\data_out_frame[10] [1]), .I1(\data_out_frame[11] [1]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n53265));
    defparam i37435_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i37342_3_lut (.I0(\data_out_frame[14] [1]), .I1(\data_out_frame[15] [1]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n53172));
    defparam i37342_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_2112_i20_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n36483), 
            .I2(\data_in_frame[1] [3]), .I3(\data_in_frame[17] [3]), .O(n7692));
    defparam mux_2112_i20_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i37341_3_lut (.I0(\data_out_frame[12] [1]), .I1(\data_out_frame[13] [1]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n53171));
    defparam i37341_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_2112_i21_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n36483), 
            .I2(\data_in_frame[1] [4]), .I3(\data_in_frame[17] [4]), .O(n7693));
    defparam mux_2112_i21_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_adj_1014 (.I0(byte_transmit_counter[6]), .I1(byte_transmit_counter[5]), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_4675));
    defparam i1_2_lut_adj_1014.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_1015 (.I0(byte_transmit_counter[4]), .I1(byte_transmit_counter[0]), 
            .I2(byte_transmit_counter[2]), .I3(byte_transmit_counter[1]), 
            .O(n4_adj_4676));
    defparam i1_4_lut_adj_1015.LUT_INIT = 16'ha8a0;
    SB_LUT4 i40666_4_lut (.I0(byte_transmit_counter[3]), .I1(byte_transmit_counter[7]), 
            .I2(n4_adj_4676), .I3(n4_adj_4675), .O(tx_transmit_N_3748));
    defparam i40666_4_lut.LUT_INIT = 16'h0013;
    SB_LUT4 i22406_2_lut (.I0(tx_active), .I1(r_SM_Main_2__N_3851[0]), .I2(GND_net), 
            .I3(GND_net), .O(n36465));
    defparam i22406_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 mux_2112_i22_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n36483), 
            .I2(\data_in_frame[1] [5]), .I3(\data_in_frame[17] [5]), .O(n7694));
    defparam mux_2112_i22_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i34131_3_lut (.I0(\FRAME_MATCHER.state[3] ), .I1(n48871), .I2(n49824), 
            .I3(GND_net), .O(n49887));
    defparam i34131_3_lut.LUT_INIT = 16'hecec;
    SB_LUT4 mux_1461_i1_4_lut (.I0(tx_transmit_N_3748), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(n7828), .I3(n8_adj_4677), .O(n6223[0]));   // verilog/coms.v(146[4] 302[11])
    defparam mux_1461_i1_4_lut.LUT_INIT = 16'h0cac;
    SB_LUT4 mux_2112_i23_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n36483), 
            .I2(\data_in_frame[1] [6]), .I3(\data_in_frame[17] [6]), .O(n7695));
    defparam mux_2112_i23_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 mux_2112_i24_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n36483), 
            .I2(\data_in_frame[1] [7]), .I3(\data_in_frame[17] [7]), .O(n7696));
    defparam mux_2112_i24_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_4_lut_adj_1016 (.I0(n49111), .I1(n49246), .I2(Kp_23__N_1602), 
            .I3(\data_in_frame[13] [2]), .O(n28406));
    defparam i1_4_lut_adj_1016.LUT_INIT = 16'h6996;
    SB_LUT4 mux_2112_i1_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n36483), 
            .I2(\data_in_frame[3] [0]), .I3(\data_in_frame[19] [0]), .O(n7673));
    defparam mux_2112_i1_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i15551_3_lut_4_lut (.I0(n37171), .I1(n48993), .I2(rx_data[7]), 
            .I3(\data_in_frame[15] [7]), .O(n29631));
    defparam i15551_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i15552_3_lut_4_lut (.I0(n37171), .I1(n48993), .I2(rx_data[6]), 
            .I3(\data_in_frame[15] [6]), .O(n29632));
    defparam i15552_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i40635_3_lut (.I0(n49824), .I1(n49911), .I2(n27235), .I3(GND_net), 
            .O(n50359));
    defparam i40635_3_lut.LUT_INIT = 16'h0101;
    SB_LUT4 i1_4_lut_adj_1017 (.I0(\FRAME_MATCHER.state[0] ), .I1(n24549), 
            .I2(\FRAME_MATCHER.state [2]), .I3(n23548), .O(n51106));
    defparam i1_4_lut_adj_1017.LUT_INIT = 16'h5040;
    SB_LUT4 i15553_3_lut_4_lut (.I0(n37171), .I1(n48993), .I2(rx_data[5]), 
            .I3(\data_in_frame[15] [5]), .O(n29633));
    defparam i15553_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 equal_333_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8_adj_4678));
    defparam equal_333_i8_2_lut_3_lut.LUT_INIT = 16'hf7f7;
    SB_LUT4 i1_4_lut_adj_1018 (.I0(n46800), .I1(n49288), .I2(n49432), 
            .I3(n52608), .O(n52614));
    defparam i1_4_lut_adj_1018.LUT_INIT = 16'h9669;
    SB_LUT4 i1_3_lut_adj_1019 (.I0(n45766), .I1(n51108), .I2(Kp_23__N_1895), 
            .I3(GND_net), .O(n51124));
    defparam i1_3_lut_adj_1019.LUT_INIT = 16'h6969;
    SB_LUT4 i40098_4_lut (.I0(n27235), .I1(n7828), .I2(n52474), .I3(n51106), 
            .O(n48905));
    defparam i40098_4_lut.LUT_INIT = 16'h1115;
    SB_LUT4 i1_4_lut_adj_1020 (.I0(n50995), .I1(\data_in_frame[23] [1]), 
            .I2(n52418), .I3(n49122), .O(n52422));
    defparam i1_4_lut_adj_1020.LUT_INIT = 16'hfdf7;
    SB_DFF \FRAME_MATCHER.rx_data_ready_prev_4012  (.Q(\FRAME_MATCHER.rx_data_ready_prev ), 
           .C(clk16MHz), .D(rx_data_ready));   // verilog/coms.v(128[12] 303[6])
    SB_DFF Kp_i8 (.Q(\Kp[8] ), .C(clk16MHz), .D(n29513));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i1_4_lut_adj_1021 (.I0(n52422), .I1(n52614), .I2(n49122), 
            .I3(n49699), .O(n31));
    defparam i1_4_lut_adj_1021.LUT_INIT = 16'hbeeb;
    SB_DFF Kp_i9 (.Q(\Kp[9] ), .C(clk16MHz), .D(n29512));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i15554_3_lut_4_lut (.I0(n37171), .I1(n48993), .I2(rx_data[4]), 
            .I3(\data_in_frame[15] [4]), .O(n29634));
    defparam i15554_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_41022 (.I0(byte_transmit_counter[3]), 
            .I1(n56715), .I2(n54596), .I3(byte_transmit_counter[4]), .O(n56898));
    defparam byte_transmit_counter_3__bdd_4_lut_41022.LUT_INIT = 16'he4aa;
    SB_DFFE setpoint__i0 (.Q(setpoint[0]), .C(clk16MHz), .E(n28716), .D(n7673));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i1_4_lut_adj_1022 (.I0(\data_in_frame[5] [0]), .I1(\data_in_frame[6] [7]), 
            .I2(\data_in_frame[4] [7]), .I3(\data_in_frame[7] [1]), .O(n52916));   // verilog/coms.v(71[16:27])
    defparam i1_4_lut_adj_1022.LUT_INIT = 16'h6996;
    SB_DFFSS \FRAME_MATCHER.i_i20  (.Q(\FRAME_MATCHER.i [20]), .C(clk16MHz), 
            .D(n2_adj_4679), .S(n3_adj_4665));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i1_3_lut_adj_1023 (.I0(n49229), .I1(n28268), .I2(n52916), 
            .I3(GND_net), .O(n27962));   // verilog/coms.v(71[16:27])
    defparam i1_3_lut_adj_1023.LUT_INIT = 16'h9696;
    SB_LUT4 i1_4_lut_adj_1024 (.I0(n49229), .I1(n27863), .I2(n49094), 
            .I3(\data_in_frame[7] [3]), .O(n46188));   // verilog/coms.v(86[17:70])
    defparam i1_4_lut_adj_1024.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1025 (.I0(n51108), .I1(n49288), .I2(n49646), 
            .I3(n52690), .O(n52696));
    defparam i1_4_lut_adj_1025.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1026 (.I0(n46188), .I1(n27962), .I2(GND_net), 
            .I3(GND_net), .O(n46727));
    defparam i1_2_lut_adj_1026.LUT_INIT = 16'h6666;
    SB_LUT4 i15555_3_lut_4_lut (.I0(n37171), .I1(n48993), .I2(rx_data[3]), 
            .I3(\data_in_frame[15] [3]), .O(n29635));
    defparam i15555_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFFSS \FRAME_MATCHER.i_i1  (.Q(\FRAME_MATCHER.i [1]), .C(clk16MHz), 
            .D(n2_adj_4680), .S(n3_adj_4660));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i15556_3_lut_4_lut (.I0(n37171), .I1(n48993), .I2(rx_data[2]), 
            .I3(\data_in_frame[15] [2]), .O(n29636));
    defparam i15556_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_adj_1027 (.I0(\data_in_frame[4] [0]), .I1(\data_in_frame[1] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n49637));   // verilog/coms.v(79[16:27])
    defparam i1_2_lut_adj_1027.LUT_INIT = 16'h6666;
    SB_LUT4 i15557_3_lut_4_lut (.I0(n37171), .I1(n48993), .I2(rx_data[1]), 
            .I3(\data_in_frame[15] [1]), .O(n29637));
    defparam i15557_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i23088_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n37171));
    defparam i23088_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 select_751_Select_1_i1_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), 
            .I1(n19836), .I2(n19602), .I3(n27218), .O(n1));
    defparam select_751_Select_1_i1_3_lut_4_lut.LUT_INIT = 16'h008f;
    SB_DFFSS \FRAME_MATCHER.i_i2  (.Q(\FRAME_MATCHER.i [2]), .C(clk16MHz), 
            .D(n2_adj_4681), .S(n3_adj_4658));   // verilog/coms.v(128[12] 303[6])
    SB_DFFSS \FRAME_MATCHER.i_i3  (.Q(\FRAME_MATCHER.i [3]), .C(clk16MHz), 
            .D(n2_adj_4682), .S(n3_adj_4657));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i1_2_lut_adj_1028 (.I0(\data_in_frame[3] [6]), .I1(\data_in_frame[6] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n28527));   // verilog/coms.v(76[16:27])
    defparam i1_2_lut_adj_1028.LUT_INIT = 16'h6666;
    SB_LUT4 i15558_3_lut_4_lut (.I0(n37171), .I1(n48993), .I2(rx_data[0]), 
            .I3(\data_in_frame[15] [0]), .O(n29638));
    defparam i15558_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_adj_1029 (.I0(\data_in_frame[8]_c [1]), .I1(n25500), 
            .I2(GND_net), .I3(GND_net), .O(n49060));
    defparam i1_2_lut_adj_1029.LUT_INIT = 16'h6666;
    SB_DFFSS \FRAME_MATCHER.i_i19  (.Q(\FRAME_MATCHER.i [19]), .C(clk16MHz), 
            .D(n2_adj_4683), .S(n3_adj_4656));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i1_3_lut_adj_1030 (.I0(\data_in_frame[6] [1]), .I1(\data_in_frame[3] [7]), 
            .I2(\data_in_frame[8][2] ), .I3(GND_net), .O(n52934));
    defparam i1_3_lut_adj_1030.LUT_INIT = 16'h9696;
    SB_LUT4 i1_4_lut_adj_1031 (.I0(n28527), .I1(n49495), .I2(n49637), 
            .I3(n52934), .O(n3_adj_4674));
    defparam i1_4_lut_adj_1031.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1032 (.I0(\FRAME_MATCHER.state[3] ), .I1(n27307), 
            .I2(GND_net), .I3(GND_net), .O(n27223));
    defparam i1_2_lut_adj_1032.LUT_INIT = 16'heeee;
    SB_DFFSS \FRAME_MATCHER.i_i4  (.Q(\FRAME_MATCHER.i [4]), .C(clk16MHz), 
            .D(n2_adj_4684), .S(n3_adj_4654));   // verilog/coms.v(128[12] 303[6])
    SB_DFFSS \FRAME_MATCHER.i_i18  (.Q(\FRAME_MATCHER.i [18]), .C(clk16MHz), 
            .D(n2_adj_4685), .S(n3_adj_4653));   // verilog/coms.v(128[12] 303[6])
    SB_DFFSS \FRAME_MATCHER.i_i17  (.Q(\FRAME_MATCHER.i [17]), .C(clk16MHz), 
            .D(n2_adj_4686), .S(n3_adj_4652));   // verilog/coms.v(128[12] 303[6])
    SB_DFFSS \FRAME_MATCHER.i_i5  (.Q(\FRAME_MATCHER.i [5]), .C(clk16MHz), 
            .D(n2_adj_4687), .S(n3_adj_4651));   // verilog/coms.v(128[12] 303[6])
    SB_DFF Kp_i10 (.Q(\Kp[10] ), .C(clk16MHz), .D(n29511));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i1_3_lut_adj_1033 (.I0(n49492), .I1(n45804), .I2(\data_in_frame[9] [7]), 
            .I3(GND_net), .O(n51163));
    defparam i1_3_lut_adj_1033.LUT_INIT = 16'h9696;
    SB_DFF Kp_i11 (.Q(\Kp[11] ), .C(clk16MHz), .D(n29510));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i1_4_lut_adj_1034 (.I0(n27223), .I1(n31), .I2(n48979), .I3(n4_adj_4688), 
            .O(n50654));
    defparam i1_4_lut_adj_1034.LUT_INIT = 16'hfffe;
    SB_DFF Kp_i12 (.Q(\Kp[12] ), .C(clk16MHz), .D(n29509));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i1_2_lut_3_lut (.I0(n27461), .I1(\data_in_frame[7] [6]), .I2(\data_in_frame[10][2] ), 
            .I3(GND_net), .O(n52728));
    defparam i1_2_lut_3_lut.LUT_INIT = 16'h9696;
    SB_DFF Kp_i13 (.Q(\Kp[13] ), .C(clk16MHz), .D(n29508));   // verilog/coms.v(128[12] 303[6])
    SB_DFF Kp_i14 (.Q(\Kp[14] ), .C(clk16MHz), .D(n29507));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i1_2_lut_adj_1035 (.I0(n28132), .I1(n28406), .I2(GND_net), 
            .I3(GND_net), .O(n49376));
    defparam i1_2_lut_adj_1035.LUT_INIT = 16'h6666;
    SB_LUT4 i24_2_lut (.I0(PWMLimit[17]), .I1(n363), .I2(GND_net), .I3(GND_net), 
            .O(n32464));
    defparam i24_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_3_lut_adj_1036 (.I0(n27461), .I1(\data_in_frame[7] [6]), 
            .I2(n27706), .I3(GND_net), .O(n27669));
    defparam i1_2_lut_3_lut_adj_1036.LUT_INIT = 16'h9696;
    SB_DFFSS \FRAME_MATCHER.i_i16  (.Q(\FRAME_MATCHER.i [16]), .C(clk16MHz), 
            .D(n2_adj_4689), .S(n3_adj_4640));   // verilog/coms.v(128[12] 303[6])
    SB_DFFSS \FRAME_MATCHER.i_i15  (.Q(\FRAME_MATCHER.i [15]), .C(clk16MHz), 
            .D(n2_adj_4690), .S(n3_adj_4639));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i1_4_lut_adj_1037 (.I0(\data_in_frame[12] [3]), .I1(\data_in_frame[10][1] ), 
            .I2(\data_in_frame[12] [4]), .I3(n51163), .O(n49543));
    defparam i1_4_lut_adj_1037.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1038 (.I0(\data_in_frame[3] [5]), .I1(\data_in_frame[1] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n49218));   // verilog/coms.v(79[16:27])
    defparam i1_2_lut_adj_1038.LUT_INIT = 16'h6666;
    SB_DFFSS \FRAME_MATCHER.i_i6  (.Q(\FRAME_MATCHER.i [6]), .C(clk16MHz), 
            .D(n2_adj_4691), .S(n3_adj_4638));   // verilog/coms.v(128[12] 303[6])
    SB_DFFSS \FRAME_MATCHER.i_i7  (.Q(\FRAME_MATCHER.i [7]), .C(clk16MHz), 
            .D(n2_adj_4692), .S(n3_adj_4637));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i38939_2_lut (.I0(n56955), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n54602));
    defparam i38939_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1_2_lut_adj_1039 (.I0(n28138), .I1(n49543), .I2(GND_net), 
            .I3(GND_net), .O(n49373));
    defparam i1_2_lut_adj_1039.LUT_INIT = 16'h6666;
    SB_DFFSS \FRAME_MATCHER.i_i8  (.Q(\FRAME_MATCHER.i [8]), .C(clk16MHz), 
            .D(n2_adj_4693), .S(n3_adj_4635));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i5_4_lut (.I0(\data_in_frame[10][1] ), .I1(n49667), .I2(\data_in_frame[12] [1]), 
            .I3(n49492), .O(n12_adj_4694));
    defparam i5_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1040 (.I0(\data_in_frame[3] [6]), .I1(\data_in_frame[6] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n49203));   // verilog/coms.v(79[16:27])
    defparam i1_2_lut_adj_1040.LUT_INIT = 16'h6666;
    SB_DFF Kp_i15 (.Q(\Kp[15] ), .C(clk16MHz), .D(n29506));   // verilog/coms.v(128[12] 303[6])
    SB_DFFSS \FRAME_MATCHER.i_i9  (.Q(\FRAME_MATCHER.i [9]), .C(clk16MHz), 
            .D(n2_adj_4695), .S(n3_adj_4634));   // verilog/coms.v(128[12] 303[6])
    SB_DFFSS \FRAME_MATCHER.i_i10  (.Q(\FRAME_MATCHER.i [10]), .C(clk16MHz), 
            .D(n2_adj_4696), .S(n3_adj_4631));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i15543_3_lut_4_lut (.I0(n8_adj_4697), .I1(n48984), .I2(rx_data[7]), 
            .I3(\data_in_frame[16] [7]), .O(n29623));
    defparam i15543_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15544_3_lut_4_lut (.I0(n8_adj_4697), .I1(n48984), .I2(rx_data[6]), 
            .I3(\data_in_frame[16] [6]), .O(n29624));
    defparam i15544_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFFSS \FRAME_MATCHER.i_i12  (.Q(\FRAME_MATCHER.i [12]), .C(clk16MHz), 
            .D(n2_adj_4698), .S(n3_adj_4630));   // verilog/coms.v(128[12] 303[6])
    SB_DFF Ki_i1 (.Q(\Ki[1] ), .C(clk16MHz), .D(n29505));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i1_4_lut_adj_1041 (.I0(n49203), .I1(n49218), .I2(\data_in_frame[5] [7]), 
            .I3(\data_in_frame[6] [1]), .O(n49021));   // verilog/coms.v(79[16:27])
    defparam i1_4_lut_adj_1041.LUT_INIT = 16'h6996;
    SB_DFFSS \FRAME_MATCHER.i_i14  (.Q(\FRAME_MATCHER.i [14]), .C(clk16MHz), 
            .D(n2_adj_4699), .S(n3_adj_4629));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i37353_3_lut (.I0(\data_out_frame[8] [0]), .I1(\data_out_frame[9] [0]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n53183));
    defparam i37353_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15545_3_lut_4_lut (.I0(n8_adj_4697), .I1(n48984), .I2(rx_data[5]), 
            .I3(\data_in_frame[16] [5]), .O(n29625));
    defparam i15545_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF Ki_i2 (.Q(\Ki[2] ), .C(clk16MHz), .D(n29504));   // verilog/coms.v(128[12] 303[6])
    SB_DFF Ki_i3 (.Q(\Ki[3] ), .C(clk16MHz), .D(n29503));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i1_2_lut_adj_1042 (.I0(\data_in_frame[2] [0]), .I1(\data_in_frame[1] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n49466));   // verilog/coms.v(79[16:27])
    defparam i1_2_lut_adj_1042.LUT_INIT = 16'h6666;
    SB_LUT4 i37354_3_lut (.I0(\data_out_frame[10] [0]), .I1(\data_out_frame[11] [0]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n53184));
    defparam i37354_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF Ki_i4 (.Q(\Ki[4] ), .C(clk16MHz), .D(n29502));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 n56898_bdd_4_lut (.I0(n56898), .I1(n56799), .I2(n7_adj_4700), 
            .I3(byte_transmit_counter[4]), .O(tx_data[0]));
    defparam n56898_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i37462_3_lut (.I0(\data_out_frame[14] [0]), .I1(\data_out_frame[15] [0]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n53292));
    defparam i37462_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i37461_3_lut (.I0(\data_out_frame[12] [0]), .I1(\data_out_frame[13] [0]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n53291));
    defparam i37461_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i37377_3_lut (.I0(\data_out_frame[8] [3]), .I1(\data_out_frame[9] [3]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n53207));
    defparam i37377_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF Ki_i5 (.Q(\Ki[5] ), .C(clk16MHz), .D(n29499));   // verilog/coms.v(128[12] 303[6])
    SB_DFF Ki_i6 (.Q(\Ki[6] ), .C(clk16MHz), .D(n29498));   // verilog/coms.v(128[12] 303[6])
    SB_DFF Ki_i7 (.Q(\Ki[7] ), .C(clk16MHz), .D(n29497));   // verilog/coms.v(128[12] 303[6])
    SB_DFF Ki_i8 (.Q(\Ki[8] ), .C(clk16MHz), .D(n29496));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i37378_3_lut (.I0(\data_out_frame[10] [3]), .I1(\data_out_frame[11] [3]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n53208));
    defparam i37378_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1043 (.I0(n49466), .I1(n49021), .I2(\data_in_frame[3] [7]), 
            .I3(\data_in_frame[4] [1]), .O(Kp_23__N_1296));   // verilog/coms.v(79[16:27])
    defparam i1_4_lut_adj_1043.LUT_INIT = 16'h6996;
    SB_DFF Ki_i9 (.Q(\Ki[9] ), .C(clk16MHz), .D(n29495));   // verilog/coms.v(128[12] 303[6])
    SB_DFF Ki_i10 (.Q(\Ki[10] ), .C(clk16MHz), .D(n29494));   // verilog/coms.v(128[12] 303[6])
    SB_DFF Ki_i11 (.Q(\Ki[11] ), .C(clk16MHz), .D(n29493));   // verilog/coms.v(128[12] 303[6])
    SB_DFF Ki_i12 (.Q(\Ki[12] ), .C(clk16MHz), .D(n29492));   // verilog/coms.v(128[12] 303[6])
    SB_DFF Ki_i13 (.Q(\Ki[13] ), .C(clk16MHz), .D(n29491));   // verilog/coms.v(128[12] 303[6])
    SB_DFF Ki_i14 (.Q(\Ki[14] ), .C(clk16MHz), .D(n29490));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i188 (.Q(\data_in_frame[23] [3]), .C(clk16MHz), 
           .D(n29487));   // verilog/coms.v(128[12] 303[6])
    SB_DFF Ki_i15 (.Q(\Ki[15] ), .C(clk16MHz), .D(n29486));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_0___i2 (.Q(\data_in[0] [1]), .C(clk16MHz), .D(n29485));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_0___i3 (.Q(\data_in[0] [2]), .C(clk16MHz), .D(n29484));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_0___i4 (.Q(\data_in[0] [3]), .C(clk16MHz), .D(n29483));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_0___i5 (.Q(\data_in[0] [4]), .C(clk16MHz), .D(n29482));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_0___i6 (.Q(\data_in[0] [5]), .C(clk16MHz), .D(n29481));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_0___i7 (.Q(\data_in[0] [6]), .C(clk16MHz), .D(n29480));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_0___i8 (.Q(\data_in[0] [7]), .C(clk16MHz), .D(n29479));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i15546_3_lut_4_lut (.I0(n8_adj_4697), .I1(n48984), .I2(rx_data[4]), 
            .I3(\data_in_frame[16] [4]), .O(n29626));
    defparam i15546_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_0___i9 (.Q(\data_in[1] [0]), .C(clk16MHz), .D(n29478));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_0___i10 (.Q(\data_in[1] [1]), .C(clk16MHz), .D(n29477));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_0___i11 (.Q(\data_in[1] [2]), .C(clk16MHz), .D(n29476));   // verilog/coms.v(128[12] 303[6])
    SB_DFFSS \FRAME_MATCHER.i_i13  (.Q(\FRAME_MATCHER.i [13]), .C(clk16MHz), 
            .D(n2_adj_4701), .S(n3_adj_4623));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i37384_3_lut (.I0(\data_out_frame[14] [3]), .I1(\data_out_frame[15] [3]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n53214));
    defparam i37384_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i37383_3_lut (.I0(\data_out_frame[12] [3]), .I1(\data_out_frame[13] [3]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n53213));
    defparam i37383_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15547_3_lut_4_lut (.I0(n8_adj_4697), .I1(n48984), .I2(rx_data[3]), 
            .I3(\data_in_frame[16] [3]), .O(n29627));
    defparam i15547_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15548_3_lut_4_lut (.I0(n8_adj_4697), .I1(n48984), .I2(rx_data[2]), 
            .I3(\data_in_frame[16] [2]), .O(n29628));
    defparam i15548_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15549_3_lut_4_lut (.I0(n8_adj_4697), .I1(n48984), .I2(rx_data[1]), 
            .I3(\data_in_frame[16] [1]), .O(n29629));
    defparam i15549_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i6_4_lut_adj_1044 (.I0(\data_in_frame[12] [2]), .I1(n12_adj_4694), 
            .I2(\data_in_frame[14] [3]), .I3(n49652), .O(n49328));
    defparam i6_4_lut_adj_1044.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1045 (.I0(\data_in_frame[16] [5]), .I1(\data_in_frame[16] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n52836));
    defparam i1_2_lut_adj_1045.LUT_INIT = 16'h6666;
    SB_LUT4 i15550_3_lut_4_lut (.I0(n8_adj_4697), .I1(n48984), .I2(rx_data[0]), 
            .I3(\data_in_frame[16] [0]), .O(n29630));
    defparam i15550_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFFESR byte_transmit_counter_i0_i1 (.Q(byte_transmit_counter[1]), .C(clk16MHz), 
            .E(n28738), .D(n9046[1]), .R(n29306));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_0___i12 (.Q(\data_in[1] [3]), .C(clk16MHz), .D(n29472));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i1_2_lut_adj_1046 (.I0(\data_in_frame[13] [1]), .I1(n26844), 
            .I2(GND_net), .I3(GND_net), .O(n49246));
    defparam i1_2_lut_adj_1046.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1047 (.I0(\data_in_frame[13] [2]), .I1(\data_in_frame[13] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n27400));
    defparam i1_2_lut_adj_1047.LUT_INIT = 16'h6666;
    SB_DFFESR byte_transmit_counter_i0_i2 (.Q(byte_transmit_counter[2]), .C(clk16MHz), 
            .E(n28738), .D(n9046[2]), .R(n29306));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i5652_2_lut_3_lut (.I0(n45364), .I1(\FRAME_MATCHER.i [31]), 
            .I2(n63_adj_6), .I3(GND_net), .O(n19602));   // verilog/coms.v(158[9:60])
    defparam i5652_2_lut_3_lut.LUT_INIT = 16'hd0d0;
    SB_LUT4 i1_4_lut_adj_1048 (.I0(n46749), .I1(n46832), .I2(n49328), 
            .I3(n52836), .O(n49249));
    defparam i1_4_lut_adj_1048.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1049 (.I0(n45364), .I1(\FRAME_MATCHER.i [31]), 
            .I2(n22875), .I3(GND_net), .O(n24251));   // verilog/coms.v(158[9:60])
    defparam i1_2_lut_3_lut_adj_1049.LUT_INIT = 16'hd0d0;
    SB_LUT4 i1_3_lut_4_lut (.I0(n45364), .I1(\FRAME_MATCHER.i [31]), .I2(n4599), 
            .I3(n27218), .O(n4));   // verilog/coms.v(158[9:60])
    defparam i1_3_lut_4_lut.LUT_INIT = 16'hf0fd;
    SB_LUT4 i1_2_lut_adj_1050 (.I0(\data_in_frame[0] [5]), .I1(\data_in_frame[0] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n49085));   // verilog/coms.v(77[16:27])
    defparam i1_2_lut_adj_1050.LUT_INIT = 16'h6666;
    SB_DFF data_in_0___i13 (.Q(\data_in[1] [4]), .C(clk16MHz), .D(n29471));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i1_2_lut_adj_1051 (.I0(\data_in_frame[0] [6]), .I1(\data_in_frame[0] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n49117));   // verilog/coms.v(71[16:27])
    defparam i1_2_lut_adj_1051.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1052 (.I0(n49117), .I1(n49032), .I2(n49085), 
            .I3(\data_in_frame[0] [1]), .O(Kp_23__N_1079));   // verilog/coms.v(71[16:27])
    defparam i1_4_lut_adj_1052.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1053 (.I0(\data_in_frame[2] [0]), .I1(n28037), 
            .I2(GND_net), .I3(GND_net), .O(n49165));   // verilog/coms.v(74[16:42])
    defparam i1_2_lut_adj_1053.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1054 (.I0(\data_in_frame[6] [7]), .I1(\data_in_frame[6] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n28066));   // verilog/coms.v(86[17:28])
    defparam i1_2_lut_adj_1054.LUT_INIT = 16'h6666;
    SB_LUT4 i1_3_lut_adj_1055 (.I0(\data_in_frame[5] [5]), .I1(n49258), 
            .I2(\data_in_frame[5] [4]), .I3(GND_net), .O(n27461));
    defparam i1_3_lut_adj_1055.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1056 (.I0(\data_in_frame[3] [7]), .I1(\data_in_frame[4] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n49074));   // verilog/coms.v(71[16:69])
    defparam i1_2_lut_adj_1056.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1057 (.I0(\data_in_frame[18] [7]), .I1(n49249), 
            .I2(\data_in_frame[19] [1]), .I3(GND_net), .O(n50429));
    defparam i2_3_lut_adj_1057.LUT_INIT = 16'h9696;
    SB_LUT4 i1_4_lut_adj_1058 (.I0(\data_in_frame[5] [3]), .I1(\data_in_frame[5] [7]), 
            .I2(\data_in_frame[4] [0]), .I3(\data_in_frame[3] [6]), .O(n52566));
    defparam i1_4_lut_adj_1058.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1059 (.I0(n49074), .I1(n49664), .I2(n49517), 
            .I3(n52566), .O(n52574));
    defparam i1_4_lut_adj_1059.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1060 (.I0(\data_in_frame[2] [1]), .I1(\data_in_frame[4] [1]), 
            .I2(\data_in_frame[1] [1]), .I3(\data_in_frame[3] [3]), .O(n52588));
    defparam i1_4_lut_adj_1060.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1061 (.I0(n27461), .I1(n52574), .I2(n49522), 
            .I3(n52572), .O(n52580));
    defparam i1_4_lut_adj_1061.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1062 (.I0(\data_in_frame[13] [7]), .I1(\data_in_frame[16] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n49042));
    defparam i1_2_lut_adj_1062.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1063 (.I0(n52592), .I1(n52580), .I2(n49540), 
            .I3(GND_net), .O(n45758));
    defparam i1_4_lut_adj_1063.LUT_INIT = 16'h9696;
    SB_LUT4 i1_4_lut_adj_1064 (.I0(\data_in_frame[6] [1]), .I1(\data_in_frame[6] [0]), 
            .I2(\data_in_frame[6] [5]), .I3(\data_in_frame[6] [2]), .O(n52552));   // verilog/coms.v(86[17:28])
    defparam i1_4_lut_adj_1064.LUT_INIT = 16'h6996;
    SB_LUT4 i1_3_lut_adj_1065 (.I0(n49206), .I1(n45758), .I2(n52552), 
            .I3(GND_net), .O(n49705));   // verilog/coms.v(86[17:28])
    defparam i1_3_lut_adj_1065.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1066 (.I0(n28268), .I1(n49705), .I2(GND_net), 
            .I3(GND_net), .O(n49221));
    defparam i1_2_lut_adj_1066.LUT_INIT = 16'h6666;
    SB_LUT4 i1_3_lut_adj_1067 (.I0(\data_in_frame[0] [1]), .I1(\data_in_frame[0] [0]), 
            .I2(\data_in_frame[2] [2]), .I3(GND_net), .O(n28037));   // verilog/coms.v(74[16:42])
    defparam i1_3_lut_adj_1067.LUT_INIT = 16'h9696;
    SB_LUT4 i1_4_lut_adj_1068 (.I0(n28303), .I1(n27954), .I2(\data_in_frame[8][6] ), 
            .I3(\data_in_frame[8] [7]), .O(n49702));   // verilog/coms.v(72[16:27])
    defparam i1_4_lut_adj_1068.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1069 (.I0(\data_in_frame[11] [7]), .I1(n46188), 
            .I2(GND_net), .I3(GND_net), .O(n49667));
    defparam i1_2_lut_adj_1069.LUT_INIT = 16'h6666;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_41062 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [0]), .I2(\data_out_frame[27] [0]), 
            .I3(byte_transmit_counter[1]), .O(n56892));
    defparam byte_transmit_counter_0__bdd_4_lut_41062.LUT_INIT = 16'he4aa;
    SB_LUT4 n56928_bdd_4_lut (.I0(n56928), .I1(n56835), .I2(n7_adj_4703), 
            .I3(byte_transmit_counter[4]), .O(tx_data[5]));
    defparam n56928_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n56922_bdd_4_lut (.I0(n56922), .I1(n56829), .I2(n7_adj_4704), 
            .I3(byte_transmit_counter[4]), .O(tx_data[4]));
    defparam n56922_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_adj_1070 (.I0(\data_in_frame[15] [5]), .I1(\data_in_frame[17] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n49475));
    defparam i1_2_lut_adj_1070.LUT_INIT = 16'h6666;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut (.I0(byte_transmit_counter[3]), 
            .I1(n56637), .I2(n54592), .I3(byte_transmit_counter[4]), .O(n56940));
    defparam byte_transmit_counter_3__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 i6_4_lut_adj_1071 (.I0(n49376), .I1(\data_in_frame[9] [3]), 
            .I2(\data_in_frame[11] [5]), .I3(n46727), .O(n15_adj_4705));
    defparam i6_4_lut_adj_1071.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1072 (.I0(\data_in_frame[7] [7]), .I1(n55901), 
            .I2(\data_in_frame[8][2] ), .I3(\data_in_frame[9] [6]), .O(n49525));
    defparam i3_4_lut_adj_1072.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1073 (.I0(\data_in_frame[4] [5]), .I1(\data_in_frame[6] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n49064));   // verilog/coms.v(76[16:43])
    defparam i1_2_lut_adj_1073.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1074 (.I0(\data_in_frame[6] [6]), .I1(n49064), 
            .I2(n28017), .I3(Kp_23__N_1209), .O(Kp_23__N_1324));   // verilog/coms.v(76[16:43])
    defparam i3_4_lut_adj_1074.LUT_INIT = 16'h6996;
    SB_DFF data_in_0___i14 (.Q(\data_in[1] [5]), .C(clk16MHz), .D(n29470));   // verilog/coms.v(128[12] 303[6])
    SB_DFFSS \FRAME_MATCHER.i_i31  (.Q(\FRAME_MATCHER.i [31]), .C(clk16MHz), 
            .D(n2_adj_4706), .S(n3_adj_4707));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i15535_3_lut_4_lut (.I0(n8_adj_4708), .I1(n48984), .I2(rx_data[7]), 
            .I3(\data_in_frame[17] [7]), .O(n29615));
    defparam i15535_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_0___i15 (.Q(\data_in[1] [6]), .C(clk16MHz), .D(n29469));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 n56916_bdd_4_lut (.I0(n56916), .I1(n56823), .I2(n7_adj_4709), 
            .I3(byte_transmit_counter[4]), .O(tx_data[3]));
    defparam n56916_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFFESR byte_transmit_counter_i0_i3 (.Q(byte_transmit_counter[3]), .C(clk16MHz), 
            .E(n28738), .D(n9046[3]), .R(n29306));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i1_4_lut_adj_1075 (.I0(DE_c), .I1(n7828), .I2(n27235), .I3(n27248), 
            .O(n48390));   // verilog/TinyFPGA_B.v(15[10:12])
    defparam i1_4_lut_adj_1075.LUT_INIT = 16'ha8ac;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_41037 (.I0(byte_transmit_counter[3]), 
            .I1(n56685), .I2(n54598), .I3(byte_transmit_counter[4]), .O(n56916));
    defparam byte_transmit_counter_3__bdd_4_lut_41037.LUT_INIT = 16'he4aa;
    SB_LUT4 i15536_3_lut_4_lut (.I0(n8_adj_4708), .I1(n48984), .I2(rx_data[6]), 
            .I3(\data_in_frame[17] [6]), .O(n29616));
    defparam i15536_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFFESR byte_transmit_counter_i0_i4 (.Q(byte_transmit_counter[4]), .C(clk16MHz), 
            .E(n28738), .D(n9046[4]), .R(n29306));   // verilog/coms.v(128[12] 303[6])
    SB_DFFESR byte_transmit_counter_i0_i5 (.Q(byte_transmit_counter[5]), .C(clk16MHz), 
            .E(n28738), .D(n9046[5]), .R(n29306));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i1_3_lut_adj_1076 (.I0(\data_in_frame[1] [2]), .I1(\data_in_frame[1] [3]), 
            .I2(\data_in_frame[3] [4]), .I3(GND_net), .O(n27706));
    defparam i1_3_lut_adj_1076.LUT_INIT = 16'h9696;
    SB_LUT4 i1_3_lut_adj_1077 (.I0(n27706), .I1(n28030), .I2(\data_in_frame[5] [5]), 
            .I3(GND_net), .O(n28050));
    defparam i1_3_lut_adj_1077.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1078 (.I0(\data_in_frame[9] [2]), .I1(Kp_23__N_1324), 
            .I2(\data_in_frame[9] [1]), .I3(GND_net), .O(n49162));   // verilog/coms.v(73[16:41])
    defparam i2_3_lut_adj_1078.LUT_INIT = 16'h9696;
    SB_LUT4 i1_4_lut_adj_1079 (.I0(\data_in_frame[8] [0]), .I1(\data_in_frame[11] [5]), 
            .I2(\data_in_frame[8]_c [1]), .I3(\data_in_frame[14] [1]), .O(n52708));
    defparam i1_4_lut_adj_1079.LUT_INIT = 16'h6996;
    SB_LUT4 i1_3_lut_adj_1080 (.I0(n52708), .I1(\data_in_frame[13] [7]), 
            .I2(\data_in_frame[9] [0]), .I3(GND_net), .O(n52710));
    defparam i1_3_lut_adj_1080.LUT_INIT = 16'h9696;
    SB_LUT4 i8_4_lut_adj_1081 (.I0(n15_adj_4705), .I1(n27680), .I2(n14_adj_4710), 
            .I3(n49246), .O(n49569));
    defparam i8_4_lut_adj_1081.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1082 (.I0(n49162), .I1(n27577), .I2(n28050), 
            .I3(n52710), .O(n52716));
    defparam i1_4_lut_adj_1082.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1083 (.I0(n46699), .I1(n49569), .I2(n49475), 
            .I3(n49042), .O(n46413));
    defparam i3_4_lut_adj_1083.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1084 (.I0(n49525), .I1(n49667), .I2(n49702), 
            .I3(n52716), .O(n52722));
    defparam i1_4_lut_adj_1084.LUT_INIT = 16'h6996;
    SB_DFFESR byte_transmit_counter_i0_i6 (.Q(byte_transmit_counter[6]), .C(clk16MHz), 
            .E(n28738), .D(n9046[6]), .R(n29306));   // verilog/coms.v(128[12] 303[6])
    SB_DFFESR byte_transmit_counter_i0_i7 (.Q(byte_transmit_counter[7]), .C(clk16MHz), 
            .E(n28738), .D(n9046[7]), .R(n29306));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i1_4_lut_adj_1085 (.I0(n49221), .I1(n50767), .I2(n52722), 
            .I3(\data_in_frame[12] [0]), .O(n46793));
    defparam i1_4_lut_adj_1085.LUT_INIT = 16'h9669;
    SB_LUT4 i15537_3_lut_4_lut (.I0(n8_adj_4708), .I1(n48984), .I2(rx_data[5]), 
            .I3(\data_in_frame[17] [5]), .O(n29617));
    defparam i15537_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_4_lut_adj_1086 (.I0(\data_in_frame[12] [5]), .I1(\data_in_frame[11] [3]), 
            .I2(\data_in_frame[11] [7]), .I3(\data_in_frame[11] [0]), .O(n52524));
    defparam i1_4_lut_adj_1086.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1087 (.I0(n52524), .I1(n49612), .I2(\data_in_frame[12] [6]), 
            .I3(\data_in_frame[9] [2]), .O(n52528));
    defparam i1_4_lut_adj_1087.LUT_INIT = 16'h6996;
    SB_DFF data_in_0___i16 (.Q(\data_in[1] [7]), .C(clk16MHz), .D(n29468));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i1_2_lut_adj_1088 (.I0(n46793), .I1(n45864), .I2(GND_net), 
            .I3(GND_net), .O(n46708));
    defparam i1_2_lut_adj_1088.LUT_INIT = 16'h9999;
    SB_DFF data_in_0___i17 (.Q(\data_in[2] [0]), .C(clk16MHz), .D(n29467));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_0___i18 (.Q(\data_in[2] [1]), .C(clk16MHz), .D(n29466));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i1_4_lut_adj_1089 (.I0(n27659), .I1(n49234), .I2(n52530), 
            .I3(n52528), .O(n52536));
    defparam i1_4_lut_adj_1089.LUT_INIT = 16'h6996;
    SB_DFF data_in_0___i19 (.Q(\data_in[2] [2]), .C(clk16MHz), .D(n29465));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i37398_3_lut (.I0(\data_out_frame[8] [4]), .I1(\data_out_frame[9] [4]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n53228));
    defparam i37398_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i37399_3_lut (.I0(\data_out_frame[10] [4]), .I1(\data_out_frame[11] [4]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n53229));
    defparam i37399_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1090 (.I0(n49335), .I1(n46727), .I2(n28403), 
            .I3(n52536), .O(n52542));
    defparam i1_4_lut_adj_1090.LUT_INIT = 16'h6996;
    SB_LUT4 i15538_3_lut_4_lut (.I0(n8_adj_4708), .I1(n48984), .I2(rx_data[4]), 
            .I3(\data_in_frame[17] [4]), .O(n29618));
    defparam i15538_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_4_lut_adj_1091 (.I0(n49446), .I1(n49582), .I2(n49373), 
            .I3(n52542), .O(n26844));
    defparam i1_4_lut_adj_1091.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1092 (.I0(\FRAME_MATCHER.state [14]), .I1(\FRAME_MATCHER.state [13]), 
            .I2(GND_net), .I3(GND_net), .O(n48));   // verilog/coms.v(128[12] 303[6])
    defparam i1_2_lut_adj_1092.LUT_INIT = 16'heeee;
    SB_LUT4 n56940_bdd_4_lut (.I0(n56940), .I1(n56847), .I2(n7_adj_4711), 
            .I3(byte_transmit_counter[4]), .O(tx_data[7]));
    defparam n56940_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF data_in_0___i20 (.Q(\data_in[2] [3]), .C(clk16MHz), .D(n29464));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_0___i21 (.Q(\data_in[2] [4]), .C(clk16MHz), .D(n29463));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_0___i22 (.Q(\data_in[2] [5]), .C(clk16MHz), .D(n29462));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_0___i23 (.Q(\data_in[2] [6]), .C(clk16MHz), .D(n29461));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_0___i24 (.Q(\data_in[2] [7]), .C(clk16MHz), .D(n29460));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_0___i25 (.Q(\data_in[3] [0]), .C(clk16MHz), .D(n29456));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_0___i26 (.Q(\data_in[3] [1]), .C(clk16MHz), .D(n29455));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_0___i27 (.Q(\data_in[3] [2]), .C(clk16MHz), .D(n29454));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_0___i28 (.Q(\data_in[3] [3]), .C(clk16MHz), .D(n29453));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_0___i29 (.Q(\data_in[3] [4]), .C(clk16MHz), .D(n29451));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i3_4_lut_adj_1093 (.I0(\FRAME_MATCHER.state [4]), .I1(\FRAME_MATCHER.state [7]), 
            .I2(\FRAME_MATCHER.state [5]), .I3(\FRAME_MATCHER.state [6]), 
            .O(n37153));
    defparam i3_4_lut_adj_1093.LUT_INIT = 16'hfffe;
    SB_LUT4 i5_4_lut_adj_1094 (.I0(\FRAME_MATCHER.state [21]), .I1(\FRAME_MATCHER.state [27]), 
            .I2(\FRAME_MATCHER.state [19]), .I3(\FRAME_MATCHER.state [20]), 
            .O(n12_adj_4712));   // verilog/coms.v(128[12] 303[6])
    defparam i5_4_lut_adj_1094.LUT_INIT = 16'hfffe;
    SB_LUT4 i3_4_lut_adj_1095 (.I0(\data_in_frame[12] [6]), .I1(n49633), 
            .I2(n27400), .I3(n27692), .O(n49696));
    defparam i3_4_lut_adj_1095.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut (.I0(n46749), .I1(n46673), .I2(\data_in_frame[16] [6]), 
            .I3(n49331), .O(n49599));
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h9669;
    SB_LUT4 i4_4_lut_adj_1096 (.I0(n49451), .I1(\data_out_frame[25] [7]), 
            .I2(\data_out_frame[25] [6]), .I3(n49578), .O(n10_adj_4713));
    defparam i4_4_lut_adj_1096.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1097 (.I0(\FRAME_MATCHER.state [24]), .I1(n12_adj_4712), 
            .I2(\FRAME_MATCHER.state [18]), .I3(\FRAME_MATCHER.state [23]), 
            .O(n48866));   // verilog/coms.v(128[12] 303[6])
    defparam i6_4_lut_adj_1097.LUT_INIT = 16'hfffe;
    SB_LUT4 i5_3_lut_adj_1098 (.I0(\data_out_frame[23] [6]), .I1(n10_adj_4713), 
            .I2(n46738), .I3(GND_net), .O(n50764));
    defparam i5_3_lut_adj_1098.LUT_INIT = 16'h6969;
    SB_LUT4 i5_4_lut_adj_1099 (.I0(n46718), .I1(n45830), .I2(n51314), 
            .I3(n25418), .O(n12_adj_4714));
    defparam i5_4_lut_adj_1099.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_1100 (.I0(\FRAME_MATCHER.state [22]), .I1(\FRAME_MATCHER.state [25]), 
            .I2(\FRAME_MATCHER.state [28]), .I3(GND_net), .O(n14_adj_4715));   // verilog/coms.v(202[5:24])
    defparam i5_3_lut_adj_1100.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_4_lut_adj_1101 (.I0(n45802), .I1(n49696), .I2(n49111), 
            .I3(\data_in_frame[17] [3]), .O(n52394));
    defparam i1_4_lut_adj_1101.LUT_INIT = 16'h6996;
    SB_DFF data_in_0___i30 (.Q(\data_in[3] [5]), .C(clk16MHz), .D(n29450));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i6_4_lut_adj_1102 (.I0(n46827), .I1(n12_adj_4714), .I2(n49412), 
            .I3(n46420), .O(n51417));
    defparam i6_4_lut_adj_1102.LUT_INIT = 16'h9669;
    SB_LUT4 i6_4_lut_adj_1103 (.I0(\FRAME_MATCHER.state [30]), .I1(\FRAME_MATCHER.state [31]), 
            .I2(\FRAME_MATCHER.state [16]), .I3(\FRAME_MATCHER.state [26]), 
            .O(n15_adj_4716));   // verilog/coms.v(202[5:24])
    defparam i6_4_lut_adj_1103.LUT_INIT = 16'hfffe;
    SB_LUT4 i8_4_lut_adj_1104 (.I0(n15_adj_4716), .I1(\FRAME_MATCHER.state [29]), 
            .I2(n14_adj_4715), .I3(\FRAME_MATCHER.state [17]), .O(n48864));   // verilog/coms.v(202[5:24])
    defparam i8_4_lut_adj_1104.LUT_INIT = 16'hfffe;
    SB_LUT4 i4_4_lut_adj_1105 (.I0(\FRAME_MATCHER.state [11]), .I1(\FRAME_MATCHER.state [8]), 
            .I2(\FRAME_MATCHER.state [10]), .I3(\FRAME_MATCHER.state [12]), 
            .O(n10_adj_4717));
    defparam i4_4_lut_adj_1105.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_adj_1106 (.I0(\data_in_frame[21] [1]), .I1(\data_in_frame[19] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n52740));
    defparam i1_2_lut_adj_1106.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1107 (.I0(n49696), .I1(n49590), .I2(GND_net), 
            .I3(GND_net), .O(n52670));
    defparam i1_2_lut_adj_1107.LUT_INIT = 16'h6666;
    SB_LUT4 i2_4_lut_adj_1108 (.I0(n48866), .I1(n37153), .I2(n48), .I3(n4_adj_4718), 
            .O(n27307));   // verilog/coms.v(202[5:24])
    defparam i2_4_lut_adj_1108.LUT_INIT = 16'hfffe;
    SB_LUT4 i15539_3_lut_4_lut (.I0(n8_adj_4708), .I1(n48984), .I2(rx_data[3]), 
            .I3(\data_in_frame[17] [3]), .O(n29619));
    defparam i15539_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_4_lut_adj_1109 (.I0(n52740), .I1(n52696), .I2(n51124), 
            .I3(\data_in_frame[20] [7]), .O(n45939));
    defparam i1_4_lut_adj_1109.LUT_INIT = 16'h9669;
    SB_LUT4 i1_4_lut_adj_1110 (.I0(\data_in_frame[15] [3]), .I1(n52670), 
            .I2(\data_in_frame[17] [4]), .I3(n46699), .O(n45874));
    defparam i1_4_lut_adj_1110.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1111 (.I0(n50279), .I1(\data_in_frame[20] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n49432));
    defparam i1_2_lut_adj_1111.LUT_INIT = 16'h9999;
    SB_LUT4 i1_2_lut_adj_1112 (.I0(\data_in_frame[1] [5]), .I1(\data_in_frame[4] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n27557));   // verilog/coms.v(79[16:27])
    defparam i1_2_lut_adj_1112.LUT_INIT = 16'h6666;
    SB_DFF data_in_0___i31 (.Q(\data_in[3] [6]), .C(clk16MHz), .D(n29449));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_0___i32 (.Q(\data_in[3] [7]), .C(clk16MHz), .D(n29448));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i33 (.Q(\data_out_frame[4] [0]), .C(clk16MHz), 
           .D(n29447));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i34 (.Q(\data_out_frame[4] [1]), .C(clk16MHz), 
           .D(n29446));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i35 (.Q(\data_out_frame[4] [2]), .C(clk16MHz), 
           .D(n29445));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i36 (.Q(\data_out_frame[4] [3]), .C(clk16MHz), 
           .D(n29444));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i37 (.Q(\data_out_frame[4] [4]), .C(clk16MHz), 
           .D(n29443));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i38 (.Q(\data_out_frame[4] [5]), .C(clk16MHz), 
           .D(n29442));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i39 (.Q(\data_out_frame[4] [6]), .C(clk16MHz), 
           .D(n29441));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i40 (.Q(\data_out_frame[4] [7]), .C(clk16MHz), 
           .D(n29440));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i41 (.Q(\data_out_frame[5] [0]), .C(clk16MHz), 
           .D(n29439));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i42 (.Q(\data_out_frame[5] [1]), .C(clk16MHz), 
           .D(n29438));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i43 (.Q(\data_out_frame[5] [2]), .C(clk16MHz), 
           .D(n29437));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i44 (.Q(\data_out_frame[5] [3]), .C(clk16MHz), 
           .D(n29436));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i45 (.Q(\data_out_frame[5] [4]), .C(clk16MHz), 
           .D(n29435));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i1_2_lut_adj_1113 (.I0(\data_in_frame[6] [3]), .I1(Kp_23__N_1203), 
            .I2(GND_net), .I3(GND_net), .O(n27577));   // verilog/coms.v(75[16:43])
    defparam i1_2_lut_adj_1113.LUT_INIT = 16'h6666;
    SB_DFF data_out_frame_0___i46 (.Q(\data_out_frame[5] [5]), .C(clk16MHz), 
           .D(n29434));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i47 (.Q(\data_out_frame[5] [6]), .C(clk16MHz), 
           .D(n29433));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i48 (.Q(\data_out_frame[5] [7]), .C(clk16MHz), 
           .D(n29432));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i49 (.Q(\data_out_frame[6] [0]), .C(clk16MHz), 
           .D(n29431));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i50 (.Q(\data_out_frame[6] [1]), .C(clk16MHz), 
           .D(n29430));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i51 (.Q(\data_out_frame[6] [2]), .C(clk16MHz), 
           .D(n29429));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i52 (.Q(\data_out_frame[6] [3]), .C(clk16MHz), 
           .D(n29428));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i53 (.Q(\data_out_frame[6] [4]), .C(clk16MHz), 
           .D(n29427));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i54 (.Q(\data_out_frame[6] [5]), .C(clk16MHz), 
           .D(n29426));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i55 (.Q(\data_out_frame[6] [6]), .C(clk16MHz), 
           .D(n29425));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i56 (.Q(\data_out_frame[6] [7]), .C(clk16MHz), 
           .D(n29424));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i57 (.Q(\data_out_frame[7] [0]), .C(clk16MHz), 
           .D(n29423));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i58 (.Q(\data_out_frame[7] [1]), .C(clk16MHz), 
           .D(n29422));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i59 (.Q(\data_out_frame[7] [2]), .C(clk16MHz), 
           .D(n29421));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i60 (.Q(\data_out_frame[7] [3]), .C(clk16MHz), 
           .D(n29420));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i1_3_lut_adj_1114 (.I0(n45811), .I1(n46666), .I2(n45874), 
            .I3(GND_net), .O(n51092));
    defparam i1_3_lut_adj_1114.LUT_INIT = 16'h6969;
    SB_DFF data_out_frame_0___i61 (.Q(\data_out_frame[7] [4]), .C(clk16MHz), 
           .D(n29419));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 n56892_bdd_4_lut (.I0(n56892), .I1(\data_out_frame[25] [0]), 
            .I2(\data_out_frame[24] [0]), .I3(byte_transmit_counter[1]), 
            .O(n56895));
    defparam n56892_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_41013 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [7]), .I2(\data_out_frame[27] [7]), 
            .I3(byte_transmit_counter[1]), .O(n56886));
    defparam byte_transmit_counter_0__bdd_4_lut_41013.LUT_INIT = 16'he4aa;
    SB_LUT4 n56886_bdd_4_lut (.I0(n56886), .I1(\data_out_frame[25] [7]), 
            .I2(\data_out_frame[24] [7]), .I3(byte_transmit_counter[1]), 
            .O(n56889));
    defparam n56886_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 equal_2277_i7_2_lut (.I0(Kp_23__N_1305), .I1(\data_in_frame[8][6] ), 
            .I2(GND_net), .I3(GND_net), .O(n7_adj_4673));   // verilog/coms.v(237[9:81])
    defparam equal_2277_i7_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_41008 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [6]), .I2(\data_out_frame[27] [6]), 
            .I3(byte_transmit_counter[1]), .O(n56880));
    defparam byte_transmit_counter_0__bdd_4_lut_41008.LUT_INIT = 16'he4aa;
    SB_LUT4 n56880_bdd_4_lut (.I0(n56880), .I1(\data_out_frame[25] [6]), 
            .I2(\data_out_frame[24] [6]), .I3(byte_transmit_counter[1]), 
            .O(n56883));
    defparam n56880_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i15540_3_lut_4_lut (.I0(n8_adj_4708), .I1(n48984), .I2(rx_data[2]), 
            .I3(\data_in_frame[17] [2]), .O(n29620));
    defparam i15540_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_adj_1115 (.I0(n45874), .I1(\data_in_frame[19] [5]), 
            .I2(n46666), .I3(GND_net), .O(n51209));
    defparam i2_3_lut_adj_1115.LUT_INIT = 16'h9696;
    SB_DFFE data_out_frame_0___i224 (.Q(\data_out_frame[27] [7]), .C(clk16MHz), 
            .E(n28807), .D(n51166));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i2_3_lut_adj_1116 (.I0(\data_in_frame[21] [6]), .I1(n51209), 
            .I2(\data_in_frame[21] [5]), .I3(GND_net), .O(n49352));
    defparam i2_3_lut_adj_1116.LUT_INIT = 16'h6969;
    SB_LUT4 i4_4_lut_adj_1117 (.I0(n27557), .I1(\data_in_frame[1] [4]), 
            .I2(n49466), .I3(n6_adj_4719), .O(n28069));   // verilog/coms.v(79[16:27])
    defparam i4_4_lut_adj_1117.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1118 (.I0(\data_in_frame[8] [3]), .I1(\data_in_frame[8][4] ), 
            .I2(GND_net), .I3(GND_net), .O(n27599));   // verilog/coms.v(76[16:43])
    defparam i1_2_lut_adj_1118.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1119 (.I0(n51092), .I1(\data_in_frame[19] [5]), 
            .I2(\data_in_frame[20] [0]), .I3(GND_net), .O(n49457));
    defparam i2_3_lut_adj_1119.LUT_INIT = 16'h6969;
    SB_LUT4 i1_2_lut_adj_1120 (.I0(\data_in_frame[1] [7]), .I1(\data_in_frame[0] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n49138));   // verilog/coms.v(71[16:69])
    defparam i1_2_lut_adj_1120.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1121 (.I0(\data_in_frame[4] [3]), .I1(\data_in_frame[4] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n49517));   // verilog/coms.v(75[16:43])
    defparam i1_2_lut_adj_1121.LUT_INIT = 16'h6666;
    SB_LUT4 i15541_3_lut_4_lut (.I0(n8_adj_4708), .I1(n48984), .I2(rx_data[1]), 
            .I3(\data_in_frame[17] [1]), .O(n29621));
    defparam i15541_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_3_lut_adj_1122 (.I0(\data_in_frame[0] [2]), .I1(\data_in_frame[0] [1]), 
            .I2(\data_in_frame[2] [3]), .I3(GND_net), .O(n28020));   // verilog/coms.v(76[16:43])
    defparam i1_3_lut_adj_1122.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1123 (.I0(\data_in_frame[15] [0]), .I1(\data_in_frame[12] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n28539));   // verilog/coms.v(72[16:27])
    defparam i1_2_lut_adj_1123.LUT_INIT = 16'h6666;
    SB_LUT4 data_in_frame_14__7__I_0_4037_2_lut (.I0(\data_in_frame[14] [7]), 
            .I1(\data_in_frame[14] [6]), .I2(GND_net), .I3(GND_net), .O(Kp_23__N_985));   // verilog/coms.v(72[16:27])
    defparam data_in_frame_14__7__I_0_4037_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1124 (.I0(\data_in_frame[12] [4]), .I1(n45762), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_4720));
    defparam i1_2_lut_adj_1124.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1125 (.I0(n28020), .I1(n49517), .I2(n49138), 
            .I3(\data_in_frame[2] [1]), .O(Kp_23__N_1209));   // verilog/coms.v(75[16:43])
    defparam i1_4_lut_adj_1125.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1126 (.I0(Kp_23__N_985), .I1(n28539), .I2(\data_in_frame[15] [1]), 
            .I3(\data_in_frame[17] [2]), .O(n52650));
    defparam i1_4_lut_adj_1126.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1127 (.I0(\data_in_frame[4] [6]), .I1(\data_in_frame[7] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n52900));   // verilog/coms.v(74[16:42])
    defparam i1_2_lut_adj_1127.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1128 (.I0(n49252), .I1(n28017), .I2(n28066), 
            .I3(n52900), .O(n27928));   // verilog/coms.v(74[16:42])
    defparam i1_4_lut_adj_1128.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1129 (.I0(Kp_23__N_1209), .I1(Kp_23__N_1206), .I2(\data_in_frame[6] [5]), 
            .I3(\data_in_frame[6] [4]), .O(Kp_23__N_1305));   // verilog/coms.v(77[16:43])
    defparam i1_4_lut_adj_1129.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1130 (.I0(\data_in_frame[9] [0]), .I1(\data_in_frame[11] [2]), 
            .I2(\data_in_frame[9] [1]), .I3(GND_net), .O(n49237));   // verilog/coms.v(72[16:27])
    defparam i2_3_lut_adj_1130.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1131 (.I0(Kp_23__N_1305), .I1(n27928), .I2(GND_net), 
            .I3(GND_net), .O(n28303));   // verilog/coms.v(72[16:27])
    defparam i1_2_lut_adj_1131.LUT_INIT = 16'h6666;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut (.I0(byte_transmit_counter[1]), 
            .I1(n53192), .I2(n53193), .I3(byte_transmit_counter[2]), .O(n56856));
    defparam byte_transmit_counter_1__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n56856_bdd_4_lut (.I0(n56856), .I1(n53190), .I2(n53189), .I3(byte_transmit_counter[2]), 
            .O(n56859));
    defparam n56856_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_40984 (.I0(byte_transmit_counter[1]), 
            .I1(n53135), .I2(n53136), .I3(byte_transmit_counter[2]), .O(n56844));
    defparam byte_transmit_counter_1__bdd_4_lut_40984.LUT_INIT = 16'he4aa;
    SB_LUT4 n56844_bdd_4_lut (.I0(n56844), .I1(n53262), .I2(n53261), .I3(byte_transmit_counter[2]), 
            .O(n56847));
    defparam n56844_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_40974 (.I0(byte_transmit_counter[1]), 
            .I1(n53177), .I2(n53178), .I3(byte_transmit_counter[2]), .O(n56838));
    defparam byte_transmit_counter_1__bdd_4_lut_40974.LUT_INIT = 16'he4aa;
    SB_LUT4 n56838_bdd_4_lut (.I0(n56838), .I1(n53244), .I2(n53243), .I3(byte_transmit_counter[2]), 
            .O(n56841));
    defparam n56838_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_adj_1132 (.I0(\data_in_frame[2] [1]), .I1(\data_in_frame[0] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n52948));   // verilog/coms.v(71[16:69])
    defparam i1_2_lut_adj_1132.LUT_INIT = 16'h6666;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_40969 (.I0(byte_transmit_counter[1]), 
            .I1(n53198), .I2(n53199), .I3(byte_transmit_counter[2]), .O(n56832));
    defparam byte_transmit_counter_1__bdd_4_lut_40969.LUT_INIT = 16'he4aa;
    SB_LUT4 n56832_bdd_4_lut (.I0(n56832), .I1(n53235), .I2(n53234), .I3(byte_transmit_counter[2]), 
            .O(n56835));
    defparam n56832_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i37408_3_lut (.I0(\data_out_frame[14] [4]), .I1(\data_out_frame[15] [4]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n53238));
    defparam i37408_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i37407_3_lut (.I0(\data_out_frame[12] [4]), .I1(\data_out_frame[13] [4]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n53237));
    defparam i37407_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_1133 (.I0(n45897), .I1(n28403), .I2(GND_net), 
            .I3(GND_net), .O(n52656));
    defparam i1_2_lut_adj_1133.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1134 (.I0(n49395), .I1(n46738), .I2(\data_out_frame[24] [0]), 
            .I3(n49605), .O(n10_adj_4721));
    defparam i4_4_lut_adj_1134.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1135 (.I0(\data_out_frame[23] [7]), .I1(n49395), 
            .I2(n49301), .I3(n28368), .O(n25418));
    defparam i3_4_lut_adj_1135.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1136 (.I0(n28138), .I1(n28272), .I2(n27811), 
            .I3(n52650), .O(n52658));
    defparam i1_4_lut_adj_1136.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1137 (.I0(n28406), .I1(n4_adj_4720), .I2(n52658), 
            .I3(n52656), .O(n52664));
    defparam i1_4_lut_adj_1137.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1138 (.I0(n25418), .I1(n49384), .I2(\data_out_frame[24] [1]), 
            .I3(GND_net), .O(n51154));
    defparam i2_3_lut_adj_1138.LUT_INIT = 16'h6969;
    SB_LUT4 i1_3_lut_adj_1139 (.I0(\data_in_frame[19] [4]), .I1(n52394), 
            .I2(n52664), .I3(GND_net), .O(n46852));
    defparam i1_3_lut_adj_1139.LUT_INIT = 16'h6969;
    SB_DFFE data_out_frame_0___i223 (.Q(\data_out_frame[27] [6]), .C(clk16MHz), 
            .E(n28807), .D(n50744));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i15542_3_lut_4_lut (.I0(n8_adj_4708), .I1(n48984), .I2(rx_data[0]), 
            .I3(\data_in_frame[17] [0]), .O(n29622));
    defparam i15542_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_4_lut_adj_1140 (.I0(n49120), .I1(n49608), .I2(n49060), 
            .I3(n52728), .O(n45762));
    defparam i1_4_lut_adj_1140.LUT_INIT = 16'h6996;
    SB_LUT4 i40068_2_lut (.I0(n28124), .I1(\data_in_frame[10] [0]), .I2(GND_net), 
            .I3(GND_net), .O(n55899));   // verilog/coms.v(97[12:25])
    defparam i40068_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_3_lut_adj_1141 (.I0(\data_in_frame[12] [3]), .I1(n49446), 
            .I2(\data_in_frame[14] [4]), .I3(GND_net), .O(n46673));
    defparam i1_3_lut_adj_1141.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_1142 (.I0(n46686), .I1(n49432), .I2(\data_in_frame[20] [4]), 
            .I3(\data_in_frame[18] [4]), .O(n45834));
    defparam i3_4_lut_adj_1142.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1143 (.I0(\data_in_frame[18] [7]), .I1(\data_in_frame[18] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n49482));   // verilog/coms.v(79[16:27])
    defparam i1_2_lut_adj_1143.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1144 (.I0(\data_in_frame[20] [7]), .I1(\data_in_frame[21] [0]), 
            .I2(n45766), .I3(GND_net), .O(n49699));
    defparam i2_3_lut_adj_1144.LUT_INIT = 16'h9696;
    SB_LUT4 i1_4_lut_adj_1145 (.I0(\data_in_frame[21] [2]), .I1(\data_in_frame[21] [3]), 
            .I2(\data_in_frame[20] [6]), .I3(\data_in_frame[21] [1]), .O(n52486));
    defparam i1_4_lut_adj_1145.LUT_INIT = 16'h6996;
    SB_LUT4 i1_3_lut_adj_1146 (.I0(n52486), .I1(\data_in_frame[21] [7]), 
            .I2(\data_in_frame[21] [4]), .I3(GND_net), .O(n52488));
    defparam i1_3_lut_adj_1146.LUT_INIT = 16'h9696;
    SB_LUT4 i1_4_lut_adj_1147 (.I0(\data_in_frame[20] [3]), .I1(n52490), 
            .I2(n49682), .I3(n52488), .O(n52494));
    defparam i1_4_lut_adj_1147.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1148 (.I0(n46682), .I1(n45512), .I2(n45834), 
            .I3(n52494), .O(n52500));
    defparam i1_4_lut_adj_1148.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1149 (.I0(n46917), .I1(n46800), .I2(n46823), 
            .I3(n52500), .O(n52506));
    defparam i1_4_lut_adj_1149.LUT_INIT = 16'h9669;
    SB_LUT4 i1_4_lut_adj_1150 (.I0(n49640), .I1(n49457), .I2(n49352), 
            .I3(n52506), .O(n52512));
    defparam i1_4_lut_adj_1150.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1151 (.I0(n46031), .I1(n51209), .I2(n25607), 
            .I3(n52362), .O(n52368));
    defparam i1_4_lut_adj_1151.LUT_INIT = 16'h9669;
    SB_LUT4 i1_4_lut_adj_1152 (.I0(n52696), .I1(n52368), .I2(n52512), 
            .I3(n49596), .O(n49122));
    defparam i1_4_lut_adj_1152.LUT_INIT = 16'h9669;
    SB_DFFE data_out_frame_0___i222 (.Q(\data_out_frame[27] [5]), .C(clk16MHz), 
            .E(n28807), .D(n50545));   // verilog/coms.v(128[12] 303[6])
    SB_DFFE data_out_frame_0___i221 (.Q(\data_out_frame[27] [4]), .C(clk16MHz), 
            .E(n28807), .D(n49180));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i1_2_lut_adj_1153 (.I0(n45874), .I1(\data_in_frame[19] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n49370));
    defparam i1_2_lut_adj_1153.LUT_INIT = 16'h6666;
    SB_DFFE data_out_frame_0___i220 (.Q(\data_out_frame[27] [3]), .C(clk16MHz), 
            .E(n28807), .D(n49340));   // verilog/coms.v(128[12] 303[6])
    SB_DFFSS \FRAME_MATCHER.i_i30  (.Q(\FRAME_MATCHER.i [30]), .C(clk16MHz), 
            .D(n2_adj_4722), .S(n3_adj_4723));   // verilog/coms.v(128[12] 303[6])
    SB_DFFE data_out_frame_0___i219 (.Q(\data_out_frame[27] [2]), .C(clk16MHz), 
            .E(n28807), .D(n50639));   // verilog/coms.v(128[12] 303[6])
    SB_DFFE data_out_frame_0___i218 (.Q(\data_out_frame[27] [1]), .C(clk16MHz), 
            .E(n28807), .D(n50933));   // verilog/coms.v(128[12] 303[6])
    SB_DFFSS \FRAME_MATCHER.i_i29  (.Q(\FRAME_MATCHER.i [29]), .C(clk16MHz), 
            .D(n2_adj_4724), .S(n3_adj_4725));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i1_2_lut_adj_1154 (.I0(\data_out_frame[21] [6]), .I1(n28368), 
            .I2(GND_net), .I3(GND_net), .O(n49605));
    defparam i1_2_lut_adj_1154.LUT_INIT = 16'h6666;
    SB_LUT4 i5_4_lut_adj_1155 (.I0(n49440), .I1(n49605), .I2(n45782), 
            .I3(n49035), .O(n12_adj_4726));
    defparam i5_4_lut_adj_1155.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1156 (.I0(n50929), .I1(n12_adj_4726), .I2(n49685), 
            .I3(n50579), .O(n51314));
    defparam i6_4_lut_adj_1156.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1157 (.I0(\data_out_frame[24] [2]), .I1(n51314), 
            .I2(GND_net), .I3(GND_net), .O(n49384));
    defparam i1_2_lut_adj_1157.LUT_INIT = 16'h9999;
    SB_LUT4 i4_4_lut_adj_1158 (.I0(n49384), .I1(n27720), .I2(\data_out_frame[24] [3]), 
            .I3(n46744), .O(n10_adj_4727));
    defparam i4_4_lut_adj_1158.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_1159 (.I0(n49379), .I1(n10_adj_4727), .I2(n46865), 
            .I3(GND_net), .O(n51110));
    defparam i5_3_lut_adj_1159.LUT_INIT = 16'h6969;
    SB_DFFSS \FRAME_MATCHER.i_i28  (.Q(\FRAME_MATCHER.i [28]), .C(clk16MHz), 
            .D(n2_adj_4728), .S(n3_adj_4729));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 data_in_frame_17__7__I_0_4040_2_lut (.I0(\data_in_frame[17] [7]), 
            .I1(\data_in_frame[17] [6]), .I2(GND_net), .I3(GND_net), .O(Kp_23__N_1720));   // verilog/coms.v(71[16:27])
    defparam data_in_frame_17__7__I_0_4040_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1160 (.I0(\data_in_frame[1] [1]), .I1(\data_in_frame[1] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n49175));   // verilog/coms.v(74[16:34])
    defparam i1_2_lut_adj_1160.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1161 (.I0(\data_in_frame[1] [5]), .I1(\data_in_frame[1] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n49071));   // verilog/coms.v(76[16:27])
    defparam i1_2_lut_adj_1161.LUT_INIT = 16'h6666;
    SB_LUT4 data_in_frame_1__7__I_0_2_lut (.I0(\data_in_frame[1] [7]), .I1(\data_in_frame[1] [6]), 
            .I2(GND_net), .I3(GND_net), .O(Kp_23__N_1103));   // verilog/coms.v(79[16:27])
    defparam data_in_frame_1__7__I_0_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_3_lut_adj_1162 (.I0(\data_in_frame[1] [0]), .I1(Kp_23__N_1098), 
            .I2(\data_in_frame[0] [5]), .I3(GND_net), .O(n26302));   // verilog/coms.v(78[16:27])
    defparam i1_3_lut_adj_1162.LUT_INIT = 16'h9696;
    SB_DFFSS \FRAME_MATCHER.i_i27  (.Q(\FRAME_MATCHER.i [27]), .C(clk16MHz), 
            .D(n2_adj_4730), .S(n3_adj_4731));   // verilog/coms.v(128[12] 303[6])
    SB_DFFSS \FRAME_MATCHER.i_i26  (.Q(\FRAME_MATCHER.i [26]), .C(clk16MHz), 
            .D(n2_adj_4732), .S(n3_adj_4733));   // verilog/coms.v(128[12] 303[6])
    SB_DFFE data_out_frame_0___i217 (.Q(\data_out_frame[27] [0]), .C(clk16MHz), 
            .E(n28807), .D(n49456));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i1_2_lut_adj_1163 (.I0(\data_in_frame[0] [3]), .I1(\data_in_frame[0] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n49032));   // verilog/coms.v(167[9:87])
    defparam i1_2_lut_adj_1163.LUT_INIT = 16'h6666;
    SB_DFFE data_out_frame_0___i216 (.Q(\data_out_frame[26] [7]), .C(clk16MHz), 
            .E(n28807), .D(n49567));   // verilog/coms.v(128[12] 303[6])
    SB_DFFE data_out_frame_0___i215 (.Q(\data_out_frame[26] [6]), .C(clk16MHz), 
            .E(n28807), .D(n51440));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i1_2_lut_adj_1164 (.I0(\data_in_frame[4] [6]), .I1(\data_in_frame[5] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n49664));
    defparam i1_2_lut_adj_1164.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1165 (.I0(Kp_23__N_1103), .I1(n49071), .I2(n49175), 
            .I3(\data_in_frame[1] [4]), .O(Kp_23__N_1098));   // verilog/coms.v(74[16:34])
    defparam i1_4_lut_adj_1165.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1166 (.I0(n7_adj_4734), .I1(\data_out_frame[21] [7]), 
            .I2(n46905), .I3(n49685), .O(n49379));
    defparam i4_4_lut_adj_1166.LUT_INIT = 16'h9669;
    SB_LUT4 i1_3_lut_adj_1167 (.I0(n49229), .I1(n26302), .I2(\data_in_frame[2] [7]), 
            .I3(GND_net), .O(n49540));   // verilog/coms.v(71[16:27])
    defparam i1_3_lut_adj_1167.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1168 (.I0(\data_in_frame[9] [2]), .I1(\data_in_frame[9] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n27352));   // verilog/coms.v(74[16:42])
    defparam i1_2_lut_adj_1168.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1169 (.I0(\data_in_frame[13] [5]), .I1(\data_in_frame[15] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n49711));   // verilog/coms.v(75[16:43])
    defparam i1_2_lut_adj_1169.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1170 (.I0(n28263), .I1(n49540), .I2(n49144), 
            .I3(n27478), .O(n27954));   // verilog/coms.v(71[16:27])
    defparam i1_4_lut_adj_1170.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1171 (.I0(n27954), .I1(n49711), .I2(n49265), 
            .I3(\data_in_frame[11] [4]), .O(n49418));   // verilog/coms.v(77[16:43])
    defparam i1_4_lut_adj_1171.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1172 (.I0(n27811), .I1(\data_in_frame[13] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n49615));   // verilog/coms.v(77[16:43])
    defparam i1_2_lut_adj_1172.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1173 (.I0(Kp_23__N_1103), .I1(n49074), .I2(n27557), 
            .I3(n52948), .O(Kp_23__N_1203));   // verilog/coms.v(71[16:69])
    defparam i1_4_lut_adj_1173.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1174 (.I0(\data_in_frame[20] [2]), .I1(\data_in_frame[18] [0]), 
            .I2(n49615), .I3(n49418), .O(n49682));   // verilog/coms.v(77[16:43])
    defparam i3_4_lut_adj_1174.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1175 (.I0(Kp_23__N_1103), .I1(n49165), .I2(\data_in_frame[4] [2]), 
            .I3(\data_in_frame[4] [3]), .O(Kp_23__N_1206));   // verilog/coms.v(74[16:42])
    defparam i1_4_lut_adj_1175.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1176 (.I0(\data_out_frame[22] [3]), .I1(n49379), 
            .I2(n46744), .I3(\data_out_frame[20] [3]), .O(n46420));
    defparam i3_4_lut_adj_1176.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1177 (.I0(n46420), .I1(n49443), .I2(GND_net), 
            .I3(GND_net), .O(n49444));
    defparam i1_2_lut_adj_1177.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1178 (.I0(\data_in_frame[6] [3]), .I1(\data_in_frame[6] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n27554));   // verilog/coms.v(86[17:28])
    defparam i1_2_lut_adj_1178.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_4_lut (.I0(n22875), .I1(n39), .I2(n48947), .I3(\FRAME_MATCHER.state [18]), 
            .O(n7_adj_4735));
    defparam i1_2_lut_4_lut.LUT_INIT = 16'hec00;
    SB_LUT4 i1_4_lut_adj_1179 (.I0(n49324), .I1(n49702), .I2(n28079), 
            .I3(Kp_23__N_1324), .O(n52382));
    defparam i1_4_lut_adj_1179.LUT_INIT = 16'h6996;
    SB_DFFE data_out_frame_0___i214 (.Q(\data_out_frame[26] [5]), .C(clk16MHz), 
            .E(n28807), .D(n49444));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i1_2_lut_4_lut_adj_1180 (.I0(n22875), .I1(n39), .I2(n48947), 
            .I3(\FRAME_MATCHER.state [20]), .O(n7_adj_4736));
    defparam i1_2_lut_4_lut_adj_1180.LUT_INIT = 16'hec00;
    SB_LUT4 i1_2_lut_4_lut_adj_1181 (.I0(n22875), .I1(n39), .I2(n48947), 
            .I3(\FRAME_MATCHER.state [24]), .O(n7_adj_4737));
    defparam i1_2_lut_4_lut_adj_1181.LUT_INIT = 16'hec00;
    SB_LUT4 i1_4_lut_adj_1182 (.I0(n52382), .I1(n49060), .I2(n46727), 
            .I3(n49688), .O(n49581));
    defparam i1_4_lut_adj_1182.LUT_INIT = 16'h9669;
    SB_LUT4 i3_4_lut_adj_1183 (.I0(n27554), .I1(Kp_23__N_1206), .I2(Kp_23__N_1203), 
            .I3(\data_in_frame[8][5] ), .O(n27604));
    defparam i3_4_lut_adj_1183.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1184 (.I0(\data_in_frame[3] [1]), .I1(\data_in_frame[7] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n52762));
    defparam i1_2_lut_adj_1184.LUT_INIT = 16'h6666;
    SB_DFFE data_out_frame_0___i213 (.Q(\data_out_frame[26] [4]), .C(clk16MHz), 
            .E(n28807), .D(n51110));   // verilog/coms.v(128[12] 303[6])
    SB_DFFE data_out_frame_0___i212 (.Q(\data_out_frame[26] [3]), .C(clk16MHz), 
            .E(n28807), .D(n51154));   // verilog/coms.v(128[12] 303[6])
    SB_DFFE data_out_frame_0___i211 (.Q(\data_out_frame[26] [2]), .C(clk16MHz), 
            .E(n28807), .D(n50862));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_40964 (.I0(byte_transmit_counter[1]), 
            .I1(n53237), .I2(n53238), .I3(byte_transmit_counter[2]), .O(n56826));
    defparam byte_transmit_counter_1__bdd_4_lut_40964.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_2_lut_4_lut_adj_1185 (.I0(n22875), .I1(n39), .I2(n48947), 
            .I3(\FRAME_MATCHER.state [26]), .O(n36478));
    defparam i1_2_lut_4_lut_adj_1185.LUT_INIT = 16'hec00;
    SB_LUT4 i1_4_lut_adj_1186 (.I0(n49172), .I1(n27863), .I2(n52762), 
            .I3(\data_in_frame[5] [4]), .O(n45804));
    defparam i1_4_lut_adj_1186.LUT_INIT = 16'h6996;
    SB_DFF data_out_frame_0___i62 (.Q(\data_out_frame[7] [5]), .C(clk16MHz), 
           .D(n29418));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i1_4_lut_adj_1187 (.I0(n45804), .I1(n49581), .I2(n49404), 
            .I3(\data_in_frame[9] [0]), .O(n50767));
    defparam i1_4_lut_adj_1187.LUT_INIT = 16'h6996;
    SB_DFFE data_out_frame_0___i210 (.Q(\data_out_frame[26] [1]), .C(clk16MHz), 
            .E(n28807), .D(n51417));   // verilog/coms.v(128[12] 303[6])
    SB_DFFE data_out_frame_0___i209 (.Q(\data_out_frame[26] [0]), .C(clk16MHz), 
            .E(n28807), .D(n50764));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 n56826_bdd_4_lut (.I0(n56826), .I1(n53229), .I2(n53228), .I3(byte_transmit_counter[2]), 
            .O(n56829));
    defparam n56826_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i37344_3_lut (.I0(\data_out_frame[16] [7]), .I1(\data_out_frame[17] [7]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n53174));
    defparam i37344_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_4114_9_lut (.I0(GND_net), .I1(byte_transmit_counter[7]), 
            .I2(GND_net), .I3(n43725), .O(n9046[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4114_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i37345_3_lut (.I0(\data_out_frame[18] [7]), .I1(\data_out_frame[19] [7]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n53175));
    defparam i37345_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_4114_8_lut (.I0(GND_net), .I1(byte_transmit_counter[6]), 
            .I2(GND_net), .I3(n43724), .O(n9046[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4114_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i3_4_lut_adj_1188 (.I0(n45884), .I1(n49460), .I2(n49010), 
            .I3(n46834), .O(n46865));
    defparam i3_4_lut_adj_1188.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1189 (.I0(\data_out_frame[24] [4]), .I1(n49415), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_4738));
    defparam i1_2_lut_adj_1189.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1190 (.I0(\data_out_frame[24] [5]), .I1(n46865), 
            .I2(\data_out_frame[20] [2]), .I3(n6_adj_4738), .O(n51440));
    defparam i4_4_lut_adj_1190.LUT_INIT = 16'h9669;
    SB_CARRY add_4114_8 (.CI(n43724), .I0(byte_transmit_counter[6]), .I1(GND_net), 
            .CO(n43725));
    SB_LUT4 add_4114_7_lut (.I0(GND_net), .I1(byte_transmit_counter[5]), 
            .I2(GND_net), .I3(n43723), .O(n9046[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4114_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i37492_3_lut (.I0(\data_out_frame[22] [7]), .I1(\data_out_frame[23] [7]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n53322));
    defparam i37492_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i37491_3_lut (.I0(\data_out_frame[20] [7]), .I1(\data_out_frame[21] [7]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n53321));
    defparam i37491_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_4114_7 (.CI(n43723), .I0(byte_transmit_counter[5]), .I1(GND_net), 
            .CO(n43724));
    SB_LUT4 select_713_Select_26_i3_2_lut (.I0(\FRAME_MATCHER.i [26]), .I1(n4623), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4733));
    defparam select_713_Select_26_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_713_Select_27_i3_2_lut (.I0(\FRAME_MATCHER.i [27]), .I1(n4623), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4731));
    defparam select_713_Select_27_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4114_6_lut (.I0(GND_net), .I1(byte_transmit_counter[4]), 
            .I2(GND_net), .I3(n43722), .O(n9046[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4114_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4114_6 (.CI(n43722), .I0(byte_transmit_counter[4]), .I1(GND_net), 
            .CO(n43723));
    SB_LUT4 add_4114_5_lut (.I0(GND_net), .I1(byte_transmit_counter[3]), 
            .I2(GND_net), .I3(n43721), .O(n9046[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4114_5_lut.LUT_INIT = 16'hC33C;
    SB_DFF driver_enable_4015 (.Q(DE_c), .C(clk16MHz), .D(n48390));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i96 (.Q(\data_out_frame[11] [7]), .C(clk16MHz), 
           .D(n30058));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i97 (.Q(\data_out_frame[12] [0]), .C(clk16MHz), 
           .D(n30057));   // verilog/coms.v(128[12] 303[6])
    SB_CARRY add_4114_5 (.CI(n43721), .I0(byte_transmit_counter[3]), .I1(GND_net), 
            .CO(n43722));
    SB_DFF data_out_frame_0___i98 (.Q(\data_out_frame[12] [1]), .C(clk16MHz), 
           .D(n30056));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i99 (.Q(\data_out_frame[12] [2]), .C(clk16MHz), 
           .D(n30055));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i100 (.Q(\data_out_frame[12] [3]), .C(clk16MHz), 
           .D(n30054));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i101 (.Q(\data_out_frame[12] [4]), .C(clk16MHz), 
           .D(n30053));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i102 (.Q(\data_out_frame[12] [5]), .C(clk16MHz), 
           .D(n30052));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i103 (.Q(\data_out_frame[12] [6]), .C(clk16MHz), 
           .D(n30051));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i104 (.Q(\data_out_frame[12] [7]), .C(clk16MHz), 
           .D(n30050));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i105 (.Q(\data_out_frame[13] [0]), .C(clk16MHz), 
           .D(n30049));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i106 (.Q(\data_out_frame[13] [1]), .C(clk16MHz), 
           .D(n30048));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i107 (.Q(\data_out_frame[13] [2]), .C(clk16MHz), 
           .D(n30047));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i108 (.Q(\data_out_frame[13] [3]), .C(clk16MHz), 
           .D(n30046));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i109 (.Q(\data_out_frame[13] [4]), .C(clk16MHz), 
           .D(n30045));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i110 (.Q(\data_out_frame[13] [5]), .C(clk16MHz), 
           .D(n30044));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i111 (.Q(\data_out_frame[13] [6]), .C(clk16MHz), 
           .D(n30043));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i112 (.Q(\data_out_frame[13] [7]), .C(clk16MHz), 
           .D(n30042));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i113 (.Q(\data_out_frame[14] [0]), .C(clk16MHz), 
           .D(n30041));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i114 (.Q(\data_out_frame[14] [1]), .C(clk16MHz), 
           .D(n30040));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i115 (.Q(\data_out_frame[14] [2]), .C(clk16MHz), 
           .D(n30039));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i116 (.Q(\data_out_frame[14] [3]), .C(clk16MHz), 
           .D(n30038));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i117 (.Q(\data_out_frame[14] [4]), .C(clk16MHz), 
           .D(n30037));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i118 (.Q(\data_out_frame[14] [5]), .C(clk16MHz), 
           .D(n30036));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i119 (.Q(\data_out_frame[14] [6]), .C(clk16MHz), 
           .D(n30035));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i120 (.Q(\data_out_frame[14] [7]), .C(clk16MHz), 
           .D(n30034));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i121 (.Q(\data_out_frame[15] [0]), .C(clk16MHz), 
           .D(n30033));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i122 (.Q(\data_out_frame[15] [1]), .C(clk16MHz), 
           .D(n30032));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i123 (.Q(\data_out_frame[15] [2]), .C(clk16MHz), 
           .D(n30031));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 add_4114_4_lut (.I0(GND_net), .I1(byte_transmit_counter[2]), 
            .I2(GND_net), .I3(n43720), .O(n9046[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4114_4_lut.LUT_INIT = 16'hC33C;
    SB_DFF data_out_frame_0___i124 (.Q(\data_out_frame[15] [3]), .C(clk16MHz), 
           .D(n30030));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i125 (.Q(\data_out_frame[15] [4]), .C(clk16MHz), 
           .D(n30029));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i126 (.Q(\data_out_frame[15] [5]), .C(clk16MHz), 
           .D(n30028));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i127 (.Q(\data_out_frame[15] [6]), .C(clk16MHz), 
           .D(n30027));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i128 (.Q(\data_out_frame[15] [7]), .C(clk16MHz), 
           .D(n30026));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i129 (.Q(\data_out_frame[16] [0]), .C(clk16MHz), 
           .D(n30025));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i130 (.Q(\data_out_frame[16] [1]), .C(clk16MHz), 
           .D(n30024));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i131 (.Q(\data_out_frame[16] [2]), .C(clk16MHz), 
           .D(n30023));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i132 (.Q(\data_out_frame[16] [3]), .C(clk16MHz), 
           .D(n30022));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i133 (.Q(\data_out_frame[16] [4]), .C(clk16MHz), 
           .D(n30021));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i134 (.Q(\data_out_frame[16] [5]), .C(clk16MHz), 
           .D(n30020));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i135 (.Q(\data_out_frame[16] [6]), .C(clk16MHz), 
           .D(n30019));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i136 (.Q(\data_out_frame[16] [7]), .C(clk16MHz), 
           .D(n30018));   // verilog/coms.v(128[12] 303[6])
    SB_CARRY add_4114_4 (.CI(n43720), .I0(byte_transmit_counter[2]), .I1(GND_net), 
            .CO(n43721));
    SB_DFF data_out_frame_0___i137 (.Q(\data_out_frame[17] [0]), .C(clk16MHz), 
           .D(n30017));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i138 (.Q(\data_out_frame[17] [1]), .C(clk16MHz), 
           .D(n30016));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i1_2_lut_adj_1191 (.I0(n27604), .I1(n49581), .I2(GND_net), 
            .I3(GND_net), .O(n49582));
    defparam i1_2_lut_adj_1191.LUT_INIT = 16'h6666;
    SB_DFF data_out_frame_0___i139 (.Q(\data_out_frame[17] [2]), .C(clk16MHz), 
           .D(n30015));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i140 (.Q(\data_out_frame[17] [3]), .C(clk16MHz), 
           .D(n30014));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i141 (.Q(\data_out_frame[17] [4]), .C(clk16MHz), 
           .D(n30013));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i142 (.Q(\data_out_frame[17] [5]), .C(clk16MHz), 
           .D(n30012));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i143 (.Q(\data_out_frame[17] [6]), .C(clk16MHz), 
           .D(n30011));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i144 (.Q(\data_out_frame[17] [7]), .C(clk16MHz), 
           .D(n30010));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i145 (.Q(\data_out_frame[18] [0]), .C(clk16MHz), 
           .D(n30009));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i146 (.Q(\data_out_frame[18] [1]), .C(clk16MHz), 
           .D(n30008));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i147 (.Q(\data_out_frame[18] [2]), .C(clk16MHz), 
           .D(n30007));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i148 (.Q(\data_out_frame[18] [3]), .C(clk16MHz), 
           .D(n30006));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i149 (.Q(\data_out_frame[18] [4]), .C(clk16MHz), 
           .D(n30005));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i150 (.Q(\data_out_frame[18] [5]), .C(clk16MHz), 
           .D(n30004));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i151 (.Q(\data_out_frame[18] [6]), .C(clk16MHz), 
           .D(n30003));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 select_713_Select_28_i3_2_lut (.I0(\FRAME_MATCHER.i [28]), .I1(n4623), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4729));
    defparam select_713_Select_28_i3_2_lut.LUT_INIT = 16'h8888;
    SB_DFF data_out_frame_0___i152 (.Q(\data_out_frame[18] [7]), .C(clk16MHz), 
           .D(n30002));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i153 (.Q(\data_out_frame[19] [0]), .C(clk16MHz), 
           .D(n30001));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i154 (.Q(\data_out_frame[19] [1]), .C(clk16MHz), 
           .D(n30000));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i155 (.Q(\data_out_frame[19] [2]), .C(clk16MHz), 
           .D(n29999));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i156 (.Q(\data_out_frame[19] [3]), .C(clk16MHz), 
           .D(n29998));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 add_4114_3_lut (.I0(GND_net), .I1(byte_transmit_counter[1]), 
            .I2(GND_net), .I3(n43719), .O(n9046[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4114_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4114_3 (.CI(n43719), .I0(byte_transmit_counter[1]), .I1(GND_net), 
            .CO(n43720));
    SB_LUT4 i15527_3_lut_4_lut (.I0(n8_adj_4739), .I1(n48984), .I2(rx_data[7]), 
            .I3(\data_in_frame[18] [7]), .O(n29607));
    defparam i15527_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_out_frame_0___i157 (.Q(\data_out_frame[19] [4]), .C(clk16MHz), 
           .D(n29997));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i158 (.Q(\data_out_frame[19] [5]), .C(clk16MHz), 
           .D(n29996));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i159 (.Q(\data_out_frame[19] [6]), .C(clk16MHz), 
           .D(n29995));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i160 (.Q(\data_out_frame[19] [7]), .C(clk16MHz), 
           .D(n29994));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i161 (.Q(\data_out_frame[20] [0]), .C(clk16MHz), 
           .D(n29993));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i162 (.Q(\data_out_frame[20] [1]), .C(clk16MHz), 
           .D(n29992));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i163 (.Q(\data_out_frame[20] [2]), .C(clk16MHz), 
           .D(n29991));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i164 (.Q(\data_out_frame[20] [3]), .C(clk16MHz), 
           .D(n29990));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i165 (.Q(\data_out_frame[20] [4]), .C(clk16MHz), 
           .D(n29989));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i166 (.Q(\data_out_frame[20] [5]), .C(clk16MHz), 
           .D(n29988));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i167 (.Q(\data_out_frame[20] [6]), .C(clk16MHz), 
           .D(n29987));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i168 (.Q(\data_out_frame[20] [7]), .C(clk16MHz), 
           .D(n29986));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i169 (.Q(\data_out_frame[21] [0]), .C(clk16MHz), 
           .D(n29985));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_40959 (.I0(byte_transmit_counter[1]), 
            .I1(n53213), .I2(n53214), .I3(byte_transmit_counter[2]), .O(n56820));
    defparam byte_transmit_counter_1__bdd_4_lut_40959.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_2_lut_adj_1192 (.I0(\data_in_frame[18] [6]), .I1(\data_in_frame[18] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n49046));   // verilog/coms.v(79[16:27])
    defparam i1_2_lut_adj_1192.LUT_INIT = 16'h6666;
    SB_DFF data_out_frame_0___i170 (.Q(\data_out_frame[21] [1]), .C(clk16MHz), 
           .D(n29984));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i171 (.Q(\data_out_frame[21] [2]), .C(clk16MHz), 
           .D(n29983));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i172 (.Q(\data_out_frame[21] [3]), .C(clk16MHz), 
           .D(n29982));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i173 (.Q(\data_out_frame[21] [4]), .C(clk16MHz), 
           .D(n29981));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i174 (.Q(\data_out_frame[21] [5]), .C(clk16MHz), 
           .D(n29980));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i175 (.Q(\data_out_frame[21] [6]), .C(clk16MHz), 
           .D(n29979));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i176 (.Q(\data_out_frame[21] [7]), .C(clk16MHz), 
           .D(n29978));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i177 (.Q(\data_out_frame[22] [0]), .C(clk16MHz), 
           .D(n29977));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i178 (.Q(\data_out_frame[22] [1]), .C(clk16MHz), 
           .D(n29976));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i15528_3_lut_4_lut (.I0(n8_adj_4739), .I1(n48984), .I2(rx_data[6]), 
            .I3(\data_in_frame[18] [6]), .O(n29608));
    defparam i15528_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 add_4114_2_lut (.I0(GND_net), .I1(byte_transmit_counter[0]), 
            .I2(tx_transmit_N_3748), .I3(GND_net), .O(n9046[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4114_2_lut.LUT_INIT = 16'hC33C;
    SB_DFF data_out_frame_0___i63 (.Q(\data_out_frame[7] [6]), .C(clk16MHz), 
           .D(n29417));   // verilog/coms.v(128[12] 303[6])
    SB_CARRY add_4114_2 (.CI(GND_net), .I0(byte_transmit_counter[0]), .I1(tx_transmit_N_3748), 
            .CO(n43719));
    SB_DFFESR byte_transmit_counter_i0_i0 (.Q(byte_transmit_counter[0]), .C(clk16MHz), 
            .E(n28738), .D(n9046[0]), .R(n29306));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 n56820_bdd_4_lut (.I0(n56820), .I1(n53208), .I2(n53207), .I3(byte_transmit_counter[2]), 
            .O(n56823));
    defparam n56820_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_4_lut_adj_1193 (.I0(n49582), .I1(n50767), .I2(n45804), 
            .I3(n52632), .O(n46699));
    defparam i1_4_lut_adj_1193.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_40954 (.I0(byte_transmit_counter[1]), 
            .I1(n53291), .I2(n53292), .I3(byte_transmit_counter[2]), .O(n56796));
    defparam byte_transmit_counter_1__bdd_4_lut_40954.LUT_INIT = 16'he4aa;
    SB_LUT4 n56796_bdd_4_lut (.I0(n56796), .I1(n53184), .I2(n53183), .I3(byte_transmit_counter[2]), 
            .O(n56799));
    defparam n56796_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF data_out_frame_0___i64 (.Q(\data_out_frame[7] [7]), .C(clk16MHz), 
           .D(n29416));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i65 (.Q(\data_out_frame[8] [0]), .C(clk16MHz), 
           .D(n29415));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i66 (.Q(\data_out_frame[8] [1]), .C(clk16MHz), 
           .D(n29414));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i67 (.Q(\data_out_frame[8] [2]), .C(clk16MHz), 
           .D(n29412));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i68 (.Q(\data_out_frame[8] [3]), .C(clk16MHz), 
           .D(n29411));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i69 (.Q(\data_out_frame[8] [4]), .C(clk16MHz), 
           .D(n29410));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i70 (.Q(\data_out_frame[8] [5]), .C(clk16MHz), 
           .D(n29408));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i71 (.Q(\data_out_frame[8] [6]), .C(clk16MHz), 
           .D(n29406));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i72 (.Q(\data_out_frame[8] [7]), .C(clk16MHz), 
           .D(n29405));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i73 (.Q(\data_out_frame[9] [0]), .C(clk16MHz), 
           .D(n29404));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i74 (.Q(\data_out_frame[9] [1]), .C(clk16MHz), 
           .D(n29403));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i75 (.Q(\data_out_frame[9] [2]), .C(clk16MHz), 
           .D(n29402));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i76 (.Q(\data_out_frame[9] [3]), .C(clk16MHz), 
           .D(n29401));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i77 (.Q(\data_out_frame[9] [4]), .C(clk16MHz), 
           .D(n29400));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i78 (.Q(\data_out_frame[9] [5]), .C(clk16MHz), 
           .D(n29397));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i79 (.Q(\data_out_frame[9] [6]), .C(clk16MHz), 
           .D(n29396));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i80 (.Q(\data_out_frame[9] [7]), .C(clk16MHz), 
           .D(n29395));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i81 (.Q(\data_out_frame[10] [0]), .C(clk16MHz), 
           .D(n29394));   // verilog/coms.v(128[12] 303[6])
    SB_DFFESR LED_4014 (.Q(LED_c), .C(clk16MHz), .E(n48905), .D(n29136), 
            .R(n50359));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i179 (.Q(\data_out_frame[22] [2]), .C(clk16MHz), 
           .D(n29975));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i15529_3_lut_4_lut (.I0(n8_adj_4739), .I1(n48984), .I2(rx_data[5]), 
            .I3(\data_in_frame[18] [5]), .O(n29609));
    defparam i15529_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_out_frame_0___i180 (.Q(\data_out_frame[22] [3]), .C(clk16MHz), 
           .D(n29974));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i181 (.Q(\data_out_frame[22] [4]), .C(clk16MHz), 
           .D(n29973));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i182 (.Q(\data_out_frame[22] [5]), .C(clk16MHz), 
           .D(n29972));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i183 (.Q(\data_out_frame[22] [6]), .C(clk16MHz), 
           .D(n29971));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i1_2_lut_adj_1194 (.I0(\data_in_frame[15] [5]), .I1(n46823), 
            .I2(GND_net), .I3(GND_net), .O(n46868));
    defparam i1_2_lut_adj_1194.LUT_INIT = 16'h6666;
    SB_DFF data_out_frame_0___i184 (.Q(\data_out_frame[22] [7]), .C(clk16MHz), 
           .D(n29970));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i185 (.Q(\data_out_frame[23] [0]), .C(clk16MHz), 
           .D(n29969));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i186 (.Q(\data_out_frame[23] [1]), .C(clk16MHz), 
           .D(n29968));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i3_4_lut_adj_1195 (.I0(\data_in_frame[15] [4]), .I1(n45897), 
            .I2(\data_in_frame[13] [2]), .I3(\data_in_frame[13] [3]), .O(n49272));
    defparam i3_4_lut_adj_1195.LUT_INIT = 16'h6996;
    SB_DFF data_out_frame_0___i187 (.Q(\data_out_frame[23] [2]), .C(clk16MHz), 
           .D(n29967));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i192 (.Q(\data_in_frame[23] [7]), .C(clk16MHz), 
           .D(n29966));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i191 (.Q(\data_in_frame[23] [6]), .C(clk16MHz), 
           .D(n29965));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i190 (.Q(\data_in_frame[23] [5]), .C(clk16MHz), 
           .D(n29964));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i189 (.Q(\data_in_frame[23] [4]), .C(clk16MHz), 
           .D(n29963));   // verilog/coms.v(128[12] 303[6])
    SB_DFF control_mode_i0_i1 (.Q(control_mode[1]), .C(clk16MHz), .D(n29962));   // verilog/coms.v(128[12] 303[6])
    SB_DFF control_mode_i0_i2 (.Q(control_mode[2]), .C(clk16MHz), .D(n29961));   // verilog/coms.v(128[12] 303[6])
    SB_DFF control_mode_i0_i3 (.Q(control_mode[3]), .C(clk16MHz), .D(n29960));   // verilog/coms.v(128[12] 303[6])
    SB_DFF control_mode_i0_i4 (.Q(control_mode[4]), .C(clk16MHz), .D(n29959));   // verilog/coms.v(128[12] 303[6])
    SB_DFF control_mode_i0_i5 (.Q(control_mode[5]), .C(clk16MHz), .D(n29958));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_40934 (.I0(byte_transmit_counter[1]), 
            .I1(n53171), .I2(n53172), .I3(byte_transmit_counter[2]), .O(n56748));
    defparam byte_transmit_counter_1__bdd_4_lut_40934.LUT_INIT = 16'he4aa;
    SB_DFF control_mode_i0_i6 (.Q(control_mode[6]), .C(clk16MHz), .D(n29957));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 n56748_bdd_4_lut (.I0(n56748), .I1(n53265), .I2(n53264), .I3(byte_transmit_counter[2]), 
            .O(n56751));
    defparam n56748_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF control_mode_i0_i7 (.Q(control_mode[7]), .C(clk16MHz), .D(n29956));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 data_in_frame_13__7__I_0_2_lut (.I0(\data_in_frame[13] [7]), .I1(\data_in_frame[13] [6]), 
            .I2(GND_net), .I3(GND_net), .O(Kp_23__N_1602));   // verilog/coms.v(86[17:28])
    defparam data_in_frame_13__7__I_0_2_lut.LUT_INIT = 16'h6666;
    SB_DFF current_limit_i0_i1 (.Q(current_limit[1]), .C(clk16MHz), .D(n29955));   // verilog/coms.v(128[12] 303[6])
    SB_DFF current_limit_i0_i2 (.Q(current_limit[2]), .C(clk16MHz), .D(n29954));   // verilog/coms.v(128[12] 303[6])
    SB_DFF current_limit_i0_i3 (.Q(current_limit[3]), .C(clk16MHz), .D(n29953));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i10_4_lut_adj_1196 (.I0(\data_in_frame[14] [2]), .I1(n49252), 
            .I2(\data_in_frame[9] [4]), .I3(n49525), .O(n28_adj_4740));
    defparam i10_4_lut_adj_1196.LUT_INIT = 16'h6996;
    SB_DFF current_limit_i0_i4 (.Q(current_limit[4]), .C(clk16MHz), .D(n29952));   // verilog/coms.v(128[12] 303[6])
    SB_DFF current_limit_i0_i5 (.Q(current_limit[5]), .C(clk16MHz), .D(n29951));   // verilog/coms.v(128[12] 303[6])
    SB_DFF current_limit_i0_i6 (.Q(current_limit[6]), .C(clk16MHz), .D(n29950));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i14_3_lut (.I0(n49226), .I1(n28_adj_4740), .I2(n49144), .I3(GND_net), 
            .O(n32));
    defparam i14_3_lut.LUT_INIT = 16'h9696;
    SB_DFF current_limit_i0_i7 (.Q(current_limit[7]), .C(clk16MHz), .D(n29949));   // verilog/coms.v(128[12] 303[6])
    SB_DFF current_limit_i0_i8 (.Q(current_limit[8]), .C(clk16MHz), .D(n29948));   // verilog/coms.v(128[12] 303[6])
    SB_DFF current_limit_i0_i9 (.Q(current_limit[9]), .C(clk16MHz), .D(n29947));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i12_4_lut_adj_1197 (.I0(n27599), .I1(n49172), .I2(\data_in_frame[4] [5]), 
            .I3(n49670), .O(n30));
    defparam i12_4_lut_adj_1197.LUT_INIT = 16'h6996;
    SB_DFF current_limit_i0_i10 (.Q(current_limit[10]), .C(clk16MHz), .D(n29946));   // verilog/coms.v(128[12] 303[6])
    SB_DFF current_limit_i0_i11 (.Q(current_limit[11]), .C(clk16MHz), .D(n29945));   // verilog/coms.v(128[12] 303[6])
    SB_DFF current_limit_i0_i12 (.Q(current_limit[12]), .C(clk16MHz), .D(n29944));   // verilog/coms.v(128[12] 303[6])
    SB_DFF current_limit_i0_i13 (.Q(current_limit[13]), .C(clk16MHz), .D(n29943));   // verilog/coms.v(128[12] 303[6])
    SB_DFF current_limit_i0_i14 (.Q(current_limit[14]), .C(clk16MHz), .D(n29942));   // verilog/coms.v(128[12] 303[6])
    SB_DFF current_limit_i0_i15 (.Q(current_limit[15]), .C(clk16MHz), .D(n29941));   // verilog/coms.v(128[12] 303[6])
    SB_DFF PWMLimit_i0_i1 (.Q(PWMLimit[1]), .C(clk16MHz), .D(n29940));   // verilog/coms.v(128[12] 303[6])
    SB_DFF PWMLimit_i0_i2 (.Q(PWMLimit[2]), .C(clk16MHz), .D(n29939));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i82 (.Q(\data_out_frame[10] [1]), .C(clk16MHz), 
           .D(n29390));   // verilog/coms.v(128[12] 303[6])
    SB_DFF PWMLimit_i0_i3 (.Q(PWMLimit[3]), .C(clk16MHz), .D(n29938));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i83 (.Q(\data_out_frame[10] [2]), .C(clk16MHz), 
           .D(n29389));   // verilog/coms.v(128[12] 303[6])
    SB_DFF PWMLimit_i0_i4 (.Q(PWMLimit[4]), .C(clk16MHz), .D(n29937));   // verilog/coms.v(128[12] 303[6])
    SB_DFF PWMLimit_i0_i5 (.Q(PWMLimit[5]), .C(clk16MHz), .D(n29936));   // verilog/coms.v(128[12] 303[6])
    SB_DFF PWMLimit_i0_i6 (.Q(PWMLimit[6]), .C(clk16MHz), .D(n29935));   // verilog/coms.v(128[12] 303[6])
    SB_DFF PWMLimit_i0_i7 (.Q(PWMLimit[7]), .C(clk16MHz), .D(n29934));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i84 (.Q(\data_out_frame[10] [3]), .C(clk16MHz), 
           .D(n29388));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i1_3_lut_adj_1198 (.I0(\data_in_frame[13] [1]), .I1(\data_in_frame[13] [2]), 
            .I2(\data_in_frame[15] [3]), .I3(GND_net), .O(n52640));
    defparam i1_3_lut_adj_1198.LUT_INIT = 16'h9696;
    SB_LUT4 i13_4_lut (.I0(\data_in_frame[5] [5]), .I1(n49478), .I2(n55899), 
            .I3(n49324), .O(n31_adj_4741));
    defparam i13_4_lut.LUT_INIT = 16'h9669;
    SB_LUT4 i1_4_lut_adj_1199 (.I0(n49335), .I1(n46699), .I2(n28272), 
            .I3(n52640), .O(n50867));
    defparam i1_4_lut_adj_1199.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1200 (.I0(\data_in_frame[15] [4]), .I1(\data_in_frame[15] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n52426));
    defparam i1_2_lut_adj_1200.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1201 (.I0(\data_in_frame[16] [4]), .I1(n52426), 
            .I2(\data_in_frame[16] [6]), .I3(\data_in_frame[15] [7]), .O(n52430));
    defparam i1_4_lut_adj_1201.LUT_INIT = 16'h6996;
    SB_DFF data_out_frame_0___i85 (.Q(\data_out_frame[10] [4]), .C(clk16MHz), 
           .D(n29387));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i86 (.Q(\data_out_frame[10] [5]), .C(clk16MHz), 
           .D(n29386));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i87 (.Q(\data_out_frame[10] [6]), .C(clk16MHz), 
           .D(n29385));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i88 (.Q(\data_out_frame[10] [7]), .C(clk16MHz), 
           .D(n29384));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i89 (.Q(\data_out_frame[11] [0]), .C(clk16MHz), 
           .D(n29383));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i90 (.Q(\data_out_frame[11] [1]), .C(clk16MHz), 
           .D(n29382));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i91 (.Q(\data_out_frame[11] [2]), .C(clk16MHz), 
           .D(n29380));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i92 (.Q(\data_out_frame[11] [3]), .C(clk16MHz), 
           .D(n29379));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i93 (.Q(\data_out_frame[11] [4]), .C(clk16MHz), 
           .D(n29378));   // verilog/coms.v(128[12] 303[6])
    SB_DFF \FRAME_MATCHER.state_i0  (.Q(\FRAME_MATCHER.state[0] ), .C(clk16MHz), 
           .D(n50741));   // verilog/coms.v(128[12] 303[6])
    SB_DFF PWMLimit_i0_i0 (.Q(PWMLimit[0]), .C(clk16MHz), .D(n29376));   // verilog/coms.v(128[12] 303[6])
    SB_DFF current_limit_i0_i0 (.Q(current_limit[0]), .C(clk16MHz), .D(n29375));   // verilog/coms.v(128[12] 303[6])
    SB_DFF control_mode_i0_i0 (.Q(control_mode[0]), .C(clk16MHz), .D(n29374));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i1 (.Q(\data_in_frame[0] [0]), .C(clk16MHz), 
           .D(n29373));   // verilog/coms.v(128[12] 303[6])
    SB_DFF neopxl_color_i0_i0 (.Q(neopxl_color[0]), .C(clk16MHz), .D(n29372));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_0___i1 (.Q(\data_in[0] [0]), .C(clk16MHz), .D(n29371));   // verilog/coms.v(128[12] 303[6])
    SB_DFF Ki_i0 (.Q(\Ki[0] ), .C(clk16MHz), .D(n29370));   // verilog/coms.v(128[12] 303[6])
    SB_DFF Kp_i0 (.Q(\Kp[0] ), .C(clk16MHz), .D(n29369));   // verilog/coms.v(128[12] 303[6])
    SB_DFF IntegralLimit_i0_i0 (.Q(IntegralLimit[0]), .C(clk16MHz), .D(n29368));   // verilog/coms.v(128[12] 303[6])
    SB_DFF PWMLimit_i0_i8 (.Q(PWMLimit[8]), .C(clk16MHz), .D(n29933));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i1_4_lut_adj_1202 (.I0(n49690), .I1(Kp_23__N_985), .I2(n52430), 
            .I3(Kp_23__N_1720), .O(n52436));
    defparam i1_4_lut_adj_1202.LUT_INIT = 16'h6996;
    SB_LUT4 i11_4_lut_adj_1203 (.I0(n49705), .I1(n25500), .I2(n49399), 
            .I3(n28069), .O(n29));
    defparam i11_4_lut_adj_1203.LUT_INIT = 16'h6996;
    SB_DFF PWMLimit_i0_i9 (.Q(PWMLimit[9]), .C(clk16MHz), .D(n29932));   // verilog/coms.v(128[12] 303[6])
    SB_DFF PWMLimit_i0_i10 (.Q(PWMLimit[10]), .C(clk16MHz), .D(n29931));   // verilog/coms.v(128[12] 303[6])
    SB_DFF PWMLimit_i0_i11 (.Q(PWMLimit[11]), .C(clk16MHz), .D(n29930));   // verilog/coms.v(128[12] 303[6])
    SB_DFF PWMLimit_i0_i12 (.Q(PWMLimit[12]), .C(clk16MHz), .D(n29929));   // verilog/coms.v(128[12] 303[6])
    SB_DFF PWMLimit_i0_i13 (.Q(PWMLimit[13]), .C(clk16MHz), .D(n29928));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 select_713_Select_29_i3_2_lut (.I0(\FRAME_MATCHER.i [29]), .I1(n4623), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4725));
    defparam select_713_Select_29_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i4_4_lut_adj_1204 (.I0(n49188), .I1(n45770), .I2(\data_out_frame[19] [7]), 
            .I3(n49364), .O(n10_adj_4742));
    defparam i4_4_lut_adj_1204.LUT_INIT = 16'h6996;
    SB_LUT4 i17_4_lut_adj_1205 (.I0(n29), .I1(n31_adj_4741), .I2(n30), 
            .I3(n32), .O(n45864));
    defparam i17_4_lut_adj_1205.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_40895 (.I0(byte_transmit_counter[1]), 
            .I1(n53279), .I2(n53280), .I3(byte_transmit_counter[2]), .O(n56712));
    defparam byte_transmit_counter_1__bdd_4_lut_40895.LUT_INIT = 16'he4aa;
    SB_LUT4 n56712_bdd_4_lut (.I0(n56712), .I1(n53202), .I2(n53201), .I3(byte_transmit_counter[2]), 
            .O(n56715));
    defparam n56712_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_40866 (.I0(byte_transmit_counter[1]), 
            .I1(n53180), .I2(n53181), .I3(byte_transmit_counter[2]), .O(n56700));
    defparam byte_transmit_counter_1__bdd_4_lut_40866.LUT_INIT = 16'he4aa;
    SB_LUT4 n56700_bdd_4_lut (.I0(n56700), .I1(n53319), .I2(n53318), .I3(byte_transmit_counter[2]), 
            .O(n56703));
    defparam n56700_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3_4_lut_adj_1206 (.I0(\data_in_frame[16] [3]), .I1(\data_in_frame[16] [2]), 
            .I2(n50453), .I3(\data_in_frame[14] [0]), .O(n49367));
    defparam i3_4_lut_adj_1206.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_40856 (.I0(byte_transmit_counter[1]), 
            .I1(n53273), .I2(n53274), .I3(byte_transmit_counter[2]), .O(n56694));
    defparam byte_transmit_counter_1__bdd_4_lut_40856.LUT_INIT = 16'he4aa;
    SB_LUT4 n56694_bdd_4_lut (.I0(n56694), .I1(n53196), .I2(n53195), .I3(byte_transmit_counter[2]), 
            .O(n56697));
    defparam n56694_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i6_4_lut_adj_1207 (.I0(n49711), .I1(n27378), .I2(n49615), 
            .I3(\data_in_frame[14] [0]), .O(n14_adj_4743));   // verilog/coms.v(75[16:43])
    defparam i6_4_lut_adj_1207.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_40851 (.I0(byte_transmit_counter[1]), 
            .I1(n53258), .I2(n53259), .I3(byte_transmit_counter[2]), .O(n56682));
    defparam byte_transmit_counter_1__bdd_4_lut_40851.LUT_INIT = 16'he4aa;
    SB_LUT4 n56682_bdd_4_lut (.I0(n56682), .I1(n53226), .I2(n53225), .I3(byte_transmit_counter[2]), 
            .O(n56685));
    defparam n56682_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i7_4_lut_adj_1208 (.I0(\data_in_frame[13] [6]), .I1(n14_adj_4743), 
            .I2(n10_adj_4744), .I3(n49478), .O(n46458));   // verilog/coms.v(75[16:43])
    defparam i7_4_lut_adj_1208.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1209 (.I0(\data_out_frame[20] [1]), .I1(n45782), 
            .I2(\data_out_frame[22] [4]), .I3(n46753), .O(n49415));
    defparam i3_4_lut_adj_1209.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1210 (.I0(\data_out_frame[22] [3]), .I1(n49415), 
            .I2(GND_net), .I3(GND_net), .O(n46718));
    defparam i1_2_lut_adj_1210.LUT_INIT = 16'h6666;
    SB_DFFE setpoint__i23 (.Q(setpoint[23]), .C(clk16MHz), .E(n28716), 
            .D(n7696));   // verilog/coms.v(128[12] 303[6])
    SB_DFFE setpoint__i22 (.Q(setpoint[22]), .C(clk16MHz), .E(n28716), 
            .D(n7695));   // verilog/coms.v(128[12] 303[6])
    SB_DFFE setpoint__i21 (.Q(setpoint[21]), .C(clk16MHz), .E(n28716), 
            .D(n7694));   // verilog/coms.v(128[12] 303[6])
    SB_DFFE setpoint__i20 (.Q(setpoint[20]), .C(clk16MHz), .E(n28716), 
            .D(n7693));   // verilog/coms.v(128[12] 303[6])
    SB_DFFE setpoint__i19 (.Q(setpoint[19]), .C(clk16MHz), .E(n28716), 
            .D(n7692));   // verilog/coms.v(128[12] 303[6])
    SB_DFFE setpoint__i18 (.Q(setpoint[18]), .C(clk16MHz), .E(n28716), 
            .D(n7691));   // verilog/coms.v(128[12] 303[6])
    SB_DFFE setpoint__i17 (.Q(setpoint[17]), .C(clk16MHz), .E(n28716), 
            .D(n7690));   // verilog/coms.v(128[12] 303[6])
    SB_DFFE setpoint__i16 (.Q(setpoint[16]), .C(clk16MHz), .E(n28716), 
            .D(n7689));   // verilog/coms.v(128[12] 303[6])
    SB_DFFE setpoint__i15 (.Q(setpoint[15]), .C(clk16MHz), .E(n28716), 
            .D(n7688));   // verilog/coms.v(128[12] 303[6])
    SB_DFFE setpoint__i14 (.Q(setpoint[14]), .C(clk16MHz), .E(n28716), 
            .D(n7687));   // verilog/coms.v(128[12] 303[6])
    SB_DFFE setpoint__i13 (.Q(setpoint[13]), .C(clk16MHz), .E(n28716), 
            .D(n7686));   // verilog/coms.v(128[12] 303[6])
    SB_DFFE setpoint__i12 (.Q(setpoint[12]), .C(clk16MHz), .E(n28716), 
            .D(n7685));   // verilog/coms.v(128[12] 303[6])
    SB_DFFE setpoint__i11 (.Q(setpoint[11]), .C(clk16MHz), .E(n28716), 
            .D(n7684));   // verilog/coms.v(128[12] 303[6])
    SB_DFFE setpoint__i10 (.Q(setpoint[10]), .C(clk16MHz), .E(n28716), 
            .D(n7683));   // verilog/coms.v(128[12] 303[6])
    SB_DFFE setpoint__i9 (.Q(setpoint[9]), .C(clk16MHz), .E(n28716), .D(n7682));   // verilog/coms.v(128[12] 303[6])
    SB_DFFE setpoint__i8 (.Q(setpoint[8]), .C(clk16MHz), .E(n28716), .D(n7681));   // verilog/coms.v(128[12] 303[6])
    SB_DFFE setpoint__i7 (.Q(setpoint[7]), .C(clk16MHz), .E(n28716), .D(n7680));   // verilog/coms.v(128[12] 303[6])
    SB_DFFE setpoint__i6 (.Q(setpoint[6]), .C(clk16MHz), .E(n28716), .D(n7679));   // verilog/coms.v(128[12] 303[6])
    SB_DFFE setpoint__i5 (.Q(setpoint[5]), .C(clk16MHz), .E(n28716), .D(n7678));   // verilog/coms.v(128[12] 303[6])
    SB_DFFE setpoint__i4 (.Q(setpoint[4]), .C(clk16MHz), .E(n28716), .D(n7677));   // verilog/coms.v(128[12] 303[6])
    SB_DFFE setpoint__i3 (.Q(setpoint[3]), .C(clk16MHz), .E(n28716), .D(n7676));   // verilog/coms.v(128[12] 303[6])
    SB_DFFE setpoint__i2 (.Q(setpoint[2]), .C(clk16MHz), .E(n28716), .D(n7675));   // verilog/coms.v(128[12] 303[6])
    SB_DFFE setpoint__i1 (.Q(setpoint[1]), .C(clk16MHz), .E(n28716), .D(n7674));   // verilog/coms.v(128[12] 303[6])
    SB_DFFSS \FRAME_MATCHER.state_i31  (.Q(\FRAME_MATCHER.state [31]), .C(clk16MHz), 
            .D(n48446), .S(n48316));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i15530_3_lut_4_lut (.I0(n8_adj_4739), .I1(n48984), .I2(rx_data[4]), 
            .I3(\data_in_frame[18] [4]), .O(n29610));
    defparam i15530_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15531_3_lut_4_lut (.I0(n8_adj_4739), .I1(n48984), .I2(rx_data[3]), 
            .I3(\data_in_frame[18] [3]), .O(n29611));
    defparam i15531_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_2_lut_adj_1211 (.I0(\data_out_frame[15] [3]), .I1(n28496), 
            .I2(GND_net), .I3(GND_net), .O(n45770));
    defparam i2_2_lut_adj_1211.LUT_INIT = 16'h6666;
    SB_LUT4 add_43_33_lut (.I0(n3746), .I1(\FRAME_MATCHER.i [31]), .I2(GND_net), 
            .I3(n43718), .O(n2_adj_4706)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_33_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i4_4_lut_adj_1212 (.I0(\data_out_frame[17] [5]), .I1(n27455), 
            .I2(\data_out_frame[17] [4]), .I3(n6_adj_4745), .O(n49016));
    defparam i4_4_lut_adj_1212.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1213 (.I0(\data_out_frame[24] [4]), .I1(\data_out_frame[24] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n49443));
    defparam i1_2_lut_adj_1213.LUT_INIT = 16'h6666;
    SB_LUT4 add_43_32_lut (.I0(n3746), .I1(\FRAME_MATCHER.i [30]), .I2(GND_net), 
            .I3(n43717), .O(n2_adj_4722)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_32_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_43_32 (.CI(n43717), .I0(\FRAME_MATCHER.i [30]), .I1(GND_net), 
            .CO(n43718));
    SB_LUT4 add_43_31_lut (.I0(n3746), .I1(\FRAME_MATCHER.i [29]), .I2(GND_net), 
            .I3(n43716), .O(n2_adj_4724)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_31_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_43_31 (.CI(n43716), .I0(\FRAME_MATCHER.i [29]), .I1(GND_net), 
            .CO(n43717));
    SB_LUT4 i6_4_lut_adj_1214 (.I0(\data_out_frame[16] [7]), .I1(\data_out_frame[13] [0]), 
            .I2(n49618), .I3(n49693), .O(n15_adj_4746));   // verilog/coms.v(76[16:43])
    defparam i6_4_lut_adj_1214.LUT_INIT = 16'h6996;
    SB_LUT4 add_43_30_lut (.I0(n3746), .I1(\FRAME_MATCHER.i [28]), .I2(GND_net), 
            .I3(n43715), .O(n2_adj_4728)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_30_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i8_4_lut_adj_1215 (.I0(n15_adj_4746), .I1(n49426), .I2(n14_adj_4747), 
            .I3(\data_out_frame[14] [6]), .O(n49395));   // verilog/coms.v(76[16:43])
    defparam i8_4_lut_adj_1215.LUT_INIT = 16'h6996;
    SB_CARRY add_43_30 (.CI(n43715), .I0(\FRAME_MATCHER.i [28]), .I1(GND_net), 
            .CO(n43716));
    SB_LUT4 i2_3_lut_adj_1216 (.I0(n49395), .I1(n27701), .I2(n50579), 
            .I3(GND_net), .O(n49578));
    defparam i2_3_lut_adj_1216.LUT_INIT = 16'h6969;
    SB_LUT4 add_43_29_lut (.I0(n3746), .I1(\FRAME_MATCHER.i [27]), .I2(GND_net), 
            .I3(n43714), .O(n2_adj_4730)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_29_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_2_lut_adj_1217 (.I0(\data_out_frame[22] [1]), .I1(n49631), 
            .I2(GND_net), .I3(GND_net), .O(n46697));
    defparam i1_2_lut_adj_1217.LUT_INIT = 16'h9999;
    SB_LUT4 i15532_3_lut_4_lut (.I0(n8_adj_4739), .I1(n48984), .I2(rx_data[2]), 
            .I3(\data_in_frame[18] [2]), .O(n29612));
    defparam i15532_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1218 (.I0(\data_out_frame[24] [1]), .I1(\data_out_frame[23] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n49355));
    defparam i1_2_lut_adj_1218.LUT_INIT = 16'h6666;
    SB_CARRY add_43_29 (.CI(n43714), .I0(\FRAME_MATCHER.i [27]), .I1(GND_net), 
            .CO(n43715));
    SB_LUT4 i3_4_lut_adj_1219 (.I0(n46172), .I1(\data_out_frame[22] [2]), 
            .I2(\data_out_frame[20] [0]), .I3(n28322), .O(n49010));
    defparam i3_4_lut_adj_1219.LUT_INIT = 16'h6996;
    SB_LUT4 add_43_28_lut (.I0(n3746), .I1(\FRAME_MATCHER.i [26]), .I2(GND_net), 
            .I3(n43713), .O(n2_adj_4732)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_28_lut.LUT_INIT = 16'h8228;
    SB_DFF PWMLimit_i0_i14 (.Q(PWMLimit[14]), .C(clk16MHz), .D(n29927));   // verilog/coms.v(128[12] 303[6])
    SB_CARRY add_43_28 (.CI(n43713), .I0(\FRAME_MATCHER.i [26]), .I1(GND_net), 
            .CO(n43714));
    SB_DFF PWMLimit_i0_i15 (.Q(PWMLimit[15]), .C(clk16MHz), .D(n29926));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 add_43_27_lut (.I0(n3746), .I1(\FRAME_MATCHER.i [25]), .I2(GND_net), 
            .I3(n43712), .O(n2_adj_4748)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_27_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i5_4_lut_adj_1220 (.I0(\data_out_frame[15] [0]), .I1(n49555), 
            .I2(\data_out_frame[13] [0]), .I3(n28448), .O(n12_adj_4749));
    defparam i5_4_lut_adj_1220.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1221 (.I0(\data_out_frame[15] [2]), .I1(n12_adj_4749), 
            .I2(\data_out_frame[19] [4]), .I3(n49332), .O(n50579));
    defparam i6_4_lut_adj_1221.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1222 (.I0(\data_out_frame[21] [7]), .I1(n1995), 
            .I2(\data_out_frame[19] [5]), .I3(n50579), .O(n49301));
    defparam i1_4_lut_adj_1222.LUT_INIT = 16'h9669;
    SB_LUT4 i40119_3_lut_4_lut (.I0(n63), .I1(n27214), .I2(tx_active), 
            .I3(r_SM_Main_2__N_3851[0]), .O(n28738));
    defparam i40119_3_lut_4_lut.LUT_INIT = 16'h5557;
    SB_LUT4 i15533_3_lut_4_lut (.I0(n8_adj_4739), .I1(n48984), .I2(rx_data[1]), 
            .I3(\data_in_frame[18] [1]), .O(n29613));
    defparam i15533_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_2_lut_3_lut (.I0(n27307), .I1(\FRAME_MATCHER.state [1]), 
            .I2(\FRAME_MATCHER.state [2]), .I3(GND_net), .O(n6));   // verilog/coms.v(202[5:24])
    defparam i2_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_DFF PWMLimit_i0_i16 (.Q(PWMLimit[16]), .C(clk16MHz), .D(n29925));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i14_4_lut_adj_1223 (.I0(\data_out_frame[19] [7]), .I1(\data_out_frame[23] [5]), 
            .I2(n46033), .I3(n49708), .O(n36));
    defparam i14_4_lut_adj_1223.LUT_INIT = 16'h6996;
    SB_CARRY add_43_27 (.CI(n43712), .I0(\FRAME_MATCHER.i [25]), .I1(GND_net), 
            .CO(n43713));
    SB_LUT4 i5_3_lut_adj_1224 (.I0(n28151), .I1(n46913), .I2(n49301), 
            .I3(GND_net), .O(n14_adj_4751));
    defparam i5_3_lut_adj_1224.LUT_INIT = 16'h6969;
    SB_LUT4 i6_4_lut_adj_1225 (.I0(n49578), .I1(n28176), .I2(\data_out_frame[21] [0]), 
            .I3(n49321), .O(n15_adj_4752));
    defparam i6_4_lut_adj_1225.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1226 (.I0(n63_adj_6), .I1(n63_adj_4650), 
            .I2(n63_adj_4644), .I3(GND_net), .O(n27180));   // verilog/coms.v(158[6] 160[9])
    defparam i1_2_lut_3_lut_adj_1226.LUT_INIT = 16'h8080;
    SB_LUT4 i8_4_lut_adj_1227 (.I0(n15_adj_4752), .I1(\data_out_frame[21] [6]), 
            .I2(n14_adj_4751), .I3(n49631), .O(n50725));
    defparam i8_4_lut_adj_1227.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_3_lut_4_lut (.I0(n27110), .I1(\FRAME_MATCHER.i [31]), 
            .I2(n22875), .I3(\FRAME_MATCHER.state [2]), .O(n3_adj_4628));   // verilog/coms.v(116[11:12])
    defparam i1_2_lut_3_lut_4_lut.LUT_INIT = 16'hd000;
    SB_LUT4 i1_2_lut_adj_1228 (.I0(\data_in_frame[20] [1]), .I1(n51346), 
            .I2(GND_net), .I3(GND_net), .O(n49640));
    defparam i1_2_lut_adj_1228.LUT_INIT = 16'h9999;
    SB_LUT4 i12_4_lut_adj_1229 (.I0(n49010), .I1(\data_out_frame[23] [7]), 
            .I2(n49673), .I3(n49355), .O(n34));
    defparam i12_4_lut_adj_1229.LUT_INIT = 16'h6996;
    SB_LUT4 i15534_3_lut_4_lut (.I0(n8_adj_4739), .I1(n48984), .I2(rx_data[0]), 
            .I3(\data_in_frame[18] [0]), .O(n29614));
    defparam i15534_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i3_3_lut_4_lut (.I0(n22875), .I1(n6_c), .I2(n27214), .I3(n63), 
            .O(n4_c));
    defparam i3_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i18_4_lut_adj_1230 (.I0(n46697), .I1(n36), .I2(n26_adj_4753), 
            .I3(\data_out_frame[24] [6]), .O(n40_adj_4754));
    defparam i18_4_lut_adj_1230.LUT_INIT = 16'h6996;
    SB_LUT4 i15519_3_lut_4_lut (.I0(n8_adj_4755), .I1(n48984), .I2(rx_data[7]), 
            .I3(\data_in_frame[19] [7]), .O(n29599));
    defparam i15519_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1231 (.I0(n27110), .I1(\FRAME_MATCHER.i [31]), 
            .I2(n22875), .I3(GND_net), .O(n24278));   // verilog/coms.v(228[6] 230[9])
    defparam i1_2_lut_3_lut_adj_1231.LUT_INIT = 16'hd0d0;
    SB_LUT4 i16_4_lut_adj_1232 (.I0(\data_out_frame[23] [1]), .I1(n50725), 
            .I2(\data_out_frame[17] [6]), .I3(n27569), .O(n38_adj_4756));
    defparam i16_4_lut_adj_1232.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1233 (.I0(\data_in_frame[16] [1]), .I1(\data_in_frame[13] [7]), 
            .I2(\data_in_frame[16] [0]), .I3(GND_net), .O(n49690));   // verilog/coms.v(75[16:43])
    defparam i1_2_lut_3_lut_adj_1233.LUT_INIT = 16'h9696;
    SB_LUT4 i17_3_lut (.I0(\data_out_frame[24] [2]), .I1(n34), .I2(\data_out_frame[23] [4]), 
            .I3(GND_net), .O(n39_adj_4757));
    defparam i17_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1234 (.I0(\data_in_frame[11] [4]), .I1(\data_in_frame[9] [5]), 
            .I2(\data_in_frame[11] [6]), .I3(GND_net), .O(n49234));   // verilog/coms.v(76[16:43])
    defparam i1_2_lut_3_lut_adj_1234.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_4_lut_adj_1235 (.I0(n28020), .I1(\data_in_frame[0] [3]), 
            .I2(\data_in_frame[2] [5]), .I3(\data_in_frame[0] [4]), .O(n49252));   // verilog/coms.v(74[16:42])
    defparam i1_2_lut_4_lut_adj_1235.LUT_INIT = 16'h6996;
    SB_LUT4 i3_1_lut_2_lut (.I0(\FRAME_MATCHER.i_31__N_2845 ), .I1(n27217), 
            .I2(GND_net), .I3(GND_net), .O(n3746));
    defparam i3_1_lut_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 i15_4_lut_adj_1236 (.I0(n49593), .I1(n49304), .I2(n49443), 
            .I3(n49016), .O(n37));
    defparam i15_4_lut_adj_1236.LUT_INIT = 16'h6996;
    SB_DFF PWMLimit_i0_i17 (.Q(PWMLimit[17]), .C(clk16MHz), .D(n29924));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i21_4_lut (.I0(n37), .I1(n39_adj_4757), .I2(n38_adj_4756), 
            .I3(n40_adj_4754), .O(n45830));
    defparam i21_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_43_26_lut (.I0(n3746), .I1(\FRAME_MATCHER.i [24]), .I2(GND_net), 
            .I3(n43711), .O(n2_adj_4758)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_26_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i37207_2_lut_4_lut (.I0(\data_in_frame[0] [3]), .I1(\data_in_frame[2] [5]), 
            .I2(\data_in_frame[0] [4]), .I3(n28037), .O(n52970));
    defparam i37207_2_lut_4_lut.LUT_INIT = 16'hff96;
    SB_LUT4 i15520_3_lut_4_lut (.I0(n8_adj_4755), .I1(n48984), .I2(rx_data[6]), 
            .I3(\data_in_frame[19] [6]), .O(n29600));
    defparam i15520_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1237 (.I0(\data_out_frame[25] [7]), .I1(\data_out_frame[24] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_4759));
    defparam i1_2_lut_adj_1237.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_4_lut_adj_1238 (.I0(\FRAME_MATCHER.state [1]), .I1(n49911), 
            .I2(\FRAME_MATCHER.state[3] ), .I3(n49824), .O(n28807));   // verilog/coms.v(128[12] 303[6])
    defparam i2_3_lut_4_lut_adj_1238.LUT_INIT = 16'h0010;
    SB_LUT4 i1_2_lut_4_lut_adj_1239 (.I0(\data_out_frame[23] [3]), .I1(\data_out_frame[20] [7]), 
            .I2(n49275), .I3(n46808), .O(n49255));
    defparam i1_2_lut_4_lut_adj_1239.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1240 (.I0(\data_out_frame[23] [5]), .I1(n46403), 
            .I2(n46738), .I3(GND_net), .O(n27715));
    defparam i1_2_lut_3_lut_adj_1240.LUT_INIT = 16'h9696;
    SB_LUT4 i4_4_lut_adj_1241 (.I0(n45830), .I1(n27715), .I2(n49552), 
            .I3(n6_adj_4759), .O(n49412));
    defparam i4_4_lut_adj_1241.LUT_INIT = 16'h6996;
    SB_DFF PWMLimit_i0_i18 (.Q(PWMLimit[18]), .C(clk16MHz), .D(n29923));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i4_4_lut_adj_1242 (.I0(\data_out_frame[25] [6]), .I1(\data_out_frame[25] [3]), 
            .I2(n49339), .I3(n6_adj_4760), .O(n46729));
    defparam i4_4_lut_adj_1242.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1243 (.I0(n50817), .I1(n50449), .I2(GND_net), 
            .I3(GND_net), .O(n6_adj_4761));
    defparam i1_2_lut_adj_1243.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_3_lut_adj_1244 (.I0(n4_c), .I1(n14_adj_4762), .I2(\FRAME_MATCHER.state [10]), 
            .I3(GND_net), .O(n48370));
    defparam i1_2_lut_3_lut_adj_1244.LUT_INIT = 16'he0e0;
    SB_LUT4 i5_3_lut_4_lut (.I0(\data_out_frame[19] [2]), .I1(n10_adj_4763), 
            .I2(\data_out_frame[15] [0]), .I3(\data_out_frame[15] [1]), 
            .O(n46738));
    defparam i5_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1245 (.I0(n4_c), .I1(n14_adj_4762), .I2(\FRAME_MATCHER.state [11]), 
            .I3(GND_net), .O(n48364));
    defparam i1_2_lut_3_lut_adj_1245.LUT_INIT = 16'he0e0;
    SB_CARRY add_43_26 (.CI(n43711), .I0(\FRAME_MATCHER.i [24]), .I1(GND_net), 
            .CO(n43712));
    SB_LUT4 add_43_25_lut (.I0(n3746), .I1(\FRAME_MATCHER.i [23]), .I2(GND_net), 
            .I3(n43710), .O(n2_adj_4764)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_25_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_2_lut_3_lut_adj_1246 (.I0(n4_c), .I1(n14_adj_4762), .I2(\FRAME_MATCHER.state [12]), 
            .I3(GND_net), .O(n48362));
    defparam i1_2_lut_3_lut_adj_1246.LUT_INIT = 16'he0e0;
    SB_CARRY add_43_25 (.CI(n43710), .I0(\FRAME_MATCHER.i [23]), .I1(GND_net), 
            .CO(n43711));
    SB_DFF PWMLimit_i0_i19 (.Q(PWMLimit[19]), .C(clk16MHz), .D(n29922));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 add_43_24_lut (.I0(n3746), .I1(\FRAME_MATCHER.i [22]), .I2(GND_net), 
            .I3(n43709), .O(n2)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_24_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_2_lut_3_lut_adj_1247 (.I0(n4_c), .I1(n14_adj_4762), .I2(\FRAME_MATCHER.state [13]), 
            .I3(GND_net), .O(n48360));
    defparam i1_2_lut_3_lut_adj_1247.LUT_INIT = 16'he0e0;
    SB_LUT4 i4_4_lut_adj_1248 (.I0(n46729), .I1(n45838), .I2(n50641), 
            .I3(n6_adj_4761), .O(n50933));
    defparam i4_4_lut_adj_1248.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1249 (.I0(n4_c), .I1(n14_adj_4762), .I2(\FRAME_MATCHER.state [14]), 
            .I3(GND_net), .O(n48358));
    defparam i1_2_lut_3_lut_adj_1249.LUT_INIT = 16'he0e0;
    SB_CARRY add_43_24 (.CI(n43709), .I0(\FRAME_MATCHER.i [22]), .I1(GND_net), 
            .CO(n43710));
    SB_LUT4 add_43_23_lut (.I0(n3746), .I1(\FRAME_MATCHER.i [21]), .I2(GND_net), 
            .I3(n43708), .O(n2_adj_4620)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_23_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_43_23 (.CI(n43708), .I0(\FRAME_MATCHER.i [21]), .I1(GND_net), 
            .CO(n43709));
    SB_LUT4 i1_2_lut_adj_1250 (.I0(\data_out_frame[15] [6]), .I1(\data_out_frame[17] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n49364));
    defparam i1_2_lut_adj_1250.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1251 (.I0(n46710), .I1(n49364), .I2(\data_out_frame[18] [0]), 
            .I3(\data_out_frame[17] [6]), .O(n10_adj_4765));
    defparam i4_4_lut_adj_1251.LUT_INIT = 16'h6996;
    SB_LUT4 add_43_22_lut (.I0(n3746), .I1(\FRAME_MATCHER.i [20]), .I2(GND_net), 
            .I3(n43707), .O(n2_adj_4679)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_22_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i4_4_lut_adj_1252 (.I0(n26774), .I1(\data_out_frame[13] [5]), 
            .I2(n50929), .I3(n49559), .O(n10_adj_4766));
    defparam i4_4_lut_adj_1252.LUT_INIT = 16'h9669;
    SB_CARRY add_43_22 (.CI(n43707), .I0(\FRAME_MATCHER.i [20]), .I1(GND_net), 
            .CO(n43708));
    SB_LUT4 add_43_21_lut (.I0(n3746), .I1(\FRAME_MATCHER.i [19]), .I2(GND_net), 
            .I3(n43706), .O(n2_adj_4683)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_21_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_2_lut_3_lut_adj_1253 (.I0(\data_out_frame[16] [7]), .I1(\data_out_frame[16] [6]), 
            .I2(n49624), .I3(GND_net), .O(n49621));
    defparam i1_2_lut_3_lut_adj_1253.LUT_INIT = 16'h9696;
    SB_CARRY add_43_21 (.CI(n43706), .I0(\FRAME_MATCHER.i [19]), .I1(GND_net), 
            .CO(n43707));
    SB_LUT4 i5_3_lut_adj_1254 (.I0(\data_out_frame[15] [7]), .I1(n10_adj_4766), 
            .I2(n46821), .I3(GND_net), .O(n45884));
    defparam i5_3_lut_adj_1254.LUT_INIT = 16'h9696;
    SB_LUT4 add_43_20_lut (.I0(n3746), .I1(\FRAME_MATCHER.i [18]), .I2(GND_net), 
            .I3(n43705), .O(n2_adj_4685)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_20_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_43_20 (.CI(n43705), .I0(\FRAME_MATCHER.i [18]), .I1(GND_net), 
            .CO(n43706));
    SB_LUT4 add_43_19_lut (.I0(n3746), .I1(\FRAME_MATCHER.i [17]), .I2(GND_net), 
            .I3(n43704), .O(n2_adj_4686)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_19_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_2_lut_3_lut_adj_1255 (.I0(n4_c), .I1(n14_adj_4762), .I2(\FRAME_MATCHER.state [15]), 
            .I3(GND_net), .O(n48356));
    defparam i1_2_lut_3_lut_adj_1255.LUT_INIT = 16'he0e0;
    SB_CARRY add_43_19 (.CI(n43704), .I0(\FRAME_MATCHER.i [17]), .I1(GND_net), 
            .CO(n43705));
    SB_LUT4 i1_2_lut_3_lut_adj_1256 (.I0(n4_c), .I1(n14_adj_4762), .I2(\FRAME_MATCHER.state [17]), 
            .I3(GND_net), .O(n48354));
    defparam i1_2_lut_3_lut_adj_1256.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1257 (.I0(n4_c), .I1(n14_adj_4762), .I2(\FRAME_MATCHER.state [25]), 
            .I3(GND_net), .O(n48350));
    defparam i1_2_lut_3_lut_adj_1257.LUT_INIT = 16'he0e0;
    SB_LUT4 add_43_18_lut (.I0(n3746), .I1(\FRAME_MATCHER.i [16]), .I2(GND_net), 
            .I3(n43703), .O(n2_adj_4689)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_18_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_2_lut_adj_1258 (.I0(\data_out_frame[20] [4]), .I1(n46804), 
            .I2(GND_net), .I3(GND_net), .O(n46905));
    defparam i1_2_lut_adj_1258.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_3_lut_adj_1259 (.I0(\data_out_frame[7] [6]), .I1(\data_out_frame[6] [0]), 
            .I2(\data_out_frame[7] [7]), .I3(GND_net), .O(n27359));   // verilog/coms.v(73[16:27])
    defparam i1_2_lut_3_lut_adj_1259.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1260 (.I0(n4_c), .I1(n14_adj_4762), .I2(\FRAME_MATCHER.state [28]), 
            .I3(GND_net), .O(n48348));
    defparam i1_2_lut_3_lut_adj_1260.LUT_INIT = 16'he0e0;
    SB_CARRY add_43_18 (.CI(n43703), .I0(\FRAME_MATCHER.i [16]), .I1(GND_net), 
            .CO(n43704));
    SB_LUT4 add_43_17_lut (.I0(n3746), .I1(\FRAME_MATCHER.i [15]), .I2(GND_net), 
            .I3(n43702), .O(n2_adj_4690)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_17_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_43_17 (.CI(n43702), .I0(\FRAME_MATCHER.i [15]), .I1(GND_net), 
            .CO(n43703));
    SB_LUT4 add_43_16_lut (.I0(n3746), .I1(\FRAME_MATCHER.i [14]), .I2(GND_net), 
            .I3(n43701), .O(n2_adj_4699)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_16_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_43_16 (.CI(n43701), .I0(\FRAME_MATCHER.i [14]), .I1(GND_net), 
            .CO(n43702));
    SB_LUT4 add_43_15_lut (.I0(n3746), .I1(\FRAME_MATCHER.i [13]), .I2(GND_net), 
            .I3(n43700), .O(n2_adj_4701)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_15_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_43_15 (.CI(n43700), .I0(\FRAME_MATCHER.i [13]), .I1(GND_net), 
            .CO(n43701));
    SB_LUT4 add_43_14_lut (.I0(n3746), .I1(\FRAME_MATCHER.i [12]), .I2(GND_net), 
            .I3(n43699), .O(n2_adj_4698)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_14_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_2_lut_3_lut_adj_1261 (.I0(n4_c), .I1(n14_adj_4762), .I2(\FRAME_MATCHER.state [30]), 
            .I3(GND_net), .O(n48346));
    defparam i1_2_lut_3_lut_adj_1261.LUT_INIT = 16'he0e0;
    SB_LUT4 i15521_3_lut_4_lut (.I0(n8_adj_4755), .I1(n48984), .I2(rx_data[5]), 
            .I3(\data_in_frame[19] [5]), .O(n29601));
    defparam i15521_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_CARRY add_43_14 (.CI(n43699), .I0(\FRAME_MATCHER.i [12]), .I1(GND_net), 
            .CO(n43700));
    SB_LUT4 i1_2_lut_3_lut_adj_1262 (.I0(n4_c), .I1(n14_adj_4762), .I2(\FRAME_MATCHER.state [31]), 
            .I3(GND_net), .O(n48316));
    defparam i1_2_lut_3_lut_adj_1262.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1263 (.I0(n39), .I1(n49), .I2(\FRAME_MATCHER.state [10]), 
            .I3(GND_net), .O(n48456));
    defparam i1_2_lut_3_lut_adj_1263.LUT_INIT = 16'he0e0;
    SB_LUT4 add_43_13_lut (.I0(n3746), .I1(\FRAME_MATCHER.i [11]), .I2(GND_net), 
            .I3(n43698), .O(n2_adj_4767)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_13_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_43_13 (.CI(n43698), .I0(\FRAME_MATCHER.i [11]), .I1(GND_net), 
            .CO(n43699));
    SB_LUT4 i1_2_lut_3_lut_adj_1264 (.I0(n39), .I1(n49), .I2(\FRAME_MATCHER.state [11]), 
            .I3(GND_net), .O(n48458));
    defparam i1_2_lut_3_lut_adj_1264.LUT_INIT = 16'he0e0;
    SB_LUT4 add_43_12_lut (.I0(n3746), .I1(\FRAME_MATCHER.i [10]), .I2(GND_net), 
            .I3(n43697), .O(n2_adj_4696)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_12_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_43_12 (.CI(n43697), .I0(\FRAME_MATCHER.i [10]), .I1(GND_net), 
            .CO(n43698));
    SB_LUT4 i1_2_lut_3_lut_adj_1265 (.I0(n39), .I1(n49), .I2(\FRAME_MATCHER.state [12]), 
            .I3(GND_net), .O(n48460));
    defparam i1_2_lut_3_lut_adj_1265.LUT_INIT = 16'he0e0;
    SB_LUT4 add_43_11_lut (.I0(n3746), .I1(\FRAME_MATCHER.i [9]), .I2(GND_net), 
            .I3(n43696), .O(n2_adj_4695)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_11_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_43_11 (.CI(n43696), .I0(\FRAME_MATCHER.i [9]), .I1(GND_net), 
            .CO(n43697));
    SB_LUT4 i1_2_lut_3_lut_adj_1266 (.I0(\data_out_frame[6] [0]), .I1(\data_out_frame[5] [7]), 
            .I2(\data_out_frame[5] [6]), .I3(GND_net), .O(n49534));   // verilog/coms.v(75[16:27])
    defparam i1_2_lut_3_lut_adj_1266.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1267 (.I0(n46033), .I1(n49552), .I2(\data_out_frame[22] [4]), 
            .I3(GND_net), .O(n46827));
    defparam i2_3_lut_adj_1267.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1268 (.I0(n39), .I1(n49), .I2(\FRAME_MATCHER.state [13]), 
            .I3(GND_net), .O(n48462));
    defparam i1_2_lut_3_lut_adj_1268.LUT_INIT = 16'he0e0;
    SB_LUT4 i15522_3_lut_4_lut (.I0(n8_adj_4755), .I1(n48984), .I2(rx_data[4]), 
            .I3(\data_in_frame[19] [4]), .O(n29602));
    defparam i15522_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 add_43_10_lut (.I0(n3746), .I1(\FRAME_MATCHER.i [8]), .I2(GND_net), 
            .I3(n43695), .O(n2_adj_4693)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_10_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_43_10 (.CI(n43695), .I0(\FRAME_MATCHER.i [8]), .I1(GND_net), 
            .CO(n43696));
    SB_LUT4 i1_2_lut_3_lut_adj_1269 (.I0(n39), .I1(n49), .I2(\FRAME_MATCHER.state [17]), 
            .I3(GND_net), .O(n48480));
    defparam i1_2_lut_3_lut_adj_1269.LUT_INIT = 16'he0e0;
    SB_LUT4 add_43_9_lut (.I0(n3746), .I1(\FRAME_MATCHER.i [7]), .I2(GND_net), 
            .I3(n43694), .O(n2_adj_4692)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_9_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_43_9 (.CI(n43694), .I0(\FRAME_MATCHER.i [7]), .I1(GND_net), 
            .CO(n43695));
    SB_LUT4 add_43_8_lut (.I0(n3746), .I1(\FRAME_MATCHER.i [6]), .I2(GND_net), 
            .I3(n43693), .O(n2_adj_4691)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_8_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i22412_2_lut_3_lut (.I0(n39), .I1(n49), .I2(\FRAME_MATCHER.state [19]), 
            .I3(GND_net), .O(n36472));
    defparam i22412_2_lut_3_lut.LUT_INIT = 16'he0e0;
    SB_LUT4 i3_4_lut_adj_1270 (.I0(\data_out_frame[25] [1]), .I1(n49454), 
            .I2(\data_out_frame[25] [0]), .I3(n50240), .O(n50639));
    defparam i3_4_lut_adj_1270.LUT_INIT = 16'h6996;
    SB_LUT4 i22413_2_lut_3_lut (.I0(n39), .I1(n49), .I2(\FRAME_MATCHER.state [21]), 
            .I3(GND_net), .O(n36474));
    defparam i22413_2_lut_3_lut.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1271 (.I0(n39), .I1(n49), .I2(\FRAME_MATCHER.state [22]), 
            .I3(GND_net), .O(n7_adj_4768));
    defparam i1_2_lut_3_lut_adj_1271.LUT_INIT = 16'he0e0;
    SB_CARRY add_43_8 (.CI(n43693), .I0(\FRAME_MATCHER.i [6]), .I1(GND_net), 
            .CO(n43694));
    SB_LUT4 add_43_7_lut (.I0(n3746), .I1(\FRAME_MATCHER.i [5]), .I2(GND_net), 
            .I3(n43692), .O(n2_adj_4687)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_7_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i22414_2_lut_3_lut (.I0(n39), .I1(n49), .I2(\FRAME_MATCHER.state [23]), 
            .I3(GND_net), .O(n36476));
    defparam i22414_2_lut_3_lut.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1272 (.I0(n39), .I1(n49), .I2(\FRAME_MATCHER.state [25]), 
            .I3(GND_net), .O(n48482));
    defparam i1_2_lut_3_lut_adj_1272.LUT_INIT = 16'he0e0;
    SB_LUT4 select_713_Select_30_i3_2_lut (.I0(\FRAME_MATCHER.i [30]), .I1(n4623), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4723));
    defparam select_713_Select_30_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_3_lut_adj_1273 (.I0(n1945), .I1(n46695), .I2(n49284), .I3(GND_net), 
            .O(n49559));
    defparam i2_3_lut_adj_1273.LUT_INIT = 16'h9696;
    SB_CARRY add_43_7 (.CI(n43692), .I0(\FRAME_MATCHER.i [5]), .I1(GND_net), 
            .CO(n43693));
    SB_LUT4 i22416_2_lut_3_lut (.I0(n39), .I1(n49), .I2(\FRAME_MATCHER.state [27]), 
            .I3(GND_net), .O(n36480));
    defparam i22416_2_lut_3_lut.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1274 (.I0(n39), .I1(n49), .I2(\FRAME_MATCHER.state [28]), 
            .I3(GND_net), .O(n48484));
    defparam i1_2_lut_3_lut_adj_1274.LUT_INIT = 16'he0e0;
    SB_LUT4 add_43_6_lut (.I0(n3746), .I1(\FRAME_MATCHER.i [4]), .I2(GND_net), 
            .I3(n43691), .O(n2_adj_4684)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_6_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_43_6 (.CI(n43691), .I0(\FRAME_MATCHER.i [4]), .I1(GND_net), 
            .CO(n43692));
    SB_LUT4 i2_3_lut_adj_1275 (.I0(n49559), .I1(n49655), .I2(n49318), 
            .I3(GND_net), .O(n46744));
    defparam i2_3_lut_adj_1275.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1276 (.I0(n39), .I1(n49), .I2(\FRAME_MATCHER.state [29]), 
            .I3(GND_net), .O(n48408));
    defparam i1_2_lut_3_lut_adj_1276.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1277 (.I0(n39), .I1(n49), .I2(\FRAME_MATCHER.state [30]), 
            .I3(GND_net), .O(n48486));
    defparam i1_2_lut_3_lut_adj_1277.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_adj_1278 (.I0(\data_out_frame[20] [3]), .I1(n46744), 
            .I2(GND_net), .I3(GND_net), .O(n46753));
    defparam i1_2_lut_adj_1278.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1279 (.I0(n49335), .I1(n27612), .I2(n49633), 
            .I3(n52436), .O(n52442));
    defparam i1_4_lut_adj_1279.LUT_INIT = 16'h6996;
    SB_LUT4 add_43_5_lut (.I0(n3746), .I1(\FRAME_MATCHER.i [3]), .I2(GND_net), 
            .I3(n43690), .O(n2_adj_4682)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_5_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_43_5 (.CI(n43690), .I0(\FRAME_MATCHER.i [3]), .I1(GND_net), 
            .CO(n43691));
    SB_LUT4 i1_2_lut_3_lut_adj_1280 (.I0(n39), .I1(n49), .I2(\FRAME_MATCHER.state [31]), 
            .I3(GND_net), .O(n48446));
    defparam i1_2_lut_3_lut_adj_1280.LUT_INIT = 16'he0e0;
    SB_LUT4 add_43_4_lut (.I0(n3746), .I1(\FRAME_MATCHER.i [2]), .I2(GND_net), 
            .I3(n43689), .O(n2_adj_4681)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_4_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_43_4 (.CI(n43689), .I0(\FRAME_MATCHER.i [2]), .I1(GND_net), 
            .CO(n43690));
    SB_LUT4 add_43_3_lut (.I0(n3746), .I1(\FRAME_MATCHER.i [1]), .I2(GND_net), 
            .I3(n43688), .O(n2_adj_4680)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_3_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i15523_3_lut_4_lut (.I0(n8_adj_4755), .I1(n48984), .I2(rx_data[3]), 
            .I3(\data_in_frame[19] [3]), .O(n29603));
    defparam i15523_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_CARRY add_43_3 (.CI(n43688), .I0(\FRAME_MATCHER.i [1]), .I1(GND_net), 
            .CO(n43689));
    SB_LUT4 i1_2_lut_adj_1281 (.I0(\data_out_frame[22] [6]), .I1(\data_out_frame[24] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n49593));
    defparam i1_2_lut_adj_1281.LUT_INIT = 16'h6666;
    SB_LUT4 add_43_2_lut (.I0(n3746), .I1(\FRAME_MATCHER.i [0]), .I2(n161), 
            .I3(GND_net), .O(n2_adj_4624)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_2_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_2_lut_4_lut_adj_1282 (.I0(n12_adj_4769), .I1(n49624), .I2(n28346), 
            .I3(GND_net), .O(n46897));
    defparam i1_2_lut_4_lut_adj_1282.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1283 (.I0(n46842), .I1(n46677), .I2(\data_out_frame[20] [5]), 
            .I3(GND_net), .O(n28176));
    defparam i2_3_lut_adj_1283.LUT_INIT = 16'h6969;
    SB_DFF data_out_frame_0___i94 (.Q(\data_out_frame[11] [5]), .C(clk16MHz), 
           .D(n29356));   // verilog/coms.v(128[12] 303[6])
    SB_CARRY add_43_2 (.CI(GND_net), .I0(\FRAME_MATCHER.i [0]), .I1(n161), 
            .CO(n43688));
    SB_DFF deadband_i0_i0 (.Q(deadband[0]), .C(clk16MHz), .D(n29355));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i1_2_lut_3_lut_adj_1284 (.I0(\data_in_frame[13] [3]), .I1(\data_in_frame[13] [4]), 
            .I2(\data_in_frame[13] [5]), .I3(GND_net), .O(n49111));   // verilog/coms.v(86[17:63])
    defparam i1_2_lut_3_lut_adj_1284.LUT_INIT = 16'h9696;
    SB_DFF PWMLimit_i0_i20 (.Q(PWMLimit[20]), .C(clk16MHz), .D(n29921));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i1_2_lut_adj_1285 (.I0(\data_out_frame[25] [2]), .I1(\data_out_frame[25] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n49339));
    defparam i1_2_lut_adj_1285.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1286 (.I0(n28176), .I1(n49593), .I2(n49347), 
            .I3(n49268), .O(n50817));
    defparam i3_4_lut_adj_1286.LUT_INIT = 16'h6996;
    SB_DFF PWMLimit_i0_i21 (.Q(PWMLimit[21]), .C(clk16MHz), .D(n29920));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i1_4_lut_adj_1287 (.I0(n49367), .I1(n52442), .I2(n49418), 
            .I3(n49240), .O(n52448));
    defparam i1_4_lut_adj_1287.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1288 (.I0(\data_in_frame[13] [3]), .I1(\data_in_frame[13] [4]), 
            .I2(n27612), .I3(GND_net), .O(n49295));   // verilog/coms.v(86[17:63])
    defparam i1_2_lut_3_lut_adj_1288.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1289 (.I0(n50817), .I1(n49339), .I2(GND_net), 
            .I3(GND_net), .O(n49340));
    defparam i1_2_lut_adj_1289.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_2_lut (.I0(n46673), .I1(\data_in_frame[16] [6]), .I2(GND_net), 
            .I3(GND_net), .O(n49646));
    defparam i1_2_lut_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i1_2_lut_adj_1290 (.I0(\data_out_frame[22] [7]), .I1(\data_out_frame[23] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n49708));
    defparam i1_2_lut_adj_1290.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_4_lut_adj_1291 (.I0(\data_out_frame[6] [3]), .I1(\data_out_frame[4] [2]), 
            .I2(\data_out_frame[4] [1]), .I3(n49534), .O(n49223));   // verilog/coms.v(75[16:43])
    defparam i1_2_lut_4_lut_adj_1291.LUT_INIT = 16'h6996;
    SB_DFF PWMLimit_i0_i22 (.Q(PWMLimit[22]), .C(clk16MHz), .D(n29919));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i1_2_lut_adj_1292 (.I0(n50375), .I1(n49350), .I2(GND_net), 
            .I3(GND_net), .O(n49630));
    defparam i1_2_lut_adj_1292.LUT_INIT = 16'h9999;
    SB_LUT4 i1_2_lut_4_lut_adj_1293 (.I0(n46673), .I1(n49052), .I2(\data_in_frame[16] [6]), 
            .I3(\data_in_frame[17] [0]), .O(n46832));
    defparam i1_2_lut_4_lut_adj_1293.LUT_INIT = 16'h9669;
    SB_DFF PWMLimit_i0_i23 (.Q(PWMLimit[23]), .C(clk16MHz), .D(n29918));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i1_2_lut_3_lut_adj_1294 (.I0(\data_out_frame[4] [0]), .I1(\data_out_frame[4] [1]), 
            .I2(\data_out_frame[6] [2]), .I3(GND_net), .O(n27319));   // verilog/coms.v(75[16:43])
    defparam i1_2_lut_3_lut_adj_1294.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1295 (.I0(\data_out_frame[10] [2]), .I1(\data_out_frame[10] [3]), 
            .I2(n49181), .I3(GND_net), .O(n6_adj_4770));   // verilog/coms.v(86[17:70])
    defparam i1_2_lut_3_lut_adj_1295.LUT_INIT = 16'h9696;
    SB_DFF \FRAME_MATCHER.state_i2  (.Q(\FRAME_MATCHER.state [2]), .C(clk16MHz), 
           .D(n57033));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i1_4_lut_adj_1296 (.I0(n46749), .I1(n28132), .I2(n52448), 
            .I3(n49272), .O(n52454));
    defparam i1_4_lut_adj_1296.LUT_INIT = 16'h9669;
    SB_DFFSS \FRAME_MATCHER.state_i30  (.Q(\FRAME_MATCHER.state [30]), .C(clk16MHz), 
            .D(n48486), .S(n48346));   // verilog/coms.v(128[12] 303[6])
    SB_DFFSS \FRAME_MATCHER.state_i29  (.Q(\FRAME_MATCHER.state [29]), .C(clk16MHz), 
            .D(n48408), .S(n37148));   // verilog/coms.v(128[12] 303[6])
    SB_DFFSS \FRAME_MATCHER.state_i28  (.Q(\FRAME_MATCHER.state [28]), .C(clk16MHz), 
            .D(n48484), .S(n48348));   // verilog/coms.v(128[12] 303[6])
    SB_DFFSS \FRAME_MATCHER.state_i27  (.Q(\FRAME_MATCHER.state [27]), .C(clk16MHz), 
            .D(n36480), .S(n37146));   // verilog/coms.v(128[12] 303[6])
    SB_DFFSS \FRAME_MATCHER.state_i26  (.Q(\FRAME_MATCHER.state [26]), .C(clk16MHz), 
            .D(n36478), .S(n48218));   // verilog/coms.v(128[12] 303[6])
    SB_DFFSS \FRAME_MATCHER.state_i25  (.Q(\FRAME_MATCHER.state [25]), .C(clk16MHz), 
            .D(n48482), .S(n48350));   // verilog/coms.v(128[12] 303[6])
    SB_DFFSS \FRAME_MATCHER.state_i24  (.Q(\FRAME_MATCHER.state [24]), .C(clk16MHz), 
            .D(n7_adj_4737), .S(n48212));   // verilog/coms.v(128[12] 303[6])
    SB_DFFSS \FRAME_MATCHER.state_i23  (.Q(\FRAME_MATCHER.state [23]), .C(clk16MHz), 
            .D(n36476), .S(n37142));   // verilog/coms.v(128[12] 303[6])
    SB_DFFSS \FRAME_MATCHER.state_i22  (.Q(\FRAME_MATCHER.state [22]), .C(clk16MHz), 
            .D(n7_adj_4768), .S(n48250));   // verilog/coms.v(128[12] 303[6])
    SB_DFFSS \FRAME_MATCHER.state_i21  (.Q(\FRAME_MATCHER.state [21]), .C(clk16MHz), 
            .D(n36474), .S(n37140));   // verilog/coms.v(128[12] 303[6])
    SB_DFFSS \FRAME_MATCHER.state_i20  (.Q(\FRAME_MATCHER.state [20]), .C(clk16MHz), 
            .D(n7_adj_4736), .S(n48214));   // verilog/coms.v(128[12] 303[6])
    SB_DFFSS \FRAME_MATCHER.state_i19  (.Q(\FRAME_MATCHER.state [19]), .C(clk16MHz), 
            .D(n36472), .S(n37136));   // verilog/coms.v(128[12] 303[6])
    SB_DFFSS \FRAME_MATCHER.state_i18  (.Q(\FRAME_MATCHER.state [18]), .C(clk16MHz), 
            .D(n7_adj_4735), .S(n48216));   // verilog/coms.v(128[12] 303[6])
    SB_DFFSS \FRAME_MATCHER.state_i17  (.Q(\FRAME_MATCHER.state [17]), .C(clk16MHz), 
            .D(n48480), .S(n48354));   // verilog/coms.v(128[12] 303[6])
    SB_DFFSS \FRAME_MATCHER.state_i16  (.Q(\FRAME_MATCHER.state [16]), .C(clk16MHz), 
            .D(n7_adj_4633), .S(n48220));   // verilog/coms.v(128[12] 303[6])
    SB_DFFSS \FRAME_MATCHER.state_i15  (.Q(\FRAME_MATCHER.state [15]), .C(clk16MHz), 
            .D(n48478), .S(n48356));   // verilog/coms.v(128[12] 303[6])
    SB_DFFSS \FRAME_MATCHER.state_i14  (.Q(\FRAME_MATCHER.state [14]), .C(clk16MHz), 
            .D(n48470), .S(n48358));   // verilog/coms.v(128[12] 303[6])
    SB_DFFSS \FRAME_MATCHER.state_i13  (.Q(\FRAME_MATCHER.state [13]), .C(clk16MHz), 
            .D(n48462), .S(n48360));   // verilog/coms.v(128[12] 303[6])
    SB_DFFSS \FRAME_MATCHER.state_i12  (.Q(\FRAME_MATCHER.state [12]), .C(clk16MHz), 
            .D(n48460), .S(n48362));   // verilog/coms.v(128[12] 303[6])
    SB_DFFSS \FRAME_MATCHER.state_i11  (.Q(\FRAME_MATCHER.state [11]), .C(clk16MHz), 
            .D(n48458), .S(n48364));   // verilog/coms.v(128[12] 303[6])
    SB_DFFSS \FRAME_MATCHER.state_i10  (.Q(\FRAME_MATCHER.state [10]), .C(clk16MHz), 
            .D(n48456), .S(n48370));   // verilog/coms.v(128[12] 303[6])
    SB_DFFSS \FRAME_MATCHER.state_i9  (.Q(\FRAME_MATCHER.state [9]), .C(clk16MHz), 
            .D(n7_adj_4771), .S(n48224));   // verilog/coms.v(128[12] 303[6])
    SB_DFFSS \FRAME_MATCHER.state_i8  (.Q(\FRAME_MATCHER.state [8]), .C(clk16MHz), 
            .D(n48454), .S(n48314));   // verilog/coms.v(128[12] 303[6])
    SB_DFFSS \FRAME_MATCHER.state_i7  (.Q(\FRAME_MATCHER.state [7]), .C(clk16MHz), 
            .D(n48452), .S(n48366));   // verilog/coms.v(128[12] 303[6])
    SB_DFFSS \FRAME_MATCHER.state_i6  (.Q(\FRAME_MATCHER.state [6]), .C(clk16MHz), 
            .D(n7_adj_4772), .S(n48222));   // verilog/coms.v(128[12] 303[6])
    SB_DFFSS \FRAME_MATCHER.state_i5  (.Q(\FRAME_MATCHER.state [5]), .C(clk16MHz), 
            .D(n48450), .S(n48368));   // verilog/coms.v(128[12] 303[6])
    SB_DFFSS \FRAME_MATCHER.state_i4  (.Q(\FRAME_MATCHER.state [4]), .C(clk16MHz), 
            .D(n48448), .S(n48310));   // verilog/coms.v(128[12] 303[6])
    SB_DFFSS \FRAME_MATCHER.state_i3  (.Q(\FRAME_MATCHER.state[3] ), .C(clk16MHz), 
            .D(n48308), .S(n48404));   // verilog/coms.v(128[12] 303[6])
    SB_DFFSS \FRAME_MATCHER.state_i1  (.Q(\FRAME_MATCHER.state [1]), .C(clk16MHz), 
            .D(n48306), .S(n57034));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i1_2_lut_4_lut_adj_1297 (.I0(n1945), .I1(n45750), .I2(n28346), 
            .I3(n28180), .O(n46695));
    defparam i1_2_lut_4_lut_adj_1297.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1298 (.I0(\data_out_frame[8] [6]), .I1(\data_out_frame[8] [3]), 
            .I2(\data_out_frame[8] [4]), .I3(\data_out_frame[8] [5]), .O(n49472));   // verilog/coms.v(77[16:43])
    defparam i1_2_lut_4_lut_adj_1298.LUT_INIT = 16'h6996;
    SB_DFFSS \FRAME_MATCHER.i_i11  (.Q(\FRAME_MATCHER.i [11]), .C(clk16MHz), 
            .D(n2_adj_4767), .S(n3_adj_4773));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i1_4_lut_adj_1299 (.I0(n49249), .I1(n45766), .I2(n45914), 
            .I3(n52454), .O(n52460));
    defparam i1_4_lut_adj_1299.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1300 (.I0(n49367), .I1(n45864), .I2(Kp_23__N_1602), 
            .I3(GND_net), .O(n50279));
    defparam i2_3_lut_adj_1300.LUT_INIT = 16'h9696;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_41032 (.I0(byte_transmit_counter[3]), 
            .I1(n56697), .I2(n54597), .I3(byte_transmit_counter[4]), .O(n56910));
    defparam byte_transmit_counter_3__bdd_4_lut_41032.LUT_INIT = 16'he4aa;
    SB_LUT4 i2_3_lut_adj_1301 (.I0(\data_out_frame[18] [2]), .I1(n28196), 
            .I2(n46172), .I3(GND_net), .O(n49318));
    defparam i2_3_lut_adj_1301.LUT_INIT = 16'h9696;
    SB_DFFSS \FRAME_MATCHER.i_i25  (.Q(\FRAME_MATCHER.i [25]), .C(clk16MHz), 
            .D(n2_adj_4748), .S(n3_adj_4774));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i3_4_lut_adj_1302 (.I0(n46842), .I1(n49318), .I2(n46821), 
            .I3(n46802), .O(n46804));
    defparam i3_4_lut_adj_1302.LUT_INIT = 16'h6996;
    SB_DFFSS \FRAME_MATCHER.i_i24  (.Q(\FRAME_MATCHER.i [24]), .C(clk16MHz), 
            .D(n2_adj_4758), .S(n3_adj_4775));   // verilog/coms.v(128[12] 303[6])
    SB_DFFSS \FRAME_MATCHER.i_i23  (.Q(\FRAME_MATCHER.i [23]), .C(clk16MHz), 
            .D(n2_adj_4764), .S(n3_adj_4776));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i95 (.Q(\data_out_frame[11] [6]), .C(clk16MHz), 
           .D(n29353));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_40841 (.I0(byte_transmit_counter[1]), 
            .I1(n53222), .I2(n53223), .I3(byte_transmit_counter[2]), .O(n56670));
    defparam byte_transmit_counter_1__bdd_4_lut_40841.LUT_INIT = 16'he4aa;
    SB_LUT4 i2_3_lut_4_lut_adj_1303 (.I0(\data_out_frame[16] [4]), .I1(n49197), 
            .I2(\data_out_frame[16] [5]), .I3(n49184), .O(n1945));
    defparam i2_3_lut_4_lut_adj_1303.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1304 (.I0(\data_out_frame[22] [6]), .I1(n27424), 
            .I2(n49679), .I3(n49537), .O(n16_adj_4777));
    defparam i6_4_lut_adj_1304.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1305 (.I0(\data_in_frame[12] [5]), .I1(n27692), 
            .I2(\data_in_frame[12] [4]), .I3(n45762), .O(n45914));
    defparam i1_2_lut_3_lut_4_lut_adj_1305.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1306 (.I0(\data_out_frame[6] [1]), .I1(\data_out_frame[5] [7]), 
            .I2(\data_out_frame[4] [0]), .I3(\data_out_frame[11] [0]), .O(n8_adj_4778));   // verilog/coms.v(77[16:43])
    defparam i1_2_lut_4_lut_adj_1306.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1307 (.I0(\data_out_frame[6] [1]), .I1(\data_out_frame[5] [7]), 
            .I2(\data_out_frame[4] [0]), .I3(GND_net), .O(n49514));
    defparam i1_2_lut_3_lut_adj_1307.LUT_INIT = 16'h9696;
    SB_LUT4 n56670_bdd_4_lut (.I0(n56670), .I1(n53232), .I2(n53231), .I3(byte_transmit_counter[2]), 
            .O(n56673));
    defparam n56670_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_3_lut_adj_1308 (.I0(\data_out_frame[11] [3]), .I1(n1168), 
            .I2(\data_out_frame[4] [7]), .I3(GND_net), .O(n49649));   // verilog/coms.v(86[17:70])
    defparam i1_2_lut_3_lut_adj_1308.LUT_INIT = 16'h9696;
    SB_LUT4 i4_4_lut_adj_1309 (.I0(n49295), .I1(n46793), .I2(\data_in_frame[16] [2]), 
            .I3(n49569), .O(n10_adj_4779));
    defparam i4_4_lut_adj_1309.LUT_INIT = 16'h6996;
    SB_LUT4 i2_2_lut_3_lut_adj_1310 (.I0(\data_out_frame[4] [4]), .I1(\data_out_frame[4] [3]), 
            .I2(\data_out_frame[6] [5]), .I3(GND_net), .O(n27584));   // verilog/coms.v(86[17:28])
    defparam i2_2_lut_3_lut_adj_1310.LUT_INIT = 16'h9696;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_40831 (.I0(byte_transmit_counter[1]), 
            .I1(n53186), .I2(n53187), .I3(byte_transmit_counter[2]), .O(n56664));
    defparam byte_transmit_counter_1__bdd_4_lut_40831.LUT_INIT = 16'he4aa;
    SB_LUT4 i7_4_lut_adj_1311 (.I0(n46913), .I1(n49630), .I2(n49708), 
            .I3(n49392), .O(n17_adj_4780));
    defparam i7_4_lut_adj_1311.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1312 (.I0(\data_out_frame[15] [2]), .I1(\data_out_frame[15] [3]), 
            .I2(\data_out_frame[13] [0]), .I3(n26802), .O(n46834));
    defparam i1_2_lut_4_lut_adj_1312.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1313 (.I0(\data_out_frame[16] [4]), .I1(n49197), 
            .I2(\data_out_frame[18] [7]), .I3(GND_net), .O(n49429));
    defparam i1_2_lut_3_lut_adj_1313.LUT_INIT = 16'h9696;
    SB_LUT4 i9_4_lut_adj_1314 (.I0(n17_adj_4780), .I1(n28170), .I2(n16_adj_4777), 
            .I3(n46804), .O(n50240));
    defparam i9_4_lut_adj_1314.LUT_INIT = 16'h6996;
    SB_LUT4 n56664_bdd_4_lut (.I0(n56664), .I1(n53241), .I2(n53240), .I3(byte_transmit_counter[2]), 
            .O(n56667));
    defparam n56664_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i2_3_lut_4_lut_adj_1315 (.I0(\data_out_frame[16] [3]), .I1(\data_out_frame[16] [2]), 
            .I2(\data_out_frame[18] [4]), .I3(n49546), .O(n46677));   // verilog/coms.v(86[17:28])
    defparam i2_3_lut_4_lut_adj_1315.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1316 (.I0(\data_out_frame[16] [3]), .I1(\data_out_frame[16] [2]), 
            .I2(\data_out_frame[16] [1]), .I3(GND_net), .O(n49197));   // verilog/coms.v(86[17:28])
    defparam i1_2_lut_3_lut_adj_1316.LUT_INIT = 16'h9696;
    SB_LUT4 i5_3_lut_adj_1317 (.I0(\data_in_frame[13] [7]), .I1(n10_adj_4779), 
            .I2(\data_in_frame[16] [1]), .I3(GND_net), .O(n46800));
    defparam i5_3_lut_adj_1317.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1318 (.I0(\data_out_frame[15] [3]), .I1(\data_out_frame[13] [0]), 
            .I2(n26802), .I3(GND_net), .O(n49280));
    defparam i1_2_lut_3_lut_adj_1318.LUT_INIT = 16'h9696;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_6_i7_3_lut_4_lut (.I0(byte_transmit_counter[2]), 
            .I1(byte_transmit_counter[1]), .I2(n53401), .I3(n53399), .O(n7_adj_4781));   // verilog/coms.v(107[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_6_i7_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_7_i7_3_lut_4_lut (.I0(byte_transmit_counter[2]), 
            .I1(byte_transmit_counter[1]), .I2(n53317), .I3(n53315), .O(n7_adj_4711));   // verilog/coms.v(107[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_7_i7_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 i1_2_lut_adj_1319 (.I0(\data_in_frame[19] [7]), .I1(n46848), 
            .I2(GND_net), .I3(GND_net), .O(n49596));
    defparam i1_2_lut_adj_1319.LUT_INIT = 16'h9999;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_3_i7_3_lut_4_lut (.I0(byte_transmit_counter[2]), 
            .I1(byte_transmit_counter[1]), .I2(n53155), .I3(n53153), .O(n7_adj_4709));   // verilog/coms.v(107[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_3_i7_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_4_i7_3_lut_4_lut (.I0(byte_transmit_counter[2]), 
            .I1(byte_transmit_counter[1]), .I2(n53149), .I3(n53147), .O(n7_adj_4704));   // verilog/coms.v(107[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_4_i7_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_5_i7_3_lut_4_lut (.I0(byte_transmit_counter[2]), 
            .I1(byte_transmit_counter[1]), .I2(n53143), .I3(n53141), .O(n7_adj_4703));   // verilog/coms.v(107[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_5_i7_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 i3_4_lut_adj_1320 (.I0(n50279), .I1(n49640), .I2(Kp_23__N_1895), 
            .I3(n46458), .O(n49358));
    defparam i3_4_lut_adj_1320.LUT_INIT = 16'h9669;
    SB_LUT4 i1_4_lut_adj_1321 (.I0(n46868), .I1(n50867), .I2(n52460), 
            .I3(n45802), .O(n52466));
    defparam i1_4_lut_adj_1321.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1322 (.I0(\data_out_frame[23] [1]), .I1(n49528), 
            .I2(n49572), .I3(\data_out_frame[20] [7]), .O(n49347));
    defparam i1_4_lut_adj_1322.LUT_INIT = 16'h9669;
    SB_LUT4 i2_4_lut_adj_1323 (.I0(n49178), .I1(n49347), .I2(\data_out_frame[25] [2]), 
            .I3(n50240), .O(n49180));
    defparam i2_4_lut_adj_1323.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_2_i7_3_lut_4_lut (.I0(byte_transmit_counter[2]), 
            .I1(byte_transmit_counter[1]), .I2(n53164), .I3(n53162), .O(n7_c));   // verilog/coms.v(107[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_2_i7_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_40826 (.I0(byte_transmit_counter[1]), 
            .I1(n53159), .I2(n53160), .I3(byte_transmit_counter[2]), .O(n56646));
    defparam byte_transmit_counter_1__bdd_4_lut_40826.LUT_INIT = 16'he4aa;
    SB_LUT4 i37422_3_lut (.I0(\data_out_frame[16] [6]), .I1(\data_out_frame[17] [6]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n53252));
    defparam i37422_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_1_i7_3_lut_4_lut (.I0(byte_transmit_counter[2]), 
            .I1(byte_transmit_counter[1]), .I2(n53170), .I3(n53168), .O(n7_adj_4622));   // verilog/coms.v(107[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_1_i7_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 n56646_bdd_4_lut (.I0(n56646), .I1(n53253), .I2(n53252), .I3(byte_transmit_counter[2]), 
            .O(n56649));
    defparam n56646_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i37423_3_lut (.I0(\data_out_frame[18] [6]), .I1(\data_out_frame[19] [6]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n53253));
    defparam i37423_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_0_i7_3_lut_4_lut (.I0(byte_transmit_counter[2]), 
            .I1(byte_transmit_counter[1]), .I2(n53308), .I3(n53306), .O(n7_adj_4700));   // verilog/coms.v(107[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_0_i7_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 i1_2_lut_adj_1324 (.I0(n49331), .I1(\data_in_frame[16] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n52556));
    defparam i1_2_lut_adj_1324.LUT_INIT = 16'h9999;
    SB_LUT4 i1_4_lut_adj_1325 (.I0(n46708), .I1(n51124), .I2(n45512), 
            .I3(n52556), .O(n46848));
    defparam i1_4_lut_adj_1325.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1326 (.I0(\data_out_frame[14] [2]), .I1(n51147), 
            .I2(n49261), .I3(GND_net), .O(n49546));   // verilog/coms.v(86[17:70])
    defparam i1_2_lut_3_lut_adj_1326.LUT_INIT = 16'h6969;
    SB_LUT4 i2_3_lut_4_lut_adj_1327 (.I0(\data_out_frame[5] [3]), .I1(\data_out_frame[9] [7]), 
            .I2(\data_out_frame[10] [0]), .I3(\data_out_frame[5] [5]), .O(n49409));
    defparam i2_3_lut_4_lut_adj_1327.LUT_INIT = 16'h6996;
    SB_LUT4 i15524_3_lut_4_lut (.I0(n8_adj_4755), .I1(n48984), .I2(rx_data[2]), 
            .I3(\data_in_frame[19] [2]), .O(n29604));
    defparam i15524_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_adj_1328 (.I0(\data_out_frame[16] [1]), .I1(n49498), 
            .I2(n28573), .I3(GND_net), .O(n49655));
    defparam i2_3_lut_adj_1328.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1329 (.I0(\data_out_frame[9] [1]), .I1(\data_out_frame[9] [3]), 
            .I2(n49661), .I3(GND_net), .O(n6_adj_4782));   // verilog/coms.v(86[17:70])
    defparam i1_2_lut_3_lut_adj_1329.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1330 (.I0(\FRAME_MATCHER.state[0] ), 
            .I1(n27223), .I2(\FRAME_MATCHER.state [1]), .I3(\FRAME_MATCHER.state [2]), 
            .O(n63_adj_4662));
    defparam i1_2_lut_3_lut_4_lut_adj_1330.LUT_INIT = 16'hefff;
    SB_LUT4 i1_4_lut_adj_1331 (.I0(\data_out_frame[18] [3]), .I1(n49261), 
            .I2(n6_adj_4783), .I3(n46802), .O(n46842));
    defparam i1_4_lut_adj_1331.LUT_INIT = 16'h9669;
    SB_LUT4 i1_4_lut_adj_1332 (.I0(n46816), .I1(n51092), .I2(n46708), 
            .I3(n52466), .O(n51346));
    defparam i1_4_lut_adj_1332.LUT_INIT = 16'h6996;
    SB_LUT4 i1_3_lut_4_lut_adj_1333 (.I0(\FRAME_MATCHER.state[0] ), .I1(n27223), 
            .I2(n2_adj_4661), .I3(n27248), .O(n4623));
    defparam i1_3_lut_4_lut_adj_1333.LUT_INIT = 16'hf0e0;
    SB_LUT4 i2_3_lut_adj_1334 (.I0(n46808), .I1(\data_out_frame[18] [5]), 
            .I2(\data_out_frame[16] [4]), .I3(GND_net), .O(n49350));
    defparam i2_3_lut_adj_1334.LUT_INIT = 16'h6969;
    SB_LUT4 i1_2_lut_adj_1335 (.I0(\data_out_frame[20] [3]), .I1(\data_out_frame[20] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n27720));
    defparam i1_2_lut_adj_1335.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1336 (.I0(\data_out_frame[15] [1]), .I1(n26802), 
            .I2(GND_net), .I3(GND_net), .O(n27894));
    defparam i1_2_lut_adj_1336.LUT_INIT = 16'h6666;
    SB_LUT4 i37330_3_lut (.I0(\data_out_frame[22] [6]), .I1(\data_out_frame[23] [6]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n53160));
    defparam i37330_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i37329_3_lut (.I0(\data_out_frame[20] [6]), .I1(\data_out_frame[21] [6]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n53159));
    defparam i37329_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1337 (.I0(\FRAME_MATCHER.state[0] ), 
            .I1(n27223), .I2(\FRAME_MATCHER.state [1]), .I3(\FRAME_MATCHER.state [2]), 
            .O(n27214));   // verilog/coms.v(128[12] 303[6])
    defparam i1_2_lut_3_lut_4_lut_adj_1337.LUT_INIT = 16'hdfff;
    SB_LUT4 i1_2_lut_4_lut_adj_1338 (.I0(\FRAME_MATCHER.state [2]), .I1(\FRAME_MATCHER.state [1]), 
            .I2(n27223), .I3(\FRAME_MATCHER.state[0] ), .O(\FRAME_MATCHER.i_31__N_2845 ));
    defparam i1_2_lut_4_lut_adj_1338.LUT_INIT = 16'h0400;
    SB_LUT4 i2_3_lut_adj_1339 (.I0(n49091), .I1(n28496), .I2(n26802), 
            .I3(GND_net), .O(n49555));
    defparam i2_3_lut_adj_1339.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_4_lut_adj_1340 (.I0(\FRAME_MATCHER.state [2]), .I1(\FRAME_MATCHER.state [1]), 
            .I2(n27223), .I3(\FRAME_MATCHER.state[0] ), .O(n60));
    defparam i1_2_lut_4_lut_adj_1340.LUT_INIT = 16'hfffb;
    SB_LUT4 i3_4_lut_adj_1341 (.I0(\data_out_frame[17] [3]), .I1(n49555), 
            .I2(n49280), .I3(n27894), .O(n49673));
    defparam i3_4_lut_adj_1341.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1342 (.I0(\data_out_frame[19] [0]), .I1(\data_out_frame[19] [1]), 
            .I2(n46370), .I3(GND_net), .O(n49392));
    defparam i1_2_lut_3_lut_adj_1342.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1343 (.I0(\data_out_frame[5] [0]), .I1(n1168), 
            .I2(\data_out_frame[7] [0]), .I3(\data_out_frame[4] [6]), .O(n28296));   // verilog/coms.v(86[17:70])
    defparam i2_3_lut_4_lut_adj_1343.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1344 (.I0(\data_out_frame[5] [0]), .I1(n1168), 
            .I2(\data_out_frame[4] [5]), .I3(\data_out_frame[6] [7]), .O(n49147));   // verilog/coms.v(86[17:70])
    defparam i2_3_lut_4_lut_adj_1344.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1345 (.I0(\data_out_frame[5] [2]), .I1(\data_out_frame[5] [1]), 
            .I2(n1191), .I3(n49200), .O(n1168));   // verilog/coms.v(74[16:34])
    defparam i2_3_lut_4_lut_adj_1345.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1346 (.I0(\data_out_frame[5] [2]), .I1(\data_out_frame[5] [1]), 
            .I2(\data_out_frame[4] [7]), .I3(GND_net), .O(n49135));   // verilog/coms.v(74[16:34])
    defparam i1_2_lut_3_lut_adj_1346.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1347 (.I0(n28318), .I1(n46834), .I2(\data_out_frame[19] [6]), 
            .I3(n49016), .O(n28368));
    defparam i2_3_lut_4_lut_adj_1347.LUT_INIT = 16'h6996;
    SB_LUT4 i13_3_lut_4_lut (.I0(n28318), .I1(n46834), .I2(n27915), .I3(\data_out_frame[11] [5]), 
            .O(n38_adj_4784));
    defparam i13_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1348 (.I0(\data_out_frame[15] [4]), .I1(\data_out_frame[15] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n28322));
    defparam i1_2_lut_adj_1348.LUT_INIT = 16'h6666;
    SB_LUT4 i2_2_lut_3_lut_4_lut (.I0(\data_in_frame[16] [1]), .I1(\data_in_frame[13] [7]), 
            .I2(\data_in_frame[16] [0]), .I3(n27954), .O(n10_adj_4744));   // verilog/coms.v(75[16:43])
    defparam i2_2_lut_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1349 (.I0(\data_out_frame[5] [1]), .I1(n28_adj_4785), 
            .I2(n28296), .I3(\data_out_frame[11] [4]), .O(n49661));   // verilog/coms.v(86[17:28])
    defparam i2_3_lut_4_lut_adj_1349.LUT_INIT = 16'h6996;
    SB_LUT4 i15525_3_lut_4_lut (.I0(n8_adj_4755), .I1(n48984), .I2(rx_data[1]), 
            .I3(\data_in_frame[19] [1]), .O(n29605));
    defparam i15525_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i5_4_lut_adj_1350 (.I0(\data_out_frame[18] [1]), .I1(n28322), 
            .I2(\data_out_frame[17] [7]), .I3(n28346), .O(n13));
    defparam i5_4_lut_adj_1350.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1351 (.I0(n13), .I1(n11_adj_4786), .I2(\data_out_frame[15] [6]), 
            .I3(n51468), .O(n49284));
    defparam i7_4_lut_adj_1351.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_3_lut_adj_1352 (.I0(\data_out_frame[5] [1]), .I1(n28_adj_4785), 
            .I2(n49107), .I3(GND_net), .O(n49502));   // verilog/coms.v(86[17:28])
    defparam i1_2_lut_3_lut_adj_1352.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1353 (.I0(n51399), .I1(\data_out_frame[12] [1]), 
            .I2(n49658), .I3(GND_net), .O(n6_adj_4787));
    defparam i1_2_lut_3_lut_adj_1353.LUT_INIT = 16'h6969;
    SB_LUT4 i1_2_lut_adj_1354 (.I0(\data_out_frame[17] [3]), .I1(\data_out_frame[17] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n49332));
    defparam i1_2_lut_adj_1354.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1355 (.I0(\data_out_frame[19] [7]), .I1(\data_out_frame[19] [6]), 
            .I2(\data_out_frame[17] [4]), .I3(\data_out_frame[17] [6]), 
            .O(n49460));
    defparam i3_4_lut_adj_1355.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1356 (.I0(\data_out_frame[17] [5]), .I1(\data_out_frame[18] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n49188));
    defparam i1_2_lut_adj_1356.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_4_lut_adj_1357 (.I0(n51399), .I1(\data_out_frame[12] [1]), 
            .I2(\data_out_frame[14] [3]), .I3(n27335), .O(n50291));
    defparam i2_3_lut_4_lut_adj_1357.LUT_INIT = 16'h9669;
    SB_LUT4 i12_4_lut_adj_1358 (.I0(n28180), .I1(\data_out_frame[18] [2]), 
            .I2(\data_out_frame[16] [0]), .I3(\data_out_frame[19] [4]), 
            .O(n28_adj_4788));   // verilog/coms.v(76[16:43])
    defparam i12_4_lut_adj_1358.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1359 (.I0(n28069), .I1(\data_in_frame[6] [3]), 
            .I2(Kp_23__N_1203), .I3(n27599), .O(n28079));   // verilog/coms.v(75[16:43])
    defparam i1_2_lut_3_lut_4_lut_adj_1359.LUT_INIT = 16'h6996;
    SB_LUT4 i3_2_lut_3_lut_4_lut (.I0(\data_out_frame[13] [5]), .I1(n26774), 
            .I2(n28180), .I3(\data_out_frame[15] [7]), .O(n11_adj_4786));
    defparam i3_2_lut_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i10_4_lut_adj_1360 (.I0(\data_out_frame[18] [3]), .I1(n49188), 
            .I2(n49460), .I3(\data_out_frame[18] [5]), .O(n26_adj_4789));   // verilog/coms.v(76[16:43])
    defparam i10_4_lut_adj_1360.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1361 (.I0(\data_out_frame[13] [5]), .I1(n26774), 
            .I2(n46172), .I3(GND_net), .O(n46710));
    defparam i1_2_lut_3_lut_adj_1361.LUT_INIT = 16'h9696;
    SB_LUT4 i5_3_lut_4_lut_adj_1362 (.I0(\data_out_frame[13] [5]), .I1(n26774), 
            .I2(n10_adj_4742), .I3(n28322), .O(n45782));
    defparam i5_3_lut_4_lut_adj_1362.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1363 (.I0(\data_out_frame[13] [5]), .I1(n26774), 
            .I2(n49655), .I3(\data_out_frame[15] [7]), .O(n46802));
    defparam i1_2_lut_3_lut_4_lut_adj_1363.LUT_INIT = 16'h6996;
    SB_LUT4 i15526_3_lut_4_lut (.I0(n8_adj_4755), .I1(n48984), .I2(rx_data[0]), 
            .I3(\data_in_frame[19] [0]), .O(n29606));
    defparam i15526_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_4_lut_adj_1364 (.I0(n1169), .I1(n10_adj_4790), .I2(n49147), 
            .I3(\data_out_frame[13] [7]), .O(n49498));
    defparam i1_2_lut_4_lut_adj_1364.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_40811 (.I0(byte_transmit_counter[1]), 
            .I1(n53321), .I2(n53322), .I3(byte_transmit_counter[2]), .O(n56634));
    defparam byte_transmit_counter_1__bdd_4_lut_40811.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_2_lut_4_lut_adj_1365 (.I0(n1169), .I1(n10_adj_4790), .I2(n49147), 
            .I3(n49298), .O(n46821));
    defparam i1_2_lut_4_lut_adj_1365.LUT_INIT = 16'h6996;
    SB_LUT4 i1_3_lut_4_lut_adj_1366 (.I0(n49331), .I1(n49046), .I2(n49562), 
            .I3(n46749), .O(n52690));
    defparam i1_3_lut_4_lut_adj_1366.LUT_INIT = 16'h9669;
    SB_LUT4 i114_3_lut_4_lut (.I0(tx_transmit_N_3748), .I1(n36465), .I2(n22875), 
            .I3(n27214), .O(n110));   // verilog/coms.v(215[11:56])
    defparam i114_3_lut_4_lut.LUT_INIT = 16'h00e0;
    SB_LUT4 i1_3_lut_adj_1367 (.I0(n49272), .I1(n50867), .I2(\data_in_frame[17] [5]), 
            .I3(GND_net), .O(n45811));
    defparam i1_3_lut_adj_1367.LUT_INIT = 16'h6969;
    SB_LUT4 i1_3_lut_4_lut_adj_1368 (.I0(tx_transmit_N_3748), .I1(n36465), 
            .I2(n27180), .I3(n27214), .O(n39));   // verilog/coms.v(215[11:56])
    defparam i1_3_lut_4_lut_adj_1368.LUT_INIT = 16'h00e0;
    SB_LUT4 n56634_bdd_4_lut (.I0(n56634), .I1(n53175), .I2(n53174), .I3(byte_transmit_counter[2]), 
            .O(n56637));
    defparam n56634_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1369 (.I0(n28069), .I1(\data_in_frame[6] [3]), 
            .I2(Kp_23__N_1203), .I3(\data_in_frame[8][4] ), .O(n28082));   // verilog/coms.v(75[16:43])
    defparam i1_2_lut_3_lut_4_lut_adj_1369.LUT_INIT = 16'h6996;
    SB_LUT4 i11_4_lut_adj_1370 (.I0(\data_out_frame[19] [3]), .I1(n49429), 
            .I2(n49531), .I3(n49284), .O(n27_adj_4791));   // verilog/coms.v(76[16:43])
    defparam i11_4_lut_adj_1370.LUT_INIT = 16'h6996;
    SB_LUT4 i9_4_lut_adj_1371 (.I0(n46897), .I1(\data_out_frame[18] [4]), 
            .I2(n6_adj_4792), .I3(n49332), .O(n25_adj_4793));   // verilog/coms.v(76[16:43])
    defparam i9_4_lut_adj_1371.LUT_INIT = 16'h9669;
    SB_LUT4 i15_4_lut_adj_1372 (.I0(n25_adj_4793), .I1(n27_adj_4791), .I2(n26_adj_4789), 
            .I3(n28_adj_4788), .O(n49679));   // verilog/coms.v(76[16:43])
    defparam i15_4_lut_adj_1372.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut_adj_1373 (.I0(n46808), .I1(n6_adj_4792), .I2(\data_out_frame[19] [5]), 
            .I3(n27747), .O(n12_adj_4794));
    defparam i5_4_lut_adj_1373.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1374 (.I0(n46894), .I1(n12_adj_4794), .I2(n49679), 
            .I3(n27785), .O(n26777));
    defparam i6_4_lut_adj_1374.LUT_INIT = 16'h9669;
    SB_LUT4 i1_3_lut_adj_1375 (.I0(n45811), .I1(n51346), .I2(\data_in_frame[18] [0]), 
            .I3(GND_net), .O(n51108));
    defparam i1_3_lut_adj_1375.LUT_INIT = 16'h6969;
    SB_LUT4 i2_3_lut_adj_1376 (.I0(n28318), .I1(n49673), .I2(\data_out_frame[17] [4]), 
            .I3(GND_net), .O(n1995));
    defparam i2_3_lut_adj_1376.LUT_INIT = 16'h9696;
    SB_LUT4 equal_330_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8_adj_4708));   // verilog/coms.v(155[7:23])
    defparam equal_330_i8_2_lut_3_lut.LUT_INIT = 16'hefef;
    SB_LUT4 i37410_3_lut (.I0(\data_out_frame[16] [5]), .I1(\data_out_frame[17] [5]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n53240));
    defparam i37410_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i37411_3_lut (.I0(\data_out_frame[18] [5]), .I1(\data_out_frame[19] [5]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n53241));
    defparam i37411_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF data_out_frame_0___i188 (.Q(\data_out_frame[23] [3]), .C(clk16MHz), 
           .D(n29874));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i189 (.Q(\data_out_frame[23] [4]), .C(clk16MHz), 
           .D(n29873));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i190 (.Q(\data_out_frame[23] [5]), .C(clk16MHz), 
           .D(n29872));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i191 (.Q(\data_out_frame[23] [6]), .C(clk16MHz), 
           .D(n29870));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i192 (.Q(\data_out_frame[23] [7]), .C(clk16MHz), 
           .D(n29868));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i193 (.Q(\data_out_frame[24] [0]), .C(clk16MHz), 
           .D(n29867));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i194 (.Q(\data_out_frame[24] [1]), .C(clk16MHz), 
           .D(n29866));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i195 (.Q(\data_out_frame[24] [2]), .C(clk16MHz), 
           .D(n29865));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i196 (.Q(\data_out_frame[24] [3]), .C(clk16MHz), 
           .D(n29864));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i197 (.Q(\data_out_frame[24] [4]), .C(clk16MHz), 
           .D(n29863));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i198 (.Q(\data_out_frame[24] [5]), .C(clk16MHz), 
           .D(n29862));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i199 (.Q(\data_out_frame[24] [6]), .C(clk16MHz), 
           .D(n29861));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i200 (.Q(\data_out_frame[24] [7]), .C(clk16MHz), 
           .D(n29834));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i201 (.Q(\data_out_frame[25] [0]), .C(clk16MHz), 
           .D(n29833));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i202 (.Q(\data_out_frame[25] [1]), .C(clk16MHz), 
           .D(n29832));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i203 (.Q(\data_out_frame[25] [2]), .C(clk16MHz), 
           .D(n29831));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i204 (.Q(\data_out_frame[25] [3]), .C(clk16MHz), 
           .D(n29830));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i205 (.Q(\data_out_frame[25] [4]), .C(clk16MHz), 
           .D(n29827));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i206 (.Q(\data_out_frame[25] [5]), .C(clk16MHz), 
           .D(n29826));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i207 (.Q(\data_out_frame[25] [6]), .C(clk16MHz), 
           .D(n29825));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i208 (.Q(\data_out_frame[25] [7]), .C(clk16MHz), 
           .D(n29824));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 equal_331_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8_adj_4697));   // verilog/coms.v(155[7:23])
    defparam equal_331_i8_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_2_lut_3_lut_adj_1377 (.I0(n28020), .I1(n27478), .I2(\data_in_frame[1] [5]), 
            .I3(GND_net), .O(n49038));   // verilog/coms.v(76[16:43])
    defparam i1_2_lut_3_lut_adj_1377.LUT_INIT = 16'h9696;
    SB_LUT4 i37357_3_lut (.I0(\data_out_frame[22] [5]), .I1(\data_out_frame[23] [5]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n53187));
    defparam i37357_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i37356_3_lut (.I0(\data_out_frame[20] [5]), .I1(\data_out_frame[21] [5]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n53186));
    defparam i37356_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3_4_lut_adj_1378 (.I0(n49350), .I1(n49440), .I2(n27569), 
            .I3(n27890), .O(n50375));
    defparam i3_4_lut_adj_1378.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1379 (.I0(n50375), .I1(n27890), .I2(\data_out_frame[22] [7]), 
            .I3(n49168), .O(n10_adj_4795));
    defparam i4_4_lut_adj_1379.LUT_INIT = 16'h9669;
    SB_DFF neopxl_color_i0_i1 (.Q(neopxl_color[1]), .C(clk16MHz), .D(n29787));   // verilog/coms.v(128[12] 303[6])
    SB_DFF neopxl_color_i0_i2 (.Q(neopxl_color[2]), .C(clk16MHz), .D(n29786));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i5_3_lut_adj_1380 (.I0(\data_out_frame[20] [4]), .I1(n10_adj_4795), 
            .I2(n46842), .I3(GND_net), .O(n49528));
    defparam i5_3_lut_adj_1380.LUT_INIT = 16'h6969;
    SB_DFF neopxl_color_i0_i3 (.Q(neopxl_color[3]), .C(clk16MHz), .D(n29781));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i1_2_lut_4_lut_adj_1381 (.I0(n46693), .I1(n49035), .I2(\data_out_frame[16] [4]), 
            .I3(\data_out_frame[21] [0]), .O(n49572));
    defparam i1_2_lut_4_lut_adj_1381.LUT_INIT = 16'h9669;
    SB_DFF neopxl_color_i0_i4 (.Q(neopxl_color[4]), .C(clk16MHz), .D(n29780));   // verilog/coms.v(128[12] 303[6])
    SB_DFF neopxl_color_i0_i5 (.Q(neopxl_color[5]), .C(clk16MHz), .D(n29779));   // verilog/coms.v(128[12] 303[6])
    SB_DFF neopxl_color_i0_i6 (.Q(neopxl_color[6]), .C(clk16MHz), .D(n29778));   // verilog/coms.v(128[12] 303[6])
    SB_DFF neopxl_color_i0_i7 (.Q(neopxl_color[7]), .C(clk16MHz), .D(n29777));   // verilog/coms.v(128[12] 303[6])
    SB_DFF neopxl_color_i0_i8 (.Q(neopxl_color[8]), .C(clk16MHz), .D(n29776));   // verilog/coms.v(128[12] 303[6])
    SB_DFF neopxl_color_i0_i9 (.Q(neopxl_color[9]), .C(clk16MHz), .D(n29775));   // verilog/coms.v(128[12] 303[6])
    SB_DFF neopxl_color_i0_i10 (.Q(neopxl_color[10]), .C(clk16MHz), .D(n29774));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i1_2_lut_4_lut_adj_1382 (.I0(n46693), .I1(n49035), .I2(\data_out_frame[16] [4]), 
            .I3(\data_out_frame[20] [6]), .O(n46913));
    defparam i1_2_lut_4_lut_adj_1382.LUT_INIT = 16'h9669;
    SB_DFF neopxl_color_i0_i11 (.Q(neopxl_color[11]), .C(clk16MHz), .D(n29773));   // verilog/coms.v(128[12] 303[6])
    SB_DFF neopxl_color_i0_i12 (.Q(neopxl_color[12]), .C(clk16MHz), .D(n29772));   // verilog/coms.v(128[12] 303[6])
    SB_DFF neopxl_color_i0_i13 (.Q(neopxl_color[13]), .C(clk16MHz), .D(n29771));   // verilog/coms.v(128[12] 303[6])
    SB_DFF neopxl_color_i0_i14 (.Q(neopxl_color[14]), .C(clk16MHz), .D(n29770));   // verilog/coms.v(128[12] 303[6])
    SB_DFF neopxl_color_i0_i15 (.Q(neopxl_color[15]), .C(clk16MHz), .D(n29769));   // verilog/coms.v(128[12] 303[6])
    SB_DFF neopxl_color_i0_i16 (.Q(neopxl_color[16]), .C(clk16MHz), .D(n29768));   // verilog/coms.v(128[12] 303[6])
    SB_DFF neopxl_color_i0_i17 (.Q(neopxl_color[17]), .C(clk16MHz), .D(n29767));   // verilog/coms.v(128[12] 303[6])
    SB_DFF neopxl_color_i0_i18 (.Q(neopxl_color[18]), .C(clk16MHz), .D(n29766));   // verilog/coms.v(128[12] 303[6])
    SB_DFF neopxl_color_i0_i19 (.Q(neopxl_color[19]), .C(clk16MHz), .D(n29765));   // verilog/coms.v(128[12] 303[6])
    SB_DFF neopxl_color_i0_i20 (.Q(neopxl_color[20]), .C(clk16MHz), .D(n29764));   // verilog/coms.v(128[12] 303[6])
    SB_DFF neopxl_color_i0_i21 (.Q(neopxl_color[21]), .C(clk16MHz), .D(n29763));   // verilog/coms.v(128[12] 303[6])
    SB_DFF neopxl_color_i0_i22 (.Q(neopxl_color[22]), .C(clk16MHz), .D(n29762));   // verilog/coms.v(128[12] 303[6])
    SB_DFF neopxl_color_i0_i23 (.Q(neopxl_color[23]), .C(clk16MHz), .D(n29761));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i2 (.Q(\data_in_frame[0] [1]), .C(clk16MHz), 
           .D(n29760));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i3 (.Q(\data_in_frame[0] [2]), .C(clk16MHz), 
           .D(n29757));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i4 (.Q(\data_in_frame[0] [3]), .C(clk16MHz), 
           .D(n29756));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i5 (.Q(\data_in_frame[0] [4]), .C(clk16MHz), 
           .D(n29755));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i6 (.Q(\data_in_frame[0] [5]), .C(clk16MHz), 
           .D(n29754));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i7 (.Q(\data_in_frame[0] [6]), .C(clk16MHz), 
           .D(n29753));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i8 (.Q(\data_in_frame[0] [7]), .C(clk16MHz), 
           .D(n29752));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i9 (.Q(\data_in_frame[1] [0]), .C(clk16MHz), 
           .D(n29751));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i10 (.Q(\data_in_frame[1] [1]), .C(clk16MHz), 
           .D(n29750));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i11 (.Q(\data_in_frame[1] [2]), .C(clk16MHz), 
           .D(n29749));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i12 (.Q(\data_in_frame[1] [3]), .C(clk16MHz), 
           .D(n29748));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i13 (.Q(\data_in_frame[1] [4]), .C(clk16MHz), 
           .D(n29747));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i14 (.Q(\data_in_frame[1] [5]), .C(clk16MHz), 
           .D(n29746));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i15 (.Q(\data_in_frame[1] [6]), .C(clk16MHz), 
           .D(n29745));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i16 (.Q(\data_in_frame[1] [7]), .C(clk16MHz), 
           .D(n29744));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i17 (.Q(\data_in_frame[2] [0]), .C(clk16MHz), 
           .D(n29743));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i18 (.Q(\data_in_frame[2] [1]), .C(clk16MHz), 
           .D(n29742));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i19 (.Q(\data_in_frame[2] [2]), .C(clk16MHz), 
           .D(n29741));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i20 (.Q(\data_in_frame[2] [3]), .C(clk16MHz), 
           .D(n29740));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i21 (.Q(\data_in_frame[2] [4]), .C(clk16MHz), 
           .D(n29739));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i22 (.Q(\data_in_frame[2] [5]), .C(clk16MHz), 
           .D(n29738));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i23 (.Q(\data_in_frame[2] [6]), .C(clk16MHz), 
           .D(n29737));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i24 (.Q(\data_in_frame[2] [7]), .C(clk16MHz), 
           .D(n29736));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i25 (.Q(\data_in_frame[3] [0]), .C(clk16MHz), 
           .D(n29735));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i26 (.Q(\data_in_frame[3] [1]), .C(clk16MHz), 
           .D(n29734));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i27 (.Q(\data_in_frame[3] [2]), .C(clk16MHz), 
           .D(n29733));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i28 (.Q(\data_in_frame[3] [3]), .C(clk16MHz), 
           .D(n29732));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i29 (.Q(\data_in_frame[3] [4]), .C(clk16MHz), 
           .D(n29731));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i30 (.Q(\data_in_frame[3] [5]), .C(clk16MHz), 
           .D(n29730));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i31 (.Q(\data_in_frame[3] [6]), .C(clk16MHz), 
           .D(n29729));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i32 (.Q(\data_in_frame[3] [7]), .C(clk16MHz), 
           .D(n29728));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i33 (.Q(\data_in_frame[4] [0]), .C(clk16MHz), 
           .D(n29727));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i34 (.Q(\data_in_frame[4] [1]), .C(clk16MHz), 
           .D(n29726));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i35 (.Q(\data_in_frame[4] [2]), .C(clk16MHz), 
           .D(n29725));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i36 (.Q(\data_in_frame[4] [3]), .C(clk16MHz), 
           .D(n29724));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i37 (.Q(\data_in_frame[4] [4]), .C(clk16MHz), 
           .D(n29723));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i38 (.Q(\data_in_frame[4] [5]), .C(clk16MHz), 
           .D(n29722));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i39 (.Q(\data_in_frame[4] [6]), .C(clk16MHz), 
           .D(n29721));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i40 (.Q(\data_in_frame[4] [7]), .C(clk16MHz), 
           .D(n29720));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i41 (.Q(\data_in_frame[5] [0]), .C(clk16MHz), 
           .D(n29719));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i42 (.Q(\data_in_frame[5] [1]), .C(clk16MHz), 
           .D(n29718));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i43 (.Q(\data_in_frame[5] [2]), .C(clk16MHz), 
           .D(n29717));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i44 (.Q(\data_in_frame[5] [3]), .C(clk16MHz), 
           .D(n29716));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i45 (.Q(\data_in_frame[5] [4]), .C(clk16MHz), 
           .D(n29715));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i46 (.Q(\data_in_frame[5] [5]), .C(clk16MHz), 
           .D(n29714));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i47 (.Q(\data_in_frame[5] [6]), .C(clk16MHz), 
           .D(n29713));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i1_2_lut_3_lut_adj_1383 (.I0(\data_out_frame[19] [5]), .I1(n26777), 
            .I2(n49537), .I3(GND_net), .O(n27890));   // verilog/coms.v(77[16:43])
    defparam i1_2_lut_3_lut_adj_1383.LUT_INIT = 16'h9696;
    SB_LUT4 i4_2_lut_3_lut (.I0(\data_out_frame[19] [5]), .I1(n26777), .I2(n49566), 
            .I3(GND_net), .O(n26_adj_4753));   // verilog/coms.v(77[16:43])
    defparam i4_2_lut_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1384 (.I0(n28020), .I1(n27478), .I2(\data_in_frame[4] [5]), 
            .I3(GND_net), .O(n28268));   // verilog/coms.v(76[16:43])
    defparam i1_2_lut_3_lut_adj_1384.LUT_INIT = 16'h9696;
    SB_DFF data_in_frame_0__i48 (.Q(\data_in_frame[5] [7]), .C(clk16MHz), 
           .D(n29712));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i49 (.Q(\data_in_frame[6] [0]), .C(clk16MHz), 
           .D(n29711));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i50 (.Q(\data_in_frame[6] [1]), .C(clk16MHz), 
           .D(n29710));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i51 (.Q(\data_in_frame[6] [2]), .C(clk16MHz), 
           .D(n29709));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1385 (.I0(\data_in_frame[18] [7]), .I1(\data_in_frame[18] [6]), 
            .I2(\data_in_frame[15] [5]), .I3(\data_in_frame[17] [7]), .O(n52490));
    defparam i1_2_lut_3_lut_4_lut_adj_1385.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0__i52 (.Q(\data_in_frame[6] [3]), .C(clk16MHz), 
           .D(n29708));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i53 (.Q(\data_in_frame[6] [4]), .C(clk16MHz), 
           .D(n29707));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i54 (.Q(\data_in_frame[6] [5]), .C(clk16MHz), 
           .D(n29706));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i55 (.Q(\data_in_frame[6] [6]), .C(clk16MHz), 
           .D(n29705));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i56 (.Q(\data_in_frame[6] [7]), .C(clk16MHz), 
           .D(n29704));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i57 (.Q(\data_in_frame[7] [0]), .C(clk16MHz), 
           .D(n29703));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i58 (.Q(\data_in_frame[7] [1]), .C(clk16MHz), 
           .D(n29702));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i59 (.Q(\data_in_frame[7] [2]), .C(clk16MHz), 
           .D(n29701));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i60 (.Q(\data_in_frame[7] [3]), .C(clk16MHz), 
           .D(n29700));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i61 (.Q(\data_in_frame[7] [4]), .C(clk16MHz), 
           .D(n29699));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i62 (.Q(\data_in_frame[7] [5]), .C(clk16MHz), 
           .D(n29698));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i63 (.Q(\data_in_frame[7] [6]), .C(clk16MHz), 
           .D(n29697));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i64 (.Q(\data_in_frame[7] [7]), .C(clk16MHz), 
           .D(n29695));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i4_4_lut_adj_1386 (.I0(n46808), .I1(\data_out_frame[23] [2]), 
            .I2(n49275), .I3(n6_adj_4796), .O(n50449));
    defparam i4_4_lut_adj_1386.LUT_INIT = 16'h9669;
    SB_DFF data_in_frame_0__i65 (.Q(\data_in_frame[8] [0]), .C(clk16MHz), 
           .D(n29694));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i66 (.Q(\data_in_frame[8]_c [1]), .C(clk16MHz), 
           .D(n29693));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i67 (.Q(\data_in_frame[8][2] ), .C(clk16MHz), 
           .D(n29692));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i68 (.Q(\data_in_frame[8] [3]), .C(clk16MHz), 
           .D(n29691));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i69 (.Q(\data_in_frame[8][4] ), .C(clk16MHz), 
           .D(n29690));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i70 (.Q(\data_in_frame[8][5] ), .C(clk16MHz), 
           .D(n29689));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i71 (.Q(\data_in_frame[8][6] ), .C(clk16MHz), 
           .D(n29688));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i72 (.Q(\data_in_frame[8] [7]), .C(clk16MHz), 
           .D(n29687));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i73 (.Q(\data_in_frame[9] [0]), .C(clk16MHz), 
           .D(n29686));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i74 (.Q(\data_in_frame[9] [1]), .C(clk16MHz), 
           .D(n29685));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i75 (.Q(\data_in_frame[9] [2]), .C(clk16MHz), 
           .D(n29684));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i76 (.Q(\data_in_frame[9] [3]), .C(clk16MHz), 
           .D(n29683));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i77 (.Q(\data_in_frame[9] [4]), .C(clk16MHz), 
           .D(n29682));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i78 (.Q(\data_in_frame[9] [5]), .C(clk16MHz), 
           .D(n29681));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i79 (.Q(\data_in_frame[9] [6]), .C(clk16MHz), 
           .D(n29680));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i80 (.Q(\data_in_frame[9] [7]), .C(clk16MHz), 
           .D(n29679));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i81 (.Q(\data_in_frame[10] [0]), .C(clk16MHz), 
           .D(n29678));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i82 (.Q(\data_in_frame[10][1] ), .C(clk16MHz), 
           .D(n29677));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i83 (.Q(\data_in_frame[10][2] ), .C(clk16MHz), 
           .D(n29676));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i84 (.Q(\data_in_frame[10][3] ), .C(clk16MHz), 
           .D(n29675));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i85 (.Q(\data_in_frame[10][4] ), .C(clk16MHz), 
           .D(n29674));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i86 (.Q(\data_in_frame[10][5] ), .C(clk16MHz), 
           .D(n29673));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i1_2_lut_adj_1387 (.I0(\data_out_frame[25] [3]), .I1(n50449), 
            .I2(GND_net), .I3(GND_net), .O(n49178));
    defparam i1_2_lut_adj_1387.LUT_INIT = 16'h9999;
    SB_DFF data_in_frame_0__i87 (.Q(\data_in_frame[10][6] ), .C(clk16MHz), 
           .D(n29672));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i88 (.Q(\data_in_frame[10][7] ), .C(clk16MHz), 
           .D(n29671));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i89 (.Q(\data_in_frame[11] [0]), .C(clk16MHz), 
           .D(n29670));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i90 (.Q(\data_in_frame[11] [1]), .C(clk16MHz), 
           .D(n29669));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i91 (.Q(\data_in_frame[11] [2]), .C(clk16MHz), 
           .D(n29668));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i92 (.Q(\data_in_frame[11] [3]), .C(clk16MHz), 
           .D(n29667));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i93 (.Q(\data_in_frame[11] [4]), .C(clk16MHz), 
           .D(n29666));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [5]), .I2(\data_out_frame[27] [5]), 
            .I3(byte_transmit_counter[1]), .O(n56976));
    defparam byte_transmit_counter_0__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_DFF data_in_frame_0__i94 (.Q(\data_in_frame[11] [5]), .C(clk16MHz), 
           .D(n29665));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i95 (.Q(\data_in_frame[11] [6]), .C(clk16MHz), 
           .D(n29664));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i96 (.Q(\data_in_frame[11] [7]), .C(clk16MHz), 
           .D(n29663));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i97 (.Q(\data_in_frame[12] [0]), .C(clk16MHz), 
           .D(n29662));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i98 (.Q(\data_in_frame[12] [1]), .C(clk16MHz), 
           .D(n29661));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i99 (.Q(\data_in_frame[12] [2]), .C(clk16MHz), 
           .D(n29660));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i100 (.Q(\data_in_frame[12] [3]), .C(clk16MHz), 
           .D(n29659));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i101 (.Q(\data_in_frame[12] [4]), .C(clk16MHz), 
           .D(n29658));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i102 (.Q(\data_in_frame[12] [5]), .C(clk16MHz), 
           .D(n29657));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i103 (.Q(\data_in_frame[12] [6]), .C(clk16MHz), 
           .D(n29656));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i104 (.Q(\data_in_frame[12] [7]), .C(clk16MHz), 
           .D(n29655));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i105 (.Q(\data_in_frame[13] [0]), .C(clk16MHz), 
           .D(n29654));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i106 (.Q(\data_in_frame[13] [1]), .C(clk16MHz), 
           .D(n29653));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i107 (.Q(\data_in_frame[13] [2]), .C(clk16MHz), 
           .D(n29652));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i108 (.Q(\data_in_frame[13] [3]), .C(clk16MHz), 
           .D(n29651));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i109 (.Q(\data_in_frame[13] [4]), .C(clk16MHz), 
           .D(n29650));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i110 (.Q(\data_in_frame[13] [5]), .C(clk16MHz), 
           .D(n29649));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i111 (.Q(\data_in_frame[13] [6]), .C(clk16MHz), 
           .D(n29648));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i112 (.Q(\data_in_frame[13] [7]), .C(clk16MHz), 
           .D(n29647));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i113 (.Q(\data_in_frame[14] [0]), .C(clk16MHz), 
           .D(n29646));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i37401_3_lut (.I0(\data_out_frame[16] [4]), .I1(\data_out_frame[17] [4]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n53231));
    defparam i37401_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF data_in_frame_0__i114 (.Q(\data_in_frame[14] [1]), .C(clk16MHz), 
           .D(n29645));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i115 (.Q(\data_in_frame[14] [2]), .C(clk16MHz), 
           .D(n29644));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i116 (.Q(\data_in_frame[14] [3]), .C(clk16MHz), 
           .D(n29643));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i37402_3_lut (.I0(\data_out_frame[18] [4]), .I1(\data_out_frame[19] [4]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n53232));
    defparam i37402_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF data_in_frame_0__i117 (.Q(\data_in_frame[14] [4]), .C(clk16MHz), 
           .D(n29642));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i118 (.Q(\data_in_frame[14] [5]), .C(clk16MHz), 
           .D(n29641));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i119 (.Q(\data_in_frame[14] [6]), .C(clk16MHz), 
           .D(n29640));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i120 (.Q(\data_in_frame[14] [7]), .C(clk16MHz), 
           .D(n29639));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i121 (.Q(\data_in_frame[15] [0]), .C(clk16MHz), 
           .D(n29638));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i122 (.Q(\data_in_frame[15] [1]), .C(clk16MHz), 
           .D(n29637));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i123 (.Q(\data_in_frame[15] [2]), .C(clk16MHz), 
           .D(n29636));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i124 (.Q(\data_in_frame[15] [3]), .C(clk16MHz), 
           .D(n29635));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i125 (.Q(\data_in_frame[15] [4]), .C(clk16MHz), 
           .D(n29634));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i126 (.Q(\data_in_frame[15] [5]), .C(clk16MHz), 
           .D(n29633));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i127 (.Q(\data_in_frame[15] [6]), .C(clk16MHz), 
           .D(n29632));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i128 (.Q(\data_in_frame[15] [7]), .C(clk16MHz), 
           .D(n29631));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i129 (.Q(\data_in_frame[16] [0]), .C(clk16MHz), 
           .D(n29630));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i130 (.Q(\data_in_frame[16] [1]), .C(clk16MHz), 
           .D(n29629));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i15511_3_lut_4_lut (.I0(n8_adj_4797), .I1(n48984), .I2(rx_data[7]), 
            .I3(\data_in_frame[20] [7]), .O(n29591));
    defparam i15511_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_frame_0__i131 (.Q(\data_in_frame[16] [2]), .C(clk16MHz), 
           .D(n29628));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i132 (.Q(\data_in_frame[16] [3]), .C(clk16MHz), 
           .D(n29627));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i133 (.Q(\data_in_frame[16] [4]), .C(clk16MHz), 
           .D(n29626));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i134 (.Q(\data_in_frame[16] [5]), .C(clk16MHz), 
           .D(n29625));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i135 (.Q(\data_in_frame[16] [6]), .C(clk16MHz), 
           .D(n29624));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i136 (.Q(\data_in_frame[16] [7]), .C(clk16MHz), 
           .D(n29623));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i137 (.Q(\data_in_frame[17] [0]), .C(clk16MHz), 
           .D(n29622));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i138 (.Q(\data_in_frame[17] [1]), .C(clk16MHz), 
           .D(n29621));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i139 (.Q(\data_in_frame[17] [2]), .C(clk16MHz), 
           .D(n29620));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i140 (.Q(\data_in_frame[17] [3]), .C(clk16MHz), 
           .D(n29619));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i141 (.Q(\data_in_frame[17] [4]), .C(clk16MHz), 
           .D(n29618));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i142 (.Q(\data_in_frame[17] [5]), .C(clk16MHz), 
           .D(n29617));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i143 (.Q(\data_in_frame[17] [6]), .C(clk16MHz), 
           .D(n29616));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i144 (.Q(\data_in_frame[17] [7]), .C(clk16MHz), 
           .D(n29615));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i145 (.Q(\data_in_frame[18] [0]), .C(clk16MHz), 
           .D(n29614));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i146 (.Q(\data_in_frame[18] [1]), .C(clk16MHz), 
           .D(n29613));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i147 (.Q(\data_in_frame[18] [2]), .C(clk16MHz), 
           .D(n29612));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i148 (.Q(\data_in_frame[18] [3]), .C(clk16MHz), 
           .D(n29611));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i149 (.Q(\data_in_frame[18] [4]), .C(clk16MHz), 
           .D(n29610));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i150 (.Q(\data_in_frame[18] [5]), .C(clk16MHz), 
           .D(n29609));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i151 (.Q(\data_in_frame[18] [6]), .C(clk16MHz), 
           .D(n29608));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i152 (.Q(\data_in_frame[18] [7]), .C(clk16MHz), 
           .D(n29607));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i153 (.Q(\data_in_frame[19] [0]), .C(clk16MHz), 
           .D(n29606));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i154 (.Q(\data_in_frame[19] [1]), .C(clk16MHz), 
           .D(n29605));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i155 (.Q(\data_in_frame[19] [2]), .C(clk16MHz), 
           .D(n29604));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i156 (.Q(\data_in_frame[19] [3]), .C(clk16MHz), 
           .D(n29603));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i157 (.Q(\data_in_frame[19] [4]), .C(clk16MHz), 
           .D(n29602));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i158 (.Q(\data_in_frame[19] [5]), .C(clk16MHz), 
           .D(n29601));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i159 (.Q(\data_in_frame[19] [6]), .C(clk16MHz), 
           .D(n29600));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i160 (.Q(\data_in_frame[19] [7]), .C(clk16MHz), 
           .D(n29599));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i161 (.Q(\data_in_frame[20] [0]), .C(clk16MHz), 
           .D(n29598));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i162 (.Q(\data_in_frame[20] [1]), .C(clk16MHz), 
           .D(n29597));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i163 (.Q(\data_in_frame[20] [2]), .C(clk16MHz), 
           .D(n29596));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i164 (.Q(\data_in_frame[20] [3]), .C(clk16MHz), 
           .D(n29595));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i1_2_lut_adj_1388 (.I0(\data_out_frame[20] [7]), .I1(\data_out_frame[20] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n27569));   // verilog/coms.v(79[16:27])
    defparam i1_2_lut_adj_1388.LUT_INIT = 16'h6666;
    SB_DFF data_in_frame_0__i165 (.Q(\data_in_frame[20] [4]), .C(clk16MHz), 
           .D(n29594));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i166 (.Q(\data_in_frame[20] [5]), .C(clk16MHz), 
           .D(n29593));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i167 (.Q(\data_in_frame[20] [6]), .C(clk16MHz), 
           .D(n29592));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i168 (.Q(\data_in_frame[20] [7]), .C(clk16MHz), 
           .D(n29591));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i169 (.Q(\data_in_frame[21] [0]), .C(clk16MHz), 
           .D(n29590));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i170 (.Q(\data_in_frame[21] [1]), .C(clk16MHz), 
           .D(n29589));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i171 (.Q(\data_in_frame[21] [2]), .C(clk16MHz), 
           .D(n29588));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i172 (.Q(\data_in_frame[21] [3]), .C(clk16MHz), 
           .D(n29587));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i173 (.Q(\data_in_frame[21] [4]), .C(clk16MHz), 
           .D(n29586));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i174 (.Q(\data_in_frame[21] [5]), .C(clk16MHz), 
           .D(n29585));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i175 (.Q(\data_in_frame[21] [6]), .C(clk16MHz), 
           .D(n29584));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i176 (.Q(\data_in_frame[21] [7]), .C(clk16MHz), 
           .D(n29583));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i177 (.Q(\data_in_frame[22] [0]), .C(clk16MHz), 
           .D(n29582));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i178 (.Q(\data_in_frame[22] [1]), .C(clk16MHz), 
           .D(n29581));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i179 (.Q(\data_in_frame[22] [2]), .C(clk16MHz), 
           .D(n29580));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i180 (.Q(\data_in_frame[22] [3]), .C(clk16MHz), 
           .D(n29579));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i181 (.Q(\data_in_frame[22] [4]), .C(clk16MHz), 
           .D(n29578));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i182 (.Q(\data_in_frame[22] [5]), .C(clk16MHz), 
           .D(n29577));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i183 (.Q(\data_in_frame[22] [6]), .C(clk16MHz), 
           .D(n29576));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i184 (.Q(\data_in_frame[22] [7]), .C(clk16MHz), 
           .D(n29575));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i185 (.Q(\data_in_frame[23] [0]), .C(clk16MHz), 
           .D(n29574));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i186 (.Q(\data_in_frame[23] [1]), .C(clk16MHz), 
           .D(n29573));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i187 (.Q(\data_in_frame[23] [2]), .C(clk16MHz), 
           .D(n29572));   // verilog/coms.v(128[12] 303[6])
    SB_DFF IntegralLimit_i0_i1 (.Q(IntegralLimit[1]), .C(clk16MHz), .D(n29571));   // verilog/coms.v(128[12] 303[6])
    SB_DFF IntegralLimit_i0_i2 (.Q(IntegralLimit[2]), .C(clk16MHz), .D(n29570));   // verilog/coms.v(128[12] 303[6])
    SB_DFF IntegralLimit_i0_i3 (.Q(IntegralLimit[3]), .C(clk16MHz), .D(n29569));   // verilog/coms.v(128[12] 303[6])
    SB_DFF IntegralLimit_i0_i4 (.Q(IntegralLimit[4]), .C(clk16MHz), .D(n29568));   // verilog/coms.v(128[12] 303[6])
    SB_DFF IntegralLimit_i0_i5 (.Q(IntegralLimit[5]), .C(clk16MHz), .D(n29567));   // verilog/coms.v(128[12] 303[6])
    SB_DFF IntegralLimit_i0_i6 (.Q(IntegralLimit[6]), .C(clk16MHz), .D(n29566));   // verilog/coms.v(128[12] 303[6])
    SB_DFF IntegralLimit_i0_i7 (.Q(IntegralLimit[7]), .C(clk16MHz), .D(n29565));   // verilog/coms.v(128[12] 303[6])
    SB_DFF IntegralLimit_i0_i8 (.Q(IntegralLimit[8]), .C(clk16MHz), .D(n29564));   // verilog/coms.v(128[12] 303[6])
    SB_DFF IntegralLimit_i0_i9 (.Q(IntegralLimit[9]), .C(clk16MHz), .D(n29563));   // verilog/coms.v(128[12] 303[6])
    SB_DFF IntegralLimit_i0_i10 (.Q(IntegralLimit[10]), .C(clk16MHz), .D(n29562));   // verilog/coms.v(128[12] 303[6])
    SB_DFF IntegralLimit_i0_i11 (.Q(IntegralLimit[11]), .C(clk16MHz), .D(n29561));   // verilog/coms.v(128[12] 303[6])
    SB_DFF IntegralLimit_i0_i12 (.Q(IntegralLimit[12]), .C(clk16MHz), .D(n29560));   // verilog/coms.v(128[12] 303[6])
    SB_DFF IntegralLimit_i0_i13 (.Q(IntegralLimit[13]), .C(clk16MHz), .D(n29559));   // verilog/coms.v(128[12] 303[6])
    SB_DFF IntegralLimit_i0_i14 (.Q(IntegralLimit[14]), .C(clk16MHz), .D(n29558));   // verilog/coms.v(128[12] 303[6])
    SB_DFF IntegralLimit_i0_i15 (.Q(IntegralLimit[15]), .C(clk16MHz), .D(n29557));   // verilog/coms.v(128[12] 303[6])
    SB_DFF IntegralLimit_i0_i16 (.Q(IntegralLimit[16]), .C(clk16MHz), .D(n29556));   // verilog/coms.v(128[12] 303[6])
    SB_DFF IntegralLimit_i0_i17 (.Q(IntegralLimit[17]), .C(clk16MHz), .D(n29555));   // verilog/coms.v(128[12] 303[6])
    SB_DFF IntegralLimit_i0_i18 (.Q(IntegralLimit[18]), .C(clk16MHz), .D(n29554));   // verilog/coms.v(128[12] 303[6])
    SB_DFF IntegralLimit_i0_i19 (.Q(IntegralLimit[19]), .C(clk16MHz), .D(n29553));   // verilog/coms.v(128[12] 303[6])
    SB_DFF IntegralLimit_i0_i20 (.Q(IntegralLimit[20]), .C(clk16MHz), .D(n29552));   // verilog/coms.v(128[12] 303[6])
    SB_DFF IntegralLimit_i0_i21 (.Q(IntegralLimit[21]), .C(clk16MHz), .D(n29551));   // verilog/coms.v(128[12] 303[6])
    SB_DFF IntegralLimit_i0_i22 (.Q(IntegralLimit[22]), .C(clk16MHz), .D(n29550));   // verilog/coms.v(128[12] 303[6])
    SB_DFF IntegralLimit_i0_i23 (.Q(IntegralLimit[23]), .C(clk16MHz), .D(n29549));   // verilog/coms.v(128[12] 303[6])
    SB_DFF deadband_i0_i1 (.Q(deadband[1]), .C(clk16MHz), .D(n29546));   // verilog/coms.v(128[12] 303[6])
    SB_DFF deadband_i0_i2 (.Q(deadband[2]), .C(clk16MHz), .D(n29545));   // verilog/coms.v(128[12] 303[6])
    SB_DFF deadband_i0_i3 (.Q(deadband[3]), .C(clk16MHz), .D(n29544));   // verilog/coms.v(128[12] 303[6])
    SB_DFF deadband_i0_i4 (.Q(deadband[4]), .C(clk16MHz), .D(n29543));   // verilog/coms.v(128[12] 303[6])
    SB_DFF deadband_i0_i5 (.Q(deadband[5]), .C(clk16MHz), .D(n29542));   // verilog/coms.v(128[12] 303[6])
    SB_DFF deadband_i0_i6 (.Q(deadband[6]), .C(clk16MHz), .D(n29541));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1389 (.I0(\data_out_frame[20] [5]), .I1(\data_out_frame[20] [1]), 
            .I2(\data_out_frame[20] [3]), .I3(\data_out_frame[20] [2]), 
            .O(n28170));   // verilog/coms.v(79[16:27])
    defparam i1_2_lut_3_lut_4_lut_adj_1389.LUT_INIT = 16'h6996;
    SB_DFF deadband_i0_i7 (.Q(deadband[7]), .C(clk16MHz), .D(n29540));   // verilog/coms.v(128[12] 303[6])
    SB_DFF deadband_i0_i8 (.Q(deadband[8]), .C(clk16MHz), .D(n29539));   // verilog/coms.v(128[12] 303[6])
    SB_DFF deadband_i0_i9 (.Q(deadband[9]), .C(clk16MHz), .D(n29538));   // verilog/coms.v(128[12] 303[6])
    SB_DFF deadband_i0_i10 (.Q(deadband[10]), .C(clk16MHz), .D(n29537));   // verilog/coms.v(128[12] 303[6])
    SB_DFF deadband_i0_i11 (.Q(deadband[11]), .C(clk16MHz), .D(n29536));   // verilog/coms.v(128[12] 303[6])
    SB_DFF deadband_i0_i12 (.Q(deadband[12]), .C(clk16MHz), .D(n29534));   // verilog/coms.v(128[12] 303[6])
    SB_DFF deadband_i0_i13 (.Q(deadband[13]), .C(clk16MHz), .D(n29533));   // verilog/coms.v(128[12] 303[6])
    SB_DFF deadband_i0_i14 (.Q(deadband[14]), .C(clk16MHz), .D(n29532));   // verilog/coms.v(128[12] 303[6])
    SB_DFF deadband_i0_i15 (.Q(deadband[15]), .C(clk16MHz), .D(n29531));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 n56976_bdd_4_lut (.I0(n56976), .I1(\data_out_frame[25] [5]), 
            .I2(\data_out_frame[24] [5]), .I3(byte_transmit_counter[1]), 
            .O(n56979));
    defparam n56976_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF deadband_i0_i16 (.Q(deadband[16]), .C(clk16MHz), .D(n29530));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i1_2_lut_adj_1390 (.I0(\data_out_frame[23] [2]), .I1(\data_out_frame[23] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n49304));
    defparam i1_2_lut_adj_1390.LUT_INIT = 16'h6666;
    SB_DFF deadband_i0_i17 (.Q(deadband[17]), .C(clk16MHz), .D(n29529));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i2_3_lut_4_lut_adj_1391 (.I0(\data_out_frame[23] [2]), .I1(\data_out_frame[23] [3]), 
            .I2(n49572), .I3(n27701), .O(n50641));
    defparam i2_3_lut_4_lut_adj_1391.LUT_INIT = 16'h6996;
    SB_DFF deadband_i0_i18 (.Q(deadband[18]), .C(clk16MHz), .D(n29527));   // verilog/coms.v(128[12] 303[6])
    SB_DFF deadband_i0_i19 (.Q(deadband[19]), .C(clk16MHz), .D(n29526));   // verilog/coms.v(128[12] 303[6])
    SB_DFF deadband_i0_i20 (.Q(deadband[20]), .C(clk16MHz), .D(n29525));   // verilog/coms.v(128[12] 303[6])
    SB_DFF deadband_i0_i21 (.Q(deadband[21]), .C(clk16MHz), .D(n29524));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i1_2_lut_adj_1392 (.I0(\data_out_frame[23] [4]), .I1(n46403), 
            .I2(GND_net), .I3(GND_net), .O(n49451));
    defparam i1_2_lut_adj_1392.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1393 (.I0(\data_out_frame[25] [5]), .I1(\data_out_frame[25] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n49082));
    defparam i1_2_lut_adj_1393.LUT_INIT = 16'h6666;
    SB_LUT4 i2_4_lut_adj_1394 (.I0(n50641), .I1(n49082), .I2(n49255), 
            .I3(n49451), .O(n50744));
    defparam i2_4_lut_adj_1394.LUT_INIT = 16'h9669;
    SB_LUT4 i37404_3_lut (.I0(\data_out_frame[8] [5]), .I1(\data_out_frame[9] [5]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n53234));
    defparam i37404_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i37405_3_lut (.I0(\data_out_frame[10] [5]), .I1(\data_out_frame[11] [5]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n53235));
    defparam i37405_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_adj_1395 (.I0(\data_out_frame[20] [7]), .I1(\data_out_frame[20] [6]), 
            .I2(n46677), .I3(GND_net), .O(n49035));
    defparam i1_2_lut_3_lut_adj_1395.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1396 (.I0(n50641), .I1(\data_out_frame[25] [3]), 
            .I2(n50449), .I3(\data_out_frame[25] [4]), .O(n50545));
    defparam i2_3_lut_4_lut_adj_1396.LUT_INIT = 16'h6996;
    SB_LUT4 i37369_3_lut (.I0(\data_out_frame[14] [5]), .I1(\data_out_frame[15] [5]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n53199));
    defparam i37369_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i37393_3_lut (.I0(\data_out_frame[22] [4]), .I1(\data_out_frame[23] [4]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n53223));
    defparam i37393_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i37368_3_lut (.I0(\data_out_frame[12] [5]), .I1(\data_out_frame[13] [5]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n53198));
    defparam i37368_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i37413_3_lut (.I0(\data_out_frame[8] [6]), .I1(\data_out_frame[9] [6]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n53243));
    defparam i37413_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i37392_3_lut (.I0(\data_out_frame[20] [4]), .I1(\data_out_frame[21] [4]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n53222));
    defparam i37392_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15512_3_lut_4_lut (.I0(n8_adj_4797), .I1(n48984), .I2(rx_data[6]), 
            .I3(\data_in_frame[20] [6]), .O(n29592));
    defparam i15512_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15513_3_lut_4_lut (.I0(n8_adj_4797), .I1(n48984), .I2(rx_data[5]), 
            .I3(\data_in_frame[20] [5]), .O(n29593));
    defparam i15513_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_4_lut_adj_1397 (.I0(\data_out_frame[23] [1]), .I1(\data_out_frame[20] [4]), 
            .I2(n10_adj_4795), .I3(n46842), .O(n6_adj_4796));
    defparam i1_2_lut_4_lut_adj_1397.LUT_INIT = 16'h9669;
    SB_LUT4 i37414_3_lut (.I0(\data_out_frame[10] [6]), .I1(\data_out_frame[11] [6]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n53244));
    defparam i37414_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i37348_3_lut (.I0(\data_out_frame[14] [6]), .I1(\data_out_frame[15] [6]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n53178));
    defparam i37348_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 select_713_Select_23_i3_2_lut (.I0(\FRAME_MATCHER.i [23]), .I1(n4623), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4776));
    defparam select_713_Select_23_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_713_Select_24_i3_2_lut (.I0(\FRAME_MATCHER.i [24]), .I1(n4623), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4775));
    defparam select_713_Select_24_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_3_lut_adj_1398 (.I0(\data_out_frame[20] [1]), .I1(\data_out_frame[20] [3]), 
            .I2(\data_out_frame[20] [2]), .I3(GND_net), .O(n49168));   // verilog/coms.v(79[16:27])
    defparam i1_2_lut_3_lut_adj_1398.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_4_lut_adj_1399 (.I0(\data_out_frame[20] [0]), .I1(n28318), 
            .I2(n49673), .I3(\data_out_frame[17] [4]), .O(n49537));   // verilog/coms.v(77[16:43])
    defparam i1_2_lut_4_lut_adj_1399.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1400 (.I0(\data_in_frame[16] [3]), .I1(n46793), 
            .I2(n45864), .I3(GND_net), .O(n49288));
    defparam i1_2_lut_3_lut_adj_1400.LUT_INIT = 16'h6969;
    SB_LUT4 i37347_3_lut (.I0(\data_out_frame[12] [6]), .I1(\data_out_frame[13] [6]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n53177));
    defparam i37347_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i37431_3_lut (.I0(\data_out_frame[8] [7]), .I1(\data_out_frame[9] [7]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n53261));
    defparam i37431_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i37432_3_lut (.I0(\data_out_frame[10] [7]), .I1(\data_out_frame[11] [7]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n53262));
    defparam i37432_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i37306_3_lut (.I0(\data_out_frame[14] [7]), .I1(\data_out_frame[15] [7]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n53136));
    defparam i37306_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1401 (.I0(tx_transmit_N_3748), .I1(tx_active), 
            .I2(r_SM_Main_2__N_3851[0]), .I3(n27214), .O(n48957));   // verilog/coms.v(215[11:56])
    defparam i1_2_lut_3_lut_4_lut_adj_1401.LUT_INIT = 16'h00fe;
    SB_LUT4 i37305_3_lut (.I0(\data_out_frame[12] [7]), .I1(\data_out_frame[13] [7]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n53135));
    defparam i37305_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1402 (.I0(\FRAME_MATCHER.state[0] ), 
            .I1(\FRAME_MATCHER.state[3] ), .I2(n27307), .I3(\FRAME_MATCHER.state [1]), 
            .O(n27217));   // verilog/coms.v(128[12] 303[6])
    defparam i1_2_lut_3_lut_4_lut_adj_1402.LUT_INIT = 16'hfffd;
    SB_LUT4 i92_2_lut_3_lut_4_lut (.I0(\FRAME_MATCHER.state[0] ), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(n27307), .I3(n4_adj_4688), .O(n75));
    defparam i92_2_lut_3_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_4_lut_adj_1403 (.I0(\data_out_frame[20] [4]), .I1(\data_out_frame[20] [5]), 
            .I2(\data_out_frame[20] [1]), .I3(n27720), .O(n49440));
    defparam i1_2_lut_4_lut_adj_1403.LUT_INIT = 16'h6996;
    SB_LUT4 i15514_3_lut_4_lut (.I0(n8_adj_4797), .I1(n48984), .I2(rx_data[4]), 
            .I3(\data_in_frame[20] [4]), .O(n29594));
    defparam i15514_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_2_lut_4_lut (.I0(n49498), .I1(n10_adj_4798), .I2(\data_out_frame[7] [6]), 
            .I3(\data_out_frame[16] [2]), .O(n6_adj_4783));
    defparam i2_2_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i37359_3_lut (.I0(\data_out_frame[8] [2]), .I1(\data_out_frame[9] [2]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n53189));
    defparam i37359_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i37360_3_lut (.I0(\data_out_frame[10] [2]), .I1(\data_out_frame[11] [2]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n53190));
    defparam i37360_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 select_713_Select_25_i3_2_lut (.I0(\FRAME_MATCHER.i [25]), .I1(n4623), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4774));
    defparam select_713_Select_25_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i37363_3_lut (.I0(\data_out_frame[14] [2]), .I1(\data_out_frame[15] [2]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n53193));
    defparam i37363_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i37362_3_lut (.I0(\data_out_frame[12] [2]), .I1(\data_out_frame[13] [2]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n53192));
    defparam i37362_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i39025_2_lut (.I0(n56961), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n54597));
    defparam i39025_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i15515_3_lut_4_lut (.I0(n8_adj_4797), .I1(n48984), .I2(rx_data[3]), 
            .I3(\data_in_frame[20] [3]), .O(n29595));
    defparam i15515_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1404 (.I0(\data_out_frame[22] [5]), .I1(\data_out_frame[20] [3]), 
            .I2(n46744), .I3(GND_net), .O(n49268));
    defparam i1_2_lut_3_lut_adj_1404.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_4_lut_adj_1405 (.I0(\data_out_frame[24] [6]), .I1(n46033), 
            .I2(n49552), .I3(\data_out_frame[22] [4]), .O(n49454));
    defparam i1_2_lut_4_lut_adj_1405.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1406 (.I0(\data_out_frame[20] [3]), .I1(\data_out_frame[20] [2]), 
            .I2(n46744), .I3(n45884), .O(n46033));
    defparam i2_3_lut_4_lut_adj_1406.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_4_lut_adj_1407 (.I0(\data_out_frame[20] [4]), .I1(n46804), 
            .I2(\data_out_frame[22] [5]), .I3(n46753), .O(n49552));
    defparam i1_2_lut_4_lut_adj_1407.LUT_INIT = 16'h9669;
    SB_LUT4 i5_3_lut_4_lut_adj_1408 (.I0(n28318), .I1(n10_adj_4765), .I2(\data_out_frame[15] [4]), 
            .I3(n49151), .O(n50929));
    defparam i5_3_lut_4_lut_adj_1408.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1409 (.I0(\data_in_frame[16] [4]), .I1(n45864), 
            .I2(\data_in_frame[16] [5]), .I3(n46673), .O(n45512));
    defparam i2_3_lut_4_lut_adj_1409.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1410 (.I0(\data_in_frame[16] [4]), .I1(n45864), 
            .I2(n49328), .I3(GND_net), .O(n49331));
    defparam i1_2_lut_3_lut_adj_1410.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1411 (.I0(\data_in_frame[18] [7]), .I1(\data_in_frame[18] [6]), 
            .I2(n49599), .I3(GND_net), .O(n46682));
    defparam i1_2_lut_3_lut_adj_1411.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_4_lut_adj_1412 (.I0(n46729), .I1(\data_out_frame[25] [0]), 
            .I2(n27715), .I3(n49454), .O(n49456));
    defparam i1_2_lut_4_lut_adj_1412.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1413 (.I0(\data_out_frame[25] [5]), .I1(\data_out_frame[25] [4]), 
            .I2(n49412), .I3(GND_net), .O(n6_adj_4760));
    defparam i1_2_lut_3_lut_adj_1413.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_4_lut_adj_1414 (.I0(n46729), .I1(\data_out_frame[25] [0]), 
            .I2(n27715), .I3(n49566), .O(n49567));
    defparam i1_2_lut_4_lut_adj_1414.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1415 (.I0(\FRAME_MATCHER.state [2]), .I1(\FRAME_MATCHER.state [1]), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_4688));   // verilog/coms.v(264[5:27])
    defparam i1_2_lut_adj_1415.LUT_INIT = 16'hdddd;
    SB_LUT4 i1_3_lut_4_lut_adj_1416 (.I0(\data_in_frame[0] [3]), .I1(\data_in_frame[2] [5]), 
            .I2(\data_in_frame[2] [6]), .I3(\data_in_frame[0] [5]), .O(n49229));   // verilog/coms.v(167[9:87])
    defparam i1_3_lut_4_lut_adj_1416.LUT_INIT = 16'h6996;
    SB_LUT4 i15516_3_lut_4_lut (.I0(n8_adj_4797), .I1(n48984), .I2(rx_data[2]), 
            .I3(\data_in_frame[20] [2]), .O(n29596));
    defparam i15516_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15517_3_lut_4_lut (.I0(n8_adj_4797), .I1(n48984), .I2(rx_data[1]), 
            .I3(\data_in_frame[20] [1]), .O(n29597));
    defparam i15517_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 select_713_Select_11_i3_2_lut (.I0(\FRAME_MATCHER.i [11]), .I1(n4623), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4773));
    defparam select_713_Select_11_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_3_lut_adj_1417 (.I0(\data_in_frame[10][6] ), .I1(n28082), 
            .I2(\data_in_frame[12] [7]), .I3(GND_net), .O(n49335));
    defparam i1_2_lut_3_lut_adj_1417.LUT_INIT = 16'h9696;
    SB_LUT4 i15518_3_lut_4_lut (.I0(n8_adj_4797), .I1(n48984), .I2(rx_data[0]), 
            .I3(\data_in_frame[20] [0]), .O(n29598));
    defparam i15518_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15672_3_lut_4_lut (.I0(n8_adj_4697), .I1(n48970), .I2(rx_data[7]), 
            .I3(\data_in_frame[0] [7]), .O(n29752));
    defparam i15672_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_4_lut_adj_1418 (.I0(\data_in_frame[10][6] ), .I1(n28082), 
            .I2(n27811), .I3(n49342), .O(n45897));
    defparam i2_3_lut_4_lut_adj_1418.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1419 (.I0(\data_out_frame[24] [5]), .I1(\data_out_frame[22] [3]), 
            .I2(n49415), .I3(GND_net), .O(n49566));
    defparam i1_2_lut_3_lut_adj_1419.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1420 (.I0(n46677), .I1(n50375), .I2(n49350), 
            .I3(GND_net), .O(n49631));
    defparam i1_2_lut_3_lut_adj_1420.LUT_INIT = 16'h6969;
    SB_LUT4 select_713_Select_0_i3_2_lut (.I0(\FRAME_MATCHER.i [0]), .I1(n4623), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4625));
    defparam select_713_Select_0_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i5_3_lut_4_lut_adj_1421 (.I0(\data_out_frame[15] [1]), .I1(n26802), 
            .I2(\data_out_frame[21] [5]), .I3(\data_out_frame[17] [1]), 
            .O(n14_adj_4747));   // verilog/coms.v(76[16:43])
    defparam i5_3_lut_4_lut_adj_1421.LUT_INIT = 16'h6996;
    SB_LUT4 i15673_3_lut_4_lut (.I0(n8_adj_4697), .I1(n48970), .I2(rx_data[6]), 
            .I3(\data_in_frame[0] [6]), .O(n29753));
    defparam i15673_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1422 (.I0(\data_in_frame[9] [7]), .I1(\data_in_frame[9] [6]), 
            .I2(n27669), .I3(n27659), .O(n28124));   // verilog/coms.v(86[17:28])
    defparam i1_2_lut_3_lut_4_lut_adj_1422.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1423 (.I0(\data_in_frame[9] [7]), .I1(\data_in_frame[9] [6]), 
            .I2(\data_in_frame[9] [5]), .I3(GND_net), .O(n49652));   // verilog/coms.v(86[17:28])
    defparam i1_2_lut_3_lut_adj_1423.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1424 (.I0(\data_out_frame[22] [0]), .I1(\data_out_frame[15] [3]), 
            .I2(n28496), .I3(GND_net), .O(n6_adj_4745));
    defparam i1_2_lut_3_lut_adj_1424.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1425 (.I0(\FRAME_MATCHER.state[0] ), .I1(n24549), 
            .I2(GND_net), .I3(GND_net), .O(n48979));
    defparam i1_2_lut_adj_1425.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1426 (.I0(n27659), .I1(n27669), .I2(n3_adj_4674), 
            .I3(Kp_23__N_1296), .O(n49324));
    defparam i1_2_lut_3_lut_4_lut_adj_1426.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1427 (.I0(Kp_23__N_1296), .I1(n28079), .I2(\data_in_frame[10][5] ), 
            .I3(n27604), .O(n28272));
    defparam i1_2_lut_4_lut_adj_1427.LUT_INIT = 16'h6996;
    SB_LUT4 i1_rep_85_2_lut (.I0(\data_in_frame[20] [3]), .I1(n49682), .I2(GND_net), 
            .I3(GND_net), .O(n57052));
    defparam i1_rep_85_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_4_lut_adj_1428 (.I0(Kp_23__N_1296), .I1(n28079), .I2(\data_in_frame[10][5] ), 
            .I3(\data_in_frame[16] [7]), .O(n49240));
    defparam i1_2_lut_4_lut_adj_1428.LUT_INIT = 16'h6996;
    SB_LUT4 i15674_3_lut_4_lut (.I0(n8_adj_4697), .I1(n48970), .I2(rx_data[5]), 
            .I3(\data_in_frame[0] [5]), .O(n29754));
    defparam i15674_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_4_lut_adj_1429 (.I0(Kp_23__N_1296), .I1(n28079), .I2(\data_in_frame[10][5] ), 
            .I3(n27692), .O(n28403));
    defparam i1_2_lut_4_lut_adj_1429.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1430 (.I0(\data_in_frame[18] [7]), .I1(\data_in_frame[18] [5]), 
            .I2(n49562), .I3(n49046), .O(Kp_23__N_1895));   // verilog/coms.v(79[16:27])
    defparam i2_3_lut_4_lut_adj_1430.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1431 (.I0(\data_out_frame[19] [0]), .I1(\data_out_frame[19] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n27785));
    defparam i1_2_lut_adj_1431.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1432 (.I0(\data_out_frame[18] [6]), .I1(\data_out_frame[16] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_4792));
    defparam i1_2_lut_adj_1432.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_4_lut_adj_1433 (.I0(\FRAME_MATCHER.state [9]), .I1(n10_adj_4717), 
            .I2(\FRAME_MATCHER.state [15]), .I3(n48), .O(n50_adj_4799));
    defparam i1_2_lut_4_lut_adj_1433.LUT_INIT = 16'hfffe;
    SB_LUT4 i4_4_lut_adj_1434 (.I0(\data_out_frame[11] [5]), .I1(\data_out_frame[7] [1]), 
            .I2(\data_out_frame[9] [3]), .I3(n49107), .O(n10_adj_4790));
    defparam i4_4_lut_adj_1434.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1435 (.I0(\FRAME_MATCHER.state [9]), .I1(n10_adj_4717), 
            .I2(\FRAME_MATCHER.state [15]), .I3(n48864), .O(n4_adj_4718));
    defparam i1_2_lut_4_lut_adj_1435.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_3_lut_4_lut_adj_1436 (.I0(\data_in_frame[11] [4]), .I1(n49478), 
            .I2(n49265), .I3(n27378), .O(n50453));   // verilog/coms.v(76[16:43])
    defparam i2_3_lut_4_lut_adj_1436.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1437 (.I0(n49272), .I1(\data_in_frame[17] [6]), 
            .I2(\data_in_frame[15] [5]), .I3(n46823), .O(n46844));
    defparam i2_3_lut_4_lut_adj_1437.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1438 (.I0(n46699), .I1(\data_in_frame[13] [3]), 
            .I2(\data_in_frame[13] [4]), .I3(n27612), .O(n46823));
    defparam i1_2_lut_4_lut_adj_1438.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_4_lut_adj_1439 (.I0(n49590), .I1(n49376), .I2(\data_in_frame[14] [7]), 
            .I3(n52664), .O(n49097));
    defparam i1_2_lut_4_lut_adj_1439.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1440 (.I0(\data_out_frame[14] [1]), .I1(n49658), 
            .I2(n49409), .I3(n51399), .O(n10_adj_4798));
    defparam i4_4_lut_adj_1440.LUT_INIT = 16'h9669;
    SB_LUT4 i5_3_lut_adj_1441 (.I0(n49498), .I1(n10_adj_4798), .I2(\data_out_frame[7] [6]), 
            .I3(GND_net), .O(n49549));
    defparam i5_3_lut_adj_1441.LUT_INIT = 16'h9696;
    SB_LUT4 i5_4_lut_adj_1442 (.I0(n49132), .I1(n49197), .I2(n46915), 
            .I3(n45836), .O(n12_adj_4800));
    defparam i5_4_lut_adj_1442.LUT_INIT = 16'h9669;
    SB_LUT4 i6_4_lut_adj_1443 (.I0(\data_out_frame[15] [1]), .I1(n12_adj_4800), 
            .I2(n46693), .I3(\data_out_frame[18] [7]), .O(n46370));
    defparam i6_4_lut_adj_1443.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1444 (.I0(\data_out_frame[18] [5]), .I1(n46370), 
            .I2(GND_net), .I3(GND_net), .O(n46894));
    defparam i1_2_lut_adj_1444.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1445 (.I0(n51147), .I1(\data_out_frame[14] [2]), 
            .I2(n27424), .I3(n6_adj_4792), .O(n46693));
    defparam i4_4_lut_adj_1445.LUT_INIT = 16'h9669;
    SB_LUT4 i2_3_lut_adj_1446 (.I0(n50291), .I1(n49549), .I2(\data_out_frame[16] [3]), 
            .I3(GND_net), .O(n46808));
    defparam i2_3_lut_adj_1446.LUT_INIT = 16'h6969;
    SB_LUT4 i15675_3_lut_4_lut (.I0(n8_adj_4697), .I1(n48970), .I2(rx_data[4]), 
            .I3(\data_in_frame[0] [4]), .O(n29755));
    defparam i15675_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i3_4_lut_adj_1447 (.I0(\data_out_frame[19] [0]), .I1(n46693), 
            .I2(n46894), .I3(\data_out_frame[21] [1]), .O(n49275));
    defparam i3_4_lut_adj_1447.LUT_INIT = 16'h9669;
    SB_LUT4 i1_3_lut_4_lut_adj_1448 (.I0(\data_in_frame[8] [7]), .I1(Kp_23__N_1324), 
            .I2(n49404), .I3(n49612), .O(n52632));
    defparam i1_3_lut_4_lut_adj_1448.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1449 (.I0(\data_in_frame[17] [7]), .I1(\data_in_frame[17] [6]), 
            .I2(n49272), .I3(GND_net), .O(n49602));
    defparam i1_2_lut_3_lut_adj_1449.LUT_INIT = 16'h6969;
    SB_LUT4 i1_2_lut_4_lut_adj_1450 (.I0(n49590), .I1(n49376), .I2(\data_in_frame[14] [7]), 
            .I3(n52394), .O(n46666));
    defparam i1_2_lut_4_lut_adj_1450.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1451 (.I0(\data_in_frame[18] [1]), .I1(\data_in_frame[18] [3]), 
            .I2(\data_in_frame[18] [2]), .I3(GND_net), .O(n49562));
    defparam i1_2_lut_3_lut_adj_1451.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1452 (.I0(\data_out_frame[19] [2]), .I1(\data_out_frame[17] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n49531));
    defparam i1_2_lut_adj_1452.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_3_lut_adj_1453 (.I0(n27928), .I1(\data_in_frame[9] [2]), 
            .I2(\data_in_frame[9] [3]), .I3(GND_net), .O(n49265));   // verilog/coms.v(76[16:43])
    defparam i1_2_lut_3_lut_adj_1453.LUT_INIT = 16'h9696;
    SB_LUT4 i4_4_lut_adj_1454 (.I0(n27584), .I1(n49126), .I2(n49649), 
            .I3(n6_adj_4782), .O(n26774));   // verilog/coms.v(86[17:70])
    defparam i4_4_lut_adj_1454.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1455 (.I0(\data_in_frame[18] [1]), .I1(\data_in_frame[18] [3]), 
            .I2(n46413), .I3(GND_net), .O(n46917));
    defparam i1_2_lut_3_lut_adj_1455.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_4_lut_adj_1456 (.I0(Kp_23__N_1098), .I1(\data_in_frame[0] [6]), 
            .I2(\data_in_frame[1] [0]), .I3(\data_in_frame[3] [0]), .O(n28263));   // verilog/coms.v(78[16:27])
    defparam i1_2_lut_4_lut_adj_1456.LUT_INIT = 16'h6996;
    SB_LUT4 i1_3_lut_4_lut_adj_1457 (.I0(\data_in_frame[5] [1]), .I1(\data_in_frame[4] [6]), 
            .I2(\data_in_frame[5] [0]), .I3(\data_in_frame[7] [2]), .O(n49144));   // verilog/coms.v(71[16:27])
    defparam i1_3_lut_4_lut_adj_1457.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1458 (.I0(\data_out_frame[11] [7]), .I1(n49409), 
            .I2(n27535), .I3(n27922), .O(n51399));
    defparam i3_4_lut_adj_1458.LUT_INIT = 16'h6996;
    SB_LUT4 i775_2_lut (.I0(\data_out_frame[11] [7]), .I1(\data_out_frame[11] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n1563));   // verilog/coms.v(72[16:27])
    defparam i775_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1459 (.I0(\data_out_frame[12] [0]), .I1(n49024), 
            .I2(\data_out_frame[5] [4]), .I3(GND_net), .O(n49658));
    defparam i2_3_lut_adj_1459.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1460 (.I0(\data_in_frame[2] [4]), .I1(\data_in_frame[0] [3]), 
            .I2(\data_in_frame[0] [2]), .I3(GND_net), .O(n27478));   // verilog/coms.v(167[9:87])
    defparam i1_2_lut_3_lut_adj_1460.LUT_INIT = 16'h9696;
    SB_LUT4 i2_2_lut_3_lut_adj_1461 (.I0(\data_out_frame[20] [7]), .I1(\data_out_frame[20] [6]), 
            .I2(n28176), .I3(GND_net), .O(n7_adj_4734));
    defparam i2_2_lut_3_lut_adj_1461.LUT_INIT = 16'h9696;
    SB_LUT4 i4_4_lut_adj_1462 (.I0(\data_out_frame[7] [5]), .I1(n1563), 
            .I2(n49502), .I3(n6_adj_4787), .O(n51147));
    defparam i4_4_lut_adj_1462.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1463 (.I0(n49135), .I1(\data_out_frame[9] [4]), 
            .I2(\data_out_frame[7] [3]), .I3(GND_net), .O(n49107));   // verilog/coms.v(74[16:34])
    defparam i2_3_lut_adj_1463.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_1464 (.I0(\data_out_frame[4] [7]), .I1(n49505), 
            .I2(n49114), .I3(\data_out_frame[5] [1]), .O(n27535));   // verilog/coms.v(74[16:34])
    defparam i3_4_lut_adj_1464.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1465 (.I0(\data_out_frame[22] [1]), .I1(n49631), 
            .I2(n26777), .I3(GND_net), .O(n49685));
    defparam i1_2_lut_3_lut_adj_1465.LUT_INIT = 16'h6969;
    SB_LUT4 i1_3_lut_4_lut_adj_1466 (.I0(n28124), .I1(\data_in_frame[10] [0]), 
            .I2(n45762), .I3(\data_in_frame[12] [2]), .O(n49446));
    defparam i1_3_lut_4_lut_adj_1466.LUT_INIT = 16'h9669;
    SB_LUT4 i4_4_lut_adj_1467 (.I0(\data_out_frame[13] [6]), .I1(n49661), 
            .I2(n49147), .I3(\data_out_frame[9] [3]), .O(n10_adj_4801));
    defparam i4_4_lut_adj_1467.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_1468 (.I0(n49511), .I1(n10_adj_4801), .I2(\data_out_frame[9] [2]), 
            .I3(GND_net), .O(n49298));
    defparam i5_3_lut_adj_1468.LUT_INIT = 16'h9696;
    SB_LUT4 i5_3_lut_4_lut_adj_1469 (.I0(\data_out_frame[24] [1]), .I1(\data_out_frame[23] [6]), 
            .I2(n10_adj_4721), .I3(\data_out_frame[21] [7]), .O(n50862));
    defparam i5_3_lut_4_lut_adj_1469.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1470 (.I0(\data_out_frame[14] [0]), .I1(n49502), 
            .I2(n27535), .I3(\data_out_frame[11] [6]), .O(n28573));
    defparam i3_4_lut_adj_1470.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1471 (.I0(n28573), .I1(n49298), .I2(\data_out_frame[13] [7]), 
            .I3(GND_net), .O(n49261));   // verilog/coms.v(86[17:70])
    defparam i2_3_lut_adj_1471.LUT_INIT = 16'h9696;
    SB_LUT4 i15676_3_lut_4_lut (.I0(n8_adj_4697), .I1(n48970), .I2(rx_data[3]), 
            .I3(\data_in_frame[0] [3]), .O(n29756));
    defparam i15676_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1472 (.I0(\data_out_frame[14] [2]), .I1(n51147), 
            .I2(GND_net), .I3(GND_net), .O(n27747));
    defparam i1_2_lut_adj_1472.LUT_INIT = 16'h9999;
    SB_LUT4 i1_3_lut_adj_1473 (.I0(\data_out_frame[6] [6]), .I1(\data_out_frame[4] [5]), 
            .I2(\data_out_frame[4] [4]), .I3(GND_net), .O(n49511));
    defparam i1_3_lut_adj_1473.LUT_INIT = 16'h9696;
    SB_LUT4 i3_3_lut_4_lut_adj_1474 (.I0(\data_in_frame[10][7] ), .I1(Kp_23__N_1305), 
            .I2(\data_in_frame[8][6] ), .I3(\data_in_frame[11] [0]), .O(n49342));
    defparam i3_3_lut_4_lut_adj_1474.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1475 (.I0(\data_out_frame[8] [5]), .I1(\data_out_frame[8] [4]), 
            .I2(\data_out_frame[11] [0]), .I3(\data_out_frame[11] [1]), 
            .O(n49129));
    defparam i1_4_lut_adj_1475.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1476 (.I0(Kp_23__N_1305), .I1(n27928), .I2(n49237), 
            .I3(\data_in_frame[8][6] ), .O(n27811));   // verilog/coms.v(97[12:25])
    defparam i2_3_lut_4_lut_adj_1476.LUT_INIT = 16'h6996;
    SB_LUT4 i2_2_lut_adj_1477 (.I0(n49129), .I1(n27319), .I2(GND_net), 
            .I3(GND_net), .O(n10_adj_4802));
    defparam i2_2_lut_adj_1477.LUT_INIT = 16'h6666;
    SB_LUT4 i1_3_lut_4_lut_adj_1478 (.I0(\data_in_frame[19] [0]), .I1(n50429), 
            .I2(n49482), .I3(n49599), .O(n52362));
    defparam i1_3_lut_4_lut_adj_1478.LUT_INIT = 16'h9669;
    SB_LUT4 i15677_3_lut_4_lut (.I0(n8_adj_4697), .I1(n48970), .I2(rx_data[2]), 
            .I3(\data_in_frame[0] [2]), .O(n29757));
    defparam i15677_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i6_4_lut_adj_1479 (.I0(n49511), .I1(\data_out_frame[10] [6]), 
            .I2(\data_out_frame[8] [6]), .I3(\data_out_frame[9] [0]), .O(n14_adj_4803));
    defparam i6_4_lut_adj_1479.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1480 (.I0(\data_out_frame[13] [2]), .I1(n14_adj_4803), 
            .I2(n10_adj_4802), .I3(\data_out_frame[8] [7]), .O(n28318));
    defparam i7_4_lut_adj_1480.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1481 (.I0(\data_in_frame[19] [0]), .I1(n50429), 
            .I2(n46682), .I3(\data_in_frame[21] [2]), .O(n49307));
    defparam i2_3_lut_4_lut_adj_1481.LUT_INIT = 16'h9669;
    SB_LUT4 i381_2_lut (.I0(n1168), .I1(\data_out_frame[4] [7]), .I2(GND_net), 
            .I3(GND_net), .O(n1169));   // verilog/coms.v(72[16:69])
    defparam i381_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_4_lut_adj_1482 (.I0(\data_in_frame[3] [6]), .I1(\data_in_frame[6] [2]), 
            .I2(\data_in_frame[4] [0]), .I3(\data_in_frame[1] [6]), .O(n6_adj_4719));   // verilog/coms.v(79[16:27])
    defparam i1_2_lut_4_lut_adj_1482.LUT_INIT = 16'h6996;
    SB_LUT4 i1_3_lut_4_lut_adj_1483 (.I0(\data_in_frame[0] [6]), .I1(\data_in_frame[1] [0]), 
            .I2(\data_in_frame[3] [2]), .I3(\data_in_frame[1] [1]), .O(n49258));   // verilog/coms.v(78[16:27])
    defparam i1_3_lut_4_lut_adj_1483.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1484 (.I0(\data_out_frame[8] [7]), .I1(\data_out_frame[8] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_4804));
    defparam i1_2_lut_adj_1484.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_3_lut_adj_1485 (.I0(\data_in_frame[0] [6]), .I1(\data_in_frame[1] [0]), 
            .I2(\data_in_frame[3] [0]), .I3(GND_net), .O(n49522));   // verilog/coms.v(78[16:27])
    defparam i1_2_lut_3_lut_adj_1485.LUT_INIT = 16'h9696;
    SB_LUT4 i15680_3_lut_4_lut (.I0(n8_adj_4697), .I1(n48970), .I2(rx_data[1]), 
            .I3(\data_in_frame[0] [1]), .O(n29760));
    defparam i15680_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i4_4_lut_adj_1486 (.I0(n28296), .I1(n27915), .I2(\data_out_frame[11] [2]), 
            .I3(n6_adj_4804), .O(n49067));
    defparam i4_4_lut_adj_1486.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1487 (.I0(\data_in_frame[3] [4]), .I1(\data_in_frame[3] [5]), 
            .I2(\data_in_frame[5] [6]), .I3(n49094), .O(n52572));
    defparam i1_2_lut_4_lut_adj_1487.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1488 (.I0(\data_in_frame[3] [4]), .I1(\data_in_frame[3] [5]), 
            .I2(\data_in_frame[5] [6]), .I3(\data_in_frame[1] [2]), .O(n49495));
    defparam i1_2_lut_4_lut_adj_1488.LUT_INIT = 16'h6996;
    SB_LUT4 i15293_3_lut_4_lut (.I0(n8_adj_4697), .I1(n48970), .I2(rx_data[0]), 
            .I3(\data_in_frame[0] [0]), .O(n29373));
    defparam i15293_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15664_3_lut_4_lut (.I0(n8_adj_4708), .I1(n48970), .I2(rx_data[7]), 
            .I3(\data_in_frame[1] [7]), .O(n29744));
    defparam i15664_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15665_3_lut_4_lut (.I0(n8_adj_4708), .I1(n48970), .I2(rx_data[6]), 
            .I3(\data_in_frame[1] [6]), .O(n29745));
    defparam i15665_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_4_lut_adj_1489 (.I0(\FRAME_MATCHER.i [4]), .I1(\FRAME_MATCHER.i [5]), 
            .I2(\FRAME_MATCHER.i [3]), .I3(n36451), .O(n48993));   // verilog/coms.v(155[7:23])
    defparam i2_3_lut_4_lut_adj_1489.LUT_INIT = 16'hefff;
    SB_LUT4 i5_4_lut_adj_1490 (.I0(\data_out_frame[10] [5]), .I1(n49472), 
            .I2(\data_out_frame[12] [7]), .I3(n27584), .O(n12_adj_4805));   // verilog/coms.v(77[16:43])
    defparam i5_4_lut_adj_1490.LUT_INIT = 16'h6996;
    SB_LUT4 i15666_3_lut_4_lut (.I0(n8_adj_4708), .I1(n48970), .I2(rx_data[5]), 
            .I3(\data_in_frame[1] [5]), .O(n29746));
    defparam i15666_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_4_lut_adj_1491 (.I0(\data_out_frame[13] [1]), .I1(\data_out_frame[10] [7]), 
            .I2(n12_adj_4805), .I3(n8_adj_4778), .O(n28496));
    defparam i1_4_lut_adj_1491.LUT_INIT = 16'h6996;
    SB_LUT4 i15667_3_lut_4_lut (.I0(n8_adj_4708), .I1(n48970), .I2(rx_data[4]), 
            .I3(\data_in_frame[1] [4]), .O(n29747));
    defparam i15667_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15668_3_lut_4_lut (.I0(n8_adj_4708), .I1(n48970), .I2(rx_data[3]), 
            .I3(\data_in_frame[1] [3]), .O(n29748));
    defparam i15668_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1492 (.I0(n49067), .I1(n49649), .I2(GND_net), 
            .I3(GND_net), .O(n6_adj_4806));   // verilog/coms.v(86[17:70])
    defparam i1_2_lut_adj_1492.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1493 (.I0(\data_out_frame[13] [4]), .I1(\data_out_frame[7] [1]), 
            .I2(n49489), .I3(n6_adj_4806), .O(n46172));   // verilog/coms.v(86[17:70])
    defparam i4_4_lut_adj_1493.LUT_INIT = 16'h6996;
    SB_LUT4 i15669_3_lut_4_lut (.I0(n8_adj_4708), .I1(n48970), .I2(rx_data[2]), 
            .I3(\data_in_frame[1] [2]), .O(n29749));
    defparam i15669_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1494 (.I0(\data_out_frame[9] [1]), .I1(\data_out_frame[9] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n49508));   // verilog/coms.v(86[17:70])
    defparam i1_2_lut_adj_1494.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1495 (.I0(\data_out_frame[5] [3]), .I1(\data_out_frame[9] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n49114));   // verilog/coms.v(74[16:34])
    defparam i1_2_lut_adj_1495.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1496 (.I0(n46686), .I1(n49602), .I2(n57052), 
            .I3(\data_in_frame[22] [4]), .O(n50853));
    defparam i3_4_lut_adj_1496.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1497 (.I0(\data_out_frame[9] [0]), .I1(\data_out_frame[9] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n49489));   // verilog/coms.v(86[17:70])
    defparam i1_2_lut_adj_1497.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1498 (.I0(n27323), .I1(n27915), .I2(\data_out_frame[8] [5]), 
            .I3(GND_net), .O(n27906));   // verilog/coms.v(76[16:43])
    defparam i2_3_lut_adj_1498.LUT_INIT = 16'h9696;
    SB_LUT4 i15670_3_lut_4_lut (.I0(n8_adj_4708), .I1(n48970), .I2(rx_data[1]), 
            .I3(\data_in_frame[1] [1]), .O(n29750));
    defparam i15670_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15671_3_lut_4_lut (.I0(n8_adj_4708), .I1(n48970), .I2(rx_data[0]), 
            .I3(\data_in_frame[1] [0]), .O(n29751));
    defparam i15671_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1499 (.I0(\data_out_frame[4] [3]), .I1(\data_out_frame[6] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_4807));   // verilog/coms.v(86[17:28])
    defparam i1_2_lut_adj_1499.LUT_INIT = 16'h6666;
    SB_LUT4 i6_3_lut (.I0(\data_out_frame[7] [2]), .I1(\data_out_frame[5] [0]), 
            .I2(\data_out_frame[4] [6]), .I3(GND_net), .O(n28_adj_4785));   // verilog/coms.v(86[17:70])
    defparam i6_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i37340_4_lut (.I0(\data_out_frame[6] [1]), .I1(byte_transmit_counter[0]), 
            .I2(byte_transmit_counter[2]), .I3(\data_out_frame[7] [1]), 
            .O(n53170));
    defparam i37340_4_lut.LUT_INIT = 16'hec2c;
    SB_LUT4 i37338_3_lut (.I0(\data_out_frame[4] [1]), .I1(\data_out_frame[5] [1]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n53168));
    defparam i37338_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_1500 (.I0(\data_out_frame[7] [3]), .I1(\data_out_frame[7] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n49505));   // verilog/coms.v(74[16:34])
    defparam i1_2_lut_adj_1500.LUT_INIT = 16'h6666;
    SB_LUT4 i2_2_lut_3_lut_adj_1501 (.I0(\data_in_frame[12] [5]), .I1(n27692), 
            .I2(n28138), .I3(GND_net), .O(n27680));
    defparam i2_2_lut_3_lut_adj_1501.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1502 (.I0(\data_out_frame[8] [7]), .I1(\data_out_frame[7] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n49126));   // verilog/coms.v(86[17:70])
    defparam i1_2_lut_adj_1502.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_4_lut_adj_1503 (.I0(\FRAME_MATCHER.i [4]), .I1(\FRAME_MATCHER.i [5]), 
            .I2(\FRAME_MATCHER.i [3]), .I3(n36451), .O(n48970));   // verilog/coms.v(155[7:23])
    defparam i2_3_lut_4_lut_adj_1503.LUT_INIT = 16'hfeff;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_41052 (.I0(byte_transmit_counter[3]), 
            .I1(n56649), .I2(n54603), .I3(byte_transmit_counter[4]), .O(n56934));
    defparam byte_transmit_counter_3__bdd_4_lut_41052.LUT_INIT = 16'he4aa;
    SB_LUT4 i2_3_lut_adj_1504 (.I0(\data_out_frame[5] [5]), .I1(\data_out_frame[5] [3]), 
            .I2(\data_out_frame[5] [4]), .I3(GND_net), .O(n49200));   // verilog/coms.v(72[16:62])
    defparam i2_3_lut_adj_1504.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1505 (.I0(\data_in_frame[22] [6]), .I1(n45834), 
            .I2(GND_net), .I3(GND_net), .O(n45980));
    defparam i1_2_lut_adj_1505.LUT_INIT = 16'h6666;
    SB_LUT4 i15656_3_lut_4_lut (.I0(n8_adj_4739), .I1(n48970), .I2(rx_data[7]), 
            .I3(\data_in_frame[2] [7]), .O(n29736));
    defparam i15656_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15657_3_lut_4_lut (.I0(n8_adj_4739), .I1(n48970), .I2(rx_data[6]), 
            .I3(\data_in_frame[2] [6]), .O(n29737));
    defparam i15657_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 select_713_Select_21_i3_2_lut (.I0(\FRAME_MATCHER.i [21]), .I1(n4623), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4621));
    defparam select_713_Select_21_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_3_lut_4_lut_adj_1506 (.I0(\data_in_frame[13] [7]), .I1(\data_in_frame[13] [6]), 
            .I2(n26844), .I3(\data_in_frame[15] [1]), .O(n45802));
    defparam i1_3_lut_4_lut_adj_1506.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut_adj_1507 (.I0(n27906), .I1(\data_out_frame[10] [7]), 
            .I2(n49067), .I3(\data_out_frame[13] [3]), .O(n12_adj_4808));
    defparam i5_4_lut_adj_1507.LUT_INIT = 16'h6996;
    SB_LUT4 i15658_3_lut_4_lut (.I0(n8_adj_4739), .I1(n48970), .I2(rx_data[5]), 
            .I3(\data_in_frame[2] [5]), .O(n29738));
    defparam i15658_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15659_3_lut_4_lut (.I0(n8_adj_4739), .I1(n48970), .I2(rx_data[4]), 
            .I3(\data_in_frame[2] [4]), .O(n29739));
    defparam i15659_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15681_3_lut_4_lut (.I0(n36483), .I1(n63_adj_4662), .I2(\data_in_frame[4] [7]), 
            .I3(neopxl_color[23]), .O(n29761));
    defparam i15681_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i6_4_lut_adj_1508 (.I0(\data_out_frame[9] [1]), .I1(n12_adj_4808), 
            .I2(n49147), .I3(\data_out_frame[11] [1]), .O(n49151));
    defparam i6_4_lut_adj_1508.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1509 (.I0(\data_out_frame[15] [7]), .I1(\data_out_frame[15] [6]), 
            .I2(\data_out_frame[16] [0]), .I3(GND_net), .O(n28196));   // verilog/coms.v(72[16:27])
    defparam i2_3_lut_adj_1509.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_4_lut_adj_1510 (.I0(\data_in_frame[9] [0]), .I1(\data_in_frame[11] [2]), 
            .I2(\data_in_frame[9] [1]), .I3(n49670), .O(n52530));
    defparam i1_2_lut_4_lut_adj_1510.LUT_INIT = 16'h6996;
    SB_LUT4 i15682_3_lut_4_lut (.I0(n36483), .I1(n63_adj_4662), .I2(\data_in_frame[4] [6]), 
            .I3(neopxl_color[22]), .O(n29762));
    defparam i15682_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1511 (.I0(\FRAME_MATCHER.i_31__N_2845 ), .I1(n27217), 
            .I2(GND_net), .I3(GND_net), .O(n2_adj_4661));
    defparam i1_2_lut_adj_1511.LUT_INIT = 16'h4444;
    SB_LUT4 i15660_3_lut_4_lut (.I0(n8_adj_4739), .I1(n48970), .I2(rx_data[3]), 
            .I3(\data_in_frame[2] [3]), .O(n29740));
    defparam i15660_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15661_3_lut_4_lut (.I0(n8_adj_4739), .I1(n48970), .I2(rx_data[2]), 
            .I3(\data_in_frame[2] [2]), .O(n29741));
    defparam i15661_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15662_3_lut_4_lut (.I0(n8_adj_4739), .I1(n48970), .I2(rx_data[1]), 
            .I3(\data_in_frame[2] [1]), .O(n29742));
    defparam i15662_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15683_3_lut_4_lut (.I0(n36483), .I1(n63_adj_4662), .I2(\data_in_frame[4] [5]), 
            .I3(neopxl_color[21]), .O(n29763));
    defparam i15683_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15663_3_lut_4_lut (.I0(n8_adj_4739), .I1(n48970), .I2(rx_data[0]), 
            .I3(\data_in_frame[2] [0]), .O(n29743));
    defparam i15663_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 equal_345_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8_adj_4739));   // verilog/coms.v(155[7:23])
    defparam equal_345_i8_2_lut_3_lut.LUT_INIT = 16'hfdfd;
    SB_LUT4 i2_3_lut_adj_1512 (.I0(\data_in_frame[23] [4]), .I1(n49307), 
            .I2(n45752), .I3(GND_net), .O(n50716));
    defparam i2_3_lut_adj_1512.LUT_INIT = 16'h9696;
    SB_LUT4 equal_336_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8_adj_4755));   // verilog/coms.v(155[7:23])
    defparam equal_336_i8_2_lut_3_lut.LUT_INIT = 16'hdfdf;
    SB_LUT4 i1_2_lut_adj_1513 (.I0(\data_out_frame[15] [4]), .I1(n49151), 
            .I2(GND_net), .I3(GND_net), .O(n27455));
    defparam i1_2_lut_adj_1513.LUT_INIT = 16'h6666;
    SB_LUT4 i13_4_lut_adj_1514 (.I0(\data_out_frame[8] [1]), .I1(n49472), 
            .I2(\data_out_frame[8] [2]), .I3(n49200), .O(n35));   // verilog/coms.v(86[17:70])
    defparam i13_4_lut_adj_1514.LUT_INIT = 16'h6996;
    SB_LUT4 i12_4_lut_adj_1515 (.I0(n49126), .I1(\data_out_frame[6] [6]), 
            .I2(n49505), .I3(n49469), .O(n34_adj_4809));   // verilog/coms.v(86[17:70])
    defparam i12_4_lut_adj_1515.LUT_INIT = 16'h6996;
    SB_LUT4 i15684_3_lut_4_lut (.I0(n36483), .I1(n63_adj_4662), .I2(\data_in_frame[4] [4]), 
            .I3(neopxl_color[20]), .O(n29764));
    defparam i15684_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i3_4_lut_adj_1516 (.I0(n45752), .I1(n25607), .I2(\data_in_frame[21] [4]), 
            .I3(\data_in_frame[23] [5]), .O(n51236));
    defparam i3_4_lut_adj_1516.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1517 (.I0(\FRAME_MATCHER.state [1]), .I1(\FRAME_MATCHER.state [2]), 
            .I2(GND_net), .I3(GND_net), .O(n27248));   // verilog/coms.v(202[5:24])
    defparam i1_2_lut_adj_1517.LUT_INIT = 16'heeee;
    SB_LUT4 i3_3_lut (.I0(n46917), .I1(n46800), .I2(\data_in_frame[22] [5]), 
            .I3(GND_net), .O(n8_adj_4810));
    defparam i3_3_lut.LUT_INIT = 16'h6969;
    SB_LUT4 i18_4_lut_adj_1518 (.I0(n35), .I1(\data_out_frame[7] [0]), .I2(n28_adj_4785), 
            .I3(\data_out_frame[7] [6]), .O(n40_adj_4811));   // verilog/coms.v(86[17:70])
    defparam i18_4_lut_adj_1518.LUT_INIT = 16'h6996;
    SB_LUT4 i1_3_lut_4_lut_adj_1519 (.I0(\data_in_frame[0] [7]), .I1(\data_in_frame[1] [1]), 
            .I2(\data_in_frame[1] [2]), .I3(\data_in_frame[3] [3]), .O(n28030));   // verilog/coms.v(74[16:34])
    defparam i1_3_lut_4_lut_adj_1519.LUT_INIT = 16'h6996;
    SB_LUT4 i16_4_lut_adj_1520 (.I0(n49223), .I1(\data_out_frame[6] [7]), 
            .I2(n49135), .I3(\data_out_frame[6] [2]), .O(n38_adj_4812));   // verilog/coms.v(86[17:70])
    defparam i16_4_lut_adj_1520.LUT_INIT = 16'h6996;
    SB_LUT4 select_713_Select_22_i3_2_lut (.I0(\FRAME_MATCHER.i [22]), .I1(n4623), 
            .I2(GND_net), .I3(GND_net), .O(n3));
    defparam select_713_Select_22_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i15648_3_lut_4_lut (.I0(n8_adj_4755), .I1(n48970), .I2(rx_data[7]), 
            .I3(\data_in_frame[3] [7]), .O(n29728));
    defparam i15648_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_3_lut_4_lut_adj_1521 (.I0(\FRAME_MATCHER.state[3] ), .I1(n48871), 
            .I2(n49824), .I3(n7828), .O(n27235));
    defparam i1_3_lut_4_lut_adj_1521.LUT_INIT = 16'hecee;
    SB_LUT4 i1_4_lut_adj_1522 (.I0(n51236), .I1(n50716), .I2(n45980), 
            .I3(n50853), .O(n52400));
    defparam i1_4_lut_adj_1522.LUT_INIT = 16'hffef;
    SB_LUT4 i20_4_lut (.I0(n4_adj_4807), .I1(n40_adj_4811), .I2(n34_adj_4809), 
            .I3(\data_out_frame[4] [5]), .O(n42_adj_4813));   // verilog/coms.v(86[17:70])
    defparam i20_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i15_4_lut_adj_1523 (.I0(\data_out_frame[5] [3]), .I1(\data_out_frame[6] [4]), 
            .I2(n49181), .I3(\data_out_frame[4] [4]), .O(n37_adj_4814));   // verilog/coms.v(86[17:70])
    defparam i15_4_lut_adj_1523.LUT_INIT = 16'h6996;
    SB_LUT4 i15649_3_lut_4_lut (.I0(n8_adj_4755), .I1(n48970), .I2(rx_data[6]), 
            .I3(\data_in_frame[3] [6]), .O(n29729));
    defparam i15649_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i4_4_lut_adj_1524 (.I0(n46832), .I1(\data_in_frame[21] [4]), 
            .I2(\data_in_frame[21] [5]), .I3(n49013), .O(n10_adj_4815));
    defparam i4_4_lut_adj_1524.LUT_INIT = 16'h9669;
    SB_LUT4 n56934_bdd_4_lut (.I0(n56934), .I1(n56841), .I2(n7_adj_4781), 
            .I3(byte_transmit_counter[4]), .O(tx_data[6]));
    defparam n56934_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i37333_3_lut (.I0(\data_out_frame[6] [2]), .I1(\data_out_frame[7] [2]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n53163));
    defparam i37333_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i6_4_lut_adj_1525 (.I0(n27906), .I1(\data_out_frame[9] [7]), 
            .I2(n49489), .I3(\data_out_frame[9] [4]), .O(n16_adj_4816));
    defparam i6_4_lut_adj_1525.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut_adj_1526 (.I0(\data_out_frame[7] [5]), .I1(n37_adj_4814), 
            .I2(n42_adj_4813), .I3(n38_adj_4812), .O(n15_adj_4817));
    defparam i5_4_lut_adj_1526.LUT_INIT = 16'h6996;
    SB_LUT4 i15650_3_lut_4_lut (.I0(n8_adj_4755), .I1(n48970), .I2(rx_data[5]), 
            .I3(\data_in_frame[3] [5]), .O(n29730));
    defparam i15650_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15651_3_lut_4_lut (.I0(n8_adj_4755), .I1(n48970), .I2(rx_data[4]), 
            .I3(\data_in_frame[3] [4]), .O(n29731));
    defparam i15651_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i7_4_lut_adj_1527 (.I0(\data_out_frame[9] [6]), .I1(n49114), 
            .I2(n49508), .I3(\data_out_frame[5] [4]), .O(n17_adj_4818));
    defparam i7_4_lut_adj_1527.LUT_INIT = 16'h6996;
    SB_LUT4 i15652_3_lut_4_lut (.I0(n8_adj_4755), .I1(n48970), .I2(rx_data[3]), 
            .I3(\data_in_frame[3] [3]), .O(n29732));
    defparam i15652_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i8_4_lut_adj_1528 (.I0(\data_out_frame[11] [4]), .I1(n17_adj_4818), 
            .I2(n15_adj_4817), .I3(n16_adj_4816), .O(n33));
    defparam i8_4_lut_adj_1528.LUT_INIT = 16'h9669;
    SB_LUT4 i15653_3_lut_4_lut (.I0(n8_adj_4755), .I1(n48970), .I2(rx_data[2]), 
            .I3(\data_in_frame[3] [2]), .O(n29733));
    defparam i15653_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15654_3_lut_4_lut (.I0(n8_adj_4755), .I1(n48970), .I2(rx_data[1]), 
            .I3(\data_in_frame[3] [1]), .O(n29734));
    defparam i15654_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15655_3_lut_4_lut (.I0(n8_adj_4755), .I1(n48970), .I2(rx_data[0]), 
            .I3(\data_in_frame[3] [0]), .O(n29735));
    defparam i15655_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15685_3_lut_4_lut (.I0(n36483), .I1(n63_adj_4662), .I2(\data_in_frame[4] [3]), 
            .I3(neopxl_color[19]), .O(n29765));
    defparam i15685_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_4_lut_adj_1529 (.I0(\data_in_frame[20] [3]), .I1(n52400), 
            .I2(n8_adj_4810), .I3(\data_in_frame[20] [4]), .O(n52402));
    defparam i1_4_lut_adj_1529.LUT_INIT = 16'hdeed;
    SB_LUT4 i15640_3_lut_4_lut (.I0(n8_adj_4797), .I1(n48970), .I2(rx_data[7]), 
            .I3(\data_in_frame[4] [7]), .O(n29720));
    defparam i15640_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15641_3_lut_4_lut (.I0(n8_adj_4797), .I1(n48970), .I2(rx_data[6]), 
            .I3(\data_in_frame[4] [6]), .O(n29721));
    defparam i15641_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16_4_lut_adj_1530 (.I0(n49151), .I1(n46172), .I2(n28496), 
            .I3(n28180), .O(n41_adj_4819));
    defparam i16_4_lut_adj_1530.LUT_INIT = 16'h6996;
    SB_LUT4 i15642_3_lut_4_lut (.I0(n8_adj_4797), .I1(n48970), .I2(rx_data[5]), 
            .I3(\data_in_frame[4] [5]), .O(n29722));
    defparam i15642_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i3_4_lut_adj_1531 (.I0(\data_out_frame[10] [1]), .I1(\data_out_frame[10] [7]), 
            .I2(n27347), .I3(n49191), .O(n51469));   // verilog/coms.v(86[17:63])
    defparam i3_4_lut_adj_1531.LUT_INIT = 16'h6996;
    SB_LUT4 i15643_3_lut_4_lut (.I0(n8_adj_4797), .I1(n48970), .I2(rx_data[4]), 
            .I3(\data_in_frame[4] [4]), .O(n29723));
    defparam i15643_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15644_3_lut_4_lut (.I0(n8_adj_4797), .I1(n48970), .I2(rx_data[3]), 
            .I3(\data_in_frame[4] [3]), .O(n29724));
    defparam i15644_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15645_3_lut_4_lut (.I0(n8_adj_4797), .I1(n48970), .I2(rx_data[2]), 
            .I3(\data_in_frame[4] [2]), .O(n29725));
    defparam i15645_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15646_3_lut_4_lut (.I0(n8_adj_4797), .I1(n48970), .I2(rx_data[1]), 
            .I3(\data_in_frame[4] [1]), .O(n29726));
    defparam i15646_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15647_3_lut_4_lut (.I0(n8_adj_4797), .I1(n48970), .I2(rx_data[0]), 
            .I3(\data_in_frame[4] [0]), .O(n29727));
    defparam i15647_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i18_4_lut_adj_1532 (.I0(n1563), .I1(n51469), .I2(n49514), 
            .I3(\data_out_frame[11] [3]), .O(n43_adj_4820));
    defparam i18_4_lut_adj_1532.LUT_INIT = 16'h6996;
    SB_LUT4 i15_4_lut_adj_1533 (.I0(\data_out_frame[14] [3]), .I1(n49243), 
            .I2(n49546), .I3(\data_out_frame[12] [5]), .O(n40_adj_4821));
    defparam i15_4_lut_adj_1533.LUT_INIT = 16'h6996;
    SB_LUT4 equal_343_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8_adj_4797));   // verilog/coms.v(155[7:23])
    defparam equal_343_i8_2_lut_3_lut.LUT_INIT = 16'hfbfb;
    SB_LUT4 i21_4_lut_adj_1534 (.I0(n41_adj_4819), .I1(n33), .I2(n49129), 
            .I3(\data_out_frame[8] [3]), .O(n46));
    defparam i21_4_lut_adj_1534.LUT_INIT = 16'h6996;
    SB_LUT4 equal_342_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8_adj_4822));   // verilog/coms.v(155[7:23])
    defparam equal_342_i8_2_lut_3_lut.LUT_INIT = 16'hbfbf;
    SB_LUT4 i15632_3_lut_4_lut (.I0(n8_adj_4822), .I1(n48970), .I2(rx_data[7]), 
            .I3(\data_in_frame[5] [7]), .O(n29712));
    defparam i15632_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15686_3_lut_4_lut (.I0(n36483), .I1(n63_adj_4662), .I2(\data_in_frame[4] [2]), 
            .I3(neopxl_color[18]), .O(n29766));
    defparam i15686_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15687_3_lut_4_lut (.I0(n36483), .I1(n63_adj_4662), .I2(\data_in_frame[4] [1]), 
            .I3(neopxl_color[17]), .O(n29767));
    defparam i15687_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14_4_lut_adj_1535 (.I0(\data_out_frame[12] [7]), .I1(n49212), 
            .I2(\data_out_frame[14] [7]), .I3(\data_out_frame[14] [1]), 
            .O(n39_adj_4823));
    defparam i14_4_lut_adj_1535.LUT_INIT = 16'h6996;
    SB_LUT4 i15633_3_lut_4_lut (.I0(n8_adj_4822), .I1(n48970), .I2(rx_data[6]), 
            .I3(\data_in_frame[5] [6]), .O(n29713));
    defparam i15633_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i37334_4_lut (.I0(n53163), .I1(byte_transmit_counter[0]), .I2(byte_transmit_counter[2]), 
            .I3(byte_transmit_counter[1]), .O(n53164));
    defparam i37334_4_lut.LUT_INIT = 16'ha0a3;
    SB_LUT4 i22_4_lut (.I0(n43_adj_4820), .I1(\data_out_frame[11] [2]), 
            .I2(n38_adj_4784), .I3(\data_out_frame[10] [0]), .O(n47));
    defparam i22_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i24_4_lut_adj_1536 (.I0(n47), .I1(n39_adj_4823), .I2(n46), 
            .I3(n40_adj_4821), .O(n51468));
    defparam i24_4_lut_adj_1536.LUT_INIT = 16'h6996;
    SB_LUT4 i3_3_lut_adj_1537 (.I0(n46844), .I1(\data_in_frame[21] [7]), 
            .I2(n49457), .I3(GND_net), .O(n8_adj_4824));
    defparam i3_3_lut_adj_1537.LUT_INIT = 16'h9696;
    SB_LUT4 i15634_3_lut_4_lut (.I0(n8_adj_4822), .I1(n48970), .I2(rx_data[5]), 
            .I3(\data_in_frame[5] [5]), .O(n29714));
    defparam i15634_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_3_lut_4_lut_adj_1538 (.I0(n28037), .I1(\data_in_frame[2] [4]), 
            .I2(n49032), .I3(\data_in_frame[4] [4]), .O(n28017));   // verilog/coms.v(76[16:43])
    defparam i1_3_lut_4_lut_adj_1538.LUT_INIT = 16'h6996;
    SB_LUT4 i37332_3_lut (.I0(\data_out_frame[4] [2]), .I1(\data_out_frame[5] [2]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n53162));
    defparam i37332_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15688_3_lut_4_lut (.I0(n36483), .I1(n63_adj_4662), .I2(\data_in_frame[4] [0]), 
            .I3(neopxl_color[16]), .O(n29768));
    defparam i15688_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15635_3_lut_4_lut (.I0(n8_adj_4822), .I1(n48970), .I2(rx_data[4]), 
            .I3(\data_in_frame[5] [4]), .O(n29715));
    defparam i15635_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15689_3_lut_4_lut (.I0(n36483), .I1(n63_adj_4662), .I2(\data_in_frame[5] [7]), 
            .I3(neopxl_color[15]), .O(n29769));
    defparam i15689_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i23065_2_lut_3_lut_4_lut (.I0(n4599), .I1(n22875), .I2(n14_adj_4762), 
            .I3(\FRAME_MATCHER.state [29]), .O(n37148));
    defparam i23065_2_lut_3_lut_4_lut.LUT_INIT = 16'hf800;
    SB_LUT4 i15690_3_lut_4_lut (.I0(n36483), .I1(n63_adj_4662), .I2(\data_in_frame[5] [6]), 
            .I3(neopxl_color[14]), .O(n29770));
    defparam i15690_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i3_4_lut_adj_1539 (.I0(n46710), .I1(n51468), .I2(n27455), 
            .I3(n28196), .O(n45750));
    defparam i3_4_lut_adj_1539.LUT_INIT = 16'h6996;
    SB_LUT4 i15636_3_lut_4_lut (.I0(n8_adj_4822), .I1(n48970), .I2(rx_data[3]), 
            .I3(\data_in_frame[5] [3]), .O(n29716));
    defparam i15636_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i23064_2_lut_3_lut_4_lut (.I0(n4599), .I1(n22875), .I2(n14_adj_4762), 
            .I3(\FRAME_MATCHER.state [27]), .O(n37146));
    defparam i23064_2_lut_3_lut_4_lut.LUT_INIT = 16'hf800;
    SB_LUT4 i15637_3_lut_4_lut (.I0(n8_adj_4822), .I1(n48970), .I2(rx_data[2]), 
            .I3(\data_in_frame[5] [2]), .O(n29717));
    defparam i15637_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i3_4_lut_adj_1540 (.I0(\data_in_frame[19] [3]), .I1(n49352), 
            .I2(n46816), .I3(\data_in_frame[23] [7]), .O(n50913));
    defparam i3_4_lut_adj_1540.LUT_INIT = 16'h9669;
    SB_LUT4 i15638_3_lut_4_lut (.I0(n8_adj_4822), .I1(n48970), .I2(rx_data[1]), 
            .I3(\data_in_frame[5] [1]), .O(n29718));
    defparam i15638_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15639_3_lut_4_lut (.I0(n8_adj_4822), .I1(n48970), .I2(rx_data[0]), 
            .I3(\data_in_frame[5] [0]), .O(n29719));
    defparam i15639_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15691_3_lut_4_lut (.I0(n36483), .I1(n63_adj_4662), .I2(\data_in_frame[5] [5]), 
            .I3(neopxl_color[13]), .O(n29771));
    defparam i15691_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i5_3_lut_4_lut_adj_1541 (.I0(\data_in_frame[13] [2]), .I1(\data_in_frame[13] [0]), 
            .I2(\data_in_frame[15] [7]), .I3(\data_in_frame[9] [4]), .O(n14_adj_4710));
    defparam i5_3_lut_4_lut_adj_1541.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1542 (.I0(n46852), .I1(n52402), .I2(n10_adj_4815), 
            .I3(\data_in_frame[23] [6]), .O(n52404));
    defparam i1_4_lut_adj_1542.LUT_INIT = 16'hdeed;
    SB_LUT4 i2_3_lut_4_lut_adj_1543 (.I0(Kp_23__N_1296), .I1(n3_adj_4674), 
            .I2(\data_in_frame[10][4] ), .I3(\data_in_frame[8] [3]), .O(n27692));   // verilog/coms.v(75[16:43])
    defparam i2_3_lut_4_lut_adj_1543.LUT_INIT = 16'h6996;
    SB_LUT4 i15624_3_lut_4_lut (.I0(n8_adj_4678), .I1(n48970), .I2(rx_data[7]), 
            .I3(\data_in_frame[6] [7]), .O(n29704));
    defparam i15624_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15625_3_lut_4_lut (.I0(n8_adj_4678), .I1(n48970), .I2(rx_data[6]), 
            .I3(\data_in_frame[6] [6]), .O(n29705));
    defparam i15625_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i23062_2_lut_3_lut_4_lut (.I0(n4599), .I1(n22875), .I2(n14_adj_4762), 
            .I3(\FRAME_MATCHER.state [23]), .O(n37142));
    defparam i23062_2_lut_3_lut_4_lut.LUT_INIT = 16'hf800;
    SB_LUT4 i15692_3_lut_4_lut (.I0(n36483), .I1(n63_adj_4662), .I2(\data_in_frame[5] [4]), 
            .I3(neopxl_color[12]), .O(n29772));
    defparam i15692_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_4_lut_adj_1544 (.I0(\data_in_frame[6] [7]), .I1(\data_in_frame[6] [6]), 
            .I2(\data_in_frame[6] [3]), .I3(\data_in_frame[6] [4]), .O(n49206));   // verilog/coms.v(86[17:28])
    defparam i1_2_lut_4_lut_adj_1544.LUT_INIT = 16'h6996;
    SB_LUT4 i15626_3_lut_4_lut (.I0(n8_adj_4678), .I1(n48970), .I2(rx_data[5]), 
            .I3(\data_in_frame[6] [5]), .O(n29706));
    defparam i15626_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15627_3_lut_4_lut (.I0(n8_adj_4678), .I1(n48970), .I2(rx_data[4]), 
            .I3(\data_in_frame[6] [4]), .O(n29707));
    defparam i15627_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15628_3_lut_4_lut (.I0(n8_adj_4678), .I1(n48970), .I2(rx_data[3]), 
            .I3(\data_in_frame[6] [3]), .O(n29708));
    defparam i15628_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15629_3_lut_4_lut (.I0(n8_adj_4678), .I1(n48970), .I2(rx_data[2]), 
            .I3(\data_in_frame[6] [2]), .O(n29709));
    defparam i15629_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_2_lut_adj_1545 (.I0(\data_in_frame[19] [7]), .I1(\data_in_frame[22] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n7_adj_4825));
    defparam i2_2_lut_adj_1545.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_4_lut_adj_1546 (.I0(n49331), .I1(n49046), .I2(n50279), 
            .I3(\data_in_frame[20] [6]), .O(n49643));
    defparam i2_3_lut_4_lut_adj_1546.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_41047 (.I0(byte_transmit_counter[3]), 
            .I1(n56667), .I2(n54601), .I3(byte_transmit_counter[4]), .O(n56928));
    defparam byte_transmit_counter_3__bdd_4_lut_41047.LUT_INIT = 16'he4aa;
    SB_LUT4 i15630_3_lut_4_lut (.I0(n8_adj_4678), .I1(n48970), .I2(rx_data[1]), 
            .I3(\data_in_frame[6] [1]), .O(n29710));
    defparam i15630_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1547 (.I0(n45750), .I1(n50291), .I2(GND_net), 
            .I3(GND_net), .O(n46915));
    defparam i1_2_lut_adj_1547.LUT_INIT = 16'h9999;
    SB_LUT4 i1_4_lut_adj_1548 (.I0(n46413), .I1(n49370), .I2(\data_in_frame[20] [0]), 
            .I3(\data_in_frame[22] [2]), .O(n52856));
    defparam i1_4_lut_adj_1548.LUT_INIT = 16'h6996;
    SB_LUT4 i15631_3_lut_4_lut (.I0(n8_adj_4678), .I1(n48970), .I2(rx_data[0]), 
            .I3(\data_in_frame[6] [0]), .O(n29711));
    defparam i15631_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1549 (.I0(\data_out_frame[14] [6]), .I1(n1519), 
            .I2(GND_net), .I3(GND_net), .O(n49212));
    defparam i1_2_lut_adj_1549.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1550 (.I0(n49212), .I1(n1516), .I2(\data_out_frame[12] [5]), 
            .I3(\data_out_frame[12] [4]), .O(n28448));   // verilog/coms.v(86[17:63])
    defparam i3_4_lut_adj_1550.LUT_INIT = 16'h6996;
    SB_LUT4 i15694_3_lut_4_lut (.I0(n36483), .I1(n63_adj_4662), .I2(\data_in_frame[5] [2]), 
            .I3(neopxl_color[10]), .O(n29774));
    defparam i15694_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i5_4_lut_adj_1551 (.I0(\data_out_frame[16] [6]), .I1(n49429), 
            .I2(n46915), .I3(n46695), .O(n12_adj_4769));
    defparam i5_4_lut_adj_1551.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1552 (.I0(n28448), .I1(n12_adj_4769), .I2(n49624), 
            .I3(n28346), .O(n46186));
    defparam i6_4_lut_adj_1552.LUT_INIT = 16'h6996;
    SB_LUT4 i1_3_lut_4_lut_adj_1553 (.I0(\data_in_frame[2] [0]), .I1(n28037), 
            .I2(Kp_23__N_1079), .I3(n52588), .O(n52592));
    defparam i1_3_lut_4_lut_adj_1553.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1554 (.I0(\data_out_frame[6] [1]), .I1(\data_out_frame[4] [0]), 
            .I2(\data_out_frame[5] [4]), .I3(GND_net), .O(n49181));   // verilog/coms.v(86[17:70])
    defparam i2_3_lut_adj_1554.LUT_INIT = 16'h9696;
    SB_LUT4 i1_4_lut_adj_1555 (.I0(n7_adj_4825), .I1(n52404), .I2(n50913), 
            .I3(n8_adj_4824), .O(n52408));
    defparam i1_4_lut_adj_1555.LUT_INIT = 16'hdfef;
    SB_LUT4 i15695_3_lut_4_lut (.I0(n36483), .I1(n63_adj_4662), .I2(\data_in_frame[5] [1]), 
            .I3(neopxl_color[9]), .O(n29775));
    defparam i15695_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15615_3_lut_4_lut (.I0(n37171), .I1(n48970), .I2(rx_data[7]), 
            .I3(\data_in_frame[7] [7]), .O(n29695));
    defparam i15615_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i15617_3_lut_4_lut (.I0(n37171), .I1(n48970), .I2(rx_data[6]), 
            .I3(\data_in_frame[7] [6]), .O(n29697));
    defparam i15617_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i15618_3_lut_4_lut (.I0(n37171), .I1(n48970), .I2(rx_data[5]), 
            .I3(\data_in_frame[7] [5]), .O(n29698));
    defparam i15618_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_adj_1556 (.I0(\data_out_frame[10] [2]), .I1(\data_out_frame[10] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n27347));   // verilog/coms.v(86[17:70])
    defparam i1_2_lut_adj_1556.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1557 (.I0(\data_out_frame[14] [5]), .I1(n27339), 
            .I2(GND_net), .I3(GND_net), .O(n49693));   // verilog/coms.v(76[16:43])
    defparam i1_2_lut_adj_1557.LUT_INIT = 16'h6666;
    SB_LUT4 i15619_3_lut_4_lut (.I0(n37171), .I1(n48970), .I2(rx_data[4]), 
            .I3(\data_in_frame[7] [4]), .O(n29699));
    defparam i15619_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i18376_3_lut (.I0(PWMLimit[17]), .I1(\data_in_frame[8]_c [1]), 
            .I2(n50654), .I3(GND_net), .O(n29924));
    defparam i18376_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i4_4_lut_adj_1558 (.I0(n27359), .I1(\data_out_frame[8] [2]), 
            .I2(\data_out_frame[8] [0]), .I3(n6_adj_4770), .O(n1516));   // verilog/coms.v(86[17:70])
    defparam i4_4_lut_adj_1558.LUT_INIT = 16'h6996;
    SB_LUT4 i15620_3_lut_4_lut (.I0(n37171), .I1(n48970), .I2(rx_data[3]), 
            .I3(\data_in_frame[7] [3]), .O(n29700));
    defparam i15620_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_41042 (.I0(byte_transmit_counter[3]), 
            .I1(n56673), .I2(n54599), .I3(byte_transmit_counter[4]), .O(n56922));
    defparam byte_transmit_counter_3__bdd_4_lut_41042.LUT_INIT = 16'he4aa;
    SB_LUT4 i15621_3_lut_4_lut (.I0(n37171), .I1(n48970), .I2(rx_data[2]), 
            .I3(\data_in_frame[7] [2]), .O(n29701));
    defparam i15621_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i15696_3_lut_4_lut (.I0(n36483), .I1(n63_adj_4662), .I2(\data_in_frame[5] [0]), 
            .I3(neopxl_color[8]), .O(n29776));
    defparam i15696_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15697_3_lut_4_lut (.I0(n36483), .I1(n63_adj_4662), .I2(\data_in_frame[6] [7]), 
            .I3(neopxl_color[7]), .O(n29777));
    defparam i15697_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i3_4_lut_adj_1559 (.I0(\data_in_frame[21] [7]), .I1(\data_in_frame[21] [6]), 
            .I2(n46031), .I3(\data_in_frame[22] [0]), .O(n51299));
    defparam i3_4_lut_adj_1559.LUT_INIT = 16'h6996;
    SB_LUT4 i15622_3_lut_4_lut (.I0(n37171), .I1(n48970), .I2(rx_data[1]), 
            .I3(\data_in_frame[7] [1]), .O(n29702));
    defparam i15622_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i15623_3_lut_4_lut (.I0(n37171), .I1(n48970), .I2(rx_data[0]), 
            .I3(\data_in_frame[7] [0]), .O(n29703));
    defparam i15623_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2_3_lut_adj_1560 (.I0(n1516), .I1(n49693), .I2(\data_out_frame[12] [4]), 
            .I3(GND_net), .O(n28180));   // verilog/coms.v(76[16:43])
    defparam i2_3_lut_adj_1560.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1561 (.I0(\data_out_frame[4] [1]), .I1(\data_out_frame[6] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n49057));   // verilog/coms.v(75[16:43])
    defparam i1_2_lut_adj_1561.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1562 (.I0(n49358), .I1(n52856), .I2(n46844), 
            .I3(n46800), .O(n52862));
    defparam i1_4_lut_adj_1562.LUT_INIT = 16'h9669;
    SB_LUT4 i2_3_lut_adj_1563 (.I0(\data_out_frame[6] [3]), .I1(\data_out_frame[4] [2]), 
            .I2(\data_out_frame[4] [1]), .I3(GND_net), .O(n27323));   // verilog/coms.v(76[16:43])
    defparam i2_3_lut_adj_1563.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1564 (.I0(\data_out_frame[5] [7]), .I1(\data_out_frame[4] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n1193));   // verilog/coms.v(86[17:70])
    defparam i1_2_lut_adj_1564.LUT_INIT = 16'h6666;
    SB_LUT4 i15607_3_lut_4_lut (.I0(n8_adj_4697), .I1(n48993), .I2(rx_data[7]), 
            .I3(\data_in_frame[8] [7]), .O(n29687));
    defparam i15607_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15608_3_lut_4_lut (.I0(n8_adj_4697), .I1(n48993), .I2(rx_data[6]), 
            .I3(\data_in_frame[8][6] ), .O(n29688));
    defparam i15608_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1565 (.I0(\data_out_frame[10] [4]), .I1(\data_out_frame[6] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n27959));   // verilog/coms.v(74[16:42])
    defparam i1_2_lut_adj_1565.LUT_INIT = 16'h6666;
    SB_LUT4 i5_3_lut_adj_1566 (.I0(\data_out_frame[8] [2]), .I1(\data_out_frame[12] [6]), 
            .I2(\data_out_frame[14] [7]), .I3(GND_net), .O(n14_adj_4826));   // verilog/coms.v(75[16:43])
    defparam i5_3_lut_adj_1566.LUT_INIT = 16'h9696;
    SB_LUT4 i15698_3_lut_4_lut (.I0(n36483), .I1(n63_adj_4662), .I2(\data_in_frame[6] [6]), 
            .I3(neopxl_color[6]), .O(n29778));
    defparam i15698_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i6_4_lut_adj_1567 (.I0(n49223), .I1(\data_out_frame[10] [5]), 
            .I2(n1193), .I3(n27319), .O(n15_adj_4827));   // verilog/coms.v(75[16:43])
    defparam i6_4_lut_adj_1567.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut_adj_1568 (.I0(n15_adj_4827), .I1(\data_out_frame[8] [4]), 
            .I2(n14_adj_4826), .I3(n27959), .O(n49618));   // verilog/coms.v(75[16:43])
    defparam i8_4_lut_adj_1568.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut_adj_1569 (.I0(\data_out_frame[8] [1]), .I1(n49057), 
            .I2(n27959), .I3(\data_out_frame[8] [3]), .O(n12_adj_4828));   // verilog/coms.v(73[16:27])
    defparam i5_4_lut_adj_1569.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1570 (.I0(\data_out_frame[5] [5]), .I1(n12_adj_4828), 
            .I2(n49101), .I3(\data_out_frame[10] [3]), .O(n1519));   // verilog/coms.v(73[16:27])
    defparam i6_4_lut_adj_1570.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_41082 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [4]), .I2(\data_out_frame[27] [4]), 
            .I3(byte_transmit_counter[1]), .O(n56970));
    defparam byte_transmit_counter_0__bdd_4_lut_41082.LUT_INIT = 16'he4aa;
    SB_LUT4 i15609_3_lut_4_lut (.I0(n8_adj_4697), .I1(n48993), .I2(rx_data[5]), 
            .I3(\data_in_frame[8][5] ), .O(n29689));
    defparam i15609_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i22453_2_lut_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n63_adj_4650), 
            .I2(n63_adj_4644), .I3(n63_adj_6), .O(\FRAME_MATCHER.state_31__N_2879 [1]));
    defparam i22453_2_lut_3_lut_4_lut.LUT_INIT = 16'h80ff;
    SB_LUT4 i15610_3_lut_4_lut (.I0(n8_adj_4697), .I1(n48993), .I2(rx_data[4]), 
            .I3(\data_in_frame[8][4] ), .O(n29690));
    defparam i15610_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15611_3_lut_4_lut (.I0(n8_adj_4697), .I1(n48993), .I2(rx_data[3]), 
            .I3(\data_in_frame[8] [3]), .O(n29691));
    defparam i15611_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_adj_1571 (.I0(n28180), .I1(\data_out_frame[15] [0]), 
            .I2(\data_out_frame[16] [7]), .I3(GND_net), .O(n49132));   // verilog/coms.v(76[16:43])
    defparam i2_3_lut_adj_1571.LUT_INIT = 16'h9696;
    SB_LUT4 i1_4_lut_adj_1572 (.I0(n52862), .I1(n51299), .I2(n46848), 
            .I3(n52408), .O(n52412));
    defparam i1_4_lut_adj_1572.LUT_INIT = 16'hff7b;
    SB_LUT4 i15612_3_lut_4_lut (.I0(n8_adj_4697), .I1(n48993), .I2(rx_data[2]), 
            .I3(\data_in_frame[8][2] ), .O(n29692));
    defparam i15612_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_adj_1573 (.I0(n1519), .I1(n49618), .I2(\data_out_frame[12] [5]), 
            .I3(GND_net), .O(n49091));
    defparam i2_3_lut_adj_1573.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1574 (.I0(\data_out_frame[15] [0]), .I1(\data_out_frame[15] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n28346));   // verilog/coms.v(77[16:43])
    defparam i1_2_lut_adj_1574.LUT_INIT = 16'h6666;
    SB_LUT4 i375_2_lut (.I0(\data_out_frame[5] [7]), .I1(\data_out_frame[5] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n1191));   // verilog/coms.v(72[16:27])
    defparam i375_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i15613_3_lut_4_lut (.I0(n8_adj_4697), .I1(n48993), .I2(rx_data[1]), 
            .I3(\data_in_frame[8]_c [1]), .O(n29693));
    defparam i15613_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15699_3_lut_4_lut (.I0(n36483), .I1(n63_adj_4662), .I2(\data_in_frame[6] [5]), 
            .I3(neopxl_color[5]), .O(n29779));
    defparam i15699_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15614_3_lut_4_lut (.I0(n8_adj_4697), .I1(n48993), .I2(rx_data[0]), 
            .I3(\data_in_frame[8] [0]), .O(n29694));
    defparam i15614_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15700_3_lut_4_lut (.I0(n36483), .I1(n63_adj_4662), .I2(\data_in_frame[6] [4]), 
            .I3(neopxl_color[4]), .O(n29780));
    defparam i15700_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i23061_2_lut_3_lut_4_lut (.I0(n4599), .I1(n22875), .I2(n14_adj_4762), 
            .I3(\FRAME_MATCHER.state [21]), .O(n37140));
    defparam i23061_2_lut_3_lut_4_lut.LUT_INIT = 16'hf800;
    SB_LUT4 i2_3_lut_adj_1575 (.I0(\data_out_frame[4] [3]), .I1(\data_out_frame[4] [2]), 
            .I2(\data_out_frame[6] [4]), .I3(GND_net), .O(n27915));   // verilog/coms.v(76[16:43])
    defparam i2_3_lut_adj_1575.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1576 (.I0(\data_out_frame[10] [6]), .I1(\data_out_frame[10] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n49191));   // verilog/coms.v(86[17:63])
    defparam i1_2_lut_adj_1576.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1577 (.I0(\data_out_frame[8] [3]), .I1(\data_out_frame[8] [4]), 
            .I2(\data_out_frame[8] [5]), .I3(GND_net), .O(n49028));   // verilog/coms.v(77[16:43])
    defparam i2_3_lut_adj_1577.LUT_INIT = 16'h9696;
    SB_LUT4 i5_4_lut_adj_1578 (.I0(n27915), .I1(\data_out_frame[12] [6]), 
            .I2(\data_out_frame[12] [7]), .I3(n49534), .O(n12_adj_4829));   // verilog/coms.v(75[16:27])
    defparam i5_4_lut_adj_1578.LUT_INIT = 16'h6996;
    SB_LUT4 i15701_3_lut_4_lut (.I0(n36483), .I1(n63_adj_4662), .I2(\data_in_frame[6] [3]), 
            .I3(neopxl_color[3]), .O(n29781));
    defparam i15701_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i6_4_lut_adj_1579 (.I0(n49028), .I1(n12_adj_4829), .I2(n49191), 
            .I3(\data_out_frame[8] [2]), .O(n26802));   // verilog/coms.v(75[16:27])
    defparam i6_4_lut_adj_1579.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1580 (.I0(\data_out_frame[7] [7]), .I1(\data_out_frame[8] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n49469));   // verilog/coms.v(75[16:27])
    defparam i1_2_lut_adj_1580.LUT_INIT = 16'h6666;
    SB_LUT4 i15706_3_lut_4_lut (.I0(n36483), .I1(n63_adj_4662), .I2(\data_in_frame[6] [2]), 
            .I3(neopxl_color[2]), .O(n29786));
    defparam i15706_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1581 (.I0(\data_out_frame[6] [0]), .I1(\data_out_frame[7] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n49101));   // verilog/coms.v(73[16:27])
    defparam i1_2_lut_adj_1581.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1582 (.I0(\data_out_frame[5] [3]), .I1(\data_out_frame[9] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n27938));   // verilog/coms.v(76[16:27])
    defparam i1_2_lut_adj_1582.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1583 (.I0(\data_out_frame[7] [5]), .I1(\data_out_frame[7] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n27922));   // verilog/coms.v(75[16:27])
    defparam i1_2_lut_adj_1583.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1584 (.I0(\data_out_frame[9] [6]), .I1(\data_out_frame[5] [2]), 
            .I2(\data_out_frame[7] [4]), .I3(GND_net), .O(n49024));   // verilog/coms.v(75[16:27])
    defparam i2_3_lut_adj_1584.LUT_INIT = 16'h9696;
    SB_LUT4 i15707_3_lut_4_lut (.I0(n36483), .I1(n63_adj_4662), .I2(\data_in_frame[6] [1]), 
            .I3(neopxl_color[1]), .O(n29787));
    defparam i15707_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i5_4_lut_adj_1585 (.I0(\data_out_frame[10] [0]), .I1(n49024), 
            .I2(\data_out_frame[12] [2]), .I3(n27922), .O(n12_adj_4830));   // verilog/coms.v(75[16:27])
    defparam i5_4_lut_adj_1585.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1586 (.I0(n49602), .I1(n49682), .I2(\data_in_frame[18] [1]), 
            .I3(\data_in_frame[22] [3]), .O(n52750));
    defparam i1_4_lut_adj_1586.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1587 (.I0(\data_out_frame[10] [1]), .I1(n12_adj_4830), 
            .I2(n49469), .I3(\data_out_frame[5] [6]), .O(n27335));   // verilog/coms.v(75[16:27])
    defparam i6_4_lut_adj_1587.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1588 (.I0(\data_out_frame[14] [4]), .I1(n27335), 
            .I2(GND_net), .I3(GND_net), .O(n49243));   // verilog/coms.v(86[17:28])
    defparam i1_2_lut_adj_1588.LUT_INIT = 16'h6666;
    SB_LUT4 i23059_2_lut_3_lut_4_lut (.I0(n4599), .I1(n22875), .I2(n14_adj_4762), 
            .I3(\FRAME_MATCHER.state [19]), .O(n37136));
    defparam i23059_2_lut_3_lut_4_lut.LUT_INIT = 16'hf800;
    SB_LUT4 i2_2_lut_adj_1589 (.I0(\data_out_frame[8] [1]), .I1(\data_out_frame[10] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n10_adj_4831));   // verilog/coms.v(76[16:27])
    defparam i2_2_lut_adj_1589.LUT_INIT = 16'h6666;
    SB_LUT4 i6_4_lut_adj_1590 (.I0(n27359), .I1(\data_out_frame[10] [2]), 
            .I2(\data_out_frame[7] [5]), .I3(n27938), .O(n14_adj_4832));   // verilog/coms.v(76[16:27])
    defparam i6_4_lut_adj_1590.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1591 (.I0(n49358), .I1(n49596), .I2(n46800), 
            .I3(n52750), .O(n51304));
    defparam i1_4_lut_adj_1591.LUT_INIT = 16'h9669;
    SB_LUT4 i7_4_lut_adj_1592 (.I0(\data_out_frame[12] [3]), .I1(n14_adj_4832), 
            .I2(n10_adj_4831), .I3(\data_out_frame[5] [7]), .O(n27339));   // verilog/coms.v(76[16:27])
    defparam i7_4_lut_adj_1592.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1593 (.I0(\data_out_frame[16] [7]), .I1(\data_out_frame[16] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n49184));   // verilog/coms.v(86[17:28])
    defparam i1_2_lut_adj_1593.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1594 (.I0(\data_out_frame[13] [0]), .I1(n26802), 
            .I2(GND_net), .I3(GND_net), .O(n45844));
    defparam i1_2_lut_adj_1594.LUT_INIT = 16'h6666;
    SB_LUT4 i15292_3_lut_4_lut (.I0(n36483), .I1(n63_adj_4662), .I2(\data_in_frame[6] [0]), 
            .I3(neopxl_color[0]), .O(n29372));
    defparam i15292_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1595 (.I0(\data_out_frame[17] [2]), .I1(\data_out_frame[19] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n49426));   // verilog/coms.v(76[16:43])
    defparam i1_2_lut_adj_1595.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1596 (.I0(n49426), .I1(n45844), .I2(\data_out_frame[21] [4]), 
            .I3(n49621), .O(n10_adj_4763));
    defparam i4_4_lut_adj_1596.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut_adj_1597 (.I0(n49621), .I1(n46897), .I2(n49091), 
            .I3(n49132), .O(n12_adj_4833));
    defparam i5_4_lut_adj_1597.LUT_INIT = 16'h9669;
    SB_LUT4 i6_4_lut_adj_1598 (.I0(\data_out_frame[19] [1]), .I1(n12_adj_4833), 
            .I2(n49531), .I3(\data_out_frame[21] [3]), .O(n46403));
    defparam i6_4_lut_adj_1598.LUT_INIT = 16'h6996;
    SB_LUT4 n56970_bdd_4_lut (.I0(n56970), .I1(\data_out_frame[25] [4]), 
            .I2(\data_out_frame[24] [4]), .I3(byte_transmit_counter[1]), 
            .O(n56973));
    defparam n56970_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i15693_3_lut_4_lut (.I0(n36483), .I1(n63_adj_4662), .I2(\data_in_frame[5] [3]), 
            .I3(neopxl_color[11]), .O(n29773));
    defparam i15693_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15503_3_lut_4_lut (.I0(n8_adj_4822), .I1(n48984), .I2(rx_data[7]), 
            .I3(\data_in_frame[21] [7]), .O(n29583));
    defparam i15503_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15504_3_lut_4_lut (.I0(n8_adj_4822), .I1(n48984), .I2(rx_data[6]), 
            .I3(\data_in_frame[21] [6]), .O(n29584));
    defparam i15504_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_4_lut_adj_1599 (.I0(n49307), .I1(n52412), .I2(n45939), 
            .I3(\data_in_frame[23] [3]), .O(n52414));
    defparam i1_4_lut_adj_1599.LUT_INIT = 16'hedde;
    SB_LUT4 i1_2_lut_adj_1600 (.I0(n46403), .I1(n46738), .I2(GND_net), 
            .I3(GND_net), .O(n49321));
    defparam i1_2_lut_adj_1600.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1601 (.I0(\data_out_frame[20] [7]), .I1(n49275), 
            .I2(n46808), .I3(GND_net), .O(n28151));
    defparam i2_3_lut_adj_1601.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1602 (.I0(n46186), .I1(n49392), .I2(\data_out_frame[21] [2]), 
            .I3(GND_net), .O(n27701));
    defparam i2_3_lut_adj_1602.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1603 (.I0(n27701), .I1(n49255), .I2(n27715), 
            .I3(GND_net), .O(n45838));
    defparam i2_3_lut_adj_1603.LUT_INIT = 16'h9696;
    SB_LUT4 i15505_3_lut_4_lut (.I0(n8_adj_4822), .I1(n48984), .I2(rx_data[5]), 
            .I3(\data_in_frame[21] [5]), .O(n29585));
    defparam i15505_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1604 (.I0(n45364), .I1(\FRAME_MATCHER.i [31]), 
            .I2(n63_adj_6), .I3(n19836), .O(n24280));   // verilog/coms.v(158[9:60])
    defparam i1_2_lut_3_lut_4_lut_adj_1604.LUT_INIT = 16'hd000;
    SB_LUT4 i2_3_lut_adj_1605 (.I0(n45838), .I1(\data_out_frame[25] [5]), 
            .I2(\data_out_frame[25] [6]), .I3(GND_net), .O(n51166));
    defparam i2_3_lut_adj_1605.LUT_INIT = 16'h9696;
    SB_LUT4 i15599_3_lut_4_lut (.I0(n8_adj_4708), .I1(n48993), .I2(rx_data[7]), 
            .I3(\data_in_frame[9] [7]), .O(n29679));
    defparam i15599_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15600_3_lut_4_lut (.I0(n8_adj_4708), .I1(n48993), .I2(rx_data[6]), 
            .I3(\data_in_frame[9] [6]), .O(n29680));
    defparam i15600_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15601_3_lut_4_lut (.I0(n8_adj_4708), .I1(n48993), .I2(rx_data[5]), 
            .I3(\data_in_frame[9] [5]), .O(n29681));
    defparam i15601_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15602_3_lut_4_lut (.I0(n8_adj_4708), .I1(n48993), .I2(rx_data[4]), 
            .I3(\data_in_frame[9] [4]), .O(n29682));
    defparam i15602_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15603_3_lut_4_lut (.I0(n8_adj_4708), .I1(n48993), .I2(rx_data[3]), 
            .I3(\data_in_frame[9] [3]), .O(n29683));
    defparam i15603_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15604_3_lut_4_lut (.I0(n8_adj_4708), .I1(n48993), .I2(rx_data[2]), 
            .I3(\data_in_frame[9] [2]), .O(n29684));
    defparam i15604_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15605_3_lut_4_lut (.I0(n8_adj_4708), .I1(n48993), .I2(rx_data[1]), 
            .I3(\data_in_frame[9] [1]), .O(n29685));
    defparam i15605_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1606 (.I0(\data_in_frame[14] [5]), .I1(n28138), 
            .I2(n49543), .I3(GND_net), .O(n46749));
    defparam i1_2_lut_3_lut_adj_1606.LUT_INIT = 16'h9696;
    SB_LUT4 i15506_3_lut_4_lut (.I0(n8_adj_4822), .I1(n48984), .I2(rx_data[4]), 
            .I3(\data_in_frame[21] [4]), .O(n29586));
    defparam i15506_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15606_3_lut_4_lut (.I0(n8_adj_4708), .I1(n48993), .I2(rx_data[0]), 
            .I3(\data_in_frame[9] [0]), .O(n29686));
    defparam i15606_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15591_3_lut_4_lut (.I0(n8_adj_4739), .I1(n48993), .I2(rx_data[7]), 
            .I3(\data_in_frame[10][7] ), .O(n29671));
    defparam i15591_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15507_3_lut_4_lut (.I0(n8_adj_4822), .I1(n48984), .I2(rx_data[3]), 
            .I3(\data_in_frame[21] [3]), .O(n29587));
    defparam i15507_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15592_3_lut_4_lut (.I0(n8_adj_4739), .I1(n48993), .I2(rx_data[6]), 
            .I3(\data_in_frame[10][6] ), .O(n29672));
    defparam i15592_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15593_3_lut_4_lut (.I0(n8_adj_4739), .I1(n48993), .I2(rx_data[5]), 
            .I3(\data_in_frame[10][5] ), .O(n29673));
    defparam i15593_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15594_3_lut_4_lut (.I0(n8_adj_4739), .I1(n48993), .I2(rx_data[4]), 
            .I3(\data_in_frame[10][4] ), .O(n29674));
    defparam i15594_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15508_3_lut_4_lut (.I0(n8_adj_4822), .I1(n48984), .I2(rx_data[2]), 
            .I3(\data_in_frame[21] [2]), .O(n29588));
    defparam i15508_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_41077 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [3]), .I2(\data_out_frame[27] [3]), 
            .I3(byte_transmit_counter[1]), .O(n56964));
    defparam byte_transmit_counter_0__bdd_4_lut_41077.LUT_INIT = 16'he4aa;
    SB_LUT4 i15509_3_lut_4_lut (.I0(n8_adj_4822), .I1(n48984), .I2(rx_data[1]), 
            .I3(\data_in_frame[21] [1]), .O(n29589));
    defparam i15509_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 n56964_bdd_4_lut (.I0(n56964), .I1(\data_out_frame[25] [3]), 
            .I2(\data_out_frame[24] [3]), .I3(byte_transmit_counter[1]), 
            .O(n56967));
    defparam n56964_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i15595_3_lut_4_lut (.I0(n8_adj_4739), .I1(n48993), .I2(rx_data[3]), 
            .I3(\data_in_frame[10][3] ), .O(n29675));
    defparam i15595_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15510_3_lut_4_lut (.I0(n8_adj_4822), .I1(n48984), .I2(rx_data[0]), 
            .I3(\data_in_frame[21] [0]), .O(n29590));
    defparam i15510_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15596_3_lut_4_lut (.I0(n8_adj_4739), .I1(n48993), .I2(rx_data[2]), 
            .I3(\data_in_frame[10][2] ), .O(n29676));
    defparam i15596_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15495_3_lut_4_lut (.I0(n8_adj_4678), .I1(n48984), .I2(rx_data[7]), 
            .I3(\data_in_frame[22] [7]), .O(n29575));
    defparam i15495_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15597_3_lut_4_lut (.I0(n8_adj_4739), .I1(n48993), .I2(rx_data[1]), 
            .I3(\data_in_frame[10][1] ), .O(n29677));
    defparam i15597_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15598_3_lut_4_lut (.I0(n8_adj_4739), .I1(n48993), .I2(rx_data[0]), 
            .I3(\data_in_frame[10] [0]), .O(n29678));
    defparam i15598_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i9_3_lut (.I0(n24549), .I1(\data_in_frame[1] [3]), .I2(\data_in_frame[1] [2]), 
            .I3(GND_net), .O(n26_adj_4834));
    defparam i9_3_lut.LUT_INIT = 16'h4040;
    SB_LUT4 i37209_4_lut (.I0(n27478), .I1(\data_in_frame[0] [6]), .I2(\data_in_frame[2] [7]), 
            .I3(\data_in_frame[0] [5]), .O(n52972));
    defparam i37209_4_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 i1_4_lut_4_lut (.I0(\FRAME_MATCHER.state[0] ), .I1(\FRAME_MATCHER.state [1]), 
            .I2(\FRAME_MATCHER.state [2]), .I3(\FRAME_MATCHER.state_31__N_2943 [3]), 
            .O(n52474));   // verilog/coms.v(146[4] 302[11])
    defparam i1_4_lut_4_lut.LUT_INIT = 16'habaf;
    SB_LUT4 i6_4_lut_adj_1607 (.I0(\data_in_frame[0] [7]), .I1(Kp_23__N_1079), 
            .I2(\data_in_frame[1] [1]), .I3(\data_in_frame[2] [1]), .O(n23));
    defparam i6_4_lut_adj_1607.LUT_INIT = 16'h2184;
    SB_LUT4 i5_4_lut_adj_1608 (.I0(\data_in_frame[1] [0]), .I1(Kp_23__N_1079), 
            .I2(n49117), .I3(n49138), .O(n22));
    defparam i5_4_lut_adj_1608.LUT_INIT = 16'h1248;
    SB_LUT4 i37211_4_lut (.I0(n4_adj_4835), .I1(\data_in_frame[2] [0]), 
            .I2(\data_in_frame[0] [0]), .I3(Kp_23__N_1079), .O(n52974));
    defparam i37211_4_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 i15_4_lut_adj_1609 (.I0(n23), .I1(n52970), .I2(n52972), .I3(n26_adj_4834), 
            .O(n32_adj_4836));
    defparam i15_4_lut_adj_1609.LUT_INIT = 16'h0200;
    SB_LUT4 i10_4_lut_adj_1610 (.I0(\data_in_frame[1] [6]), .I1(\data_in_frame[1] [4]), 
            .I2(n28020), .I3(\data_in_frame[1] [5]), .O(n27_adj_4837));
    defparam i10_4_lut_adj_1610.LUT_INIT = 16'h0800;
    SB_LUT4 i16_4_lut_adj_1611 (.I0(n27_adj_4837), .I1(n32_adj_4836), .I2(n52974), 
            .I3(n22), .O(\FRAME_MATCHER.state_31__N_2943 [3]));
    defparam i16_4_lut_adj_1611.LUT_INIT = 16'h0800;
    SB_LUT4 i1_2_lut_adj_1612 (.I0(\FRAME_MATCHER.state[3] ), .I1(n49824), 
            .I2(GND_net), .I3(GND_net), .O(n48882));
    defparam i1_2_lut_adj_1612.LUT_INIT = 16'h2222;
    SB_LUT4 i1_3_lut_adj_1613 (.I0(n49643), .I1(n49699), .I2(\data_in_frame[23] [2]), 
            .I3(GND_net), .O(n52744));
    defparam i1_3_lut_adj_1613.LUT_INIT = 16'h9696;
    SB_LUT4 i37277_2_lut (.I0(\FRAME_MATCHER.state[3] ), .I1(\FRAME_MATCHER.state [2]), 
            .I2(GND_net), .I3(GND_net), .O(n53040));
    defparam i37277_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_1614 (.I0(\FRAME_MATCHER.state [1]), .I1(n48882), 
            .I2(n53040), .I3(\FRAME_MATCHER.state[0] ), .O(n24055));
    defparam i1_4_lut_adj_1614.LUT_INIT = 16'hccce;
    SB_LUT4 i3_4_lut_adj_1615 (.I0(\FRAME_MATCHER.state [1]), .I1(\FRAME_MATCHER.state_31__N_2943 [3]), 
            .I2(n24055), .I3(n48871), .O(n24210));
    defparam i3_4_lut_adj_1615.LUT_INIT = 16'h0080;
    SB_LUT4 i15496_3_lut_4_lut (.I0(n8_adj_4678), .I1(n48984), .I2(rx_data[6]), 
            .I3(\data_in_frame[22] [6]), .O(n29576));
    defparam i15496_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1616 (.I0(n27339), .I1(\data_out_frame[14] [4]), 
            .I2(n27335), .I3(GND_net), .O(n27424));   // verilog/coms.v(86[17:28])
    defparam i1_2_lut_3_lut_adj_1616.LUT_INIT = 16'h9696;
    SB_LUT4 i15497_3_lut_4_lut (.I0(n8_adj_4678), .I1(n48984), .I2(rx_data[5]), 
            .I3(\data_in_frame[22] [5]), .O(n29577));
    defparam i15497_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15498_3_lut_4_lut (.I0(n8_adj_4678), .I1(n48984), .I2(rx_data[4]), 
            .I3(\data_in_frame[22] [4]), .O(n29578));
    defparam i15498_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15499_3_lut_4_lut (.I0(n8_adj_4678), .I1(n48984), .I2(rx_data[3]), 
            .I3(\data_in_frame[22] [3]), .O(n29579));
    defparam i15499_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15500_3_lut_4_lut (.I0(n8_adj_4678), .I1(n48984), .I2(rx_data[2]), 
            .I3(\data_in_frame[22] [2]), .O(n29580));
    defparam i15500_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15583_3_lut_4_lut (.I0(n8_adj_4755), .I1(n48993), .I2(rx_data[7]), 
            .I3(\data_in_frame[11] [7]), .O(n29663));
    defparam i15583_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15584_3_lut_4_lut (.I0(n8_adj_4755), .I1(n48993), .I2(rx_data[6]), 
            .I3(\data_in_frame[11] [6]), .O(n29664));
    defparam i15584_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15585_3_lut_4_lut (.I0(n8_adj_4755), .I1(n48993), .I2(rx_data[5]), 
            .I3(\data_in_frame[11] [5]), .O(n29665));
    defparam i15585_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15586_3_lut_4_lut (.I0(n8_adj_4755), .I1(n48993), .I2(rx_data[4]), 
            .I3(\data_in_frame[11] [4]), .O(n29666));
    defparam i15586_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15587_3_lut_4_lut (.I0(n8_adj_4755), .I1(n48993), .I2(rx_data[3]), 
            .I3(\data_in_frame[11] [3]), .O(n29667));
    defparam i15587_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15588_3_lut_4_lut (.I0(n8_adj_4755), .I1(n48993), .I2(rx_data[2]), 
            .I3(\data_in_frame[11] [2]), .O(n29668));
    defparam i15588_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15501_3_lut_4_lut (.I0(n8_adj_4678), .I1(n48984), .I2(rx_data[1]), 
            .I3(\data_in_frame[22] [1]), .O(n29581));
    defparam i15501_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15589_3_lut_4_lut (.I0(n8_adj_4755), .I1(n48993), .I2(rx_data[1]), 
            .I3(\data_in_frame[11] [1]), .O(n29669));
    defparam i15589_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_4_lut_adj_1617 (.I0(n1945), .I1(n45750), .I2(\data_out_frame[15] [0]), 
            .I3(\data_out_frame[15] [1]), .O(n45836));
    defparam i2_3_lut_4_lut_adj_1617.LUT_INIT = 16'h6996;
    SB_LUT4 i15590_3_lut_4_lut (.I0(n8_adj_4755), .I1(n48993), .I2(rx_data[0]), 
            .I3(\data_in_frame[11] [0]), .O(n29670));
    defparam i15590_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15575_3_lut_4_lut (.I0(n8_adj_4797), .I1(n48993), .I2(rx_data[7]), 
            .I3(\data_in_frame[12] [7]), .O(n29655));
    defparam i15575_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15502_3_lut_4_lut (.I0(n8_adj_4678), .I1(n48984), .I2(rx_data[0]), 
            .I3(\data_in_frame[22] [0]), .O(n29582));
    defparam i15502_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15576_3_lut_4_lut (.I0(n8_adj_4797), .I1(n48993), .I2(rx_data[6]), 
            .I3(\data_in_frame[12] [6]), .O(n29656));
    defparam i15576_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15577_3_lut_4_lut (.I0(n8_adj_4797), .I1(n48993), .I2(rx_data[5]), 
            .I3(\data_in_frame[12] [5]), .O(n29657));
    defparam i15577_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15578_3_lut_4_lut (.I0(n8_adj_4797), .I1(n48993), .I2(rx_data[4]), 
            .I3(\data_in_frame[12] [4]), .O(n29658));
    defparam i15578_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15579_3_lut_4_lut (.I0(n8_adj_4797), .I1(n48993), .I2(rx_data[3]), 
            .I3(\data_in_frame[12] [3]), .O(n29659));
    defparam i15579_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15580_3_lut_4_lut (.I0(n8_adj_4797), .I1(n48993), .I2(rx_data[2]), 
            .I3(\data_in_frame[12] [2]), .O(n29660));
    defparam i15580_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15581_3_lut_4_lut (.I0(n8_adj_4797), .I1(n48993), .I2(rx_data[1]), 
            .I3(\data_in_frame[12] [1]), .O(n29661));
    defparam i15581_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i37487_4_lut (.I0(\data_out_frame[6] [7]), .I1(byte_transmit_counter[0]), 
            .I2(byte_transmit_counter[2]), .I3(\data_out_frame[7] [7]), 
            .O(n53317));
    defparam i37487_4_lut.LUT_INIT = 16'hec2c;
    SB_LUT4 i37485_3_lut (.I0(\data_out_frame[4] [7]), .I1(\data_out_frame[5] [7]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n53315));
    defparam i37485_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15582_3_lut_4_lut (.I0(n8_adj_4797), .I1(n48993), .I2(rx_data[0]), 
            .I3(\data_in_frame[12] [0]), .O(n29662));
    defparam i15582_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i37313_3_lut_4_lut (.I0(byte_transmit_counter[0]), .I1(byte_transmit_counter[1]), 
            .I2(byte_transmit_counter[2]), .I3(n53142), .O(n53143));   // verilog/coms.v(107[34:55])
    defparam i37313_3_lut_4_lut.LUT_INIT = 16'hf202;
    SB_LUT4 i2_3_lut_4_lut_adj_1618 (.I0(\FRAME_MATCHER.state [1]), .I1(\FRAME_MATCHER.state[0] ), 
            .I2(n48871), .I3(\FRAME_MATCHER.state [2]), .O(n7828));
    defparam i2_3_lut_4_lut_adj_1618.LUT_INIT = 16'hfffe;
    SB_LUT4 i34072_2_lut_3_lut (.I0(\FRAME_MATCHER.state [1]), .I1(\FRAME_MATCHER.state[0] ), 
            .I2(\FRAME_MATCHER.state [2]), .I3(GND_net), .O(n49824));
    defparam i34072_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i3_3_lut_4_lut_adj_1619 (.I0(\FRAME_MATCHER.state [2]), .I1(\FRAME_MATCHER.state [1]), 
            .I2(n36465), .I3(\FRAME_MATCHER.state[0] ), .O(n8_adj_4677));
    defparam i3_3_lut_4_lut_adj_1619.LUT_INIT = 16'hf7ff;
    SB_LUT4 i2_3_lut_4_lut_adj_1620 (.I0(n48866), .I1(n48864), .I2(n37153), 
            .I3(n50_adj_4799), .O(n49911));
    defparam i2_3_lut_4_lut_adj_1620.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_3_lut_4_lut_adj_1621 (.I0(n48866), .I1(n48864), .I2(n50_adj_4799), 
            .I3(n37153), .O(n48871));
    defparam i2_3_lut_4_lut_adj_1621.LUT_INIT = 16'hfffe;
    SB_LUT4 i15567_3_lut_4_lut (.I0(n8_adj_4822), .I1(n48993), .I2(rx_data[7]), 
            .I3(\data_in_frame[13] [7]), .O(n29647));
    defparam i15567_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i37478_3_lut_4_lut (.I0(byte_transmit_counter[0]), .I1(byte_transmit_counter[1]), 
            .I2(byte_transmit_counter[2]), .I3(n53307), .O(n53308));   // verilog/coms.v(107[34:55])
    defparam i37478_3_lut_4_lut.LUT_INIT = 16'hf202;
    SB_LUT4 i15568_3_lut_4_lut (.I0(n8_adj_4822), .I1(n48993), .I2(rx_data[6]), 
            .I3(\data_in_frame[13] [6]), .O(n29648));
    defparam i15568_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1622 (.I0(n27339), .I1(\data_out_frame[14] [4]), 
            .I2(n27335), .I3(\data_out_frame[17] [0]), .O(n49624));
    defparam i1_2_lut_3_lut_4_lut_adj_1622.LUT_INIT = 16'h6996;
    SB_LUT4 i1_3_lut_4_lut_adj_1623 (.I0(n3_adj_4674), .I1(\data_in_frame[8]_c [1]), 
            .I2(n25500), .I3(\data_in_frame[10][3] ), .O(n28138));
    defparam i1_3_lut_4_lut_adj_1623.LUT_INIT = 16'h6996;
    SB_LUT4 i15569_3_lut_4_lut (.I0(n8_adj_4822), .I1(n48993), .I2(rx_data[5]), 
            .I3(\data_in_frame[13] [5]), .O(n29649));
    defparam i15569_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15570_3_lut_4_lut (.I0(n8_adj_4822), .I1(n48993), .I2(rx_data[4]), 
            .I3(\data_in_frame[13] [4]), .O(n29650));
    defparam i15570_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1624 (.I0(n110), .I1(n49), .I2(\FRAME_MATCHER.state [4]), 
            .I3(GND_net), .O(n48448));   // verilog/coms.v(116[11:12])
    defparam i1_2_lut_3_lut_adj_1624.LUT_INIT = 16'he0e0;
    SB_LUT4 i15571_3_lut_4_lut (.I0(n8_adj_4822), .I1(n48993), .I2(rx_data[3]), 
            .I3(\data_in_frame[13] [3]), .O(n29651));
    defparam i15571_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15572_3_lut_4_lut (.I0(n8_adj_4822), .I1(n48993), .I2(rx_data[2]), 
            .I3(\data_in_frame[13] [2]), .O(n29652));
    defparam i15572_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15573_3_lut_4_lut (.I0(n8_adj_4822), .I1(n48993), .I2(rx_data[1]), 
            .I3(\data_in_frame[13] [1]), .O(n29653));
    defparam i15573_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15574_3_lut_4_lut (.I0(n8_adj_4822), .I1(n48993), .I2(rx_data[0]), 
            .I3(\data_in_frame[13] [0]), .O(n29654));
    defparam i15574_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i38945_2_lut (.I0(n56967), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n54598));
    defparam i38945_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1_2_lut_3_lut_adj_1625 (.I0(n110), .I1(n49), .I2(\FRAME_MATCHER.state [5]), 
            .I3(GND_net), .O(n48450));   // verilog/coms.v(116[11:12])
    defparam i1_2_lut_3_lut_adj_1625.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1626 (.I0(n110), .I1(n49), .I2(\FRAME_MATCHER.state [6]), 
            .I3(GND_net), .O(n7_adj_4772));   // verilog/coms.v(116[11:12])
    defparam i1_2_lut_3_lut_adj_1626.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1627 (.I0(n110), .I1(n49), .I2(\FRAME_MATCHER.state [7]), 
            .I3(GND_net), .O(n48452));   // verilog/coms.v(116[11:12])
    defparam i1_2_lut_3_lut_adj_1627.LUT_INIT = 16'he0e0;
    SB_LUT4 i15559_3_lut_4_lut (.I0(n8_adj_4678), .I1(n48993), .I2(rx_data[7]), 
            .I3(\data_in_frame[14] [7]), .O(n29639));
    defparam i15559_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15560_3_lut_4_lut (.I0(n8_adj_4678), .I1(n48993), .I2(rx_data[6]), 
            .I3(\data_in_frame[14] [6]), .O(n29640));
    defparam i15560_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1628 (.I0(n110), .I1(n49), .I2(\FRAME_MATCHER.state [8]), 
            .I3(GND_net), .O(n48454));   // verilog/coms.v(116[11:12])
    defparam i1_2_lut_3_lut_adj_1628.LUT_INIT = 16'he0e0;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_41072 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [2]), .I2(\data_out_frame[27] [2]), 
            .I3(byte_transmit_counter[1]), .O(n56958));
    defparam byte_transmit_counter_0__bdd_4_lut_41072.LUT_INIT = 16'he4aa;
    SB_LUT4 i15561_3_lut_4_lut (.I0(n8_adj_4678), .I1(n48993), .I2(rx_data[5]), 
            .I3(\data_in_frame[14] [5]), .O(n29641));
    defparam i15561_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15562_3_lut_4_lut (.I0(n8_adj_4678), .I1(n48993), .I2(rx_data[4]), 
            .I3(\data_in_frame[14] [4]), .O(n29642));
    defparam i15562_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i37324_3_lut (.I0(\data_out_frame[6] [3]), .I1(\data_out_frame[7] [3]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n53154));
    defparam i37324_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i37325_4_lut (.I0(n53154), .I1(byte_transmit_counter[1]), .I2(byte_transmit_counter[2]), 
            .I3(byte_transmit_counter[0]), .O(n53155));
    defparam i37325_4_lut.LUT_INIT = 16'hafa3;
    SB_LUT4 i37323_3_lut (.I0(\data_out_frame[4] [3]), .I1(\data_out_frame[5] [3]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n53153));
    defparam i37323_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15563_3_lut_4_lut (.I0(n8_adj_4678), .I1(n48993), .I2(rx_data[3]), 
            .I3(\data_in_frame[14] [3]), .O(n29643));
    defparam i15563_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i40773_2_lut_3_lut (.I0(\FRAME_MATCHER.state [1]), .I1(\FRAME_MATCHER.state [2]), 
            .I2(\FRAME_MATCHER.state[0] ), .I3(GND_net), .O(n29136));
    defparam i40773_2_lut_3_lut.LUT_INIT = 16'h0e0e;
    SB_LUT4 i1_2_lut_3_lut_adj_1629 (.I0(n110), .I1(n49), .I2(\FRAME_MATCHER.state [9]), 
            .I3(GND_net), .O(n7_adj_4771));   // verilog/coms.v(116[11:12])
    defparam i1_2_lut_3_lut_adj_1629.LUT_INIT = 16'he0e0;
    SB_LUT4 select_713_Select_31_i3_2_lut (.I0(\FRAME_MATCHER.i [31]), .I1(n4623), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4707));
    defparam select_713_Select_31_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i40070_2_lut_3_lut (.I0(n28124), .I1(\data_in_frame[8] [3]), 
            .I2(\data_in_frame[8][4] ), .I3(GND_net), .O(n55901));
    defparam i40070_2_lut_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i15564_3_lut_4_lut (.I0(n8_adj_4678), .I1(n48993), .I2(rx_data[2]), 
            .I3(\data_in_frame[14] [2]), .O(n29644));
    defparam i15564_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15565_3_lut_4_lut (.I0(n8_adj_4678), .I1(n48993), .I2(rx_data[1]), 
            .I3(\data_in_frame[14] [1]), .O(n29645));
    defparam i15565_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15566_3_lut_4_lut (.I0(n8_adj_4678), .I1(n48993), .I2(rx_data[0]), 
            .I3(\data_in_frame[14] [0]), .O(n29646));
    defparam i15566_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15492_3_lut_4_lut (.I0(n37171), .I1(n48984), .I2(rx_data[2]), 
            .I3(\data_in_frame[23] [2]), .O(n29572));
    defparam i15492_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i15493_3_lut_4_lut (.I0(n37171), .I1(n48984), .I2(rx_data[1]), 
            .I3(\data_in_frame[23] [1]), .O(n29573));
    defparam i15493_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i15494_3_lut_4_lut (.I0(n37171), .I1(n48984), .I2(rx_data[0]), 
            .I3(\data_in_frame[23] [0]), .O(n29574));
    defparam i15494_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i38989_2_lut (.I0(n56889), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n54592));
    defparam i38989_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1_2_lut_4_lut_adj_1630 (.I0(\data_in_frame[13] [0]), .I1(\data_in_frame[12] [5]), 
            .I2(n27692), .I3(n28138), .O(n28132));
    defparam i1_2_lut_4_lut_adj_1630.LUT_INIT = 16'h6996;
    SB_LUT4 n56958_bdd_4_lut (.I0(n56958), .I1(\data_out_frame[25] [2]), 
            .I2(\data_out_frame[24] [2]), .I3(byte_transmit_counter[1]), 
            .O(n56961));
    defparam n56958_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i15883_3_lut_4_lut (.I0(n37171), .I1(n48984), .I2(rx_data[4]), 
            .I3(\data_in_frame[23] [4]), .O(n29963));
    defparam i15883_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_adj_1631 (.I0(\data_in_frame[12] [7]), .I1(n49342), 
            .I2(GND_net), .I3(GND_net), .O(n49590));
    defparam i1_2_lut_adj_1631.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1632 (.I0(n27604), .I1(\data_in_frame[15] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n49633));
    defparam i1_2_lut_adj_1632.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1633 (.I0(n49328), .I1(\data_in_frame[16] [5]), 
            .I2(n46673), .I3(GND_net), .O(n45766));
    defparam i2_3_lut_adj_1633.LUT_INIT = 16'h9696;
    SB_LUT4 i37318_3_lut (.I0(\data_out_frame[6] [4]), .I1(\data_out_frame[7] [4]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n53148));
    defparam i37318_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1634 (.I0(n49495), .I1(n28382), .I2(\data_in_frame[1] [4]), 
            .I3(\data_in_frame[8] [0]), .O(n49492));
    defparam i1_4_lut_adj_1634.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1635 (.I0(\state[0] ), .I1(\state[2] ), .I2(\state[3] ), 
            .I3(GND_net), .O(n7936));
    defparam i1_2_lut_3_lut_adj_1635.LUT_INIT = 16'h0202;
    SB_LUT4 i37319_4_lut (.I0(n53148), .I1(byte_transmit_counter[1]), .I2(byte_transmit_counter[2]), 
            .I3(byte_transmit_counter[0]), .O(n53149));
    defparam i37319_4_lut.LUT_INIT = 16'haca3;
    SB_LUT4 i1_3_lut_adj_1636 (.I0(\data_in_frame[16] [7]), .I1(n45914), 
            .I2(\data_in_frame[14] [6]), .I3(GND_net), .O(n49052));
    defparam i1_3_lut_adj_1636.LUT_INIT = 16'h9696;
    SB_LUT4 i37317_3_lut (.I0(\data_out_frame[4] [4]), .I1(\data_out_frame[5] [4]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n53147));
    defparam i37317_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3_4_lut_adj_1637 (.I0(\data_in_frame[11] [3]), .I1(n49162), 
            .I2(\data_in_frame[8] [7]), .I3(n27962), .O(n27612));   // verilog/coms.v(73[16:41])
    defparam i3_4_lut_adj_1637.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1638 (.I0(n28382), .I1(n28268), .I2(n49705), 
            .I3(GND_net), .O(n49120));
    defparam i1_2_lut_3_lut_adj_1638.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1639 (.I0(\data_in_frame[10][7] ), .I1(\data_in_frame[11] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n49612));
    defparam i1_2_lut_adj_1639.LUT_INIT = 16'h6666;
    SB_LUT4 i2_4_lut_adj_1640 (.I0(n49652), .I1(\data_in_frame[9] [4]), 
            .I2(\data_in_frame[9] [1]), .I3(n27352), .O(n49404));
    defparam i2_4_lut_adj_1640.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1641 (.I0(\data_in_frame[12] [0]), .I1(\data_in_frame[9] [7]), 
            .I2(\data_in_frame[12] [1]), .I3(GND_net), .O(n49670));
    defparam i2_3_lut_adj_1641.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1642 (.I0(\data_in_frame[5] [3]), .I1(n28030), 
            .I2(GND_net), .I3(GND_net), .O(n49172));
    defparam i1_2_lut_adj_1642.LUT_INIT = 16'h6666;
    SB_LUT4 i37312_3_lut (.I0(\data_out_frame[6] [5]), .I1(\data_out_frame[7] [5]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n53142));
    defparam i37312_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_adj_1643 (.I0(\data_in_frame[2] [6]), .I1(\data_in_frame[0] [5]), 
            .I2(\data_in_frame[0] [4]), .I3(\data_in_frame[5] [3]), .O(n52864));
    defparam i1_2_lut_4_lut_adj_1643.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1644 (.I0(\data_in_frame[2] [6]), .I1(\data_in_frame[0] [5]), 
            .I2(\data_in_frame[0] [4]), .I3(GND_net), .O(n4_adj_4835));   // verilog/coms.v(77[16:27])
    defparam i1_2_lut_3_lut_adj_1644.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1645 (.I0(\data_in_frame[3] [5]), .I1(\data_in_frame[5] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n52774));   // verilog/coms.v(76[16:27])
    defparam i1_2_lut_adj_1645.LUT_INIT = 16'h6666;
    SB_LUT4 i37311_3_lut (.I0(\data_out_frame[4] [5]), .I1(\data_out_frame[5] [5]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n53141));
    defparam i37311_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_adj_1646 (.I0(\data_in_frame[7] [7]), .I1(n27706), 
            .I2(n28030), .I3(\data_in_frame[5] [5]), .O(n28382));   // verilog/coms.v(76[16:27])
    defparam i1_2_lut_4_lut_adj_1646.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1647 (.I0(n28527), .I1(n28382), .I2(n49071), 
            .I3(n52774), .O(n25500));   // verilog/coms.v(76[16:27])
    defparam i1_4_lut_adj_1647.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1648 (.I0(n27706), .I1(\data_in_frame[8] [0]), 
            .I2(n49399), .I3(GND_net), .O(n49688));
    defparam i1_2_lut_3_lut_adj_1648.LUT_INIT = 16'h9696;
    SB_LUT4 i22461_3_lut_4_lut (.I0(n122), .I1(n27110), .I2(\FRAME_MATCHER.i [31]), 
            .I3(n63_adj_6), .O(\FRAME_MATCHER.state_31__N_3007[2] ));   // verilog/coms.v(228[6] 230[9])
    defparam i22461_3_lut_4_lut.LUT_INIT = 16'hae0c;
    SB_LUT4 i2_4_lut_adj_1649 (.I0(n60), .I1(n75), .I2(n2_adj_4661), .I3(n63_adj_4662), 
            .O(n6_c));
    defparam i2_4_lut_adj_1649.LUT_INIT = 16'h8000;
    SB_LUT4 i1_2_lut_adj_1650 (.I0(\data_in_frame[9] [4]), .I1(n27659), 
            .I2(GND_net), .I3(GND_net), .O(n27378));
    defparam i1_2_lut_adj_1650.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_4_lut_adj_1651 (.I0(\FRAME_MATCHER.state[0] ), .I1(n27223), 
            .I2(n4_adj_4688), .I3(n36546), .O(n6_adj_4663));
    defparam i1_2_lut_4_lut_adj_1651.LUT_INIT = 16'hfe00;
    SB_LUT4 i1_2_lut_adj_1652 (.I0(\data_in_frame[9] [5]), .I1(\data_in_frame[11] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n49478));   // verilog/coms.v(75[16:43])
    defparam i1_2_lut_adj_1652.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1653 (.I0(\data_in_frame[18] [2]), .I1(n46458), 
            .I2(GND_net), .I3(GND_net), .O(n46686));
    defparam i1_2_lut_adj_1653.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1654 (.I0(n27217), .I1(n24280), .I2(n24278), 
            .I3(\FRAME_MATCHER.state [2]), .O(n14_adj_4762));
    defparam i1_4_lut_adj_1654.LUT_INIT = 16'h5044;
    SB_LUT4 i1_4_lut_adj_1655 (.I0(n46832), .I1(\data_in_frame[21] [3]), 
            .I2(n49013), .I3(n50429), .O(n45752));
    defparam i1_4_lut_adj_1655.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1656 (.I0(\data_in_frame[19] [2]), .I1(n46100), 
            .I2(GND_net), .I3(GND_net), .O(n49013));
    defparam i1_2_lut_adj_1656.LUT_INIT = 16'h6666;
    SB_LUT4 i5842_2_lut (.I0(n63_adj_4650), .I1(n63_adj_4644), .I2(GND_net), 
            .I3(GND_net), .O(n19836));   // verilog/coms.v(140[4] 142[7])
    defparam i5842_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i5_4_lut_adj_1657 (.I0(\data_in_frame[12] [5]), .I1(n49240), 
            .I2(\data_in_frame[17] [1]), .I3(\data_in_frame[14] [5]), .O(n12_adj_4838));
    defparam i5_4_lut_adj_1657.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1658 (.I0(n28539), .I1(n12_adj_4838), .I2(n49543), 
            .I3(\data_in_frame[14] [7]), .O(n46100));
    defparam i6_4_lut_adj_1658.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1659 (.I0(n46100), .I1(n49097), .I2(GND_net), 
            .I3(GND_net), .O(n46816));
    defparam i1_2_lut_adj_1659.LUT_INIT = 16'h6666;
    SB_LUT4 i1_3_lut_adj_1660 (.I0(\FRAME_MATCHER.i_31__N_2845 ), .I1(n22875), 
            .I2(n4452), .I3(GND_net), .O(n49));
    defparam i1_3_lut_adj_1660.LUT_INIT = 16'h0808;
    SB_LUT4 i15884_3_lut_4_lut (.I0(n37171), .I1(n48984), .I2(rx_data[5]), 
            .I3(\data_in_frame[23] [5]), .O(n29964));
    defparam i15884_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i15885_3_lut_4_lut (.I0(n37171), .I1(n48984), .I2(rx_data[6]), 
            .I3(\data_in_frame[23] [6]), .O(n29965));
    defparam i15885_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i38943_2_lut (.I0(n56973), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n54599));
    defparam i38943_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i39023_2_lut (.I0(n56979), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n54601));
    defparam i39023_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1_2_lut_4_lut_adj_1661 (.I0(n3303), .I1(n22875), .I2(\FRAME_MATCHER.state [2]), 
            .I3(n27217), .O(n5_adj_4626));
    defparam i1_2_lut_4_lut_adj_1661.LUT_INIT = 16'h0040;
    SB_LUT4 i15886_3_lut_4_lut (.I0(n37171), .I1(n48984), .I2(rx_data[7]), 
            .I3(\data_in_frame[23] [7]), .O(n29966));
    defparam i15886_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_4_lut_adj_1662 (.I0(n49046), .I1(\data_in_frame[18] [5]), 
            .I2(\data_in_frame[18] [3]), .I3(\data_in_frame[22] [7]), .O(n52608));
    defparam i1_4_lut_adj_1662.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_41067 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [1]), .I2(\data_out_frame[27] [1]), 
            .I3(byte_transmit_counter[1]), .O(n56952));
    defparam byte_transmit_counter_0__bdd_4_lut_41067.LUT_INIT = 16'he4aa;
    SB_LUT4 i37571_4_lut (.I0(\data_out_frame[6] [6]), .I1(byte_transmit_counter[0]), 
            .I2(byte_transmit_counter[2]), .I3(\data_out_frame[7] [6]), 
            .O(n53401));
    defparam i37571_4_lut.LUT_INIT = 16'hec2c;
    SB_LUT4 i37569_3_lut (.I0(\data_out_frame[4] [6]), .I1(\data_out_frame[5] [6]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n53399));
    defparam i37569_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut_4_lut_adj_1663 (.I0(n8_adj_4697), .I1(\FRAME_MATCHER.i [4]), 
            .I2(n27304), .I3(\FRAME_MATCHER.i [3]), .O(n27110));
    defparam i1_3_lut_4_lut_adj_1663.LUT_INIT = 16'hfefc;
    SB_LUT4 i38949_2_lut (.I0(n56883), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n54603));
    defparam i38949_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1_2_lut_4_lut_adj_1664 (.I0(\FRAME_MATCHER.state [2]), .I1(n45364), 
            .I2(\FRAME_MATCHER.i [31]), .I3(n22875), .O(n3_adj_4627));
    defparam i1_2_lut_4_lut_adj_1664.LUT_INIT = 16'h5100;
    SB_LUT4 mux_2112_i2_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n36483), 
            .I2(\data_in_frame[3] [1]), .I3(\data_in_frame[19] [1]), .O(n7674));
    defparam mux_2112_i2_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 mux_2112_i3_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n36483), 
            .I2(\data_in_frame[3] [2]), .I3(\data_in_frame[19] [2]), .O(n7675));
    defparam mux_2112_i3_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 mux_2112_i4_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n36483), 
            .I2(\data_in_frame[3] [3]), .I3(\data_in_frame[19] [3]), .O(n7676));
    defparam mux_2112_i4_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i22482_2_lut (.I0(n27214), .I1(n63), .I2(GND_net), .I3(GND_net), 
            .O(n36546));
    defparam i22482_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i3_3_lut_adj_1665 (.I0(\FRAME_MATCHER.state[0] ), .I1(n6), .I2(\FRAME_MATCHER.state[3] ), 
            .I3(GND_net), .O(n63));   // verilog/coms.v(202[5:24])
    defparam i3_3_lut_adj_1665.LUT_INIT = 16'hefef;
    SB_LUT4 i22392_2_lut_4_lut (.I0(\FRAME_MATCHER.i_31__N_2845 ), .I1(n27217), 
            .I2(rx_data_ready), .I3(\FRAME_MATCHER.rx_data_ready_prev ), 
            .O(n36451));
    defparam i22392_2_lut_4_lut.LUT_INIT = 16'h00b0;
    SB_LUT4 i15231_2_lut (.I0(n28738), .I1(n27214), .I2(GND_net), .I3(GND_net), 
            .O(n29306));   // verilog/coms.v(128[12] 303[6])
    defparam i15231_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 n56952_bdd_4_lut (.I0(n56952), .I1(\data_out_frame[25] [1]), 
            .I2(\data_out_frame[24] [1]), .I3(byte_transmit_counter[1]), 
            .O(n56955));
    defparam n56952_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_4_lut_adj_1666 (.I0(n52744), .I1(n52414), .I2(n45939), 
            .I3(n51304), .O(n52418));
    defparam i1_4_lut_adj_1666.LUT_INIT = 16'hffed;
    SB_LUT4 i1_4_lut_adj_1667 (.I0(n49643), .I1(n49122), .I2(\data_in_frame[23] [0]), 
            .I3(n49699), .O(n50995));
    defparam i1_4_lut_adj_1667.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1668 (.I0(\data_in_frame[1] [0]), .I1(Kp_23__N_1098), 
            .I2(\data_in_frame[0] [5]), .I3(\data_in_frame[2] [7]), .O(n27862));
    defparam i1_2_lut_4_lut_adj_1668.LUT_INIT = 16'h6996;
    SB_LUT4 i1_3_lut_4_lut_adj_1669 (.I0(n45874), .I1(\data_in_frame[19] [6]), 
            .I2(n46852), .I3(n45811), .O(n46031));
    defparam i1_3_lut_4_lut_adj_1669.LUT_INIT = 16'h9669;
    SB_LUT4 mux_2112_i5_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n36483), 
            .I2(\data_in_frame[3] [4]), .I3(\data_in_frame[19] [4]), .O(n7677));
    defparam mux_2112_i5_3_lut_4_lut.LUT_INIT = 16'hfd20;
    uart_tx tx (.n28848(n28848), .clk16MHz(clk16MHz), .n29280(n29280), 
            .\r_SM_Main_2__N_3851[0] (r_SM_Main_2__N_3851[0]), .r_SM_Main({r_SM_Main}), 
            .\r_SM_Main_2__N_3848[1] (\r_SM_Main_2__N_3848[1] ), .GND_net(GND_net), 
            .\r_Bit_Index[0] (\r_Bit_Index[0] ), .VCC_net(VCC_net), .tx_o(tx_o), 
            .tx_data({tx_data}), .n19728(n19728), .n29842(n29842), .n29413(n29413), 
            .tx_active(tx_active), .n57032(n57032), .n4(n4_adj_7), .tx_enable(tx_enable)) /* synthesis syn_module_defined=1 */ ;   // verilog/coms.v(108[10:70])
    uart_rx rx (.r_SM_Main({r_SM_Main_adj_15}), .\r_SM_Main_2__N_3777[2] (\r_SM_Main_2__N_3777[2] ), 
            .GND_net(GND_net), .r_Rx_Data(r_Rx_Data), .n28852(n28852), 
            .clk16MHz(clk16MHz), .n29282(n29282), .VCC_net(VCC_net), .RX_N_10(RX_N_10), 
            .\r_Bit_Index[0] (\r_Bit_Index[0]_adj_11 ), .n4(n4_adj_12), 
            .n36556(n36556), .n4_adj_4(n4_adj_13), .n4_adj_5(n4_adj_14), 
            .n29845(n29845), .n48522(n48522), .rx_data_ready(rx_data_ready), 
            .n48878(n48878), .n29880(n29880), .rx_data({rx_data}), .n29878(n29878), 
            .n29877(n29877), .n29871(n29871), .n29860(n29860), .n29849(n29849), 
            .n29759(n29759), .n29528(n29528), .n27208(n27208), .n27203(n27203)) /* synthesis syn_module_defined=1 */ ;   // verilog/coms.v(94[10:44])
    
endmodule
//
// Verilog Description of module uart_tx
//

module uart_tx (n28848, clk16MHz, n29280, \r_SM_Main_2__N_3851[0] , 
            r_SM_Main, \r_SM_Main_2__N_3848[1] , GND_net, \r_Bit_Index[0] , 
            VCC_net, tx_o, tx_data, n19728, n29842, n29413, tx_active, 
            n57032, n4, tx_enable) /* synthesis syn_module_defined=1 */ ;
    output n28848;
    input clk16MHz;
    output n29280;
    input \r_SM_Main_2__N_3851[0] ;
    output [2:0]r_SM_Main;
    output \r_SM_Main_2__N_3848[1] ;
    input GND_net;
    output \r_Bit_Index[0] ;
    input VCC_net;
    output tx_o;
    input [7:0]tx_data;
    output n19728;
    input n29842;
    input n29413;
    output tx_active;
    input n57032;
    output n4;
    output tx_enable;
    
    wire clk16MHz /* synthesis SET_AS_NETWORK=clk16MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    wire [2:0]n307;
    wire [2:0]r_Bit_Index;   // verilog/uart_tx.v(33[16:27])
    wire [8:0]n41;
    
    wire n1;
    wire [8:0]r_Clock_Count;   // verilog/uart_tx.v(32[16:29])
    
    wire n29180, n37070, n21944, n21945, o_Tx_Serial_N_3879, n3;
    wire [7:0]r_Tx_Data;   // verilog/uart_tx.v(34[16:25])
    
    wire n53246, n53247, n53250, n53249, n44622, n44621, n44620, 
        n44619, n44618, n44617, n44616, n44615, n26719, n56742, 
        n3_adj_4619, n50990, n10;
    
    SB_DFFESR r_Bit_Index_i1 (.Q(r_Bit_Index[1]), .C(clk16MHz), .E(n28848), 
            .D(n307[1]), .R(n29280));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFESR r_Bit_Index_i2 (.Q(r_Bit_Index[2]), .C(clk16MHz), .E(n28848), 
            .D(n307[2]), .R(n29280));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFESR r_Clock_Count_2292__i0 (.Q(r_Clock_Count[0]), .C(clk16MHz), 
            .E(n1), .D(n41[0]), .R(n29180));   // verilog/uart_tx.v(118[34:51])
    SB_LUT4 i7985_4_lut (.I0(\r_SM_Main_2__N_3851[0] ), .I1(n37070), .I2(r_SM_Main[1]), 
            .I3(\r_SM_Main_2__N_3848[1] ), .O(n21944));   // verilog/uart_tx.v(43[7] 142[14])
    defparam i7985_4_lut.LUT_INIT = 16'hca0a;
    SB_LUT4 i7986_3_lut (.I0(n21944), .I1(\r_SM_Main_2__N_3848[1] ), .I2(r_SM_Main[0]), 
            .I3(GND_net), .O(n21945));   // verilog/uart_tx.v(43[7] 142[14])
    defparam i7986_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 r_SM_Main_2__I_0_56_i3_3_lut (.I0(r_SM_Main[0]), .I1(o_Tx_Serial_N_3879), 
            .I2(r_SM_Main[1]), .I3(GND_net), .O(n3));   // verilog/uart_tx.v(43[7] 142[14])
    defparam r_SM_Main_2__I_0_56_i3_3_lut.LUT_INIT = 16'he5e5;
    SB_LUT4 i37416_3_lut (.I0(r_Tx_Data[0]), .I1(r_Tx_Data[1]), .I2(\r_Bit_Index[0] ), 
            .I3(GND_net), .O(n53246));
    defparam i37416_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i37417_3_lut (.I0(r_Tx_Data[2]), .I1(r_Tx_Data[3]), .I2(\r_Bit_Index[0] ), 
            .I3(GND_net), .O(n53247));
    defparam i37417_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i37420_3_lut (.I0(r_Tx_Data[6]), .I1(r_Tx_Data[7]), .I2(\r_Bit_Index[0] ), 
            .I3(GND_net), .O(n53250));
    defparam i37420_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i37419_3_lut (.I0(r_Tx_Data[4]), .I1(r_Tx_Data[5]), .I2(\r_Bit_Index[0] ), 
            .I3(GND_net), .O(n53249));
    defparam i37419_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 r_Clock_Count_2292_add_4_10_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[8]), .I3(n44622), .O(n41[8])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2292_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 r_Clock_Count_2292_add_4_9_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[7]), .I3(n44621), .O(n41[7])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2292_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2292_add_4_9 (.CI(n44621), .I0(GND_net), .I1(r_Clock_Count[7]), 
            .CO(n44622));
    SB_LUT4 r_Clock_Count_2292_add_4_8_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[6]), .I3(n44620), .O(n41[6])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2292_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2292_add_4_8 (.CI(n44620), .I0(GND_net), .I1(r_Clock_Count[6]), 
            .CO(n44621));
    SB_LUT4 r_Clock_Count_2292_add_4_7_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[5]), .I3(n44619), .O(n41[5])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2292_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2292_add_4_7 (.CI(n44619), .I0(GND_net), .I1(r_Clock_Count[5]), 
            .CO(n44620));
    SB_LUT4 r_Clock_Count_2292_add_4_6_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[4]), .I3(n44618), .O(n41[4])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2292_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2292_add_4_6 (.CI(n44618), .I0(GND_net), .I1(r_Clock_Count[4]), 
            .CO(n44619));
    SB_LUT4 r_Clock_Count_2292_add_4_5_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[3]), .I3(n44617), .O(n41[3])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2292_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2292_add_4_5 (.CI(n44617), .I0(GND_net), .I1(r_Clock_Count[3]), 
            .CO(n44618));
    SB_LUT4 r_Clock_Count_2292_add_4_4_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[2]), .I3(n44616), .O(n41[2])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2292_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2292_add_4_4 (.CI(n44616), .I0(GND_net), .I1(r_Clock_Count[2]), 
            .CO(n44617));
    SB_LUT4 r_Clock_Count_2292_add_4_3_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[1]), .I3(n44615), .O(n41[1])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2292_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2292_add_4_3 (.CI(n44615), .I0(GND_net), .I1(r_Clock_Count[1]), 
            .CO(n44616));
    SB_LUT4 r_Clock_Count_2292_add_4_2_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[0]), .I3(VCC_net), .O(n41[0])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2292_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2292_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(r_Clock_Count[0]), 
            .CO(n44615));
    SB_DFFE o_Tx_Serial_45 (.Q(tx_o), .C(clk16MHz), .E(n1), .D(n3));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i0 (.Q(r_Tx_Data[0]), .C(clk16MHz), .E(n26719), 
            .D(tx_data[0]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFSR r_SM_Main_i0 (.Q(r_SM_Main[0]), .C(clk16MHz), .D(n21945), 
            .R(r_SM_Main[2]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_LUT4 i5778_2_lut (.I0(\r_SM_Main_2__N_3851[0] ), .I1(r_SM_Main[0]), 
            .I2(GND_net), .I3(GND_net), .O(n19728));   // verilog/uart_tx.v(43[7] 142[14])
    defparam i5778_2_lut.LUT_INIT = 16'h2222;
    SB_DFFESR r_Clock_Count_2292__i1 (.Q(r_Clock_Count[1]), .C(clk16MHz), 
            .E(n1), .D(n41[1]), .R(n29180));   // verilog/uart_tx.v(118[34:51])
    SB_DFFESR r_Clock_Count_2292__i2 (.Q(r_Clock_Count[2]), .C(clk16MHz), 
            .E(n1), .D(n41[2]), .R(n29180));   // verilog/uart_tx.v(118[34:51])
    SB_DFFESR r_Clock_Count_2292__i3 (.Q(r_Clock_Count[3]), .C(clk16MHz), 
            .E(n1), .D(n41[3]), .R(n29180));   // verilog/uart_tx.v(118[34:51])
    SB_DFFESR r_Clock_Count_2292__i4 (.Q(r_Clock_Count[4]), .C(clk16MHz), 
            .E(n1), .D(n41[4]), .R(n29180));   // verilog/uart_tx.v(118[34:51])
    SB_DFFESR r_Clock_Count_2292__i5 (.Q(r_Clock_Count[5]), .C(clk16MHz), 
            .E(n1), .D(n41[5]), .R(n29180));   // verilog/uart_tx.v(118[34:51])
    SB_DFFESR r_Clock_Count_2292__i6 (.Q(r_Clock_Count[6]), .C(clk16MHz), 
            .E(n1), .D(n41[6]), .R(n29180));   // verilog/uart_tx.v(118[34:51])
    SB_DFFESR r_Clock_Count_2292__i7 (.Q(r_Clock_Count[7]), .C(clk16MHz), 
            .E(n1), .D(n41[7]), .R(n29180));   // verilog/uart_tx.v(118[34:51])
    SB_DFFESR r_Clock_Count_2292__i8 (.Q(r_Clock_Count[8]), .C(clk16MHz), 
            .E(n1), .D(n41[8]), .R(n29180));   // verilog/uart_tx.v(118[34:51])
    SB_DFF r_Bit_Index_i0 (.Q(\r_Bit_Index[0] ), .C(clk16MHz), .D(n29842));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Tx_Active_47 (.Q(tx_active), .C(clk16MHz), .D(n29413));   // verilog/uart_tx.v(40[10] 143[8])
    SB_LUT4 r_Bit_Index_1__bdd_4_lut (.I0(r_Bit_Index[1]), .I1(n53249), 
            .I2(n53250), .I3(r_Bit_Index[2]), .O(n56742));
    defparam r_Bit_Index_1__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n56742_bdd_4_lut (.I0(n56742), .I1(n53247), .I2(n53246), .I3(r_Bit_Index[2]), 
            .O(o_Tx_Serial_N_3879));
    defparam n56742_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFFSR r_SM_Main_i1 (.Q(r_SM_Main[1]), .C(clk16MHz), .D(n3_adj_4619), 
            .R(r_SM_Main[2]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i7 (.Q(r_Tx_Data[7]), .C(clk16MHz), .E(n26719), 
            .D(tx_data[7]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i6 (.Q(r_Tx_Data[6]), .C(clk16MHz), .E(n26719), 
            .D(tx_data[6]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i5 (.Q(r_Tx_Data[5]), .C(clk16MHz), .E(n26719), 
            .D(tx_data[5]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i4 (.Q(r_Tx_Data[4]), .C(clk16MHz), .E(n26719), 
            .D(tx_data[4]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i3 (.Q(r_Tx_Data[3]), .C(clk16MHz), .E(n26719), 
            .D(tx_data[3]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i2 (.Q(r_Tx_Data[2]), .C(clk16MHz), .E(n26719), 
            .D(tx_data[2]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i1 (.Q(r_Tx_Data[1]), .C(clk16MHz), .E(n26719), 
            .D(tx_data[1]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_SM_Main_i2 (.Q(r_SM_Main[2]), .C(clk16MHz), .D(n57032));   // verilog/uart_tx.v(40[10] 143[8])
    SB_LUT4 i40116_4_lut (.I0(r_SM_Main[2]), .I1(\r_SM_Main_2__N_3848[1] ), 
            .I2(r_SM_Main[1]), .I3(r_SM_Main[0]), .O(n29180));
    defparam i40116_4_lut.LUT_INIT = 16'h4445;
    SB_LUT4 i1_1_lut (.I0(r_SM_Main[2]), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n1));
    defparam i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_3_lut_4_lut_4_lut (.I0(\r_SM_Main_2__N_3848[1] ), .I1(r_SM_Main[0]), 
            .I2(r_SM_Main[1]), .I3(r_SM_Main[2]), .O(n4));
    defparam i1_3_lut_4_lut_4_lut.LUT_INIT = 16'h008f;
    SB_LUT4 i2471_3_lut (.I0(r_Bit_Index[2]), .I1(r_Bit_Index[1]), .I2(\r_Bit_Index[0] ), 
            .I3(GND_net), .O(n307[2]));   // verilog/uart_tx.v(98[36:51])
    defparam i2471_3_lut.LUT_INIT = 16'h6a6a;
    SB_LUT4 i3_4_lut (.I0(r_Clock_Count[0]), .I1(r_Clock_Count[3]), .I2(r_Clock_Count[1]), 
            .I3(r_Clock_Count[2]), .O(n50990));
    defparam i3_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i4_4_lut (.I0(r_Clock_Count[4]), .I1(r_Clock_Count[5]), .I2(n50990), 
            .I3(r_Clock_Count[8]), .O(n10));
    defparam i4_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i5_3_lut (.I0(r_Clock_Count[6]), .I1(n10), .I2(r_Clock_Count[7]), 
            .I3(GND_net), .O(\r_SM_Main_2__N_3848[1] ));
    defparam i5_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i2_3_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), .I2(\r_Bit_Index[0] ), 
            .I3(GND_net), .O(n37070));
    defparam i2_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i15200_3_lut (.I0(n28848), .I1(n37070), .I2(r_SM_Main[1]), 
            .I3(GND_net), .O(n29280));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i15200_3_lut.LUT_INIT = 16'h8a8a;
    SB_LUT4 i2464_2_lut (.I0(r_Bit_Index[1]), .I1(\r_Bit_Index[0] ), .I2(GND_net), 
            .I3(GND_net), .O(n307[1]));   // verilog/uart_tx.v(98[36:51])
    defparam i2464_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_4_lut (.I0(r_SM_Main[2]), .I1(r_SM_Main[0]), .I2(\r_SM_Main_2__N_3851[0] ), 
            .I3(r_SM_Main[1]), .O(n26719));
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h0010;
    SB_LUT4 i1_3_lut_4_lut (.I0(r_SM_Main[2]), .I1(r_SM_Main[0]), .I2(r_SM_Main[1]), 
            .I3(\r_SM_Main_2__N_3848[1] ), .O(n28848));
    defparam i1_3_lut_4_lut.LUT_INIT = 16'h1101;
    SB_LUT4 i9998_2_lut_3_lut (.I0(\r_SM_Main_2__N_3848[1] ), .I1(r_SM_Main[0]), 
            .I2(r_SM_Main[1]), .I3(GND_net), .O(n3_adj_4619));
    defparam i9998_2_lut_3_lut.LUT_INIT = 16'h7878;
    SB_LUT4 o_Tx_Serial_I_0_1_lut (.I0(tx_o), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(tx_enable));   // verilog/uart_tx.v(38[24:36])
    defparam o_Tx_Serial_I_0_1_lut.LUT_INIT = 16'h5555;
    
endmodule
//
// Verilog Description of module uart_rx
//

module uart_rx (r_SM_Main, \r_SM_Main_2__N_3777[2] , GND_net, r_Rx_Data, 
            n28852, clk16MHz, n29282, VCC_net, RX_N_10, \r_Bit_Index[0] , 
            n4, n36556, n4_adj_4, n4_adj_5, n29845, n48522, rx_data_ready, 
            n48878, n29880, rx_data, n29878, n29877, n29871, n29860, 
            n29849, n29759, n29528, n27208, n27203) /* synthesis syn_module_defined=1 */ ;
    output [2:0]r_SM_Main;
    output \r_SM_Main_2__N_3777[2] ;
    input GND_net;
    output r_Rx_Data;
    output n28852;
    input clk16MHz;
    output n29282;
    input VCC_net;
    input RX_N_10;
    output \r_Bit_Index[0] ;
    output n4;
    output n36556;
    output n4_adj_4;
    output n4_adj_5;
    input n29845;
    input n48522;
    output rx_data_ready;
    input n48878;
    input n29880;
    output [7:0]rx_data;
    input n29878;
    input n29877;
    input n29871;
    input n29860;
    input n29849;
    input n29759;
    input n29528;
    output n27208;
    output n27203;
    
    wire clk16MHz /* synthesis SET_AS_NETWORK=clk16MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    
    wire n28, n33112, n48602;
    wire [2:0]n326;
    wire [2:0]r_Bit_Index;   // verilog/uart_rx.v(33[17:28])
    wire [7:0]n37;
    
    wire n28800;
    wire [7:0]r_Clock_Count;   // verilog/uart_rx.v(32[17:30])
    
    wire n29188, n37072, n31, n48875, n29, n33, n44614, n44613, 
        n44612, n44611, n44610, n44609, n44608, r_Rx_Data_R, n27091, 
        n48936, n54612, n6;
    
    SB_LUT4 i1_2_lut (.I0(r_SM_Main[0]), .I1(\r_SM_Main_2__N_3777[2] ), 
            .I2(GND_net), .I3(GND_net), .O(n28));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i1_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i13_4_lut (.I0(n33112), .I1(n28), .I2(r_SM_Main[1]), .I3(r_Rx_Data), 
            .O(n48602));   // verilog/uart_rx.v(30[17:26])
    defparam i13_4_lut.LUT_INIT = 16'h303a;
    SB_DFFESR r_Bit_Index_i2 (.Q(r_Bit_Index[2]), .C(clk16MHz), .E(n28852), 
            .D(n326[2]), .R(n29282));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFFESR r_Clock_Count_2290__i0 (.Q(r_Clock_Count[0]), .C(clk16MHz), 
            .E(n28800), .D(n37[0]), .R(n29188));   // verilog/uart_rx.v(120[34:51])
    SB_DFFESR r_Clock_Count_2290__i1 (.Q(r_Clock_Count[1]), .C(clk16MHz), 
            .E(n28800), .D(n37[1]), .R(n29188));   // verilog/uart_rx.v(120[34:51])
    SB_LUT4 i33_3_lut (.I0(n37072), .I1(\r_SM_Main_2__N_3777[2] ), .I2(r_SM_Main[0]), 
            .I3(GND_net), .O(n31));   // verilog/uart_rx.v(30[17:26])
    defparam i33_3_lut.LUT_INIT = 16'hc7c7;
    SB_LUT4 i34_3_lut (.I0(r_Rx_Data), .I1(n48875), .I2(r_SM_Main[0]), 
            .I3(GND_net), .O(n29));   // verilog/uart_rx.v(30[17:26])
    defparam i34_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i32_3_lut (.I0(n29), .I1(n31), .I2(r_SM_Main[1]), .I3(GND_net), 
            .O(n33));   // verilog/uart_rx.v(30[17:26])
    defparam i32_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 r_Clock_Count_2290_add_4_9_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[7]), .I3(n44614), .O(n37[7])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2290_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 r_Clock_Count_2290_add_4_8_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[6]), .I3(n44613), .O(n37[6])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2290_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2290_add_4_8 (.CI(n44613), .I0(GND_net), .I1(r_Clock_Count[6]), 
            .CO(n44614));
    SB_LUT4 r_Clock_Count_2290_add_4_7_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[5]), .I3(n44612), .O(n37[5])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2290_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2290_add_4_7 (.CI(n44612), .I0(GND_net), .I1(r_Clock_Count[5]), 
            .CO(n44613));
    SB_LUT4 r_Clock_Count_2290_add_4_6_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[4]), .I3(n44611), .O(n37[4])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2290_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2290_add_4_6 (.CI(n44611), .I0(GND_net), .I1(r_Clock_Count[4]), 
            .CO(n44612));
    SB_LUT4 r_Clock_Count_2290_add_4_5_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[3]), .I3(n44610), .O(n37[3])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2290_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2290_add_4_5 (.CI(n44610), .I0(GND_net), .I1(r_Clock_Count[3]), 
            .CO(n44611));
    SB_LUT4 r_Clock_Count_2290_add_4_4_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[2]), .I3(n44609), .O(n37[2])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2290_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_DFFESR r_Clock_Count_2290__i2 (.Q(r_Clock_Count[2]), .C(clk16MHz), 
            .E(n28800), .D(n37[2]), .R(n29188));   // verilog/uart_rx.v(120[34:51])
    SB_CARRY r_Clock_Count_2290_add_4_4 (.CI(n44609), .I0(GND_net), .I1(r_Clock_Count[2]), 
            .CO(n44610));
    SB_DFFESR r_Clock_Count_2290__i3 (.Q(r_Clock_Count[3]), .C(clk16MHz), 
            .E(n28800), .D(n37[3]), .R(n29188));   // verilog/uart_rx.v(120[34:51])
    SB_LUT4 r_Clock_Count_2290_add_4_3_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[1]), .I3(n44608), .O(n37[1])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2290_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2290_add_4_3 (.CI(n44608), .I0(GND_net), .I1(r_Clock_Count[1]), 
            .CO(n44609));
    SB_LUT4 r_Clock_Count_2290_add_4_2_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[0]), .I3(VCC_net), .O(n37[0])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2290_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2290_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(r_Clock_Count[0]), 
            .CO(n44608));
    SB_DFFSR r_SM_Main_i0 (.Q(r_SM_Main[0]), .C(clk16MHz), .D(n33), .R(r_SM_Main[2]));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Data_50 (.Q(r_Rx_Data), .C(clk16MHz), .D(r_Rx_Data_R));   // verilog/uart_rx.v(41[10] 45[8])
    SB_DFF r_Rx_Data_R_49 (.Q(r_Rx_Data_R), .C(clk16MHz), .D(RX_N_10));   // verilog/uart_rx.v(41[10] 45[8])
    SB_DFFESR r_Clock_Count_2290__i4 (.Q(r_Clock_Count[4]), .C(clk16MHz), 
            .E(n28800), .D(n37[4]), .R(n29188));   // verilog/uart_rx.v(120[34:51])
    SB_DFFESR r_Clock_Count_2290__i5 (.Q(r_Clock_Count[5]), .C(clk16MHz), 
            .E(n28800), .D(n37[5]), .R(n29188));   // verilog/uart_rx.v(120[34:51])
    SB_DFFESR r_Clock_Count_2290__i6 (.Q(r_Clock_Count[6]), .C(clk16MHz), 
            .E(n28800), .D(n37[6]), .R(n29188));   // verilog/uart_rx.v(120[34:51])
    SB_DFFESR r_Clock_Count_2290__i7 (.Q(r_Clock_Count[7]), .C(clk16MHz), 
            .E(n28800), .D(n37[7]), .R(n29188));   // verilog/uart_rx.v(120[34:51])
    SB_LUT4 i2442_2_lut (.I0(r_Bit_Index[1]), .I1(\r_Bit_Index[0] ), .I2(GND_net), 
            .I3(GND_net), .O(n326[1]));   // verilog/uart_rx.v(102[36:51])
    defparam i2442_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 equal_379_i4_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(GND_net), .I3(GND_net), .O(n4));   // verilog/uart_rx.v(97[17:39])
    defparam equal_379_i4_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i22492_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), .I2(GND_net), 
            .I3(GND_net), .O(n36556));
    defparam i22492_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 equal_377_i4_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_4));   // verilog/uart_rx.v(97[17:39])
    defparam equal_377_i4_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 equal_375_i4_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_5));   // verilog/uart_rx.v(97[17:39])
    defparam equal_375_i4_2_lut.LUT_INIT = 16'hbbbb;
    SB_DFF r_Bit_Index_i0 (.Q(\r_Bit_Index[0] ), .C(clk16MHz), .D(n29845));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_DV_52 (.Q(rx_data_ready), .C(clk16MHz), .D(n48522));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFFESR r_Bit_Index_i1 (.Q(r_Bit_Index[1]), .C(clk16MHz), .E(n28852), 
            .D(n326[1]), .R(n29282));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_SM_Main_i2 (.Q(r_SM_Main[2]), .C(clk16MHz), .D(n48878));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFFSR r_SM_Main_i1 (.Q(r_SM_Main[1]), .C(clk16MHz), .D(n48602), 
            .R(r_SM_Main[2]));   // verilog/uart_rx.v(49[10] 144[8])
    SB_LUT4 i2_3_lut (.I0(n27091), .I1(r_Clock_Count[3]), .I2(n48936), 
            .I3(GND_net), .O(n48875));
    defparam i2_3_lut.LUT_INIT = 16'h1010;
    SB_LUT4 i1_2_lut_adj_951 (.I0(r_SM_Main[0]), .I1(n48875), .I2(GND_net), 
            .I3(GND_net), .O(n33112));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i1_2_lut_adj_951.LUT_INIT = 16'h8888;
    SB_LUT4 i39516_3_lut (.I0(r_Rx_Data), .I1(r_SM_Main[0]), .I2(n48875), 
            .I3(GND_net), .O(n54612));
    defparam i39516_3_lut.LUT_INIT = 16'h7373;
    SB_LUT4 i1_4_lut (.I0(r_SM_Main[2]), .I1(n54612), .I2(\r_SM_Main_2__N_3777[2] ), 
            .I3(r_SM_Main[1]), .O(n29188));
    defparam i1_4_lut.LUT_INIT = 16'h5044;
    SB_LUT4 i40771_4_lut (.I0(r_Rx_Data), .I1(r_SM_Main[2]), .I2(r_SM_Main[1]), 
            .I3(n33112), .O(n28800));
    defparam i40771_4_lut.LUT_INIT = 16'h3133;
    SB_LUT4 i2_3_lut_adj_952 (.I0(r_Clock_Count[0]), .I1(r_Clock_Count[1]), 
            .I2(r_Clock_Count[2]), .I3(GND_net), .O(n48936));
    defparam i2_3_lut_adj_952.LUT_INIT = 16'h8080;
    SB_LUT4 i3_4_lut (.I0(r_Clock_Count[4]), .I1(r_Clock_Count[7]), .I2(r_Clock_Count[6]), 
            .I3(r_Clock_Count[5]), .O(n27091));   // verilog/uart_rx.v(118[17:47])
    defparam i3_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_2_lut (.I0(r_SM_Main[0]), .I1(r_SM_Main[2]), .I2(GND_net), 
            .I3(GND_net), .O(n6));
    defparam i2_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i22991_3_lut (.I0(r_Clock_Count[3]), .I1(n27091), .I2(n48936), 
            .I3(GND_net), .O(\r_SM_Main_2__N_3777[2] ));
    defparam i22991_3_lut.LUT_INIT = 16'hecec;
    SB_LUT4 i2_3_lut_adj_953 (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(\r_Bit_Index[0] ), .I3(GND_net), .O(n37072));
    defparam i2_3_lut_adj_953.LUT_INIT = 16'h8080;
    SB_LUT4 i15202_3_lut (.I0(n28852), .I1(n37072), .I2(r_SM_Main[1]), 
            .I3(GND_net), .O(n29282));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i15202_3_lut.LUT_INIT = 16'h8a8a;
    SB_LUT4 i2449_3_lut (.I0(r_Bit_Index[2]), .I1(r_Bit_Index[1]), .I2(\r_Bit_Index[0] ), 
            .I3(GND_net), .O(n326[2]));   // verilog/uart_rx.v(102[36:51])
    defparam i2449_3_lut.LUT_INIT = 16'h6a6a;
    SB_DFF r_Rx_Byte_i5 (.Q(rx_data[5]), .C(clk16MHz), .D(n29880));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i4 (.Q(rx_data[4]), .C(clk16MHz), .D(n29878));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i3 (.Q(rx_data[3]), .C(clk16MHz), .D(n29877));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i2 (.Q(rx_data[2]), .C(clk16MHz), .D(n29871));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i7 (.Q(rx_data[7]), .C(clk16MHz), .D(n29860));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i0 (.Q(rx_data[0]), .C(clk16MHz), .D(n29849));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i1 (.Q(rx_data[1]), .C(clk16MHz), .D(n29759));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i6 (.Q(rx_data[6]), .C(clk16MHz), .D(n29528));   // verilog/uart_rx.v(49[10] 144[8])
    SB_LUT4 i1_3_lut_4_lut (.I0(\r_SM_Main_2__N_3777[2] ), .I1(r_SM_Main[0]), 
            .I2(r_SM_Main[2]), .I3(r_SM_Main[1]), .O(n28852));
    defparam i1_3_lut_4_lut.LUT_INIT = 16'h0203;
    SB_LUT4 i1_2_lut_4_lut (.I0(n6), .I1(\r_SM_Main_2__N_3777[2] ), .I2(r_SM_Main[1]), 
            .I3(\r_Bit_Index[0] ), .O(n27208));
    defparam i1_2_lut_4_lut.LUT_INIT = 16'hffbf;
    SB_LUT4 i1_2_lut_4_lut_adj_954 (.I0(n6), .I1(\r_SM_Main_2__N_3777[2] ), 
            .I2(r_SM_Main[1]), .I3(\r_Bit_Index[0] ), .O(n27203));
    defparam i1_2_lut_4_lut_adj_954.LUT_INIT = 16'hbfff;
    
endmodule
//
// Verilog Description of module pwm
//

module pwm (pwm_out, clk32MHz, GND_net, VCC_net, pwm_setpoint) /* synthesis syn_module_defined=1 */ ;
    output pwm_out;
    input clk32MHz;
    input GND_net;
    input VCC_net;
    input [23:0]pwm_setpoint;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[16:24])
    
    wire pwm_out_N_908;
    wire [23:0]n101;
    wire [23:0]pwm_counter;   // verilog/pwm.v(11[19:30])
    
    wire n44532, n44531, n44530, pwm_counter_23__N_906, n44529, n44528, 
        n44527, n44526, n44525, n44524, n44523, n44522, n44521, 
        n44520, n44519, n44518, n44517, n44516, n44515, n44514, 
        n44513, n44512, n44511, n44510, n8, n54937, n16, n54971, 
        n6, n10, n54948, n12, n41, n39, n45, n37, n43, n29, 
        n31, n23, n25, n35, n33, n11, n13, n15, n27, n9, 
        n17, n19, n21, n54960, n54954, n30, n55343, n55339, 
        n55764, n55528, n55804, n55598, n55599, n24, n54939, n55456, 
        n55167, n4, n55596, n55597, n54950, n55774, n55169, n55858, 
        n55859, n55833, n54941, n55708, n55175, n55792, n51426, 
        n22, n15_adj_4614, n20, n24_adj_4615, n19_adj_4616;
    
    SB_DFF pwm_out_12 (.Q(pwm_out), .C(clk32MHz), .D(pwm_out_N_908));   // verilog/pwm.v(16[12] 26[6])
    SB_LUT4 pwm_counter_2282_add_4_25_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[23]), 
            .I3(n44532), .O(n101[23])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2282_add_4_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 pwm_counter_2282_add_4_24_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[22]), 
            .I3(n44531), .O(n101[22])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2282_add_4_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_2282_add_4_24 (.CI(n44531), .I0(GND_net), .I1(pwm_counter[22]), 
            .CO(n44532));
    SB_LUT4 pwm_counter_2282_add_4_23_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[21]), 
            .I3(n44530), .O(n101[21])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2282_add_4_23_lut.LUT_INIT = 16'hC33C;
    SB_DFFSR pwm_counter_2282__i23 (.Q(pwm_counter[23]), .C(clk32MHz), .D(n101[23]), 
            .R(pwm_counter_23__N_906));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_2282__i22 (.Q(pwm_counter[22]), .C(clk32MHz), .D(n101[22]), 
            .R(pwm_counter_23__N_906));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_2282__i21 (.Q(pwm_counter[21]), .C(clk32MHz), .D(n101[21]), 
            .R(pwm_counter_23__N_906));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_2282__i20 (.Q(pwm_counter[20]), .C(clk32MHz), .D(n101[20]), 
            .R(pwm_counter_23__N_906));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_2282__i19 (.Q(pwm_counter[19]), .C(clk32MHz), .D(n101[19]), 
            .R(pwm_counter_23__N_906));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_2282__i18 (.Q(pwm_counter[18]), .C(clk32MHz), .D(n101[18]), 
            .R(pwm_counter_23__N_906));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_2282__i17 (.Q(pwm_counter[17]), .C(clk32MHz), .D(n101[17]), 
            .R(pwm_counter_23__N_906));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_2282__i16 (.Q(pwm_counter[16]), .C(clk32MHz), .D(n101[16]), 
            .R(pwm_counter_23__N_906));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_2282__i15 (.Q(pwm_counter[15]), .C(clk32MHz), .D(n101[15]), 
            .R(pwm_counter_23__N_906));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_2282__i14 (.Q(pwm_counter[14]), .C(clk32MHz), .D(n101[14]), 
            .R(pwm_counter_23__N_906));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_2282__i13 (.Q(pwm_counter[13]), .C(clk32MHz), .D(n101[13]), 
            .R(pwm_counter_23__N_906));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_2282__i12 (.Q(pwm_counter[12]), .C(clk32MHz), .D(n101[12]), 
            .R(pwm_counter_23__N_906));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_2282__i11 (.Q(pwm_counter[11]), .C(clk32MHz), .D(n101[11]), 
            .R(pwm_counter_23__N_906));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_2282__i10 (.Q(pwm_counter[10]), .C(clk32MHz), .D(n101[10]), 
            .R(pwm_counter_23__N_906));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_2282__i9 (.Q(pwm_counter[9]), .C(clk32MHz), .D(n101[9]), 
            .R(pwm_counter_23__N_906));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_2282__i8 (.Q(pwm_counter[8]), .C(clk32MHz), .D(n101[8]), 
            .R(pwm_counter_23__N_906));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_2282__i7 (.Q(pwm_counter[7]), .C(clk32MHz), .D(n101[7]), 
            .R(pwm_counter_23__N_906));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_2282__i6 (.Q(pwm_counter[6]), .C(clk32MHz), .D(n101[6]), 
            .R(pwm_counter_23__N_906));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_2282__i5 (.Q(pwm_counter[5]), .C(clk32MHz), .D(n101[5]), 
            .R(pwm_counter_23__N_906));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_2282__i4 (.Q(pwm_counter[4]), .C(clk32MHz), .D(n101[4]), 
            .R(pwm_counter_23__N_906));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_2282__i3 (.Q(pwm_counter[3]), .C(clk32MHz), .D(n101[3]), 
            .R(pwm_counter_23__N_906));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_2282__i2 (.Q(pwm_counter[2]), .C(clk32MHz), .D(n101[2]), 
            .R(pwm_counter_23__N_906));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_2282__i1 (.Q(pwm_counter[1]), .C(clk32MHz), .D(n101[1]), 
            .R(pwm_counter_23__N_906));   // verilog/pwm.v(17[20:33])
    SB_CARRY pwm_counter_2282_add_4_23 (.CI(n44530), .I0(GND_net), .I1(pwm_counter[21]), 
            .CO(n44531));
    SB_LUT4 pwm_counter_2282_add_4_22_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[20]), 
            .I3(n44529), .O(n101[20])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2282_add_4_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_2282_add_4_22 (.CI(n44529), .I0(GND_net), .I1(pwm_counter[20]), 
            .CO(n44530));
    SB_LUT4 pwm_counter_2282_add_4_21_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[19]), 
            .I3(n44528), .O(n101[19])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2282_add_4_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_2282_add_4_21 (.CI(n44528), .I0(GND_net), .I1(pwm_counter[19]), 
            .CO(n44529));
    SB_LUT4 pwm_counter_2282_add_4_20_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[18]), 
            .I3(n44527), .O(n101[18])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2282_add_4_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_2282_add_4_20 (.CI(n44527), .I0(GND_net), .I1(pwm_counter[18]), 
            .CO(n44528));
    SB_LUT4 pwm_counter_2282_add_4_19_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[17]), 
            .I3(n44526), .O(n101[17])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2282_add_4_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_2282_add_4_19 (.CI(n44526), .I0(GND_net), .I1(pwm_counter[17]), 
            .CO(n44527));
    SB_LUT4 pwm_counter_2282_add_4_18_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[16]), 
            .I3(n44525), .O(n101[16])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2282_add_4_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_2282_add_4_18 (.CI(n44525), .I0(GND_net), .I1(pwm_counter[16]), 
            .CO(n44526));
    SB_LUT4 pwm_counter_2282_add_4_17_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[15]), 
            .I3(n44524), .O(n101[15])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2282_add_4_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_2282_add_4_17 (.CI(n44524), .I0(GND_net), .I1(pwm_counter[15]), 
            .CO(n44525));
    SB_LUT4 pwm_counter_2282_add_4_16_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[14]), 
            .I3(n44523), .O(n101[14])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2282_add_4_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_2282_add_4_16 (.CI(n44523), .I0(GND_net), .I1(pwm_counter[14]), 
            .CO(n44524));
    SB_LUT4 pwm_counter_2282_add_4_15_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[13]), 
            .I3(n44522), .O(n101[13])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2282_add_4_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_2282_add_4_15 (.CI(n44522), .I0(GND_net), .I1(pwm_counter[13]), 
            .CO(n44523));
    SB_LUT4 pwm_counter_2282_add_4_14_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[12]), 
            .I3(n44521), .O(n101[12])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2282_add_4_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_2282_add_4_14 (.CI(n44521), .I0(GND_net), .I1(pwm_counter[12]), 
            .CO(n44522));
    SB_LUT4 pwm_counter_2282_add_4_13_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[11]), 
            .I3(n44520), .O(n101[11])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2282_add_4_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_2282_add_4_13 (.CI(n44520), .I0(GND_net), .I1(pwm_counter[11]), 
            .CO(n44521));
    SB_LUT4 pwm_counter_2282_add_4_12_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[10]), 
            .I3(n44519), .O(n101[10])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2282_add_4_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_2282_add_4_12 (.CI(n44519), .I0(GND_net), .I1(pwm_counter[10]), 
            .CO(n44520));
    SB_LUT4 pwm_counter_2282_add_4_11_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[9]), 
            .I3(n44518), .O(n101[9])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2282_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_2282_add_4_11 (.CI(n44518), .I0(GND_net), .I1(pwm_counter[9]), 
            .CO(n44519));
    SB_LUT4 pwm_counter_2282_add_4_10_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[8]), 
            .I3(n44517), .O(n101[8])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2282_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_2282_add_4_10 (.CI(n44517), .I0(GND_net), .I1(pwm_counter[8]), 
            .CO(n44518));
    SB_LUT4 pwm_counter_2282_add_4_9_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[7]), 
            .I3(n44516), .O(n101[7])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2282_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_2282_add_4_9 (.CI(n44516), .I0(GND_net), .I1(pwm_counter[7]), 
            .CO(n44517));
    SB_LUT4 pwm_counter_2282_add_4_8_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[6]), 
            .I3(n44515), .O(n101[6])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2282_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_2282_add_4_8 (.CI(n44515), .I0(GND_net), .I1(pwm_counter[6]), 
            .CO(n44516));
    SB_LUT4 pwm_counter_2282_add_4_7_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[5]), 
            .I3(n44514), .O(n101[5])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2282_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_2282_add_4_7 (.CI(n44514), .I0(GND_net), .I1(pwm_counter[5]), 
            .CO(n44515));
    SB_LUT4 pwm_counter_2282_add_4_6_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[4]), 
            .I3(n44513), .O(n101[4])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2282_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_2282_add_4_6 (.CI(n44513), .I0(GND_net), .I1(pwm_counter[4]), 
            .CO(n44514));
    SB_LUT4 pwm_counter_2282_add_4_5_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[3]), 
            .I3(n44512), .O(n101[3])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2282_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_2282_add_4_5 (.CI(n44512), .I0(GND_net), .I1(pwm_counter[3]), 
            .CO(n44513));
    SB_LUT4 pwm_counter_2282_add_4_4_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[2]), 
            .I3(n44511), .O(n101[2])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2282_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_2282_add_4_4 (.CI(n44511), .I0(GND_net), .I1(pwm_counter[2]), 
            .CO(n44512));
    SB_LUT4 pwm_counter_2282_add_4_3_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[1]), 
            .I3(n44510), .O(n101[1])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2282_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_2282_add_4_3 (.CI(n44510), .I0(GND_net), .I1(pwm_counter[1]), 
            .CO(n44511));
    SB_LUT4 pwm_counter_2282_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[0]), 
            .I3(VCC_net), .O(n101[0])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2282_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_2282_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(pwm_counter[0]), 
            .CO(n44510));
    SB_DFFSR pwm_counter_2282__i0 (.Q(pwm_counter[0]), .C(clk32MHz), .D(n101[0]), 
            .R(pwm_counter_23__N_906));   // verilog/pwm.v(17[20:33])
    SB_LUT4 duty_23__I_0_i8_3_lut_3_lut (.I0(pwm_setpoint[4]), .I1(pwm_setpoint[8]), 
            .I2(pwm_counter[8]), .I3(GND_net), .O(n8));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i8_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i39107_2_lut_4_lut (.I0(pwm_counter[21]), .I1(pwm_setpoint[21]), 
            .I2(pwm_counter[9]), .I3(pwm_setpoint[9]), .O(n54937));
    defparam i39107_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 duty_23__I_0_i16_3_lut_3_lut (.I0(pwm_setpoint[9]), .I1(pwm_setpoint[21]), 
            .I2(pwm_counter[21]), .I3(GND_net), .O(n16));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i16_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i39141_3_lut_4_lut (.I0(pwm_counter[3]), .I1(pwm_setpoint[3]), 
            .I2(pwm_setpoint[2]), .I3(pwm_counter[2]), .O(n54971));   // verilog/pwm.v(21[8:24])
    defparam i39141_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 duty_23__I_0_i6_3_lut_3_lut (.I0(pwm_counter[3]), .I1(pwm_setpoint[3]), 
            .I2(pwm_setpoint[2]), .I3(GND_net), .O(n6));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 duty_23__I_0_i10_3_lut_3_lut (.I0(pwm_setpoint[5]), .I1(pwm_setpoint[6]), 
            .I2(pwm_counter[6]), .I3(GND_net), .O(n10));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i10_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i39118_2_lut_4_lut (.I0(pwm_counter[16]), .I1(pwm_setpoint[16]), 
            .I2(pwm_counter[7]), .I3(pwm_setpoint[7]), .O(n54948));
    defparam i39118_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 duty_23__I_0_i12_3_lut_3_lut (.I0(pwm_setpoint[7]), .I1(pwm_setpoint[16]), 
            .I2(pwm_counter[16]), .I3(GND_net), .O(n12));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i12_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 duty_23__I_0_i41_2_lut (.I0(pwm_counter[20]), .I1(pwm_setpoint[20]), 
            .I2(GND_net), .I3(GND_net), .O(n41));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i39_2_lut (.I0(pwm_counter[19]), .I1(pwm_setpoint[19]), 
            .I2(GND_net), .I3(GND_net), .O(n39));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i45_2_lut (.I0(pwm_counter[22]), .I1(pwm_setpoint[22]), 
            .I2(GND_net), .I3(GND_net), .O(n45));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i45_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i37_2_lut (.I0(pwm_counter[18]), .I1(pwm_setpoint[18]), 
            .I2(GND_net), .I3(GND_net), .O(n37));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i43_2_lut (.I0(pwm_counter[21]), .I1(pwm_setpoint[21]), 
            .I2(GND_net), .I3(GND_net), .O(n43));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i29_2_lut (.I0(pwm_counter[14]), .I1(pwm_setpoint[14]), 
            .I2(GND_net), .I3(GND_net), .O(n29));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i31_2_lut (.I0(pwm_counter[15]), .I1(pwm_setpoint[15]), 
            .I2(GND_net), .I3(GND_net), .O(n31));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i23_2_lut (.I0(pwm_counter[11]), .I1(pwm_setpoint[11]), 
            .I2(GND_net), .I3(GND_net), .O(n23));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i25_2_lut (.I0(pwm_counter[12]), .I1(pwm_setpoint[12]), 
            .I2(GND_net), .I3(GND_net), .O(n25));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i35_2_lut (.I0(pwm_counter[17]), .I1(pwm_setpoint[17]), 
            .I2(GND_net), .I3(GND_net), .O(n35));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i33_2_lut (.I0(pwm_counter[16]), .I1(pwm_setpoint[16]), 
            .I2(GND_net), .I3(GND_net), .O(n33));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i11_2_lut (.I0(pwm_counter[5]), .I1(pwm_setpoint[5]), 
            .I2(GND_net), .I3(GND_net), .O(n11));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i13_2_lut (.I0(pwm_counter[6]), .I1(pwm_setpoint[6]), 
            .I2(GND_net), .I3(GND_net), .O(n13));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i15_2_lut (.I0(pwm_counter[7]), .I1(pwm_setpoint[7]), 
            .I2(GND_net), .I3(GND_net), .O(n15));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i27_2_lut (.I0(pwm_counter[13]), .I1(pwm_setpoint[13]), 
            .I2(GND_net), .I3(GND_net), .O(n27));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i9_2_lut (.I0(pwm_counter[4]), .I1(pwm_setpoint[4]), 
            .I2(GND_net), .I3(GND_net), .O(n9));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i17_2_lut (.I0(pwm_counter[8]), .I1(pwm_setpoint[8]), 
            .I2(GND_net), .I3(GND_net), .O(n17));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i19_2_lut (.I0(pwm_counter[9]), .I1(pwm_setpoint[9]), 
            .I2(GND_net), .I3(GND_net), .O(n19));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i21_2_lut (.I0(pwm_counter[10]), .I1(pwm_setpoint[10]), 
            .I2(GND_net), .I3(GND_net), .O(n21));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i39130_4_lut (.I0(n21), .I1(n19), .I2(n17), .I3(n9), .O(n54960));
    defparam i39130_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i39124_4_lut (.I0(n27), .I1(n15), .I2(n13), .I3(n11), .O(n54954));
    defparam i39124_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 duty_23__I_0_i30_3_lut (.I0(n12), .I1(pwm_setpoint[17]), .I2(n35), 
            .I3(GND_net), .O(n30));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i39512_4_lut (.I0(n13), .I1(n11), .I2(n9), .I3(n54971), 
            .O(n55343));
    defparam i39512_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i39508_4_lut (.I0(n19), .I1(n17), .I2(n15), .I3(n55343), 
            .O(n55339));
    defparam i39508_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i39933_4_lut (.I0(n25), .I1(n23), .I2(n21), .I3(n55339), 
            .O(n55764));
    defparam i39933_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i39697_4_lut (.I0(n31), .I1(n29), .I2(n27), .I3(n55764), 
            .O(n55528));
    defparam i39697_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i39973_4_lut (.I0(n37), .I1(n35), .I2(n33), .I3(n55528), 
            .O(n55804));
    defparam i39973_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i39767_3_lut (.I0(n6), .I1(pwm_setpoint[10]), .I2(n21), .I3(GND_net), 
            .O(n55598));   // verilog/pwm.v(21[8:24])
    defparam i39767_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i39768_3_lut (.I0(n55598), .I1(pwm_setpoint[11]), .I2(n23), 
            .I3(GND_net), .O(n55599));   // verilog/pwm.v(21[8:24])
    defparam i39768_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i24_3_lut (.I0(n16), .I1(pwm_setpoint[22]), .I2(n45), 
            .I3(GND_net), .O(n24));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i39109_4_lut (.I0(n43), .I1(n25), .I2(n23), .I3(n54960), 
            .O(n54939));
    defparam i39109_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i39625_4_lut (.I0(n24), .I1(n8), .I2(n45), .I3(n54937), 
            .O(n55456));   // verilog/pwm.v(21[8:24])
    defparam i39625_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i39336_3_lut (.I0(n55599), .I1(pwm_setpoint[12]), .I2(n25), 
            .I3(GND_net), .O(n55167));   // verilog/pwm.v(21[8:24])
    defparam i39336_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i4_4_lut (.I0(pwm_counter[0]), .I1(pwm_setpoint[1]), 
            .I2(pwm_counter[1]), .I3(pwm_setpoint[0]), .O(n4));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i4_4_lut.LUT_INIT = 16'h4d0c;
    SB_LUT4 i39765_3_lut (.I0(n4), .I1(pwm_setpoint[13]), .I2(n27), .I3(GND_net), 
            .O(n55596));   // verilog/pwm.v(21[8:24])
    defparam i39765_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i39766_3_lut (.I0(n55596), .I1(pwm_setpoint[14]), .I2(n29), 
            .I3(GND_net), .O(n55597));   // verilog/pwm.v(21[8:24])
    defparam i39766_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i39120_4_lut (.I0(n33), .I1(n31), .I2(n29), .I3(n54954), 
            .O(n54950));
    defparam i39120_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i39943_4_lut (.I0(n30), .I1(n10), .I2(n35), .I3(n54948), 
            .O(n55774));   // verilog/pwm.v(21[8:24])
    defparam i39943_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i39338_3_lut (.I0(n55597), .I1(pwm_setpoint[15]), .I2(n31), 
            .I3(GND_net), .O(n55169));   // verilog/pwm.v(21[8:24])
    defparam i39338_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i40027_4_lut (.I0(n55169), .I1(n55774), .I2(n35), .I3(n54950), 
            .O(n55858));   // verilog/pwm.v(21[8:24])
    defparam i40027_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i40028_3_lut (.I0(n55858), .I1(pwm_setpoint[18]), .I2(n37), 
            .I3(GND_net), .O(n55859));   // verilog/pwm.v(21[8:24])
    defparam i40028_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i40002_3_lut (.I0(n55859), .I1(pwm_setpoint[19]), .I2(n39), 
            .I3(GND_net), .O(n55833));   // verilog/pwm.v(21[8:24])
    defparam i40002_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i39111_4_lut (.I0(n43), .I1(n41), .I2(n39), .I3(n55804), 
            .O(n54941));
    defparam i39111_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i39877_4_lut (.I0(n55167), .I1(n55456), .I2(n45), .I3(n54939), 
            .O(n55708));   // verilog/pwm.v(21[8:24])
    defparam i39877_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i39344_3_lut (.I0(n55833), .I1(pwm_setpoint[20]), .I2(n41), 
            .I3(GND_net), .O(n55175));   // verilog/pwm.v(21[8:24])
    defparam i39344_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i39961_4_lut (.I0(n55175), .I1(n55708), .I2(n45), .I3(n54941), 
            .O(n55792));   // verilog/pwm.v(21[8:24])
    defparam i39961_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i39962_3_lut (.I0(n55792), .I1(pwm_counter[23]), .I2(pwm_setpoint[23]), 
            .I3(GND_net), .O(pwm_out_N_908));   // verilog/pwm.v(21[8:24])
    defparam i39962_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i2_3_lut (.I0(pwm_counter[6]), .I1(pwm_counter[8]), .I2(pwm_counter[7]), 
            .I3(GND_net), .O(n51426));
    defparam i2_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i9_4_lut (.I0(pwm_counter[17]), .I1(pwm_counter[18]), .I2(pwm_counter[13]), 
            .I3(pwm_counter[16]), .O(n22));
    defparam i9_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_4_lut (.I0(n51426), .I1(pwm_counter[22]), .I2(pwm_counter[10]), 
            .I3(pwm_counter[9]), .O(n15_adj_4614));
    defparam i2_4_lut.LUT_INIT = 16'heccc;
    SB_LUT4 i7_3_lut (.I0(pwm_counter[20]), .I1(pwm_counter[21]), .I2(pwm_counter[11]), 
            .I3(GND_net), .O(n20));
    defparam i7_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i11_4_lut (.I0(n15_adj_4614), .I1(n22), .I2(pwm_counter[15]), 
            .I3(pwm_counter[14]), .O(n24_adj_4615));
    defparam i11_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i6_2_lut (.I0(pwm_counter[19]), .I1(pwm_counter[12]), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_4616));
    defparam i6_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i40781_4_lut (.I0(pwm_counter[23]), .I1(n19_adj_4616), .I2(n24_adj_4615), 
            .I3(n20), .O(pwm_counter_23__N_906));   // verilog/pwm.v(18[8:40])
    defparam i40781_4_lut.LUT_INIT = 16'h5554;
    
endmodule
//
// Verilog Description of module TLI4970
//

module TLI4970 (\state[0] , GND_net, \data[12] , n5, \state[1] , \data[15] , 
            n28729, clk16MHz, VCC_net, n15, n5_adj_1, n36554, n36528, 
            n6, n30067, n30066, \data[11] , n30059, \data[10] , 
            n29407, n9, clk_out, n29398, CS_c, n29391, \current[0] , 
            \current[15] , n7, n29916, \data[9] , n29892, \data[8] , 
            n29891, \current[1] , n29890, \current[2] , n29889, \current[3] , 
            n29888, \current[4] , n29887, \current[5] , n29886, \current[6] , 
            n29885, \current[7] , n29884, \current[8] , n29883, \current[9] , 
            n29882, \current[10] , n29881, \current[11] , n29879, 
            \data[7] , n29876, \data[6] , n29869, \data[5] , n29850, 
            \data[0] , n29839, \data[4] , n29838, \data[3] , n29823, 
            \data[2] , n29758, \data[1] , CS_CLK_c, n27258, n27271, 
            n27232, n27198, n6_adj_2, n5_adj_3, n27264, state_7__N_4499) /* synthesis syn_noprune=1, syn_module_defined=1 */ ;
    output \state[0] ;
    input GND_net;
    output \data[12] ;
    output n5;
    output \state[1] ;
    output \data[15] ;
    output n28729;
    input clk16MHz;
    input VCC_net;
    output n15;
    output n5_adj_1;
    output n36554;
    output n36528;
    output n6;
    input n30067;
    input n30066;
    output \data[11] ;
    input n30059;
    output \data[10] ;
    input n29407;
    input n9;
    output clk_out;
    input n29398;
    output CS_c;
    input n29391;
    output \current[0] ;
    output \current[15] ;
    output n7;
    input n29916;
    output \data[9] ;
    input n29892;
    output \data[8] ;
    input n29891;
    output \current[1] ;
    input n29890;
    output \current[2] ;
    input n29889;
    output \current[3] ;
    input n29888;
    output \current[4] ;
    input n29887;
    output \current[5] ;
    input n29886;
    output \current[6] ;
    input n29885;
    output \current[7] ;
    input n29884;
    output \current[8] ;
    input n29883;
    output \current[9] ;
    input n29882;
    output \current[10] ;
    input n29881;
    output \current[11] ;
    input n29879;
    output \data[7] ;
    input n29876;
    output \data[6] ;
    input n29869;
    output \data[5] ;
    input n29850;
    output \data[0] ;
    input n29839;
    output \data[4] ;
    input n29838;
    output \data[3] ;
    input n29823;
    output \data[2] ;
    input n29758;
    output \data[1] ;
    output CS_CLK_c;
    output n27258;
    output n27271;
    output n27232;
    output n27198;
    output n6_adj_2;
    output n5_adj_3;
    output n27264;
    output state_7__N_4499;
    
    wire clk_slow /* synthesis is_clock=1, SET_AS_NETWORK=\tli/clk_slow */ ;   // verilog/tli4970.v(11[7:15])
    wire clk16MHz /* synthesis SET_AS_NETWORK=clk16MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    
    wire n7796;
    wire [13:0]n241;
    wire [7:0]counter;   // verilog/tli4970.v(12[13:20])
    
    wire clk_slow_N_4413;
    wire [7:0]bit_counter;   // verilog/tli4970.v(26[13:24])
    
    wire clk_slow_N_4412, n54587, n24130;
    wire [2:0]n17;
    
    wire n44607, n44606;
    wire [11:0]n53;
    wire [15:0]delay_counter;   // verilog/tli4970.v(28[14:27])
    
    wire n44605, n44604, n44603, n44602, n44601, n44600, n44599, 
        n44598, n44597, n44596, n44595, n36977;
    wire [7:0]n37;
    
    wire n28797, n29175, n10895, n28875, n29156, n24107, n24109, 
        n24111, delay_counter_15__N_4494, n44665, n44664, n44663, 
        n44662, n54546, n44661, n54538, n44660, n54537, n44659, 
        n6_adj_4613, n8, n12, n10;
    
    SB_LUT4 i2151_1_lut (.I0(\state[0] ), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n7796));   // verilog/tli4970.v(35[10] 68[6])
    defparam i2151_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i2416_1_lut (.I0(\data[12] ), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n241[13]));
    defparam i2416_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i2388_3_lut (.I0(counter[0]), .I1(counter[2]), .I2(counter[1]), 
            .I3(GND_net), .O(clk_slow_N_4413));
    defparam i2388_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 equal_358_i5_2_lut (.I0(bit_counter[0]), .I1(bit_counter[1]), 
            .I2(GND_net), .I3(GND_net), .O(n5));   // verilog/tli4970.v(54[9:26])
    defparam equal_358_i5_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 clk_slow_I_0_72_2_lut (.I0(clk_slow), .I1(clk_slow_N_4413), 
            .I2(GND_net), .I3(GND_net), .O(clk_slow_N_4412));   // verilog/tli4970.v(15[5] 18[8])
    defparam clk_slow_I_0_72_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i10080_3_lut (.I0(\state[0] ), .I1(n54587), .I2(\state[1] ), 
            .I3(GND_net), .O(n24130));   // verilog/tli4970.v(55[24:39])
    defparam i10080_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i40088_3_lut (.I0(\data[15] ), .I1(\state[1] ), .I2(\state[0] ), 
            .I3(GND_net), .O(n28729));
    defparam i40088_3_lut.LUT_INIT = 16'h4040;
    SB_DFF clk_slow_63 (.Q(clk_slow), .C(clk16MHz), .D(clk_slow_N_4412));   // verilog/tli4970.v(13[10] 19[6])
    SB_LUT4 counter_2287_2288_add_4_4_lut (.I0(GND_net), .I1(GND_net), .I2(counter[2]), 
            .I3(n44607), .O(n17[2])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2287_2288_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 counter_2287_2288_add_4_3_lut (.I0(GND_net), .I1(GND_net), .I2(counter[1]), 
            .I3(n44606), .O(n17[1])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2287_2288_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_2287_2288_add_4_3 (.CI(n44606), .I0(GND_net), .I1(counter[1]), 
            .CO(n44607));
    SB_LUT4 counter_2287_2288_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(counter[0]), 
            .I3(VCC_net), .O(n17[0])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2287_2288_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_2287_2288_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(counter[0]), 
            .CO(n44606));
    SB_LUT4 delay_counter_2285_2286_add_4_13_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[11]), .I3(n44605), .O(n53[11])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_2285_2286_add_4_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 delay_counter_2285_2286_add_4_12_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[10]), .I3(n44604), .O(n53[10])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_2285_2286_add_4_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_2285_2286_add_4_12 (.CI(n44604), .I0(GND_net), 
            .I1(delay_counter[10]), .CO(n44605));
    SB_LUT4 delay_counter_2285_2286_add_4_11_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[9]), .I3(n44603), .O(n53[9])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_2285_2286_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_2285_2286_add_4_11 (.CI(n44603), .I0(GND_net), 
            .I1(delay_counter[9]), .CO(n44604));
    SB_LUT4 delay_counter_2285_2286_add_4_10_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[8]), .I3(n44602), .O(n53[8])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_2285_2286_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_2285_2286_add_4_10 (.CI(n44602), .I0(GND_net), 
            .I1(delay_counter[8]), .CO(n44603));
    SB_LUT4 delay_counter_2285_2286_add_4_9_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[7]), .I3(n44601), .O(n53[7])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_2285_2286_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_2285_2286_add_4_9 (.CI(n44601), .I0(GND_net), 
            .I1(delay_counter[7]), .CO(n44602));
    SB_LUT4 delay_counter_2285_2286_add_4_8_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[6]), .I3(n44600), .O(n53[6])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_2285_2286_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_2285_2286_add_4_8 (.CI(n44600), .I0(GND_net), 
            .I1(delay_counter[6]), .CO(n44601));
    SB_LUT4 delay_counter_2285_2286_add_4_7_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[5]), .I3(n44599), .O(n53[5])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_2285_2286_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_2285_2286_add_4_7 (.CI(n44599), .I0(GND_net), 
            .I1(delay_counter[5]), .CO(n44600));
    SB_LUT4 delay_counter_2285_2286_add_4_6_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[4]), .I3(n44598), .O(n53[4])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_2285_2286_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_2285_2286_add_4_6 (.CI(n44598), .I0(GND_net), 
            .I1(delay_counter[4]), .CO(n44599));
    SB_LUT4 delay_counter_2285_2286_add_4_5_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[3]), .I3(n44597), .O(n53[3])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_2285_2286_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_2285_2286_add_4_5 (.CI(n44597), .I0(GND_net), 
            .I1(delay_counter[3]), .CO(n44598));
    SB_LUT4 delay_counter_2285_2286_add_4_4_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[2]), .I3(n44596), .O(n53[2])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_2285_2286_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_2285_2286_add_4_4 (.CI(n44596), .I0(GND_net), 
            .I1(delay_counter[2]), .CO(n44597));
    SB_LUT4 delay_counter_2285_2286_add_4_3_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[1]), .I3(n44595), .O(n53[1])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_2285_2286_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_2285_2286_add_4_3 (.CI(n44595), .I0(GND_net), 
            .I1(delay_counter[1]), .CO(n44596));
    SB_LUT4 delay_counter_2285_2286_add_4_2_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[0]), .I3(VCC_net), .O(n53[0])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_2285_2286_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_2285_2286_add_4_2 (.CI(VCC_net), .I0(GND_net), 
            .I1(delay_counter[0]), .CO(n44595));
    SB_LUT4 i40658_2_lut (.I0(n15), .I1(\state[0] ), .I2(GND_net), .I3(GND_net), 
            .O(n36977));
    defparam i40658_2_lut.LUT_INIT = 16'h1111;
    SB_DFFNESR bit_counter_2296__i4 (.Q(bit_counter[4]), .C(clk_slow), .E(n28797), 
            .D(n37[4]), .R(n29175));   // verilog/tli4970.v(55[24:39])
    SB_DFFNESR bit_counter_2296__i5 (.Q(bit_counter[5]), .C(clk_slow), .E(n28797), 
            .D(n37[5]), .R(n29175));   // verilog/tli4970.v(55[24:39])
    SB_DFFNESR bit_counter_2296__i6 (.Q(bit_counter[6]), .C(clk_slow), .E(n28797), 
            .D(n37[6]), .R(n29175));   // verilog/tli4970.v(55[24:39])
    SB_LUT4 equal_361_i5_2_lut (.I0(bit_counter[0]), .I1(bit_counter[1]), 
            .I2(GND_net), .I3(GND_net), .O(n5_adj_1));   // verilog/tli4970.v(54[9:26])
    defparam equal_361_i5_2_lut.LUT_INIT = 16'hbbbb;
    SB_DFFNESR bit_counter_2296__i7 (.Q(bit_counter[7]), .C(clk_slow), .E(n28797), 
            .D(n37[7]), .R(n29175));   // verilog/tli4970.v(55[24:39])
    SB_LUT4 i22490_2_lut (.I0(bit_counter[0]), .I1(bit_counter[1]), .I2(GND_net), 
            .I3(GND_net), .O(n36554));
    defparam i22490_2_lut.LUT_INIT = 16'h8888;
    SB_DFFNESR state_i1 (.Q(\state[1] ), .C(clk_slow), .E(n28875), .D(n10895), 
            .R(n29156));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFNE bit_counter_2296__i3 (.Q(bit_counter[3]), .C(clk_slow), .E(n28797), 
            .D(n24107));   // verilog/tli4970.v(55[24:39])
    SB_LUT4 i22464_2_lut (.I0(bit_counter[2]), .I1(bit_counter[3]), .I2(GND_net), 
            .I3(GND_net), .O(n36528));
    defparam i22464_2_lut.LUT_INIT = 16'h8888;
    SB_DFFNE bit_counter_2296__i2 (.Q(bit_counter[2]), .C(clk_slow), .E(n28797), 
            .D(n24109));   // verilog/tli4970.v(55[24:39])
    SB_DFFNE bit_counter_2296__i1 (.Q(bit_counter[1]), .C(clk_slow), .E(n28797), 
            .D(n24111));   // verilog/tli4970.v(55[24:39])
    SB_DFFSR counter_2287_2288__i3 (.Q(counter[2]), .C(clk16MHz), .D(n17[2]), 
            .R(clk_slow_N_4413));   // verilog/tli4970.v(14[16:27])
    SB_DFFSR counter_2287_2288__i2 (.Q(counter[1]), .C(clk16MHz), .D(n17[1]), 
            .R(clk_slow_N_4413));   // verilog/tli4970.v(14[16:27])
    SB_DFFNSR delay_counter_2285_2286__i12 (.Q(delay_counter[11]), .C(clk_slow), 
            .D(n53[11]), .R(delay_counter_15__N_4494));   // verilog/tli4970.v(40[24:39])
    SB_DFFNSR delay_counter_2285_2286__i11 (.Q(delay_counter[10]), .C(clk_slow), 
            .D(n53[10]), .R(delay_counter_15__N_4494));   // verilog/tli4970.v(40[24:39])
    SB_DFFNSR delay_counter_2285_2286__i10 (.Q(delay_counter[9]), .C(clk_slow), 
            .D(n53[9]), .R(delay_counter_15__N_4494));   // verilog/tli4970.v(40[24:39])
    SB_DFFNSR delay_counter_2285_2286__i9 (.Q(delay_counter[8]), .C(clk_slow), 
            .D(n53[8]), .R(delay_counter_15__N_4494));   // verilog/tli4970.v(40[24:39])
    SB_DFFNSR delay_counter_2285_2286__i8 (.Q(delay_counter[7]), .C(clk_slow), 
            .D(n53[7]), .R(delay_counter_15__N_4494));   // verilog/tli4970.v(40[24:39])
    SB_DFFNSR delay_counter_2285_2286__i7 (.Q(delay_counter[6]), .C(clk_slow), 
            .D(n53[6]), .R(delay_counter_15__N_4494));   // verilog/tli4970.v(40[24:39])
    SB_DFFNSR delay_counter_2285_2286__i6 (.Q(delay_counter[5]), .C(clk_slow), 
            .D(n53[5]), .R(delay_counter_15__N_4494));   // verilog/tli4970.v(40[24:39])
    SB_DFFNSR delay_counter_2285_2286__i5 (.Q(delay_counter[4]), .C(clk_slow), 
            .D(n53[4]), .R(delay_counter_15__N_4494));   // verilog/tli4970.v(40[24:39])
    SB_DFFNSR delay_counter_2285_2286__i4 (.Q(delay_counter[3]), .C(clk_slow), 
            .D(n53[3]), .R(delay_counter_15__N_4494));   // verilog/tli4970.v(40[24:39])
    SB_DFFNSR delay_counter_2285_2286__i3 (.Q(delay_counter[2]), .C(clk_slow), 
            .D(n53[2]), .R(delay_counter_15__N_4494));   // verilog/tli4970.v(40[24:39])
    SB_DFFNSR delay_counter_2285_2286__i2 (.Q(delay_counter[1]), .C(clk_slow), 
            .D(n53[1]), .R(delay_counter_15__N_4494));   // verilog/tli4970.v(40[24:39])
    SB_LUT4 equal_364_i6_2_lut (.I0(bit_counter[2]), .I1(bit_counter[3]), 
            .I2(GND_net), .I3(GND_net), .O(n6));   // verilog/tli4970.v(54[9:26])
    defparam equal_364_i6_2_lut.LUT_INIT = 16'hdddd;
    SB_DFFN data_i12 (.Q(\data[12] ), .C(clk_slow), .D(n30067));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i11 (.Q(\data[11] ), .C(clk_slow), .D(n30066));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i10 (.Q(\data[10] ), .C(clk_slow), .D(n30059));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFNESS state_i0 (.Q(\state[0] ), .C(clk_slow), .E(n28875), .D(n36977), 
            .S(n29156));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i15 (.Q(\data[15] ), .C(clk_slow), .D(n29407));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN clk_out_67 (.Q(clk_out), .C(clk_slow), .D(n9));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN slave_select_66 (.Q(CS_c), .C(clk_slow), .D(n29398));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i1 (.Q(\current[0] ), .C(clk_slow), .D(n29391));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFNSR delay_counter_2285_2286__i1 (.Q(delay_counter[0]), .C(clk_slow), 
            .D(n53[0]), .R(delay_counter_15__N_4494));   // verilog/tli4970.v(40[24:39])
    SB_DFFSR counter_2287_2288__i1 (.Q(counter[0]), .C(clk16MHz), .D(n17[0]), 
            .R(clk_slow_N_4413));   // verilog/tli4970.v(14[16:27])
    SB_DFFNE bit_counter_2296__i0 (.Q(bit_counter[0]), .C(clk_slow), .E(n28797), 
            .D(n24130));   // verilog/tli4970.v(55[24:39])
    SB_DFFNE current__i13 (.Q(\current[15] ), .C(clk_slow), .E(n28729), 
            .D(n241[13]));   // verilog/tli4970.v(35[10] 68[6])
    SB_LUT4 i15096_2_lut_2_lut (.I0(\state[1] ), .I1(\state[0] ), .I2(GND_net), 
            .I3(GND_net), .O(n29175));   // verilog/tli4970.v(55[24:39])
    defparam i15096_2_lut_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 equal_371_i7_2_lut_4_lut (.I0(bit_counter[0]), .I1(bit_counter[1]), 
            .I2(bit_counter[2]), .I3(bit_counter[3]), .O(n7));   // verilog/tli4970.v(54[9:26])
    defparam equal_371_i7_2_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_DFFN data_i9 (.Q(\data[9] ), .C(clk_slow), .D(n29916));   // verilog/tli4970.v(35[10] 68[6])
    SB_LUT4 i1_2_lut_4_lut (.I0(n15), .I1(\state[1] ), .I2(\state[0] ), 
            .I3(delay_counter_15__N_4494), .O(n28875));
    defparam i1_2_lut_4_lut.LUT_INIT = 16'hfff4;
    SB_LUT4 i15076_2_lut_4_lut (.I0(n15), .I1(\state[1] ), .I2(\state[0] ), 
            .I3(delay_counter_15__N_4494), .O(n29156));
    defparam i15076_2_lut_4_lut.LUT_INIT = 16'h0b00;
    SB_DFFN data_i8 (.Q(\data[8] ), .C(clk_slow), .D(n29892));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i2 (.Q(\current[1] ), .C(clk_slow), .D(n29891));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i3 (.Q(\current[2] ), .C(clk_slow), .D(n29890));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i4 (.Q(\current[3] ), .C(clk_slow), .D(n29889));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i5 (.Q(\current[4] ), .C(clk_slow), .D(n29888));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i6 (.Q(\current[5] ), .C(clk_slow), .D(n29887));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i7 (.Q(\current[6] ), .C(clk_slow), .D(n29886));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i8 (.Q(\current[7] ), .C(clk_slow), .D(n29885));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i9 (.Q(\current[8] ), .C(clk_slow), .D(n29884));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i10 (.Q(\current[9] ), .C(clk_slow), .D(n29883));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i11 (.Q(\current[10] ), .C(clk_slow), .D(n29882));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i12 (.Q(\current[11] ), .C(clk_slow), .D(n29881));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i7 (.Q(\data[7] ), .C(clk_slow), .D(n29879));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i6 (.Q(\data[6] ), .C(clk_slow), .D(n29876));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i5 (.Q(\data[5] ), .C(clk_slow), .D(n29869));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i0 (.Q(\data[0] ), .C(clk_slow), .D(n29850));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i4 (.Q(\data[4] ), .C(clk_slow), .D(n29839));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i3 (.Q(\data[3] ), .C(clk_slow), .D(n29838));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i2 (.Q(\data[2] ), .C(clk_slow), .D(n29823));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i1 (.Q(\data[1] ), .C(clk_slow), .D(n29758));   // verilog/tli4970.v(35[10] 68[6])
    SB_LUT4 bit_counter_2296_add_4_9_lut (.I0(GND_net), .I1(VCC_net), .I2(bit_counter[7]), 
            .I3(n44665), .O(n37[7])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_counter_2296_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 bit_counter_2296_add_4_8_lut (.I0(GND_net), .I1(VCC_net), .I2(bit_counter[6]), 
            .I3(n44664), .O(n37[6])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_counter_2296_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY bit_counter_2296_add_4_8 (.CI(n44664), .I0(VCC_net), .I1(bit_counter[6]), 
            .CO(n44665));
    SB_LUT4 bit_counter_2296_add_4_7_lut (.I0(GND_net), .I1(VCC_net), .I2(bit_counter[5]), 
            .I3(n44663), .O(n37[5])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_counter_2296_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY bit_counter_2296_add_4_7 (.CI(n44663), .I0(VCC_net), .I1(bit_counter[5]), 
            .CO(n44664));
    SB_LUT4 bit_counter_2296_add_4_6_lut (.I0(GND_net), .I1(VCC_net), .I2(bit_counter[4]), 
            .I3(n44662), .O(n37[4])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_counter_2296_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY bit_counter_2296_add_4_6 (.CI(n44662), .I0(VCC_net), .I1(bit_counter[4]), 
            .CO(n44663));
    SB_LUT4 bit_counter_2296_add_4_5_lut (.I0(n7796), .I1(VCC_net), .I2(bit_counter[3]), 
            .I3(n44661), .O(n54546)) /* synthesis syn_instantiated=1 */ ;
    defparam bit_counter_2296_add_4_5_lut.LUT_INIT = 16'h8228;
    SB_CARRY bit_counter_2296_add_4_5 (.CI(n44661), .I0(VCC_net), .I1(bit_counter[3]), 
            .CO(n44662));
    SB_LUT4 bit_counter_2296_add_4_4_lut (.I0(n7796), .I1(VCC_net), .I2(bit_counter[2]), 
            .I3(n44660), .O(n54538)) /* synthesis syn_instantiated=1 */ ;
    defparam bit_counter_2296_add_4_4_lut.LUT_INIT = 16'h8228;
    SB_CARRY bit_counter_2296_add_4_4 (.CI(n44660), .I0(VCC_net), .I1(bit_counter[2]), 
            .CO(n44661));
    SB_LUT4 bit_counter_2296_add_4_3_lut (.I0(n7796), .I1(VCC_net), .I2(bit_counter[1]), 
            .I3(n44659), .O(n54537)) /* synthesis syn_instantiated=1 */ ;
    defparam bit_counter_2296_add_4_3_lut.LUT_INIT = 16'h8228;
    SB_CARRY bit_counter_2296_add_4_3 (.CI(n44659), .I0(VCC_net), .I1(bit_counter[1]), 
            .CO(n44660));
    SB_LUT4 bit_counter_2296_add_4_2_lut (.I0(n7796), .I1(GND_net), .I2(bit_counter[0]), 
            .I3(VCC_net), .O(n54587)) /* synthesis syn_instantiated=1 */ ;
    defparam bit_counter_2296_add_4_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY bit_counter_2296_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(bit_counter[0]), 
            .CO(n44659));
    SB_LUT4 spi_clk_I_0_i1_3_lut (.I0(clk_slow), .I1(clk_out), .I2(CS_c), 
            .I3(GND_net), .O(CS_CLK_c));   // verilog/tli4970.v(23[20:53])
    defparam spi_clk_I_0_i1_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i1_2_lut_4_lut_adj_946 (.I0(\state[0] ), .I1(\state[1] ), .I2(bit_counter[0]), 
            .I3(bit_counter[1]), .O(n27258));   // verilog/tli4970.v(43[5] 67[12])
    defparam i1_2_lut_4_lut_adj_946.LUT_INIT = 16'hfbff;
    SB_LUT4 i1_2_lut_4_lut_adj_947 (.I0(\state[0] ), .I1(\state[1] ), .I2(bit_counter[0]), 
            .I3(bit_counter[1]), .O(n27271));   // verilog/tli4970.v(43[5] 67[12])
    defparam i1_2_lut_4_lut_adj_947.LUT_INIT = 16'hffbf;
    SB_LUT4 i1_2_lut_4_lut_adj_948 (.I0(\state[0] ), .I1(\state[1] ), .I2(bit_counter[0]), 
            .I3(bit_counter[1]), .O(n27232));   // verilog/tli4970.v(43[5] 67[12])
    defparam i1_2_lut_4_lut_adj_948.LUT_INIT = 16'hfffb;
    SB_LUT4 i2_3_lut_4_lut (.I0(bit_counter[2]), .I1(bit_counter[3]), .I2(\state[0] ), 
            .I3(\state[1] ), .O(n27198));   // verilog/tli4970.v(43[5] 67[12])
    defparam i2_3_lut_4_lut.LUT_INIT = 16'hfbff;
    SB_LUT4 i10068_3_lut (.I0(\state[0] ), .I1(n54537), .I2(\state[1] ), 
            .I3(GND_net), .O(n24111));   // verilog/tli4970.v(55[24:39])
    defparam i10068_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10066_3_lut (.I0(\state[0] ), .I1(n54538), .I2(\state[1] ), 
            .I3(GND_net), .O(n24109));   // verilog/tli4970.v(55[24:39])
    defparam i10066_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10064_3_lut (.I0(\state[0] ), .I1(n54546), .I2(\state[1] ), 
            .I3(GND_net), .O(n24107));   // verilog/tli4970.v(55[24:39])
    defparam i10064_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 equal_371_i6_2_lut (.I0(bit_counter[2]), .I1(bit_counter[3]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_2));   // verilog/tli4970.v(54[9:26])
    defparam equal_371_i6_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 equal_363_i5_2_lut (.I0(bit_counter[0]), .I1(bit_counter[1]), 
            .I2(GND_net), .I3(GND_net), .O(n5_adj_3));   // verilog/tli4970.v(54[9:26])
    defparam equal_363_i5_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut (.I0(bit_counter[5]), .I1(bit_counter[4]), .I2(GND_net), 
            .I3(GND_net), .O(n6_adj_4613));   // verilog/tli4970.v(56[12:26])
    defparam i1_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i4_4_lut (.I0(bit_counter[6]), .I1(bit_counter[7]), .I2(n7), 
            .I3(n6_adj_4613), .O(n15));   // verilog/tli4970.v(56[12:26])
    defparam i4_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_4_lut_adj_949 (.I0(\state[0] ), .I1(\state[1] ), .I2(bit_counter[0]), 
            .I3(bit_counter[1]), .O(n27264));   // verilog/tli4970.v(43[5] 67[12])
    defparam i1_2_lut_4_lut_adj_949.LUT_INIT = 16'hbfff;
    SB_LUT4 i3_3_lut (.I0(delay_counter[1]), .I1(delay_counter[2]), .I2(delay_counter[4]), 
            .I3(GND_net), .O(n8));
    defparam i3_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i2389_4_lut (.I0(delay_counter[3]), .I1(delay_counter[5]), .I2(n8), 
            .I3(delay_counter[0]), .O(n12));
    defparam i2389_4_lut.LUT_INIT = 16'hccc8;
    SB_LUT4 i4_4_lut_adj_950 (.I0(delay_counter[11]), .I1(delay_counter[7]), 
            .I2(delay_counter[8]), .I3(delay_counter[9]), .O(n10));
    defparam i4_4_lut_adj_950.LUT_INIT = 16'h8000;
    SB_LUT4 i5_4_lut (.I0(delay_counter[10]), .I1(n10), .I2(n12), .I3(delay_counter[6]), 
            .O(delay_counter_15__N_4494));
    defparam i5_4_lut.LUT_INIT = 16'h8880;
    SB_LUT4 mux_2384_i2_3_lut (.I0(n15), .I1(\state[1] ), .I2(\state[0] ), 
            .I3(GND_net), .O(n10895));
    defparam mux_2384_i2_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 state_7__I_0_77_i9_2_lut (.I0(\state[0] ), .I1(\state[1] ), 
            .I2(GND_net), .I3(GND_net), .O(state_7__N_4499));   // verilog/tli4970.v(53[7:17])
    defparam state_7__I_0_77_i9_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 i14977_2_lut (.I0(\state[1] ), .I1(\state[0] ), .I2(GND_net), 
            .I3(GND_net), .O(n28797));
    defparam i14977_2_lut.LUT_INIT = 16'h6666;
    
endmodule
