// Verilog netlist produced by program LSE :  version Diamond Version 0.0.0
// Netlist written on Mon Feb 17 17:50:09 2020
//
// Verilog Description of module TinyFPGA_B
//

module TinyFPGA_B (CLK, LED, USBPU, ENCODER0_A, ENCODER0_B, ENCODER1_A, 
            ENCODER1_B, HALL1, HALL2, HALL3, FAULT_N, NEOPXL, DE, 
            TX, RX, CS_CLK, CS, CS_MISO, SCL, SDA, INLC, INHC, 
            INLB, INHB, INLA, INHA) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(2[8:18])
    input CLK;   // verilog/TinyFPGA_B.v(3[9:12])
    output LED;   // verilog/TinyFPGA_B.v(4[10:13])
    output USBPU;   // verilog/TinyFPGA_B.v(5[10:15])
    input ENCODER0_A;   // verilog/TinyFPGA_B.v(6[9:19])
    input ENCODER0_B;   // verilog/TinyFPGA_B.v(7[9:19])
    input ENCODER1_A;   // verilog/TinyFPGA_B.v(8[9:19])
    input ENCODER1_B;   // verilog/TinyFPGA_B.v(9[9:19])
    input HALL1 /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(10[9:14])
    input HALL2 /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(11[9:14])
    input HALL3 /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(12[9:14])
    input FAULT_N;   // verilog/TinyFPGA_B.v(13[9:16])
    output NEOPXL;   // verilog/TinyFPGA_B.v(14[10:16])
    output DE;   // verilog/TinyFPGA_B.v(15[10:12])
    output TX /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(16[10:12])
    input RX;   // verilog/TinyFPGA_B.v(17[9:11])
    output CS_CLK;   // verilog/TinyFPGA_B.v(18[10:16])
    output CS;   // verilog/TinyFPGA_B.v(19[10:12])
    input CS_MISO;   // verilog/TinyFPGA_B.v(20[9:16])
    inout SCL /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(21[9:12])
    inout SDA /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(22[9:12])
    output INLC;   // verilog/TinyFPGA_B.v(23[10:14])
    output INHC;   // verilog/TinyFPGA_B.v(24[10:14])
    output INLB;   // verilog/TinyFPGA_B.v(25[10:14])
    output INHB;   // verilog/TinyFPGA_B.v(26[10:14])
    output INLA;   // verilog/TinyFPGA_B.v(27[10:14])
    output INHA;   // verilog/TinyFPGA_B.v(28[10:14])
    
    wire CLK_c /* synthesis SET_AS_NETWORK=CLK_c, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(3[9:12])
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    
    wire GND_net, VCC_net, LED_c, ENCODER0_A_N, ENCODER0_B_N, ENCODER1_A_N, 
        ENCODER1_B_N, NEOPXL_c, DE_c, RX_c, CS_CLK_c, CS_c, CS_MISO_c, 
        INLC_c_0, INHC_c_0, INLB_c_0, INHB_c_0, INLA_c_0, INHA_c_0;
    wire [7:0]ID;   // verilog/TinyFPGA_B.v(39[11:13])
    wire [23:0]neopxl_color;   // verilog/TinyFPGA_B.v(41[13:25])
    
    wire hall1, hall2, hall3, pwm_out, dir, GHA, GHB, GHC;
    wire [23:0]pwm_setpoint;   // verilog/TinyFPGA_B.v(87[20:32])
    wire [23:0]duty;   // verilog/TinyFPGA_B.v(88[21:25])
    
    wire h1, h2, h3;
    wire [7:0]commutation_state;   // verilog/TinyFPGA_B.v(132[12:29])
    wire [7:0]commutation_state_prev;   // verilog/TinyFPGA_B.v(133[12:34])
    
    wire dti;
    wire [7:0]dti_counter;   // verilog/TinyFPGA_B.v(142[12:23])
    
    wire tx_o, tx_enable;
    wire [23:0]encoder0_position_scaled;   // verilog/TinyFPGA_B.v(239[21:45])
    wire [23:0]encoder1_position_scaled;   // verilog/TinyFPGA_B.v(241[21:45])
    wire [23:0]displacement;   // verilog/TinyFPGA_B.v(242[21:33])
    wire [23:0]setpoint;   // verilog/TinyFPGA_B.v(243[22:30])
    
    wire n50202;
    wire [23:0]Kp;   // verilog/TinyFPGA_B.v(244[22:24])
    wire [23:0]Ki;   // verilog/TinyFPGA_B.v(245[22:24])
    wire [7:0]control_mode;   // verilog/TinyFPGA_B.v(247[14:26])
    wire [23:0]PWMLimit;   // verilog/TinyFPGA_B.v(248[22:30])
    wire [23:0]IntegralLimit;   // verilog/TinyFPGA_B.v(249[22:35])
    
    wire n38535, n38883;
    wire [15:0]current;   // verilog/TinyFPGA_B.v(251[22:29])
    
    wire n38534;
    wire [15:0]current_limit;   // verilog/TinyFPGA_B.v(252[22:35])
    wire [23:0]motor_state;   // verilog/TinyFPGA_B.v(281[22:33])
    wire [7:0]data;   // verilog/TinyFPGA_B.v(344[14:18])
    
    wire data_ready, sda_out, sda_enable, scl, scl_enable;
    wire [31:0]delay_counter;   // verilog/TinyFPGA_B.v(368[11:24])
    
    wire read;
    wire [2:0]\ID_READOUT_FSM.state ;   // verilog/TinyFPGA_B.v(376[15:20])
    
    wire pwm_setpoint_23__N_239, n38882, n287, n34648, n321, n325, 
        n326, n327, n328, n329, n330, n331, n332, n333, n334, 
        n335, n336, n340, n341, n342, n343, n344, n345, n346, 
        n347, n348, n349, n350, n351, n352, n353, n354, n355, 
        n356, n357, n358, n359, n360, n361, n362, n363, n6, 
        n23, n50240, n17, n15, n6_adj_5242, n39053, n38881, n35468, 
        n38880, n38533, n35466;
    wire [23:0]pwm_setpoint_23__N_11;
    
    wire n4, n44933;
    wire [7:0]commutation_state_7__N_240;
    
    wire commutation_state_7__N_248, n29167;
    wire [31:0]encoder0_position;   // verilog/TinyFPGA_B.v(238[11:28])
    
    wire n39052, n38879, GHA_N_391, GLA_N_408, GHB_N_413, GLB_N_422, 
        GHC_N_427, GLC_N_436, dti_N_440, n29164, n29162, n29161, 
        n29160, RX_N_10, n1855;
    wire [31:0]motor_state_23__N_123;
    wire [32:0]encoder0_position_scaled_23__N_51;
    
    wire encoder1_position_scaled_23__N_303;
    wire [31:0]encoder1_position_scaled_23__N_75;
    wire [23:0]displacement_23__N_99;
    
    wire n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, 
        n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, 
        n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, 
        n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, 
        read_N_445, n1415, n50020, n38532, n38878, n38877, n38876, 
        n4_adj_5243, n38531, n15_adj_5244, n14, n38469, n38875, 
        n1896;
    wire [31:0]encoder1_position;   // verilog/TinyFPGA_B.v(240[11:28])
    
    wire n29159, n29158;
    wire [31:0]timer;   // verilog/neopixel.v(9[12:17])
    wire [3:0]state;   // verilog/neopixel.v(16[20:25])
    wire [31:0]\neo_pixel_transmitter.t0 ;   // verilog/neopixel.v(28[14:16])
    
    wire n35458, n38468, n39051, n38874, n623, n622, n621;
    wire [3:0]state_3__N_552;
    
    wire n44987, n51402, n51396, n51390, n51673, n51384, n51378, 
        n8, n50356, n4208, n29157, n29156, n39050, n38873, n39049, 
        n39048, n29155, n29154, n38872, n29153, n29152, n4_adj_5245, 
        n29151, n7494, n38871, n39047, n38870, n39046, n17_adj_5246, 
        n16, n39045, n38869, n38868, n4508, n4507, n4506, n4505, 
        n4504, n4503, n4502, n4501, n4500, n4499, n4498, n15_adj_5247, 
        n38867, n38866, n38865, n39044, n39043, n29150, n29149, 
        n43326, n29148, n38864, n39042, n35432, n29147, n29146, 
        n39041, n38863, n29145, n39040, n29144, n4_adj_5248, n29143, 
        n29142, n39039, n38862, n29141;
    wire [2:0]reg_B;   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(142[19:24])
    
    wire n39038, n11, n15_adj_5249, n2, n544, n543, n542, n541, 
        n540, n539, n538, n14_adj_5250, n15_adj_5251, n16_adj_5252, 
        n17_adj_5253, n18, n19, n20, n21, n22, n23_adj_5254, n24, 
        n29140, n29139, n3, n4_adj_5255, n5, n6_adj_5256, n7, 
        n8_adj_5257, n9, n10, n11_adj_5258, n12, n13, n14_adj_5259, 
        n15_adj_5260, n16_adj_5261, n17_adj_5262, n18_adj_5263, n19_adj_5264, 
        n20_adj_5265, n21_adj_5266, n22_adj_5267, n23_adj_5268, n24_adj_5269, 
        n25, n29138, n29137, n29136, n29135, rx_data_ready;
    wire [7:0]rx_data;   // verilog/coms.v(92[13:20])
    wire [7:0]\data_in[3] ;   // verilog/coms.v(96[12:19])
    wire [7:0]\data_in[2] ;   // verilog/coms.v(96[12:19])
    wire [7:0]\data_in[1] ;   // verilog/coms.v(96[12:19])
    wire [7:0]\data_in[0] ;   // verilog/coms.v(96[12:19])
    
    wire n39037, n39036, n39035, n39034, n38861, n38860;
    wire [7:0]\data_in_frame[22] ;   // verilog/coms.v(97[12:25])
    wire [7:0]\data_in_frame[21] ;   // verilog/coms.v(97[12:25])
    wire [7:0]\data_in_frame[20] ;   // verilog/coms.v(97[12:25])
    wire [7:0]\data_in_frame[14] ;   // verilog/coms.v(97[12:25])
    wire [7:0]\data_in_frame[13] ;   // verilog/coms.v(97[12:25])
    wire [7:0]\data_in_frame[12] ;   // verilog/coms.v(97[12:25])
    wire [7:0]\data_in_frame[11] ;   // verilog/coms.v(97[12:25])
    wire [7:0]\data_in_frame[10] ;   // verilog/coms.v(97[12:25])
    wire [7:0]\data_in_frame[9] ;   // verilog/coms.v(97[12:25])
    wire [7:0]\data_in_frame[8] ;   // verilog/coms.v(97[12:25])
    wire [7:0]\data_in_frame[6] ;   // verilog/coms.v(97[12:25])
    wire [7:0]\data_in_frame[5] ;   // verilog/coms.v(97[12:25])
    wire [7:0]\data_in_frame[4] ;   // verilog/coms.v(97[12:25])
    wire [7:0]\data_in_frame[3] ;   // verilog/coms.v(97[12:25])
    wire [7:0]\data_in_frame[2] ;   // verilog/coms.v(97[12:25])
    wire [7:0]\data_in_frame[1] ;   // verilog/coms.v(97[12:25])
    wire [7:0]\data_out_frame[25] ;   // verilog/coms.v(98[12:26])
    wire [7:0]\data_out_frame[24] ;   // verilog/coms.v(98[12:26])
    wire [7:0]\data_out_frame[23] ;   // verilog/coms.v(98[12:26])
    wire [7:0]\data_out_frame[22] ;   // verilog/coms.v(98[12:26])
    wire [7:0]\data_out_frame[21] ;   // verilog/coms.v(98[12:26])
    wire [7:0]\data_out_frame[20] ;   // verilog/coms.v(98[12:26])
    wire [7:0]\data_out_frame[19] ;   // verilog/coms.v(98[12:26])
    wire [7:0]\data_out_frame[18] ;   // verilog/coms.v(98[12:26])
    wire [7:0]\data_out_frame[17] ;   // verilog/coms.v(98[12:26])
    wire [7:0]\data_out_frame[16] ;   // verilog/coms.v(98[12:26])
    wire [7:0]\data_out_frame[15] ;   // verilog/coms.v(98[12:26])
    wire [7:0]\data_out_frame[14] ;   // verilog/coms.v(98[12:26])
    wire [7:0]\data_out_frame[13] ;   // verilog/coms.v(98[12:26])
    wire [7:0]\data_out_frame[12] ;   // verilog/coms.v(98[12:26])
    wire [7:0]\data_out_frame[11] ;   // verilog/coms.v(98[12:26])
    wire [7:0]\data_out_frame[10] ;   // verilog/coms.v(98[12:26])
    wire [7:0]\data_out_frame[9] ;   // verilog/coms.v(98[12:26])
    wire [7:0]\data_out_frame[8] ;   // verilog/coms.v(98[12:26])
    wire [7:0]\data_out_frame[7] ;   // verilog/coms.v(98[12:26])
    wire [7:0]\data_out_frame[6] ;   // verilog/coms.v(98[12:26])
    wire [7:0]\data_out_frame[5] ;   // verilog/coms.v(98[12:26])
    wire [7:0]\data_out_frame[4] ;   // verilog/coms.v(98[12:26])
    
    wire n44972, tx_active, n50022, n46128, n39033, n39032, n38859, 
        n50024, n42724, n25_adj_5270, n17_adj_5271, n38858, n4486, 
        n4485, n4497, n4496, n38857, n4488, n39031, n38856, n38855, 
        n50376, n39030, n38854, n38853, n39029, n39028, n4_adj_5272, 
        n51372, n51366, n51360, n51354, n51348, n51342, n51336, 
        n51330, n7_adj_5273, n38852, n39027, n38851, n537, n535, 
        n534, n533, n532, n7417, n35428, n531, n38850, n39026, 
        n35426, n39025, n38849, n38848, n39024, n39023, n39022, 
        n39021, n39020, n39019, n39018, n38847, n39017, n39016, 
        n38846, n38845, n39015, n39014, n38844, n39013, n39012, 
        n39011, n39010, n38843, n39009, n39008, n35424, n38842, 
        n39007, n39006, n39005, n38841, n38840, n38839, n38838, 
        n39004, n39003, n39002, n38837, n38836, n39001, n35420, 
        n34664, n34660, n35418, n38835, n35416, n35414, n39000, 
        n35410, n35408, n38467, n38999, n38998, n38997, n35402, 
        n38834, n38996, n38995, n38833, n35400, n38994, n35398, 
        n38832, n38993, n38831, n38830, n38992, n38829, n38466, 
        n35394, n38991, n38990, n38989, n38988, n38828, n35392, 
        n38987, n38986, n38985, n38984, n38983, n38982, n35388, 
        n38465, n38453, n38981, n35450, n38452, n38980, n6_adj_5274, 
        n38979, n38978, n38977, n38976, n38975, n38974, n35456, 
        n38973, n38972, n38971, n38970, n38811, n38810, n38969, 
        n38809, n38968, n38967, n38966, n38965, n38808, n38964, 
        n38963, n38962, n38807, n38961, n38960, n38959, n38958, 
        n38957, n38956, n38955, n38954, n38953, n38806, n38952, 
        n38805, n38951, n38950, n38804, n38803, n38949, n38948, 
        n38464, n46053, n10_adj_5275, n12_adj_5276, n19_adj_5277, 
        n2_adj_5278, n21_adj_5279, n530, n529, n528, n46084, n527, 
        n526, n525, n522, n521, n520, n38802, n38947, n38675, 
        n38674, n8_adj_5280, n38801, n38463, n7_adj_5281, n38800, 
        n38799, n519, n49719, n14_adj_5282, n38798, n38673, n10_adj_5283, 
        n49526, n44835, n38672, n51159, n38671, n38797, n38796, 
        n38795, n38946, n38794, n38945, n38944, n38499, n38498, 
        n38793, n38792, n45290, n50084, n44694, n5_adj_5284, n517, 
        n516, n43386, n44670, n38670, n4_adj_5285, n44668, n49518, 
        n12_adj_5286, n44748, n43380, n44666, n44664, n44661, n38943, 
        n4_adj_5287, n13_adj_5288, n38942, n44637, n49513, n44924, 
        n50463, n50455, n50454, n50451, n50544, n9_adj_5289, n27152, 
        n50635, n33, n32, n31, n30, n29, n28, n27, n26, n25_adj_5290, 
        n24_adj_5291, n23_adj_5292, n22_adj_5293, n21_adj_5294, n20_adj_5295, 
        n19_adj_5296, n18_adj_5297, n17_adj_5298, n16_adj_5299, n15_adj_5300, 
        n14_adj_5301, n13_adj_5302, n12_adj_5303, n11_adj_5304, n10_adj_5305, 
        n9_adj_5306, n8_adj_5307, n7_adj_5308, n6_adj_5309, n5_adj_5310, 
        n4_adj_5311, n3_adj_5312, n2_adj_5313, n25_adj_5314, n24_adj_5315, 
        n23_adj_5316, n22_adj_5317, n11_adj_5318, n50238, n21_adj_5319, 
        n20_adj_5320, n15_adj_5321, n19_adj_5322, n18_adj_5323, n17_adj_5324, 
        n16_adj_5325, n15_adj_5326, n14_adj_5327, n13_adj_5328, n12_adj_5329, 
        n11_adj_5330, n10_adj_5331, n9_adj_5332, n8_adj_5333, n7_adj_5334, 
        n6_adj_5335, n5_adj_5336, n4_adj_5337, n3_adj_5338, n50004, 
        n15_adj_5339, n38497, n50010, n24462, n6130, n6_adj_5340, 
        n29679, n29678, n29677, n29676, n29675, n29674, n29673, 
        n29672, n29671, n29670, n29669, n29668, n29667, n29666, 
        n29665, n29664, n29663, n29662, n29661, n29660, n29659, 
        n29658, n29657, n29656, n29655, n38791, n29654, n29653, 
        n29652, n29651, n29650, n29649, n29648, n29647, n29646, 
        n29645, n29644, n29643, n29642, n29641, n29640, n29639, 
        n29638, n10_adj_5341, n29637, n29636, n29635, n29634, n29633, 
        n29632, n29631, n29630, n8_adj_5342, n29629, n29628, n29627, 
        n29626, n29625, n29624, n29623, n29622, n29621, n29620, 
        n29619, n29618, n29617, n29616, n29615, n29614, n29134, 
        n29613, n29612, n50784, n29611, n29610, n29609, n29608, 
        n29607, n29606, n29605, n29604, n29133;
    wire [1:0]a_new;   // vhdl/quadrature_decoder.vhd(40[9:14])
    
    wire b_prev, n29602, n29599, n29598, n29597, n29596, n29595, 
        n29594, n29593, n29592, n29591, n29590, n29589, direction_N_4071, 
        n38451, n29588, n29587, n29586, n29585, n27143, n29584, 
        n29583, n29582, n29581, n29580, n29579, n29578, n29577, 
        n29576, n29575, n29574, n29573, n29572, n29571, n29570, 
        n29569, n29568, n49501, n29567, n4495, n4494, n29566, 
        n29565, n50386, n29564, n29563, n29562, n29561, n29560, 
        n29559, n29558, n29557, n29556, n29555, n29553, n29552, 
        n29551, n29550, n29549, n29548, n29547, n29546, n29545, 
        n29132;
    wire [1:0]a_new_adj_5490;   // vhdl/quadrature_decoder.vhd(40[9:14])
    
    wire b_prev_adj_5344, n2204, n2195, n38669, n29544, n29543, 
        n29542, n29541, n29540, n29539, n49819, n38790, n38462, 
        n38668, direction_N_4071_adj_5345, n38667, n29538, n29537, 
        n29536, n29535, n29534, n29533, n29532, n29531, n29530, 
        n29529, n29528, n29527, n29526, n29525, n29524, n29523, 
        n29522, n29521, n29520, n29519, n29518, n29517, n4493, 
        n4492, n4491, n4490, n4489, n29516, n29510, n29508, n43822, 
        n29506, n4_adj_5346, n29131, n29130, n29129, n29128, n29127, 
        n29126, n29125, n29124, n29123, n29122, n29121, n29120, 
        n29119, n29118, n29117, n29116, n29115, n29114, n44662, 
        n29505, n29504, n29503, n5_adj_5347, n29502, n29501, n29500, 
        n29113, n29499, n29498, n29497, rw;
    wire [7:0]state_adj_5510;   // verilog/eeprom.v(23[11:16])
    
    wire n51192, n51414, n29496, n29495, n29494, n29493, n29492, 
        n29491, n29490, n29489, n29488, n29487, n29486, n29485, 
        n29484, n29483, n29482, n9_adj_5349, n8_adj_5350, n29481, 
        n29480, n29479, n16_adj_5351, n29112, n29111, clk_out;
    wire [15:0]data_adj_5514;   // verilog/tli4970.v(27[14:18])
    wire [7:0]state_adj_5516;   // verilog/tli4970.v(29[13:18])
    
    wire n29478, n29477, n29476, n29475, n4_adj_5362, n7_adj_5363, 
        n6_adj_5364, n5_adj_5365, n4_adj_5366, n29474, n27013, n27167, 
        n29473, n29472, n29471, n29470, n11_adj_5367, n29469, n29468, 
        n29467, n29466, n29465, n29464, n29463, n29462, n29461, 
        n29460, n29459, n29458, n29457, n29456, n29455, n29454, 
        n29453, n5_adj_5368, n29110, n27015, n29452, n29451, n29450, 
        n30_adj_5369, n29449, state_7__N_4460, n29448, n45982, n29109, 
        n29108, n29447, n29446, n29445, n29444, n12_adj_5370, n10_adj_5371, 
        n8_adj_5372, n6_adj_5373, n4_adj_5374, n45800, n29107, r_Rx_Data;
    wire [2:0]r_Bit_Index;   // verilog/uart_rx.v(33[17:28])
    wire [2:0]r_SM_Main;   // verilog/uart_rx.v(36[17:26])
    
    wire n38496, n9_adj_5375, n13_adj_5376, n24_adj_5377, n29106, 
        n38941, n38666, n38940, n29105, n29104, n38665, n38450, 
        n4723, n4722, n4721, n4720;
    wire [2:0]r_SM_Main_2__N_3706;
    
    wire n38939, n29103, n50256;
    wire [2:0]r_SM_Main_adj_5525;   // verilog/uart_tx.v(31[16:25])
    wire [2:0]r_Bit_Index_adj_5527;   // verilog/uart_tx.v(33[16:27])
    
    wire n38789, n38788;
    wire [2:0]r_SM_Main_2__N_3777;
    
    wire n29102, n29101, n4719, n4718, n4717, n4716, n4715, n4714, 
        n4713, n4712, n4711, n4487, n29404, n29403, n29402, n29401, 
        n29400, n29399, n29398, n29397, n29396, n29395, n29394, 
        n29393, n29392, n29391, n29390, n29389, n29388;
    wire [7:0]state_adj_5537;   // verilog/i2c_controller.v(33[12:17])
    wire [7:0]saved_addr;   // verilog/i2c_controller.v(34[12:22])
    
    wire n29100, enable_slow_N_4354, n7754, n29099, n38495;
    wire [7:0]state_7__N_4251;
    
    wire n4710, n4709, n4708, n4707, n4706, n4705, n4704, n4703, 
        n4702, n4701, n4700, n4698, n29098, n7210, n29097;
    wire [7:0]state_7__N_4267;
    
    wire n38664, n38787, n38786, n38785, n38938, n38937, n29096, 
        n49837, n28_adj_5383, n26_adj_5384, n38663, n29095, n29094, 
        n29093, n29092, n29091, n29090, n29089, n29088, n19_adj_5385, 
        n28_adj_5386, n38936, n29087, n29086, n29085, n29084, n29083, 
        n29082, n29081, n29080, n29079, n29078, n29077, n29076, 
        n29075, n29074, n29073, n29069, n29067, n29066, n29065, 
        n29064, n29063, n29062, n29061, n29060, n29059, n29057, 
        n29056, n29055, n45989, n29054, n39523, n38935, n39522, 
        n7_adj_5387, n731, n39521, n38494, n38449, n38662, n8413, 
        n8412, n8411, n8410, n8409, n8408, n50754, n828, n829, 
        n830, n831, n832, n833, n39520, n861, n896, n897, n898, 
        n899, n900, n901, n927, n928, n929, n930, n931, n932, 
        n933, n38493, n937, n938, n38784, n28666, n950, n39519, 
        n960, n45056, n995, n996, n997, n998, n999, n1000, n1001, 
        n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, 
        n29019, n1059, n39518, n38934, n39517, n45028, n39516, 
        n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, 
        n1101, n35558, n38783, n38782, n1125, n1126, n1127, n1128, 
        n1129, n1130, n1131, n1132, n1133, n38933, n38932, n28662, 
        n1158, n28933, n39515, n39514, n39513, n1193, n1194, n1195, 
        n1196, n1197, n1198, n1199, n1200, n1201, n1224, n1225, 
        n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, 
        n1257, n1292, n1293, n1294, n1295, n1296, n1297_adj_5388, 
        n1298_adj_5389, n1299_adj_5390, n1300_adj_5391, n1301_adj_5392, 
        n51468, n1323_adj_5393, n1324_adj_5394, n1325_adj_5395, n1326_adj_5396, 
        n1327_adj_5397, n1328_adj_5398, n1329, n1330, n1331, n1332, 
        n1333, n45355, n1356, n38931, n51462, n1391, n1392, n1393, 
        n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, 
        n38930, n1422, n1423, n1424, n1425, n1426, n1427, n1428, 
        n1429, n1430, n1431, n1432, n1433, n1455, n51112, n1490, 
        n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, 
        n1499, n1500, n1501, n1521, n1522, n1523, n1524, n1525, 
        n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, 
        n1554, n39512, n39511, n39510, n39509, n39508, n1589, 
        n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, 
        n1598, n1599, n1600, n1601, n39507, n38492, n1620, n1621, 
        n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, 
        n1630, n1631, n1632, n1633, n1653, n39506, n39505, n39504, 
        n24278, n1688, n1689, n1690, n1691, n1692, n1693, n1694, 
        n1695, n1696, n1697, n1698, n1699, n1700, n1701, n38929, 
        n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, 
        n1727, n1728, n1729, n1730, n1731, n1732, n1733, n51099, 
        n1752, n49745, n1787, n1788, n1789, n1790, n1791, n1792, 
        n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, 
        n1801, n1818, n1819, n1820, n1821, n1822, n1823, n1824, 
        n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, 
        n1833, n38928, n38491, n38781, n1851, n39503, n39502, 
        n39501, n44993, n38780, n1886, n1887, n1888, n1889, n1890, 
        n1891_adj_5399, n1892, n1893, n1894, n1895, n1896_adj_5400, 
        n1897, n1898, n1899, n1900, n1901, n27180, n27171, n1917, 
        n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, 
        n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, 
        n39500, n1950, n39499, n49736, n39498, n39497, n39496, 
        n51602, n1985, n1986, n1987, n1988, n1989, n1990, n1991, 
        n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, 
        n2000, n2001, n46250, n2016, n2017, n2018, n2019, n2020, 
        n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, 
        n2029, n2030, n2031, n2032, n2033, n49732, n2049, n51727, 
        n39495, n43848, n51084, n2084, n2085, n2086, n2087, n2088, 
        n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, 
        n2097, n2098, n2099, n2100, n2101, n43847, n2115, n2116, 
        n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, 
        n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, 
        n2133, n2148, n43724, n2183, n2184, n2185, n2186, n2187, 
        n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195_adj_5401, 
        n2196, n2197, n2198, n2199, n2200, n2201, n45016, n2214, 
        n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, 
        n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, 
        n2231, n2232, n2233, n2247, n39494, n2281, n2282, n2283, 
        n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, 
        n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, 
        n2300, n2301, n2313, n2314, n2315, n2316, n2317, n2318, 
        n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, 
        n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2346, 
        n43839, n39493, n43838, n2381, n2382, n2383, n2384, n2385, 
        n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, 
        n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, 
        n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, 
        n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, 
        n2428, n2429, n2430, n2431, n2432, n2433, n51456, n2445, 
        n49722, n38461, n29052, n46347, n2480, n2481, n2482, n2483, 
        n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, 
        n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, 
        n2500, n2501, n2511, n2512, n2513, n2514, n2515, n2516, 
        n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524, 
        n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, 
        n2533, n46081, n2544, n2579, n2580, n2581, n2582, n2583, 
        n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, 
        n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, 
        n2600, n2601, n47201, n2610, n2611, n2612, n2613, n2614, 
        n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, 
        n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, 
        n2631, n2632, n2633, n5_adj_5402, n2643, n50462, n47195, 
        n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685, 
        n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, 
        n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, 
        n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716, 
        n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, 
        n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, 
        n2733, n50702, n2742, n47189, n38460, n49713, n2776, n2777, 
        n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785, 
        n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, 
        n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, 
        n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815, 
        n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, 
        n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, 
        n2832, n2833, n2841, n51069, n29339, n47183, n2876, n2877, 
        n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885, 
        n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, 
        n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, 
        n29338, n2907, n2908, n2909, n2910, n2911, n2912, n2913, 
        n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, 
        n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929, 
        n2930, n2931, n2932, n2933, n2940, n27147, n2975, n2976, 
        n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984, 
        n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, 
        n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, 
        n3001, n3006, n3007, n3008, n3009, n3010, n3011, n3012, 
        n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, 
        n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, 
        n3029, n3030, n3031, n3032, n3033, n3039, n29336, n28592, 
        n47177, n3074, n3075, n3076, n3077, n3078, n3079, n3080, 
        n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, 
        n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, 
        n3097, n3098, n3099, n3100, n3101, n3105, n3106, n3107, 
        n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115, 
        n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, 
        n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, 
        n3132, n3133, n38490, n29335, n3138, n27177, n47173, n3173, 
        n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, 
        n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189, 
        n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, 
        n3198, n3199, n3200, n3201, n3204, n3205, n3206, n3207, 
        n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215, 
        n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, 
        n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, 
        n3232, n3233, n29334, n3237, n3271, n3272, n3273, n3274, 
        n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, 
        n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, 
        n3291, n3292, n3293, n3294, n3295, n3296, n3298, n3299, 
        n3300, n3301, n50002, n27034, n47161, n47159, n47157, 
        n51053, n29333, n28562, n51709, n43824, n29332, n29331, 
        n43506, n29330, n24_adj_5403, n28537, n29329, n28522, n28521, 
        n29328, n62, n29327, n42404, n29326, n27037, n47145, n29325, 
        n29051, n29324, n47139, n47133, n44929, n29323, n28482, 
        n29322, n29321, n28835, n28458, n47127, n51450, n47121, 
        n47119, n47117, n51036, n46354, n47095, n51705, n27028, 
        n47089, n51018, n7_adj_5404, n38661, n47083, n47081, n29050, 
        n38927, n47075, n47071, n47069, n51444, n51703, n50593, 
        n50697, n38459, n38779, n38778, n38777, n38458, n38776, 
        n38489, n44913, n38488, n38457, n50427, n38487, n44908, 
        n47051, n47045, n47039, n38660, n47033, n47031, n38659, 
        n29049, n47023, n38926, n50241, n47011, n51438, n38925, 
        n38924, n47005, n38658, n38456, n47001, n50319, n38486, 
        n50999, n46995, n50365, n46993, n38448, n29047, n29046, 
        n38923, n38922, n51700, n48, n49, n50, n51, n52, n53, 
        n54, n55, n38485, n38657, n38656, n38921, n29045, n38484, 
        n29043, n29042, n38920, n38919, n38918, n38655, n38654, 
        n46979, n46975, n10621, n46969, n46967, n51697, n16_adj_5405, 
        n15_adj_5406, n14_adj_5407, n13_adj_5408, n12_adj_5409, n51692, 
        n49452, n38483, n46961, n38447, n38917, n39313, n38482, 
        n38916, n39312, n39311, n39310, n49357, n38915, n49422, 
        n38653, n39309, n35277, n46953, n39308, n38446, n39307, 
        n38914, n39306, n39305, n39304, n29290, n29288, n39303, 
        n39302, n39301, n38913, n39300, n50979, n39299, n39298, 
        n39297, n39296, n39295, n29270, n29269, n29268, n29267, 
        n29266, n29265, n29264, n29263, n29262, n29261, n29260, 
        n29259, n29258, n29257, n29256, n29255, n39294, n46941, 
        n46935, n46933, n39293, n39292, n39291, n29249, n29245, 
        n29244, n29243, n29242, n29241, n29240, n29239, n29238, 
        n29237, n50374, n39290, n46925, n38912, n39289, n39288, 
        n39287, n29233, n39286, n39285, n39284, n39283, n39282, 
        n39281, n29041, n29040, n29230, n29225, n29224, n29223, 
        n39280, n38911, n46923, n39279, n50364, n29033, n29032, 
        n29031, n29030, n29029, n29028, n29027, n29026, n29025, 
        n29221, n29220, n29219, n29218, n29217, n29216, n29215, 
        n29214, n39278, n39277, n46913, n38481, n39276, n46907, 
        n46903, n39275, n39274, n29213, n29212, n29211, n29210, 
        n29209, n29208, n29207, n29206, n29205, n29204, n29203, 
        n29202, n29201, n29200, n29199, n29198, n29197, n29196, 
        n29195, n29194, n29193, n29192, n29191, n29190, n29189, 
        n29188, n29187, n29184, n29183, n29182, n39273, n38910, 
        n39272, n39271, n39270, n29024, n29023, n29022, n29181, 
        n29180, n29179, n29178, n29177, n29176, n29175, n29174, 
        n38553, n39269, n28972, n29018, n29173, n29172, n29171, 
        n29170, n29169, n29168, n10_adj_5410, n39268, n49415, n50958, 
        n29021, n39267, n39266, n39265, n39264, n39263, n39262, 
        n39261, n49339, n46887, n39260, n27174, n39259, n46881, 
        n39258, n39257, n39256, n50426, n49335, n2_adj_5411, n3_adj_5412, 
        n4_adj_5413, n5_adj_5414, n6_adj_5415, n7_adj_5416, n8_adj_5417, 
        n9_adj_5418, n10_adj_5419, n11_adj_5420, n12_adj_5421, n13_adj_5422, 
        n14_adj_5423, n15_adj_5424, n16_adj_5425, n17_adj_5426, n18_adj_5427, 
        n19_adj_5428, n20_adj_5429, n21_adj_5430, n22_adj_5431, n23_adj_5432, 
        n24_adj_5433, n25_adj_5434, n26_adj_5435, n27_adj_5436, n28_adj_5437, 
        n29_adj_5438, n30_adj_5439, n31_adj_5440, n32_adj_5441, n33_adj_5442, 
        n49334, n46863, n39255, n38480, n39254, n39253, n46857, 
        n39252, n39251, n39250, n39249, n39248, n50937, n46849, 
        n27126, n47975, n39247, n39246, n39245, n39244, n39243, 
        n39242, n29020, n39241, n39240, n39239, n39238, n39237, 
        n45933, n39236, n27131, n39235, n39234, n39233, n46837, 
        n39232, n39231, n39230, n39229, n39228, n46833, n39227, 
        n39226, n50315, n39225, n39224, n39223, n39222, n39221, 
        n39220, n51432, n39219, n39218, n39217, n39216, n39215, 
        n39214, n46821, n46815, n39213, n39212, n39211, n39210, 
        n39209, n39208, n46807, n39207, n39206, n39205, n39204, 
        n39203, n39202, n46801, n39201, n38909, n46440, n39200, 
        n14_adj_5443, n45203, n38908, n28970, n39199, n39198, n39197, 
        n39196, n39195, n38907, n39194, n39193, n38906, n10_adj_5444, 
        n38905, n38552, n46793, n39192, n44998, n39191, n39190, 
        n34717, n39189, n39188, n39187, n38551, n39186, n39185, 
        n39184, n39183, n39182, n39181, n39180, n38550, n38479, 
        n38478, n39179, n6_adj_5445, n39178, n39177, n39176, n39175, 
        n39174, n38549, n39173, n39172, n46783, n39171, n39170, 
        n39169, n39168, n39167, n38477, n38548, n39166, n39165, 
        n39164, n39163, n39162, n38904, n39161, n39160, n39159, 
        n46777, n38903, n39158, n39157, n39156, n39155, n38902, 
        n39154, n46773, n38547, n38901, n39153, n39152, n19541, 
        n39151, n39150, n39149, n39148, n46767, n39147, n39146, 
        n39145, n35498, n39144, n39143, n38546, n39142, n35496, 
        n39141, n39140, n39139, n39138, n39137, n46765, n38900, 
        n39136, n38899, n39135, n39134, n39133, n38545, n38898, 
        n38897, n39132, n35492, n38896, n39131, n46757, n39130, 
        n39129, n39128, n39127, n39126, n39125, n39124, n39123, 
        n39122, n39121, n38544, n38895, n39120, n38543, n39119, 
        n39118, n39117, n39116, n39115, n38542, n39114, n39113, 
        n38894, n39112, n39111, n35484, n39110, n38476, n39109, 
        n38475, n39108, n39107, n39106, n39105, n39104, n46743, 
        n38474, n38541, n38473, n39103, n38540, n39102, n49374, 
        n34695, n39101, n39100, n39099, n39098, n39097, n39096, 
        n38893, n38892, n39095, n39094, n39093, n39092, n38539, 
        n39091, n39090, n39089, n39088, n39087, n39086, n34690, 
        n39085, n38891, n39084, n38472, n39083, n39082, n39081, 
        n38471, n46737, n39080, n35474, n39079, n34688, n39078, 
        n39077, n39076, n39075, n39074, n39073, n38538, n38537, 
        n39072, n39071, n38890, n39070, n39069, n39068, n38889, 
        n39067, n39066, n39065, n39064, n38455, n39063, n27014, 
        n39062, n46731, n38888, n38454, n38536, n39061, n39060, 
        n39059, n39058, n39057, n39056, n7_adj_5446, n39055, n39054, 
        n13_adj_5447, n38887, n38886, n17_adj_5448, n19_adj_5449, 
        n21_adj_5450, n27_adj_5451, n31_adj_5452, n46725, n37, n38885, 
        n38884, n38470, n50914, n46719, n46717, n46703, n46697, 
        n46691, n46689, n50384, n46683, n46679, n44970, n46677, 
        n50668, n50217, n46665, n46663, n46661, n46659, n46657, 
        n46655, n46653, n46651, n46649, n46647, n46645, n46643, 
        n46641, n44955, n46412, n46410, n46639, n46635, n51408, 
        n10_adj_5453, n46627, n46625, n50214, n46623, n46621, n46619, 
        n46617, n46611, n46609, n46603, n46599, n46591, n51426, 
        n49302, n50161, n46585, n50890, n50452, n46579, n46577, 
        n46569, n49298, n49297, n49296, n49295, n46563, n46561, 
        n49294, n49293, n50312, n49292, n49289, n50865, n46551, 
        n46545, n50029, n46539, n46533, n43630, n44905, n46531, 
        n50160, n50242, n51420, n6_adj_5454, n50221;
    
    VCC i2 (.Y(VCC_net));
    SB_IO hall2_input (.PACKAGE_PIN(HALL2), .LATCH_INPUT_VALUE(GND_net), 
          .INPUT_CLK(GND_net), .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_1(GND_net), .D_OUT_0(GND_net), .D_IN_0(hall2)) /* synthesis syn_instantiated=1, IO_FF_IN=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam hall2_input.PIN_TYPE = 6'b000001;
    defparam hall2_input.PULLUP = 1'b1;
    defparam hall2_input.NEG_TRIGGER = 1'b0;
    defparam hall2_input.IO_STANDARD = "SB_LVCMOS";
    SB_IO hall3_input (.PACKAGE_PIN(HALL3), .LATCH_INPUT_VALUE(GND_net), 
          .INPUT_CLK(GND_net), .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_1(GND_net), .D_OUT_0(GND_net), .D_IN_0(hall3)) /* synthesis syn_instantiated=1, IO_FF_IN=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam hall3_input.PIN_TYPE = 6'b000001;
    defparam hall3_input.PULLUP = 1'b1;
    defparam hall3_input.NEG_TRIGGER = 1'b0;
    defparam hall3_input.IO_STANDARD = "SB_LVCMOS";
    SB_IO tx_output (.PACKAGE_PIN(TX), .LATCH_INPUT_VALUE(GND_net), .INPUT_CLK(GND_net), 
          .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(tx_enable), .D_OUT_1(GND_net), 
          .D_OUT_0(tx_o)) /* synthesis syn_instantiated=1 */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam tx_output.PIN_TYPE = 6'b101001;
    defparam tx_output.PULLUP = 1'b1;
    defparam tx_output.NEG_TRIGGER = 1'b0;
    defparam tx_output.IO_STANDARD = "SB_LVCMOS";
    SB_DFF commutation_state_prev_i0 (.Q(commutation_state_prev[0]), .C(CLK_c), 
           .D(commutation_state[0]));   // verilog/TinyFPGA_B.v(144[9] 223[5])
    SB_DFF dir_187 (.Q(dir), .C(CLK_c), .D(pwm_setpoint_23__N_239));   // verilog/TinyFPGA_B.v(104[9] 130[5])
    SB_LUT4 unary_minus_19_inv_0_i12_1_lut (.I0(duty[11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n14_adj_5259));   // verilog/TinyFPGA_B.v(123[25:30])
    defparam unary_minus_19_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_19_inv_0_i13_1_lut (.I0(duty[12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n13));   // verilog/TinyFPGA_B.v(123[25:30])
    defparam unary_minus_19_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_DFFE dti_189 (.Q(dti), .C(CLK_c), .E(n28458), .D(dti_N_440));   // verilog/TinyFPGA_B.v(144[9] 223[5])
    SB_LUT4 i1_3_lut (.I0(n1226), .I1(n1227), .I2(n1228), .I3(GND_net), 
            .O(n46837));
    defparam i1_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_4_lut (.I0(n1229), .I1(n35428), .I2(n1230), .I3(n1231), 
            .O(n44908));
    defparam i1_4_lut.LUT_INIT = 16'ha080;
    SB_LUT4 i35500_4_lut (.I0(n1225), .I1(n1224), .I2(n44908), .I3(n46837), 
            .O(n1257));
    defparam i35500_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i15207_3_lut (.I0(IntegralLimit[4]), .I1(\data_in_frame[13] [4]), 
            .I2(n28521), .I3(GND_net), .O(n29155));   // verilog/coms.v(128[12] 303[6])
    defparam i15207_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15593_3_lut (.I0(\data_out_frame[23] [0]), .I1(neopxl_color[16]), 
            .I2(n24278), .I3(GND_net), .O(n29541));   // verilog/coms.v(128[12] 303[6])
    defparam i15593_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF encoder0_position_scaled_i0 (.Q(encoder0_position_scaled[0]), .C(CLK_c), 
           .D(encoder0_position_scaled_23__N_51[0]));   // verilog/TinyFPGA_B.v(337[10] 341[6])
    SB_DFF encoder1_position_scaled_i0 (.Q(encoder1_position_scaled[0]), .C(CLK_c), 
           .D(encoder1_position_scaled_23__N_75[0]));   // verilog/TinyFPGA_B.v(337[10] 341[6])
    SB_LUT4 encoder0_position_31__I_0_i701_3_lut (.I0(n1026), .I1(n1093), 
            .I2(n1059), .I3(GND_net), .O(n1125));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i701_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i706_3_lut (.I0(n1031), .I1(n1098), 
            .I2(n1059), .I3(GND_net), .O(n1130));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i706_3_lut.LUT_INIT = 16'hacac;
    SB_IO sda_output (.PACKAGE_PIN(SDA), .LATCH_INPUT_VALUE(GND_net), .INPUT_CLK(GND_net), 
          .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(sda_enable), .D_OUT_1(GND_net), 
          .D_OUT_0(sda_out), .D_IN_0(state_7__N_4267[3])) /* synthesis syn_instantiated=1 */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam sda_output.PIN_TYPE = 6'b101001;
    defparam sda_output.PULLUP = 1'b1;
    defparam sda_output.NEG_TRIGGER = 1'b0;
    defparam sda_output.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 encoder0_position_31__I_0_i705_3_lut (.I0(n1030), .I1(n1097), 
            .I2(n1059), .I3(GND_net), .O(n1129));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i705_3_lut.LUT_INIT = 16'hacac;
    SB_DFF displacement_i0 (.Q(displacement[0]), .C(CLK_c), .D(displacement_23__N_99[0]));   // verilog/TinyFPGA_B.v(337[10] 341[6])
    SB_IO CS_pad (.PACKAGE_PIN(CS), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(CS_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam CS_pad.PIN_TYPE = 6'b011001;
    defparam CS_pad.PULLUP = 1'b0;
    defparam CS_pad.NEG_TRIGGER = 1'b0;
    defparam CS_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO scl_output (.PACKAGE_PIN(SCL), .LATCH_INPUT_VALUE(GND_net), .INPUT_CLK(GND_net), 
          .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(scl_enable), .D_OUT_1(GND_net), 
          .D_OUT_0(scl)) /* synthesis syn_instantiated=1 */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam scl_output.PIN_TYPE = 6'b101001;
    defparam scl_output.PULLUP = 1'b1;
    defparam scl_output.NEG_TRIGGER = 1'b0;
    defparam scl_output.IO_STANDARD = "SB_LVCMOS";
    SB_IO hall1_input (.PACKAGE_PIN(HALL1), .LATCH_INPUT_VALUE(GND_net), 
          .INPUT_CLK(GND_net), .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_1(GND_net), .D_OUT_0(GND_net), .D_IN_0(hall1)) /* synthesis syn_instantiated=1, IO_FF_IN=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam hall1_input.PIN_TYPE = 6'b000001;
    defparam hall1_input.PULLUP = 1'b1;
    defparam hall1_input.NEG_TRIGGER = 1'b0;
    defparam hall1_input.IO_STANDARD = "SB_LVCMOS";
    \neopixel(CLOCK_SPEED_HZ=16000000)  nx (.GND_net(GND_net), .timer({timer}), 
            .CLK_c(CLK_c), .\neo_pixel_transmitter.t0 ({\neo_pixel_transmitter.t0 }), 
            .neopxl_color({neopxl_color}), .VCC_net(VCC_net), .\state[1] (state[1]), 
            .n42404(n42404), .\state_3__N_552[1] (state_3__N_552[1]), .LED_c(LED_c), 
            .n29069(n29069), .n28592(n28592), .n44637(n44637), .n29022(n29022), 
            .n29498(n29498), .n29497(n29497), .n29496(n29496), .n29495(n29495), 
            .n29494(n29494), .n29493(n29493), .n29492(n29492), .n29491(n29491), 
            .n29490(n29490), .n29489(n29489), .n29488(n29488), .n29487(n29487), 
            .n29486(n29486), .n29485(n29485), .n29484(n29484), .n29483(n29483), 
            .n29482(n29482), .n29481(n29481), .n29480(n29480), .n29479(n29479), 
            .n29478(n29478), .n29477(n29477), .n29476(n29476), .n29475(n29475), 
            .n29474(n29474), .n29473(n29473), .n29472(n29472), .n29471(n29471), 
            .n29470(n29470), .n29469(n29469), .n29468(n29468), .NEOPXL_c(NEOPXL_c)) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(43[24] 49[2])
    SB_LUT4 mux_1005_i23_3_lut (.I0(duty[22]), .I1(n341), .I2(duty[23]), 
            .I3(GND_net), .O(n4701));   // verilog/TinyFPGA_B.v(118[13] 129[7])
    defparam mux_1005_i23_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i35166_1_lut (.I0(n2544), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n50754));
    defparam i35166_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 inv_1004_i24_1_lut (.I0(current[15]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2));   // verilog/TinyFPGA_B.v(118[13] 129[7])
    defparam inv_1004_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i4933_2_lut (.I0(n340), .I1(duty[23]), .I2(GND_net), .I3(GND_net), 
            .O(n4700));
    defparam i4933_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i35114_1_lut (.I0(n2643), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n50702));
    defparam i35114_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_19_inv_0_i14_1_lut (.I0(duty[13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n12));   // verilog/TinyFPGA_B.v(123[25:30])
    defparam unary_minus_19_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i28_3_lut (.I0(encoder0_position[27]), 
            .I1(n6_adj_5309), .I2(encoder0_position[31]), .I3(GND_net), 
            .O(n517));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_mux_3_i28_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1005_i9_3_lut (.I0(duty[8]), .I1(n355), .I2(duty[23]), 
            .I3(GND_net), .O(n4715));   // verilog/TinyFPGA_B.v(118[13] 129[7])
    defparam mux_1005_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_19_inv_0_i2_1_lut (.I0(duty[1]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n24_adj_5269));   // verilog/TinyFPGA_B.v(123[25:30])
    defparam unary_minus_19_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_1005_i10_3_lut (.I0(duty[9]), .I1(n354), .I2(duty[23]), 
            .I3(GND_net), .O(n4714));   // verilog/TinyFPGA_B.v(118[13] 129[7])
    defparam mux_1005_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i1_1_lut (.I0(encoder0_position[0]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n33_adj_5442));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i29_3_lut (.I0(encoder0_position[28]), 
            .I1(n5_adj_5310), .I2(encoder0_position[31]), .I3(GND_net), 
            .O(n516));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_mux_3_i29_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i30_3_lut (.I0(encoder0_position[29]), 
            .I1(n4_adj_5311), .I2(encoder0_position[31]), .I3(GND_net), 
            .O(n623));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_mux_3_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i2_1_lut (.I0(encoder0_position[1]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n32_adj_5441));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i31_3_lut (.I0(encoder0_position[30]), 
            .I1(n3_adj_5312), .I2(encoder0_position[31]), .I3(GND_net), 
            .O(n622));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_mux_3_i31_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i3_1_lut (.I0(encoder0_position[2]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n31_adj_5440));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_i704_3_lut (.I0(n1029), .I1(n1096), 
            .I2(n1059), .I3(GND_net), .O(n1128));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i704_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i703_3_lut (.I0(n1028), .I1(n1095), 
            .I2(n1059), .I3(GND_net), .O(n1127));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i703_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i702_3_lut (.I0(n1027), .I1(n1094), 
            .I2(n1059), .I3(GND_net), .O(n1126));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i702_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i709_3_lut (.I0(n521), .I1(n1101), 
            .I2(n1059), .I3(GND_net), .O(n1133));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i709_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i4930_2_lut (.I0(n2_adj_5313), .I1(encoder0_position[31]), .I2(GND_net), 
            .I3(GND_net), .O(n621));
    defparam i4930_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 encoder0_position_31__I_0_i708_3_lut (.I0(n1033), .I1(n1100), 
            .I2(n1059), .I3(GND_net), .O(n1132));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i708_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i707_3_lut (.I0(n1032), .I1(n1099), 
            .I2(n1059), .I3(GND_net), .O(n1131));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i707_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i23_3_lut (.I0(encoder0_position[22]), 
            .I1(n11_adj_5304), .I2(encoder0_position[31]), .I3(GND_net), 
            .O(n522));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_mux_3_i23_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i35511_1_lut (.I0(n1158), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n51099));
    defparam i35511_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i15594_3_lut (.I0(\data_out_frame[22] [7]), .I1(current[7]), 
            .I2(n24278), .I3(GND_net), .O(n29542));   // verilog/coms.v(128[12] 303[6])
    defparam i15594_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i21543_4_lut (.I0(n522), .I1(n1131), .I2(n1132), .I3(n1133), 
            .O(n35492));
    defparam i21543_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 i1_3_lut_adj_1742 (.I0(n1126), .I1(n1127), .I2(n1128), .I3(GND_net), 
            .O(n46599));
    defparam i1_3_lut_adj_1742.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_2_lut (.I0(n1129), .I1(n1130), .I2(GND_net), .I3(GND_net), 
            .O(n46833));
    defparam i1_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i35514_4_lut (.I0(n46833), .I1(n1125), .I2(n46599), .I3(n35492), 
            .O(n1158));
    defparam i35514_4_lut.LUT_INIT = 16'h0103;
    SB_LUT4 encoder0_position_31__I_0_i636_3_lut (.I0(n929), .I1(n996), 
            .I2(n960), .I3(GND_net), .O(n1028));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i636_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i635_rep_63_3_lut (.I0(n928), .I1(n995), 
            .I2(n960), .I3(GND_net), .O(n1027));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i635_rep_63_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i639_3_lut (.I0(n932), .I1(n999), 
            .I2(n960), .I3(GND_net), .O(n1031));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i639_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i638_3_lut (.I0(n931), .I1(n998), 
            .I2(n960), .I3(GND_net), .O(n1030));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i638_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i4_1_lut (.I0(encoder0_position[3]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n30_adj_5439));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_19_inv_0_i15_1_lut (.I0(duty[14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_5258));   // verilog/TinyFPGA_B.v(123[25:30])
    defparam unary_minus_19_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_i637_3_lut (.I0(n930), .I1(n997), 
            .I2(n960), .I3(GND_net), .O(n1029));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i637_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i570_3_lut (.I0(n831), .I1(n898), 
            .I2(n861), .I3(GND_net), .O(n930));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i570_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i569_3_lut (.I0(n830), .I1(n897), 
            .I2(n861), .I3(GND_net), .O(n929));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i569_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i568_3_lut (.I0(n829), .I1(n896), 
            .I2(n861), .I3(GND_net), .O(n928));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i568_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29152_3_lut (.I0(n4_adj_5311), .I1(n8410), .I2(n44661), .I3(GND_net), 
            .O(n44664));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam i29152_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29153_3_lut (.I0(encoder0_position[29]), .I1(n44664), .I2(encoder0_position[31]), 
            .I3(GND_net), .O(n830));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam i29153_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut_adj_1743 (.I0(n5_adj_5284), .I1(n3_adj_5312), .I2(encoder0_position[31]), 
            .I3(GND_net), .O(n46933));
    defparam i1_3_lut_adj_1743.LUT_INIT = 16'h8080;
    SB_LUT4 unary_minus_19_inv_0_i16_1_lut (.I0(duty[15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n10));   // verilog/TinyFPGA_B.v(123[25:30])
    defparam unary_minus_19_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_i500_4_lut (.I0(n2_adj_5313), .I1(n8408), 
            .I2(n46933), .I3(encoder0_position[31]), .O(n828));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i500_4_lut.LUT_INIT = 16'h8a80;
    SB_LUT4 i29150_3_lut (.I0(n3_adj_5312), .I1(n8409), .I2(n44661), .I3(GND_net), 
            .O(n44662));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam i29150_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29151_3_lut (.I0(encoder0_position[30]), .I1(n44662), .I2(encoder0_position[31]), 
            .I3(GND_net), .O(n829));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam i29151_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i27_3_lut (.I0(encoder0_position[26]), 
            .I1(n7_adj_5308), .I2(encoder0_position[31]), .I3(GND_net), 
            .O(n731));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_mux_3_i27_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1744 (.I0(n4_adj_5311), .I1(n5_adj_5310), .I2(n731), 
            .I3(n6_adj_5309), .O(n5_adj_5284));
    defparam i1_4_lut_adj_1744.LUT_INIT = 16'heeea;
    SB_LUT4 i1_3_lut_adj_1745 (.I0(n3_adj_5312), .I1(n2_adj_5313), .I2(n5_adj_5284), 
            .I3(GND_net), .O(n44661));
    defparam i1_3_lut_adj_1745.LUT_INIT = 16'h8080;
    SB_LUT4 i29159_3_lut (.I0(encoder0_position[26]), .I1(n44670), .I2(encoder0_position[31]), 
            .I3(GND_net), .O(n833));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam i29159_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29156_3_lut (.I0(n6_adj_5309), .I1(n8412), .I2(n44661), .I3(GND_net), 
            .O(n44668));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam i29156_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29157_3_lut (.I0(encoder0_position[27]), .I1(n44668), .I2(encoder0_position[31]), 
            .I3(GND_net), .O(n832));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam i29157_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29154_3_lut (.I0(n5_adj_5310), .I1(n8411), .I2(n44661), .I3(GND_net), 
            .O(n44666));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam i29154_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29155_3_lut (.I0(encoder0_position[28]), .I1(n44666), .I2(encoder0_position[31]), 
            .I3(GND_net), .O(n831));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam i29155_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i21549_4_lut (.I0(n519), .I1(n831), .I2(n832), .I3(n833), 
            .O(n35498));
    defparam i21549_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 i21625_4_lut (.I0(n829), .I1(n828), .I2(n35498), .I3(n830), 
            .O(n861));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam i21625_4_lut.LUT_INIT = 16'heccc;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i26_3_lut (.I0(encoder0_position[25]), 
            .I1(n8_adj_5307), .I2(encoder0_position[31]), .I3(GND_net), 
            .O(n519));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_mux_3_i26_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29158_3_lut (.I0(n7_adj_5308), .I1(n8413), .I2(n44661), .I3(GND_net), 
            .O(n44670));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam i29158_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i573_3_lut (.I0(n519), .I1(n901), 
            .I2(n861), .I3(GND_net), .O(n933));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i573_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i572_3_lut (.I0(n833), .I1(n900), 
            .I2(n861), .I3(GND_net), .O(n932));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i572_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i571_3_lut (.I0(n832), .I1(n899), 
            .I2(n861), .I3(GND_net), .O(n931));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i571_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i21547_4_lut (.I0(n520), .I1(n931), .I2(n932), .I3(n933), 
            .O(n35496));
    defparam i21547_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 i15595_3_lut (.I0(current[11]), .I1(data_adj_5514[11]), .I2(n28537), 
            .I3(GND_net), .O(n29543));   // verilog/tli4970.v(35[10] 68[6])
    defparam i15595_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_19_inv_0_i17_1_lut (.I0(duty[16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n9));   // verilog/TinyFPGA_B.v(123[25:30])
    defparam unary_minus_19_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_2_lut_adj_1746 (.I0(n929), .I1(n930), .I2(GND_net), .I3(GND_net), 
            .O(n46757));
    defparam i1_2_lut_adj_1746.LUT_INIT = 16'h8888;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i5_1_lut (.I0(encoder0_position[4]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n29_adj_5438));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_4_lut_adj_1747 (.I0(n927), .I1(n46757), .I2(n928), .I3(n35496), 
            .O(n960));
    defparam i1_4_lut_adj_1747.LUT_INIT = 16'hfefa;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i6_1_lut (.I0(encoder0_position[5]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n28_adj_5437));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i25_3_lut (.I0(encoder0_position[24]), 
            .I1(n9_adj_5306), .I2(encoder0_position[31]), .I3(GND_net), 
            .O(n520));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_mux_3_i25_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i641_3_lut (.I0(n520), .I1(n1001), 
            .I2(n960), .I3(GND_net), .O(n1033));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i641_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i640_3_lut (.I0(n933), .I1(n1000), 
            .I2(n960), .I3(GND_net), .O(n1032));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i640_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15596_3_lut (.I0(current[10]), .I1(data_adj_5514[10]), .I2(n28537), 
            .I3(GND_net), .O(n29544));   // verilog/tli4970.v(35[10] 68[6])
    defparam i15596_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i24_3_lut (.I0(encoder0_position[23]), 
            .I1(n10_adj_5305), .I2(encoder0_position[31]), .I3(GND_net), 
            .O(n521));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_mux_3_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i35524_1_lut (.I0(n1059), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n51112));
    defparam i35524_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i21484_3_lut (.I0(n521), .I1(n1032), .I2(n1033), .I3(GND_net), 
            .O(n35432));
    defparam i21484_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i1_4_lut_adj_1748 (.I0(n1029), .I1(n35432), .I2(n1030), .I3(n1031), 
            .O(n44913));
    defparam i1_4_lut_adj_1748.LUT_INIT = 16'ha080;
    SB_LUT4 i35527_4_lut (.I0(n1026), .I1(n44913), .I2(n1027), .I3(n1028), 
            .O(n1059));
    defparam i35527_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i32_1_lut (.I0(encoder0_position[31]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n2_adj_5411));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i32_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i15072_3_lut (.I0(\data_out_frame[12] [7]), .I1(setpoint[23]), 
            .I2(n24278), .I3(GND_net), .O(n29020));   // verilog/coms.v(128[12] 303[6])
    defparam i15072_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i7_1_lut (.I0(encoder0_position[6]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n27_adj_5436));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 LessThan_15_i15_2_lut (.I0(current[7]), .I1(current_limit[7]), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_5247));   // verilog/TinyFPGA_B.v(119[9:30])
    defparam LessThan_15_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i13_2_lut (.I0(current[6]), .I1(current_limit[6]), 
            .I2(GND_net), .I3(GND_net), .O(n13_adj_5288));   // verilog/TinyFPGA_B.v(119[9:30])
    defparam LessThan_15_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i19_2_lut (.I0(current[9]), .I1(current_limit[9]), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_5385));   // verilog/TinyFPGA_B.v(119[9:30])
    defparam LessThan_15_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i17_2_lut (.I0(current[8]), .I1(current_limit[8]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_5246));   // verilog/TinyFPGA_B.v(119[9:30])
    defparam LessThan_15_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i7_2_lut (.I0(current[3]), .I1(current_limit[3]), 
            .I2(GND_net), .I3(GND_net), .O(n7_adj_5363));   // verilog/TinyFPGA_B.v(119[9:30])
    defparam LessThan_15_i7_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i9_2_lut (.I0(current[4]), .I1(current_limit[4]), 
            .I2(GND_net), .I3(GND_net), .O(n9_adj_5349));   // verilog/TinyFPGA_B.v(119[9:30])
    defparam LessThan_15_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i11_2_lut (.I0(current[5]), .I1(current_limit[5]), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_5318));   // verilog/TinyFPGA_B.v(119[9:30])
    defparam LessThan_15_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 unary_minus_19_inv_0_i18_1_lut (.I0(duty[17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n8_adj_5257));   // verilog/TinyFPGA_B.v(123[25:30])
    defparam unary_minus_19_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 LessThan_15_i5_2_lut (.I0(current[2]), .I1(current_limit[2]), 
            .I2(GND_net), .I3(GND_net), .O(n5_adj_5365));   // verilog/TinyFPGA_B.v(119[9:30])
    defparam LessThan_15_i5_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i8_1_lut (.I0(encoder0_position[7]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n26_adj_5435));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i9_1_lut (.I0(encoder0_position[8]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n25_adj_5434));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i33865_4_lut (.I0(n11_adj_5318), .I1(n9_adj_5349), .I2(n7_adj_5363), 
            .I3(n5_adj_5365), .O(n49452));
    defparam i33865_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 LessThan_15_i16_3_lut (.I0(n8_adj_5350), .I1(current_limit[9]), 
            .I2(n19_adj_5385), .I3(GND_net), .O(n16));   // verilog/TinyFPGA_B.v(119[9:30])
    defparam LessThan_15_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_15_i4_4_lut (.I0(current_limit[0]), .I1(current_limit[1]), 
            .I2(current[1]), .I3(current[0]), .O(n4_adj_5366));   // verilog/TinyFPGA_B.v(119[9:30])
    defparam LessThan_15_i4_4_lut.LUT_INIT = 16'h0c8e;
    SB_LUT4 i34572_3_lut (.I0(n4_adj_5366), .I1(current_limit[5]), .I2(n11_adj_5318), 
            .I3(GND_net), .O(n50160));   // verilog/TinyFPGA_B.v(119[9:30])
    defparam i34572_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34573_3_lut (.I0(n50160), .I1(current_limit[6]), .I2(n13_adj_5288), 
            .I3(GND_net), .O(n50161));   // verilog/TinyFPGA_B.v(119[9:30])
    defparam i34573_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_19_inv_0_i19_1_lut (.I0(duty[18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n7));   // verilog/TinyFPGA_B.v(123[25:30])
    defparam unary_minus_19_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i33835_4_lut (.I0(n17_adj_5246), .I1(n15_adj_5247), .I2(n13_adj_5288), 
            .I3(n49452), .O(n49422));
    defparam i33835_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i10_1_lut (.I0(encoder0_position[9]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n24_adj_5433));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i34798_4_lut (.I0(n16), .I1(n6_adj_5364), .I2(n19_adj_5385), 
            .I3(n49415), .O(n50386));   // verilog/TinyFPGA_B.v(119[9:30])
    defparam i34798_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i11_1_lut (.I0(encoder0_position[10]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n23_adj_5432));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i34157_3_lut (.I0(n50161), .I1(current_limit[7]), .I2(n15_adj_5247), 
            .I3(GND_net), .O(n49745));   // verilog/TinyFPGA_B.v(119[9:30])
    defparam i34157_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34866_4_lut (.I0(n49745), .I1(n50386), .I2(n19_adj_5385), 
            .I3(n49422), .O(n50454));   // verilog/TinyFPGA_B.v(119[9:30])
    defparam i34866_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i34867_3_lut (.I0(n50454), .I1(current_limit[10]), .I2(current[10]), 
            .I3(GND_net), .O(n50455));   // verilog/TinyFPGA_B.v(119[9:30])
    defparam i34867_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i34863_3_lut (.I0(n50455), .I1(current_limit[11]), .I2(current[11]), 
            .I3(GND_net), .O(n50451));   // verilog/TinyFPGA_B.v(119[9:30])
    defparam i34863_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i34837_3_lut (.I0(n50451), .I1(current_limit[12]), .I2(current[15]), 
            .I3(GND_net), .O(n26_adj_5384));   // verilog/TinyFPGA_B.v(119[9:30])
    defparam i34837_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 LessThan_15_i28_3_lut (.I0(n26_adj_5384), .I1(current_limit[13]), 
            .I2(current[15]), .I3(GND_net), .O(n28_adj_5383));   // verilog/TinyFPGA_B.v(119[9:30])
    defparam LessThan_15_i28_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i34621_4_lut (.I0(n28_adj_5383), .I1(current[15]), .I2(current_limit[15]), 
            .I3(current_limit[14]), .O(n287));   // verilog/TinyFPGA_B.v(119[9:30])
    defparam i34621_4_lut.LUT_INIT = 16'h8f0e;
    SB_LUT4 LessThan_11_i17_2_lut (.I0(current[8]), .I1(duty[8]), .I2(GND_net), 
            .I3(GND_net), .O(n17));   // verilog/TinyFPGA_B.v(111[10:22])
    defparam LessThan_11_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_11_i19_2_lut (.I0(current[9]), .I1(duty[9]), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_5277));   // verilog/TinyFPGA_B.v(111[10:22])
    defparam LessThan_11_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_11_i21_2_lut (.I0(current[10]), .I1(duty[10]), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_5279));   // verilog/TinyFPGA_B.v(111[10:22])
    defparam LessThan_11_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_11_i23_2_lut (.I0(current[11]), .I1(duty[11]), .I2(GND_net), 
            .I3(GND_net), .O(n23));   // verilog/TinyFPGA_B.v(111[10:22])
    defparam LessThan_11_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_11_i7_2_lut (.I0(current[3]), .I1(duty[3]), .I2(GND_net), 
            .I3(GND_net), .O(n7_adj_5387));   // verilog/TinyFPGA_B.v(111[10:22])
    defparam LessThan_11_i7_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_11_i9_2_lut (.I0(current[4]), .I1(duty[4]), .I2(GND_net), 
            .I3(GND_net), .O(n9_adj_5375));   // verilog/TinyFPGA_B.v(111[10:22])
    defparam LessThan_11_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_11_i11_2_lut (.I0(current[5]), .I1(duty[5]), .I2(GND_net), 
            .I3(GND_net), .O(n11));   // verilog/TinyFPGA_B.v(111[10:22])
    defparam LessThan_11_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_11_i13_2_lut (.I0(current[6]), .I1(duty[6]), .I2(GND_net), 
            .I3(GND_net), .O(n13_adj_5376));   // verilog/TinyFPGA_B.v(111[10:22])
    defparam LessThan_11_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_11_i15_2_lut (.I0(current[7]), .I1(duty[7]), .I2(GND_net), 
            .I3(GND_net), .O(n15));   // verilog/TinyFPGA_B.v(111[10:22])
    defparam LessThan_11_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut (.I0(duty[15]), .I1(duty[20]), .I2(n321), .I3(GND_net), 
            .O(n12_adj_5409));   // verilog/TinyFPGA_B.v(122[11:24])
    defparam i2_3_lut.LUT_INIT = 16'h7e7e;
    SB_LUT4 i33939_4_lut (.I0(duty[3]), .I1(duty[2]), .I2(n334), .I3(n335), 
            .O(n49526));
    defparam i33939_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 LessThan_18_i9_rep_162_2_lut (.I0(duty[4]), .I1(n333), .I2(GND_net), 
            .I3(GND_net), .O(n51703));   // verilog/TinyFPGA_B.v(122[11:24])
    defparam LessThan_18_i9_rep_162_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i33931_4_lut (.I0(duty[5]), .I1(n51703), .I2(n332), .I3(n49526), 
            .O(n49518));
    defparam i33931_4_lut.LUT_INIT = 16'h5a7b;
    SB_LUT4 LessThan_18_i13_rep_186_2_lut (.I0(duty[6]), .I1(n331), .I2(GND_net), 
            .I3(GND_net), .O(n51727));   // verilog/TinyFPGA_B.v(122[11:24])
    defparam LessThan_18_i13_rep_186_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i34496_4_lut (.I0(duty[7]), .I1(n51727), .I2(n330), .I3(n49518), 
            .O(n50084));
    defparam i34496_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 LessThan_18_i17_rep_168_2_lut (.I0(duty[8]), .I1(n329), .I2(GND_net), 
            .I3(GND_net), .O(n51709));   // verilog/TinyFPGA_B.v(122[11:24])
    defparam LessThan_18_i17_rep_168_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i34249_4_lut (.I0(duty[9]), .I1(n51709), .I2(n328), .I3(n50084), 
            .O(n49837));
    defparam i34249_4_lut.LUT_INIT = 16'hdeff;
    SB_LUT4 LessThan_18_i21_rep_159_2_lut (.I0(duty[10]), .I1(n327), .I2(GND_net), 
            .I3(GND_net), .O(n51700));   // verilog/TinyFPGA_B.v(122[11:24])
    defparam LessThan_18_i21_rep_159_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 unary_minus_19_inv_0_i20_1_lut (.I0(duty[19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_5256));   // verilog/TinyFPGA_B.v(123[25:30])
    defparam unary_minus_19_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 LessThan_18_i10_3_lut (.I0(n332), .I1(n331), .I2(duty[6]), 
            .I3(GND_net), .O(n10_adj_5371));   // verilog/TinyFPGA_B.v(122[11:24])
    defparam LessThan_18_i10_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i33926_4_lut (.I0(duty[6]), .I1(duty[5]), .I2(n331), .I3(n332), 
            .O(n49513));
    defparam i33926_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 LessThan_18_i15_rep_151_2_lut (.I0(duty[7]), .I1(n330), .I2(GND_net), 
            .I3(GND_net), .O(n51692));   // verilog/TinyFPGA_B.v(122[11:24])
    defparam LessThan_18_i15_rep_151_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i12_1_lut (.I0(encoder0_position[11]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n22_adj_5431));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i13_1_lut (.I0(encoder0_position[12]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n21_adj_5430));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i14_1_lut (.I0(encoder0_position[13]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n20_adj_5429));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_DFFESR delay_counter_i0_i11 (.Q(delay_counter[11]), .C(CLK_c), .E(n7417), 
            .D(n1317), .R(n28933));   // verilog/TinyFPGA_B.v(375[10] 403[6])
    SB_DFFESR delay_counter_i0_i12 (.Q(delay_counter[12]), .C(CLK_c), .E(n7417), 
            .D(n1316), .R(n28933));   // verilog/TinyFPGA_B.v(375[10] 403[6])
    SB_DFFESR delay_counter_i0_i13 (.Q(delay_counter[13]), .C(CLK_c), .E(n7417), 
            .D(n1315), .R(n28933));   // verilog/TinyFPGA_B.v(375[10] 403[6])
    SB_DFFESR delay_counter_i0_i14 (.Q(delay_counter[14]), .C(CLK_c), .E(n7417), 
            .D(n1314), .R(n28933));   // verilog/TinyFPGA_B.v(375[10] 403[6])
    SB_DFFESR delay_counter_i0_i15 (.Q(delay_counter[15]), .C(CLK_c), .E(n7417), 
            .D(n1313), .R(n28933));   // verilog/TinyFPGA_B.v(375[10] 403[6])
    SB_DFFESR delay_counter_i0_i16 (.Q(delay_counter[16]), .C(CLK_c), .E(n7417), 
            .D(n1312), .R(n28933));   // verilog/TinyFPGA_B.v(375[10] 403[6])
    SB_DFFESR delay_counter_i0_i17 (.Q(delay_counter[17]), .C(CLK_c), .E(n7417), 
            .D(n1311), .R(n28933));   // verilog/TinyFPGA_B.v(375[10] 403[6])
    SB_DFFESR delay_counter_i0_i18 (.Q(delay_counter[18]), .C(CLK_c), .E(n7417), 
            .D(n1310), .R(n28933));   // verilog/TinyFPGA_B.v(375[10] 403[6])
    SB_DFFESR delay_counter_i0_i19 (.Q(delay_counter[19]), .C(CLK_c), .E(n7417), 
            .D(n1309), .R(n28933));   // verilog/TinyFPGA_B.v(375[10] 403[6])
    SB_DFFESR delay_counter_i0_i20 (.Q(delay_counter[20]), .C(CLK_c), .E(n7417), 
            .D(n1308), .R(n28933));   // verilog/TinyFPGA_B.v(375[10] 403[6])
    SB_DFFESR delay_counter_i0_i21 (.Q(delay_counter[21]), .C(CLK_c), .E(n7417), 
            .D(n1307), .R(n28933));   // verilog/TinyFPGA_B.v(375[10] 403[6])
    SB_DFFESR delay_counter_i0_i22 (.Q(delay_counter[22]), .C(CLK_c), .E(n7417), 
            .D(n1306), .R(n28933));   // verilog/TinyFPGA_B.v(375[10] 403[6])
    SB_DFFESR delay_counter_i0_i23 (.Q(delay_counter[23]), .C(CLK_c), .E(n7417), 
            .D(n1305), .R(n28933));   // verilog/TinyFPGA_B.v(375[10] 403[6])
    SB_DFFESR delay_counter_i0_i24 (.Q(delay_counter[24]), .C(CLK_c), .E(n7417), 
            .D(n1304), .R(n28933));   // verilog/TinyFPGA_B.v(375[10] 403[6])
    SB_DFFESR delay_counter_i0_i25 (.Q(delay_counter[25]), .C(CLK_c), .E(n7417), 
            .D(n1303), .R(n28933));   // verilog/TinyFPGA_B.v(375[10] 403[6])
    SB_DFFESR delay_counter_i0_i26 (.Q(delay_counter[26]), .C(CLK_c), .E(n7417), 
            .D(n1302), .R(n28933));   // verilog/TinyFPGA_B.v(375[10] 403[6])
    SB_DFFESR delay_counter_i0_i27 (.Q(delay_counter[27]), .C(CLK_c), .E(n7417), 
            .D(n1301), .R(n28933));   // verilog/TinyFPGA_B.v(375[10] 403[6])
    SB_DFFESR delay_counter_i0_i28 (.Q(delay_counter[28]), .C(CLK_c), .E(n7417), 
            .D(n1300), .R(n28933));   // verilog/TinyFPGA_B.v(375[10] 403[6])
    SB_LUT4 LessThan_18_i4_3_lut (.I0(n49289), .I1(n336), .I2(duty[1]), 
            .I3(GND_net), .O(n4_adj_5374));   // verilog/TinyFPGA_B.v(122[11:24])
    defparam LessThan_18_i4_3_lut.LUT_INIT = 16'h8e8e;
    SB_DFFESR delay_counter_i0_i29 (.Q(delay_counter[29]), .C(CLK_c), .E(n7417), 
            .D(n1299), .R(n28933));   // verilog/TinyFPGA_B.v(375[10] 403[6])
    SB_DFFESR delay_counter_i0_i30 (.Q(delay_counter[30]), .C(CLK_c), .E(n7417), 
            .D(n1298), .R(n28933));   // verilog/TinyFPGA_B.v(375[10] 403[6])
    SB_DFFESR delay_counter_i0_i31 (.Q(delay_counter[31]), .C(CLK_c), .E(n7417), 
            .D(n1297), .R(n28933));   // verilog/TinyFPGA_B.v(375[10] 403[6])
    SB_LUT4 LessThan_18_i12_3_lut (.I0(n10_adj_5371), .I1(n330), .I2(duty[7]), 
            .I3(GND_net), .O(n12_adj_5370));   // verilog/TinyFPGA_B.v(122[11:24])
    defparam LessThan_18_i12_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i15_1_lut (.I0(encoder0_position[14]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n19_adj_5428));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i16_1_lut (.I0(encoder0_position[15]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n18_adj_5427));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i34144_3_lut (.I0(n15), .I1(n13_adj_5376), .I2(n11), .I3(GND_net), 
            .O(n49732));
    defparam i34144_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i34131_4_lut (.I0(current[15]), .I1(duty[13]), .I2(duty[14]), 
            .I3(n49732), .O(n49719));
    defparam i34131_4_lut.LUT_INIT = 16'h7eff;
    SB_LUT4 i34422_4_lut (.I0(current[15]), .I1(duty[16]), .I2(duty[17]), 
            .I3(n15), .O(n50010));
    defparam i34422_4_lut.LUT_INIT = 16'hff7e;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i17_1_lut (.I0(encoder0_position[16]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n17_adj_5426));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 LessThan_11_i30_4_lut (.I0(duty[7]), .I1(duty[17]), .I2(current[15]), 
            .I3(duty[16]), .O(n30_adj_5369));   // verilog/TinyFPGA_B.v(111[10:22])
    defparam LessThan_11_i30_4_lut.LUT_INIT = 16'h8f0e;
    SB_LUT4 i34148_4_lut (.I0(n9_adj_5375), .I1(n7_adj_5387), .I2(current[2]), 
            .I3(duty[2]), .O(n49736));
    defparam i34148_4_lut.LUT_INIT = 16'heffe;
    SB_LUT4 unary_minus_19_inv_0_i21_1_lut (.I0(duty[20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n5));   // verilog/TinyFPGA_B.v(123[25:30])
    defparam unary_minus_19_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i34436_4_lut (.I0(n15), .I1(n13_adj_5376), .I2(n11), .I3(n49736), 
            .O(n50024));
    defparam i34436_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i34434_4_lut (.I0(n21_adj_5279), .I1(n19_adj_5277), .I2(n17), 
            .I3(n50024), .O(n50022));
    defparam i34434_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i34724_4_lut (.I0(current[15]), .I1(n23), .I2(duty[12]), .I3(n50022), 
            .O(n50312));
    defparam i34724_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i18_1_lut (.I0(encoder0_position[17]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n16_adj_5425));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i19_1_lut (.I0(encoder0_position[18]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n15_adj_5424));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i34134_4_lut (.I0(current[15]), .I1(duty[13]), .I2(duty[14]), 
            .I3(n50312), .O(n49722));
    defparam i34134_4_lut.LUT_INIT = 16'h7eff;
    SB_LUT4 i34614_4_lut (.I0(current[15]), .I1(duty[15]), .I2(duty[16]), 
            .I3(n49722), .O(n50202));
    defparam i34614_4_lut.LUT_INIT = 16'hff7e;
    SB_LUT4 i34786_4_lut (.I0(current[15]), .I1(duty[17]), .I2(duty[18]), 
            .I3(n50202), .O(n50374));
    defparam i34786_4_lut.LUT_INIT = 16'hff7e;
    SB_LUT4 i15219_3_lut (.I0(Ki[15]), .I1(\data_in_frame[4] [7]), .I2(n28521), 
            .I3(GND_net), .O(n29167));   // verilog/coms.v(128[12] 303[6])
    defparam i15219_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34864_4_lut (.I0(current[15]), .I1(duty[19]), .I2(duty[20]), 
            .I3(n50374), .O(n50452));
    defparam i34864_4_lut.LUT_INIT = 16'hff7e;
    SB_LUT4 i15220_3_lut (.I0(Ki[14]), .I1(\data_in_frame[4] [6]), .I2(n28521), 
            .I3(GND_net), .O(n29168));   // verilog/coms.v(128[12] 303[6])
    defparam i15220_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15221_3_lut (.I0(Ki[13]), .I1(\data_in_frame[4] [5]), .I2(n28521), 
            .I3(GND_net), .O(n29169));   // verilog/coms.v(128[12] 303[6])
    defparam i15221_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5502_3_lut_4_lut (.I0(commutation_state[2]), .I1(commutation_state[1]), 
            .I2(commutation_state[0]), .I3(dir), .O(GHC_N_427));   // verilog/TinyFPGA_B.v(201[7] 220[14])
    defparam i5502_3_lut_4_lut.LUT_INIT = 16'h21cc;
    SB_LUT4 i15222_3_lut (.I0(Ki[12]), .I1(\data_in_frame[4] [4]), .I2(n28521), 
            .I3(GND_net), .O(n29170));   // verilog/coms.v(128[12] 303[6])
    defparam i15222_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i33787_4_lut (.I0(n21_adj_5279), .I1(n19_adj_5277), .I2(n17), 
            .I3(n9_adj_5375), .O(n49374));
    defparam i33787_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i34231_4_lut (.I0(current[15]), .I1(duty[21]), .I2(duty[22]), 
            .I3(n19_adj_5277), .O(n49819));
    defparam i34231_4_lut.LUT_INIT = 16'hff7e;
    SB_LUT4 i5504_3_lut_4_lut (.I0(commutation_state[2]), .I1(commutation_state[1]), 
            .I2(commutation_state[0]), .I3(dir), .O(GLC_N_436));   // verilog/TinyFPGA_B.v(201[7] 220[14])
    defparam i5504_3_lut_4_lut.LUT_INIT = 16'hcc21;
    SB_LUT4 LessThan_11_i24_4_lut (.I0(duty[9]), .I1(duty[22]), .I2(current[15]), 
            .I3(duty[21]), .O(n24_adj_5377));   // verilog/TinyFPGA_B.v(111[10:22])
    defparam LessThan_11_i24_4_lut.LUT_INIT = 16'h8f0e;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i20_1_lut (.I0(encoder0_position[19]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n14_adj_5423));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i15071_3_lut (.I0(\data_out_frame[13] [0]), .I1(setpoint[8]), 
            .I2(n24278), .I3(GND_net), .O(n29019));   // verilog/coms.v(128[12] 303[6])
    defparam i15071_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i21_1_lut (.I0(encoder0_position[20]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n13_adj_5422));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i34652_3_lut (.I0(n6_adj_5242), .I1(duty[10]), .I2(n21_adj_5279), 
            .I3(GND_net), .O(n50240));   // verilog/TinyFPGA_B.v(111[10:22])
    defparam i34652_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34653_3_lut (.I0(n50240), .I1(duty[11]), .I2(n23), .I3(GND_net), 
            .O(n50241));   // verilog/TinyFPGA_B.v(111[10:22])
    defparam i34653_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15159_3_lut (.I0(\data_out_frame[7] [0]), .I1(encoder0_position_scaled[8]), 
            .I2(n24278), .I3(GND_net), .O(n29107));   // verilog/coms.v(128[12] 303[6])
    defparam i15159_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15223_3_lut (.I0(Ki[11]), .I1(\data_in_frame[4] [3]), .I2(n28521), 
            .I3(GND_net), .O(n29171));   // verilog/coms.v(128[12] 303[6])
    defparam i15223_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34432_4_lut (.I0(current[15]), .I1(n23), .I2(duty[12]), .I3(n49374), 
            .O(n50020));
    defparam i34432_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 i34414_4_lut (.I0(current[15]), .I1(duty[21]), .I2(duty[22]), 
            .I3(n50020), .O(n50002));
    defparam i34414_4_lut.LUT_INIT = 16'h7eff;
    SB_LUT4 i34626_3_lut (.I0(n24_adj_5377), .I1(n8_adj_5342), .I2(n49819), 
            .I3(GND_net), .O(n50214));   // verilog/TinyFPGA_B.v(111[10:22])
    defparam i34626_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i34633_3_lut (.I0(n50241), .I1(duty[12]), .I2(current[15]), 
            .I3(GND_net), .O(n50221));   // verilog/TinyFPGA_B.v(111[10:22])
    defparam i34633_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 dti_counter_2244_add_4_9_lut (.I0(n49292), .I1(n34648), .I2(dti_counter[7]), 
            .I3(n39313), .O(n48)) /* synthesis syn_instantiated=1 */ ;
    defparam dti_counter_2244_add_4_9_lut.LUT_INIT = 16'hE22E;
    SB_LUT4 LessThan_18_i8_3_lut (.I0(n333), .I1(n329), .I2(duty[8]), 
            .I3(GND_net), .O(n8_adj_5372));   // verilog/TinyFPGA_B.v(122[11:24])
    defparam LessThan_18_i8_3_lut.LUT_INIT = 16'h8e8e;
    SB_DFFESR delay_counter_i0_i5 (.Q(delay_counter[5]), .C(CLK_c), .E(n7417), 
            .D(n1323), .R(n28933));   // verilog/TinyFPGA_B.v(375[10] 403[6])
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i22_1_lut (.I0(encoder0_position[21]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n12_adj_5421));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i23_1_lut (.I0(encoder0_position[22]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n11_adj_5420));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i15160_3_lut (.I0(\data_out_frame[6] [7]), .I1(encoder0_position_scaled[23]), 
            .I2(n24278), .I3(GND_net), .O(n29108));   // verilog/coms.v(128[12] 303[6])
    defparam i15160_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i24_1_lut (.I0(encoder0_position[23]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n10_adj_5419));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i15224_3_lut (.I0(Ki[10]), .I1(\data_in_frame[4] [2]), .I2(n28521), 
            .I3(GND_net), .O(n29172));   // verilog/coms.v(128[12] 303[6])
    defparam i15224_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15161_3_lut (.I0(\data_out_frame[6] [6]), .I1(encoder0_position_scaled[22]), 
            .I2(n24278), .I3(GND_net), .O(n29109));   // verilog/coms.v(128[12] 303[6])
    defparam i15161_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i25_1_lut (.I0(encoder0_position[24]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n9_adj_5418));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i25_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i15225_3_lut (.I0(Ki[9]), .I1(\data_in_frame[4] [1]), .I2(n28521), 
            .I3(GND_net), .O(n29173));   // verilog/coms.v(128[12] 303[6])
    defparam i15225_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 dti_counter_2244_add_4_8_lut (.I0(n49293), .I1(n34648), .I2(dti_counter[6]), 
            .I3(n39312), .O(n49)) /* synthesis syn_instantiated=1 */ ;
    defparam dti_counter_2244_add_4_8_lut.LUT_INIT = 16'hE22E;
    SB_LUT4 i15226_3_lut (.I0(Ki[8]), .I1(\data_in_frame[4] [0]), .I2(n28521), 
            .I3(GND_net), .O(n29174));   // verilog/coms.v(128[12] 303[6])
    defparam i15226_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15162_3_lut (.I0(\data_out_frame[6] [5]), .I1(encoder0_position_scaled[21]), 
            .I2(n24278), .I3(GND_net), .O(n29110));   // verilog/coms.v(128[12] 303[6])
    defparam i15162_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i33914_4_lut (.I0(duty[8]), .I1(duty[4]), .I2(n329), .I3(n333), 
            .O(n49501));
    defparam i33914_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 i15163_3_lut (.I0(\data_out_frame[6] [4]), .I1(encoder0_position_scaled[20]), 
            .I2(n24278), .I3(GND_net), .O(n29111));   // verilog/coms.v(128[12] 303[6])
    defparam i15163_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15164_3_lut (.I0(\data_out_frame[6] [3]), .I1(encoder0_position_scaled[19]), 
            .I2(n24278), .I3(GND_net), .O(n29112));   // verilog/coms.v(128[12] 303[6])
    defparam i15164_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY dti_counter_2244_add_4_8 (.CI(n39312), .I0(n34648), .I1(dti_counter[6]), 
            .CO(n39313));
    SB_LUT4 dti_counter_2244_add_4_7_lut (.I0(n49294), .I1(n34648), .I2(dti_counter[5]), 
            .I3(n39311), .O(n50)) /* synthesis syn_instantiated=1 */ ;
    defparam dti_counter_2244_add_4_7_lut.LUT_INIT = 16'hE22E;
    SB_LUT4 LessThan_18_i19_rep_164_2_lut (.I0(duty[9]), .I1(n328), .I2(GND_net), 
            .I3(GND_net), .O(n51705));   // verilog/TinyFPGA_B.v(122[11:24])
    defparam LessThan_18_i19_rep_164_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i15165_3_lut (.I0(\data_out_frame[6] [2]), .I1(encoder0_position_scaled[18]), 
            .I2(n24278), .I3(GND_net), .O(n29113));   // verilog/coms.v(128[12] 303[6])
    defparam i15165_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15227_3_lut (.I0(Ki[7]), .I1(\data_in_frame[5] [7]), .I2(n28521), 
            .I3(GND_net), .O(n29175));   // verilog/coms.v(128[12] 303[6])
    defparam i15227_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15166_3_lut (.I0(\data_out_frame[6] [1]), .I1(encoder0_position_scaled[17]), 
            .I2(n24278), .I3(GND_net), .O(n29114));   // verilog/coms.v(128[12] 303[6])
    defparam i15166_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15167_3_lut (.I0(\data_out_frame[6] [0]), .I1(encoder0_position_scaled[16]), 
            .I2(n24278), .I3(GND_net), .O(n29115));   // verilog/coms.v(128[12] 303[6])
    defparam i15167_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15168_3_lut (.I0(\data_out_frame[5] [7]), .I1(control_mode[7]), 
            .I2(n24278), .I3(GND_net), .O(n29116));   // verilog/coms.v(128[12] 303[6])
    defparam i15168_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i35496_1_lut (.I0(n1257), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n51084));
    defparam i35496_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_19_inv_0_i22_1_lut (.I0(duty[21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_5255));   // verilog/TinyFPGA_B.v(123[25:30])
    defparam unary_minus_19_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i15228_3_lut (.I0(Ki[6]), .I1(\data_in_frame[5] [6]), .I2(n28521), 
            .I3(GND_net), .O(n29176));   // verilog/coms.v(128[12] 303[6])
    defparam i15228_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15229_3_lut (.I0(Ki[5]), .I1(\data_in_frame[5] [5]), .I2(n28521), 
            .I3(GND_net), .O(n29177));   // verilog/coms.v(128[12] 303[6])
    defparam i15229_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15169_3_lut (.I0(\data_out_frame[5] [6]), .I1(control_mode[6]), 
            .I2(n24278), .I3(GND_net), .O(n29117));   // verilog/coms.v(128[12] 303[6])
    defparam i15169_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15170_3_lut (.I0(\data_out_frame[5] [5]), .I1(control_mode[5]), 
            .I2(n24278), .I3(GND_net), .O(n29118));   // verilog/coms.v(128[12] 303[6])
    defparam i15170_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15171_3_lut (.I0(\data_out_frame[5] [4]), .I1(control_mode[4]), 
            .I2(n24278), .I3(GND_net), .O(n29119));   // verilog/coms.v(128[12] 303[6])
    defparam i15171_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i26_1_lut (.I0(encoder0_position[25]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n8_adj_5417));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i26_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i15172_3_lut (.I0(\data_out_frame[5] [3]), .I1(control_mode[3]), 
            .I2(n24278), .I3(GND_net), .O(n29120));   // verilog/coms.v(128[12] 303[6])
    defparam i15172_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15173_3_lut (.I0(\data_out_frame[5] [2]), .I1(control_mode[2]), 
            .I2(n24278), .I3(GND_net), .O(n29121));   // verilog/coms.v(128[12] 303[6])
    defparam i15173_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15174_3_lut (.I0(\data_out_frame[5] [1]), .I1(control_mode[1]), 
            .I2(n24278), .I3(GND_net), .O(n29122));   // verilog/coms.v(128[12] 303[6])
    defparam i15174_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15175_3_lut (.I0(\data_out_frame[5] [0]), .I1(control_mode[0]), 
            .I2(n24278), .I3(GND_net), .O(n29123));   // verilog/coms.v(128[12] 303[6])
    defparam i15175_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_18_i6_3_lut (.I0(n335), .I1(n334), .I2(duty[3]), 
            .I3(GND_net), .O(n6_adj_5373));   // verilog/TinyFPGA_B.v(122[11:24])
    defparam LessThan_18_i6_3_lut.LUT_INIT = 16'h8e8e;
    SB_CARRY dti_counter_2244_add_4_7 (.CI(n39311), .I0(n34648), .I1(dti_counter[5]), 
            .CO(n39312));
    SB_LUT4 dti_counter_2244_add_4_6_lut (.I0(n49295), .I1(n34648), .I2(dti_counter[4]), 
            .I3(n39310), .O(n51)) /* synthesis syn_instantiated=1 */ ;
    defparam dti_counter_2244_add_4_6_lut.LUT_INIT = 16'hE22E;
    SB_CARRY dti_counter_2244_add_4_6 (.CI(n39310), .I0(n34648), .I1(dti_counter[4]), 
            .CO(n39311));
    SB_LUT4 i15176_3_lut (.I0(\data_out_frame[4] [7]), .I1(ID[7]), .I2(n24278), 
            .I3(GND_net), .O(n29124));   // verilog/coms.v(128[12] 303[6])
    defparam i15176_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15230_3_lut (.I0(Ki[4]), .I1(\data_in_frame[5] [4]), .I2(n28521), 
            .I3(GND_net), .O(n29178));   // verilog/coms.v(128[12] 303[6])
    defparam i15230_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_18_i16_3_lut (.I0(n8_adj_5372), .I1(n328), .I2(duty[9]), 
            .I3(GND_net), .O(n16_adj_5351));   // verilog/TinyFPGA_B.v(122[11:24])
    defparam LessThan_18_i16_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i34776_4_lut (.I0(n16_adj_5351), .I1(n6_adj_5373), .I2(n51705), 
            .I3(n49501), .O(n50364));   // verilog/TinyFPGA_B.v(122[11:24])
    defparam i34776_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i34777_3_lut (.I0(n50364), .I1(n327), .I2(duty[10]), .I3(GND_net), 
            .O(n50365));   // verilog/TinyFPGA_B.v(122[11:24])
    defparam i34777_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i34727_3_lut (.I0(n50365), .I1(n326), .I2(duty[11]), .I3(GND_net), 
            .O(n50315));   // verilog/TinyFPGA_B.v(122[11:24])
    defparam i34727_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i6_4_lut (.I0(duty[13]), .I1(n12_adj_5409), .I2(duty[21]), 
            .I3(n321), .O(n16_adj_5405));   // verilog/TinyFPGA_B.v(122[11:24])
    defparam i6_4_lut.LUT_INIT = 16'hdffe;
    SB_LUT4 i4_3_lut (.I0(duty[19]), .I1(duty[16]), .I2(n321), .I3(GND_net), 
            .O(n14_adj_5407));   // verilog/TinyFPGA_B.v(122[11:24])
    defparam i4_3_lut.LUT_INIT = 16'h7e7e;
    SB_LUT4 i5_3_lut (.I0(duty[14]), .I1(duty[18]), .I2(n321), .I3(GND_net), 
            .O(n15_adj_5406));   // verilog/TinyFPGA_B.v(122[11:24])
    defparam i5_3_lut.LUT_INIT = 16'h7e7e;
    SB_LUT4 i3_3_lut (.I0(duty[22]), .I1(duty[17]), .I2(n321), .I3(GND_net), 
            .O(n13_adj_5408));   // verilog/TinyFPGA_B.v(122[11:24])
    defparam i3_3_lut.LUT_INIT = 16'h7e7e;
    SB_LUT4 i34668_4_lut (.I0(duty[11]), .I1(n51700), .I2(n326), .I3(n49837), 
            .O(n50256));
    defparam i34668_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 dti_counter_2244_add_4_5_lut (.I0(n49296), .I1(n34648), .I2(dti_counter[3]), 
            .I3(n39309), .O(n52)) /* synthesis syn_instantiated=1 */ ;
    defparam dti_counter_2244_add_4_5_lut.LUT_INIT = 16'hE22E;
    SB_LUT4 i15597_3_lut (.I0(current[9]), .I1(data_adj_5514[9]), .I2(n28537), 
            .I3(GND_net), .O(n29545));   // verilog/tli4970.v(35[10] 68[6])
    defparam i15597_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_18_i25_rep_156_2_lut (.I0(duty[12]), .I1(n325), .I2(GND_net), 
            .I3(GND_net), .O(n51697));   // verilog/TinyFPGA_B.v(122[11:24])
    defparam LessThan_18_i25_rep_156_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i15231_3_lut (.I0(Ki[3]), .I1(\data_in_frame[5] [3]), .I2(n28521), 
            .I3(GND_net), .O(n29179));   // verilog/coms.v(128[12] 303[6])
    defparam i15231_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14_3_lut (.I0(h2), .I1(h3), .I2(h1), .I3(GND_net), .O(n6_adj_5454));
    defparam i14_3_lut.LUT_INIT = 16'h7e7e;
    SB_LUT4 i1_3_lut_adj_1749 (.I0(h3), .I1(h2), .I2(h1), .I3(GND_net), 
            .O(commutation_state_7__N_240[0]));   // verilog/TinyFPGA_B.v(164[4] 166[7])
    defparam i1_3_lut_adj_1749.LUT_INIT = 16'h1414;
    SB_LUT4 i15440_3_lut (.I0(\data_in_frame[6] [7]), .I1(rx_data[7]), .I2(n43839), 
            .I3(GND_net), .O(n29388));   // verilog/coms.v(128[12] 303[6])
    defparam i15440_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15441_3_lut (.I0(\data_in_frame[6] [6]), .I1(rx_data[6]), .I2(n43839), 
            .I3(GND_net), .O(n29389));   // verilog/coms.v(128[12] 303[6])
    defparam i15441_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15232_3_lut (.I0(Ki[2]), .I1(\data_in_frame[5] [2]), .I2(n28521), 
            .I3(GND_net), .O(n29180));   // verilog/coms.v(128[12] 303[6])
    defparam i15232_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY dti_counter_2244_add_4_5 (.CI(n39309), .I0(n34648), .I1(dti_counter[3]), 
            .CO(n39310));
    SB_LUT4 dti_counter_2244_add_4_4_lut (.I0(n49297), .I1(n34648), .I2(dti_counter[2]), 
            .I3(n39308), .O(n53)) /* synthesis syn_instantiated=1 */ ;
    defparam dti_counter_2244_add_4_4_lut.LUT_INIT = 16'hE22E;
    SB_LUT4 i35080_1_lut (.I0(n2841), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n50668));
    defparam i35080_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i34650_4_lut (.I0(n12_adj_5370), .I1(n4_adj_5374), .I2(n51692), 
            .I3(n49513), .O(n50238));   // verilog/TinyFPGA_B.v(122[11:24])
    defparam i34650_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i15442_3_lut (.I0(\data_in_frame[6] [5]), .I1(rx_data[5]), .I2(n43839), 
            .I3(GND_net), .O(n29390));   // verilog/coms.v(128[12] 303[6])
    defparam i15442_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15233_3_lut (.I0(Ki[1]), .I1(\data_in_frame[5] [1]), .I2(n28521), 
            .I3(GND_net), .O(n29181));   // verilog/coms.v(128[12] 303[6])
    defparam i15233_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34441_3_lut (.I0(n50315), .I1(n325), .I2(duty[12]), .I3(GND_net), 
            .O(n50029));   // verilog/TinyFPGA_B.v(122[11:24])
    defparam i34441_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i15443_3_lut (.I0(\data_in_frame[6] [4]), .I1(rx_data[4]), .I2(n43839), 
            .I3(GND_net), .O(n29391));   // verilog/coms.v(128[12] 303[6])
    defparam i15443_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i9_4_lut (.I0(n13_adj_5408), .I1(n15_adj_5406), .I2(n14_adj_5407), 
            .I3(n16_adj_5405), .O(n45203));   // verilog/TinyFPGA_B.v(122[11:24])
    defparam i9_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i34768_4_lut (.I0(n50029), .I1(n50238), .I2(n51697), .I3(n50256), 
            .O(n50356));   // verilog/TinyFPGA_B.v(122[11:24])
    defparam i34768_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 mux_250_i1_4_lut (.I0(encoder1_position_scaled[0]), .I1(displacement[0]), 
            .I2(n15_adj_5249), .I3(n15_adj_5321), .O(motor_state_23__N_123[0]));   // verilog/TinyFPGA_B.v(285[5] 287[10])
    defparam mux_250_i1_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_250_i2_4_lut (.I0(encoder1_position_scaled[1]), .I1(displacement[1]), 
            .I2(n15_adj_5249), .I3(n15_adj_5321), .O(motor_state_23__N_123[1]));   // verilog/TinyFPGA_B.v(285[5] 287[10])
    defparam mux_250_i2_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 LessThan_11_i4_4_lut (.I0(duty[0]), .I1(duty[1]), .I2(current[1]), 
            .I3(current[0]), .O(n4_adj_5285));   // verilog/TinyFPGA_B.v(111[10:22])
    defparam LessThan_11_i4_4_lut.LUT_INIT = 16'h0c8e;
    SB_DFFESR delay_counter_i0_i6 (.Q(delay_counter[6]), .C(CLK_c), .E(n7417), 
            .D(n1322), .R(n28933));   // verilog/TinyFPGA_B.v(375[10] 403[6])
    SB_LUT4 mux_1005_i1_3_lut (.I0(duty[0]), .I1(n363), .I2(duty[23]), 
            .I3(GND_net), .O(n4723));   // verilog/TinyFPGA_B.v(118[13] 129[7])
    defparam mux_1005_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34654_3_lut (.I0(n4_adj_5285), .I1(duty[13]), .I2(current[15]), 
            .I3(GND_net), .O(n50242));   // verilog/TinyFPGA_B.v(111[10:22])
    defparam i34654_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i15444_3_lut (.I0(\data_in_frame[6] [3]), .I1(rx_data[3]), .I2(n43839), 
            .I3(GND_net), .O(n29392));   // verilog/coms.v(128[12] 303[6])
    defparam i15444_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i34126_4_lut (.I0(current[15]), .I1(duty[15]), .I2(duty[16]), 
            .I3(n49719), .O(n49713));
    defparam i34126_4_lut.LUT_INIT = 16'h5adb;
    SB_LUT4 i15234_3_lut (.I0(Kp[15]), .I1(\data_in_frame[2] [7]), .I2(n28521), 
            .I3(GND_net), .O(n29182));   // verilog/coms.v(128[12] 303[6])
    defparam i15234_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15445_3_lut (.I0(\data_in_frame[6] [2]), .I1(rx_data[2]), .I2(n43839), 
            .I3(GND_net), .O(n29393));   // verilog/coms.v(128[12] 303[6])
    defparam i15445_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 LessThan_11_i35_rep_132_2_lut (.I0(current[15]), .I1(duty[17]), 
            .I2(GND_net), .I3(GND_net), .O(n51673));   // verilog/TinyFPGA_B.v(111[10:22])
    defparam LessThan_11_i35_rep_132_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i15235_3_lut (.I0(Kp[14]), .I1(\data_in_frame[2] [6]), .I2(n28521), 
            .I3(GND_net), .O(n29183));   // verilog/coms.v(128[12] 303[6])
    defparam i15235_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15236_4_lut (.I0(CS_MISO_c), .I1(data_adj_5514[9]), .I2(n6), 
            .I3(n27167), .O(n29184));   // verilog/tli4970.v(35[10] 68[6])
    defparam i15236_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 mux_1005_i11_3_lut (.I0(duty[10]), .I1(n353), .I2(duty[23]), 
            .I3(GND_net), .O(n4713));   // verilog/TinyFPGA_B.v(118[13] 129[7])
    defparam mux_1005_i11_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15446_3_lut (.I0(\data_in_frame[6] [1]), .I1(rx_data[1]), .I2(n43839), 
            .I3(GND_net), .O(n29394));   // verilog/coms.v(128[12] 303[6])
    defparam i15446_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i34796_3_lut (.I0(n30_adj_5369), .I1(n10_adj_5275), .I2(n50010), 
            .I3(GND_net), .O(n50384));   // verilog/TinyFPGA_B.v(111[10:22])
    defparam i34796_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i34631_4_lut (.I0(n50242), .I1(duty[15]), .I2(current[15]), 
            .I3(duty[14]), .O(n28_adj_5386));   // verilog/TinyFPGA_B.v(111[10:22])
    defparam i34631_4_lut.LUT_INIT = 16'h8f0e;
    SB_LUT4 i34874_4_lut (.I0(n28_adj_5386), .I1(n50384), .I2(n51673), 
            .I3(n49713), .O(n50462));   // verilog/TinyFPGA_B.v(111[10:22])
    defparam i34874_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i34875_3_lut (.I0(n50462), .I1(duty[18]), .I2(current[15]), 
            .I3(GND_net), .O(n50463));   // verilog/TinyFPGA_B.v(111[10:22])
    defparam i34875_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i34416_4_lut (.I0(current[15]), .I1(duty[21]), .I2(duty[22]), 
            .I3(n50452), .O(n50004));
    defparam i34416_4_lut.LUT_INIT = 16'h7eff;
    SB_LUT4 i34788_3_lut (.I0(n50221), .I1(n50214), .I2(n50002), .I3(GND_net), 
            .O(n50376));   // verilog/TinyFPGA_B.v(111[10:22])
    defparam i34788_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34629_4_lut (.I0(n50463), .I1(duty[20]), .I2(current[15]), 
            .I3(duty[19]), .O(n50217));   // verilog/TinyFPGA_B.v(111[10:22])
    defparam i34629_4_lut.LUT_INIT = 16'h8f0e;
    SB_LUT4 i34838_3_lut (.I0(n50217), .I1(n50376), .I2(n50004), .I3(GND_net), 
            .O(n50426));   // verilog/TinyFPGA_B.v(111[10:22])
    defparam i34838_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34731_4_lut (.I0(n50356), .I1(duty[23]), .I2(n321), .I3(n45203), 
            .O(n50319));   // verilog/TinyFPGA_B.v(122[11:24])
    defparam i34731_4_lut.LUT_INIT = 16'hcc8e;
    SB_LUT4 i34839_3_lut (.I0(n50426), .I1(current[15]), .I2(duty[23]), 
            .I3(GND_net), .O(n50427));   // verilog/TinyFPGA_B.v(111[10:22])
    defparam i34839_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i15447_3_lut (.I0(\data_in_frame[6] [0]), .I1(rx_data[0]), .I2(n43839), 
            .I3(GND_net), .O(n29395));   // verilog/coms.v(128[12] 303[6])
    defparam i15447_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14877_4_lut (.I0(n50427), .I1(n50319), .I2(duty[23]), .I3(n287), 
            .O(n4208));
    defparam i14877_4_lut.LUT_INIT = 16'h0f35;
    SB_LUT4 i3_4_lut (.I0(\ID_READOUT_FSM.state [1]), .I1(n62), .I2(delay_counter[31]), 
            .I3(\ID_READOUT_FSM.state [0]), .O(n46412));
    defparam i3_4_lut.LUT_INIT = 16'h0004;
    SB_LUT4 i15239_3_lut (.I0(Kp[13]), .I1(\data_in_frame[2] [5]), .I2(n28521), 
            .I3(GND_net), .O(n29187));   // verilog/coms.v(128[12] 303[6])
    defparam i15239_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15240_3_lut (.I0(Kp[12]), .I1(\data_in_frame[2] [4]), .I2(n28521), 
            .I3(GND_net), .O(n29188));   // verilog/coms.v(128[12] 303[6])
    defparam i15240_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15448_3_lut (.I0(\data_in_frame[5] [7]), .I1(rx_data[7]), .I2(n43838), 
            .I3(GND_net), .O(n29396));   // verilog/coms.v(128[12] 303[6])
    defparam i15448_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15449_3_lut (.I0(\data_in_frame[5] [6]), .I1(rx_data[6]), .I2(n43838), 
            .I3(GND_net), .O(n29397));   // verilog/coms.v(128[12] 303[6])
    defparam i15449_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15241_3_lut (.I0(Kp[11]), .I1(\data_in_frame[2] [3]), .I2(n28521), 
            .I3(GND_net), .O(n29189));   // verilog/coms.v(128[12] 303[6])
    defparam i15241_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15242_3_lut (.I0(Kp[10]), .I1(\data_in_frame[2] [2]), .I2(n28521), 
            .I3(GND_net), .O(n29190));   // verilog/coms.v(128[12] 303[6])
    defparam i15242_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15243_3_lut (.I0(Kp[9]), .I1(\data_in_frame[2] [1]), .I2(n28521), 
            .I3(GND_net), .O(n29191));   // verilog/coms.v(128[12] 303[6])
    defparam i15243_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15450_3_lut (.I0(\data_in_frame[5] [5]), .I1(rx_data[5]), .I2(n43838), 
            .I3(GND_net), .O(n29398));   // verilog/coms.v(128[12] 303[6])
    defparam i15450_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15451_3_lut (.I0(\data_in_frame[5] [4]), .I1(rx_data[4]), .I2(n43838), 
            .I3(GND_net), .O(n29399));   // verilog/coms.v(128[12] 303[6])
    defparam i15451_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15244_3_lut (.I0(Kp[8]), .I1(\data_in_frame[2] [0]), .I2(n28521), 
            .I3(GND_net), .O(n29192));   // verilog/coms.v(128[12] 303[6])
    defparam i15244_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15245_3_lut (.I0(Kp[7]), .I1(\data_in_frame[3] [7]), .I2(n28521), 
            .I3(GND_net), .O(n29193));   // verilog/coms.v(128[12] 303[6])
    defparam i15245_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15246_3_lut (.I0(Kp[6]), .I1(\data_in_frame[3] [6]), .I2(n28521), 
            .I3(GND_net), .O(n29194));   // verilog/coms.v(128[12] 303[6])
    defparam i15246_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15452_3_lut (.I0(\data_in_frame[5] [3]), .I1(rx_data[3]), .I2(n43838), 
            .I3(GND_net), .O(n29400));   // verilog/coms.v(128[12] 303[6])
    defparam i15452_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15247_3_lut (.I0(Kp[5]), .I1(\data_in_frame[3] [5]), .I2(n28521), 
            .I3(GND_net), .O(n29195));   // verilog/coms.v(128[12] 303[6])
    defparam i15247_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY dti_counter_2244_add_4_4 (.CI(n39308), .I0(n34648), .I1(dti_counter[2]), 
            .CO(n39309));
    SB_LUT4 i15248_3_lut (.I0(Kp[4]), .I1(\data_in_frame[3] [4]), .I2(n28521), 
            .I3(GND_net), .O(n29196));   // verilog/coms.v(128[12] 303[6])
    defparam i15248_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15249_3_lut (.I0(Kp[3]), .I1(\data_in_frame[3] [3]), .I2(n28521), 
            .I3(GND_net), .O(n29197));   // verilog/coms.v(128[12] 303[6])
    defparam i15249_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15453_3_lut (.I0(\data_in_frame[5] [2]), .I1(rx_data[2]), .I2(n43838), 
            .I3(GND_net), .O(n29401));   // verilog/coms.v(128[12] 303[6])
    defparam i15453_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15250_3_lut (.I0(Kp[2]), .I1(\data_in_frame[3] [2]), .I2(n28521), 
            .I3(GND_net), .O(n29198));   // verilog/coms.v(128[12] 303[6])
    defparam i15250_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15251_3_lut (.I0(Kp[1]), .I1(\data_in_frame[3] [1]), .I2(n28521), 
            .I3(GND_net), .O(n29199));   // verilog/coms.v(128[12] 303[6])
    defparam i15251_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_250_i3_4_lut (.I0(encoder1_position_scaled[2]), .I1(displacement[2]), 
            .I2(n15_adj_5249), .I3(n15_adj_5321), .O(motor_state_23__N_123[2]));   // verilog/TinyFPGA_B.v(285[5] 287[10])
    defparam mux_250_i3_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i15252_3_lut (.I0(\data_in[3] [7]), .I1(rx_data[7]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n29200));   // verilog/coms.v(128[12] 303[6])
    defparam i15252_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n10621_bdd_4_lut_35824 (.I0(n10621), .I1(current[15]), .I2(duty[20]), 
            .I3(n4208), .O(n51450));
    defparam n10621_bdd_4_lut_35824.LUT_INIT = 16'he4aa;
    SB_LUT4 i15454_3_lut (.I0(\data_in_frame[5] [1]), .I1(rx_data[1]), .I2(n43838), 
            .I3(GND_net), .O(n29402));   // verilog/coms.v(128[12] 303[6])
    defparam i15454_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15253_3_lut (.I0(\data_in[3] [6]), .I1(rx_data[6]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n29201));   // verilog/coms.v(128[12] 303[6])
    defparam i15253_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15254_3_lut (.I0(\data_in[3] [5]), .I1(rx_data[5]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n29202));   // verilog/coms.v(128[12] 303[6])
    defparam i15254_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1005_i2_3_lut (.I0(duty[1]), .I1(n362), .I2(duty[23]), 
            .I3(GND_net), .O(n4722));   // verilog/TinyFPGA_B.v(118[13] 129[7])
    defparam mux_1005_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15255_3_lut (.I0(\data_in[3] [4]), .I1(rx_data[4]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n29203));   // verilog/coms.v(128[12] 303[6])
    defparam i15255_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 dti_counter_2244_add_4_3_lut (.I0(n49298), .I1(n34648), .I2(dti_counter[1]), 
            .I3(n39307), .O(n54)) /* synthesis syn_instantiated=1 */ ;
    defparam dti_counter_2244_add_4_3_lut.LUT_INIT = 16'hE22E;
    SB_CARRY dti_counter_2244_add_4_3 (.CI(n39307), .I0(n34648), .I1(dti_counter[1]), 
            .CO(n39308));
    SB_LUT4 dti_counter_2244_add_4_2_lut (.I0(n49334), .I1(n2195), .I2(dti_counter[0]), 
            .I3(VCC_net), .O(n55)) /* synthesis syn_instantiated=1 */ ;
    defparam dti_counter_2244_add_4_2_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 i15256_3_lut (.I0(\data_in[3] [3]), .I1(rx_data[3]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n29204));   // verilog/coms.v(128[12] 303[6])
    defparam i15256_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15257_3_lut (.I0(\data_in[3] [2]), .I1(rx_data[2]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n29205));   // verilog/coms.v(128[12] 303[6])
    defparam i15257_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15455_3_lut (.I0(\data_in_frame[5] [0]), .I1(rx_data[0]), .I2(n43838), 
            .I3(GND_net), .O(n29403));   // verilog/coms.v(128[12] 303[6])
    defparam i15455_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15258_3_lut (.I0(\data_in[3] [1]), .I1(rx_data[1]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n29206));   // verilog/coms.v(128[12] 303[6])
    defparam i15258_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_250_i4_4_lut (.I0(encoder1_position_scaled[3]), .I1(displacement[3]), 
            .I2(n15_adj_5249), .I3(n15_adj_5321), .O(motor_state_23__N_123[3]));   // verilog/TinyFPGA_B.v(285[5] 287[10])
    defparam mux_250_i4_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i15259_3_lut (.I0(\data_in[3] [0]), .I1(rx_data[0]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n29207));   // verilog/coms.v(128[12] 303[6])
    defparam i15259_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15260_3_lut (.I0(\data_in[2] [7]), .I1(\data_in[3] [7]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n29208));   // verilog/coms.v(128[12] 303[6])
    defparam i15260_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15456_4_lut (.I0(r_Rx_Data), .I1(rx_data[1]), .I2(n4_adj_5287), 
            .I3(n27126), .O(n29404));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i15456_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 mux_250_i5_4_lut (.I0(encoder1_position_scaled[4]), .I1(displacement[4]), 
            .I2(n15_adj_5249), .I3(n15_adj_5321), .O(motor_state_23__N_123[4]));   // verilog/TinyFPGA_B.v(285[5] 287[10])
    defparam mux_250_i5_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i15261_3_lut (.I0(\data_in[2] [6]), .I1(\data_in[3] [6]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n29209));   // verilog/coms.v(128[12] 303[6])
    defparam i15261_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15262_3_lut (.I0(\data_in[2] [5]), .I1(\data_in[3] [5]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n29210));   // verilog/coms.v(128[12] 303[6])
    defparam i15262_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15263_3_lut (.I0(\data_in[2] [4]), .I1(\data_in[3] [4]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n29211));   // verilog/coms.v(128[12] 303[6])
    defparam i15263_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15264_3_lut (.I0(\data_in[2] [3]), .I1(\data_in[3] [3]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n29212));   // verilog/coms.v(128[12] 303[6])
    defparam i15264_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15265_3_lut (.I0(\data_in[2] [2]), .I1(\data_in[3] [2]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n29213));   // verilog/coms.v(128[12] 303[6])
    defparam i15265_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1005_i3_3_lut (.I0(duty[2]), .I1(n361), .I2(duty[23]), 
            .I3(GND_net), .O(n4721));   // verilog/TinyFPGA_B.v(118[13] 129[7])
    defparam mux_1005_i3_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY dti_counter_2244_add_4_2 (.CI(VCC_net), .I0(n2195), .I1(dti_counter[0]), 
            .CO(n39307));
    SB_LUT4 add_2773_25_lut (.I0(n51112), .I1(n2_adj_5411), .I2(n1059), 
            .I3(n39306), .O(encoder0_position_scaled_23__N_51[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2773_25_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 i15266_3_lut (.I0(\data_in[2] [1]), .I1(\data_in[3] [1]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n29214));   // verilog/coms.v(128[12] 303[6])
    defparam i15266_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15267_3_lut (.I0(\data_in[2] [0]), .I1(\data_in[3] [0]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n29215));   // verilog/coms.v(128[12] 303[6])
    defparam i15267_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15268_3_lut (.I0(\data_in[1] [7]), .I1(\data_in[2] [7]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n29216));   // verilog/coms.v(128[12] 303[6])
    defparam i15268_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_250_i6_4_lut (.I0(encoder1_position_scaled[5]), .I1(displacement[5]), 
            .I2(n15_adj_5249), .I3(n15_adj_5321), .O(motor_state_23__N_123[5]));   // verilog/TinyFPGA_B.v(285[5] 287[10])
    defparam mux_250_i6_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i15269_3_lut (.I0(\data_in[1] [6]), .I1(\data_in[2] [6]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n29217));   // verilog/coms.v(128[12] 303[6])
    defparam i15269_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2773_24_lut (.I0(n51099), .I1(n2_adj_5411), .I2(n1158), 
            .I3(n39305), .O(encoder0_position_scaled_23__N_51[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2773_24_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2773_24 (.CI(n39305), .I0(n2_adj_5411), .I1(n1158), .CO(n39306));
    SB_LUT4 i15270_3_lut (.I0(\data_in[1] [5]), .I1(\data_in[2] [5]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n29218));   // verilog/coms.v(128[12] 303[6])
    defparam i15270_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15271_3_lut (.I0(\data_in[1] [4]), .I1(\data_in[2] [4]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n29219));   // verilog/coms.v(128[12] 303[6])
    defparam i15271_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15272_3_lut (.I0(\data_in[1] [3]), .I1(\data_in[2] [3]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n29220));   // verilog/coms.v(128[12] 303[6])
    defparam i15272_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15273_3_lut (.I0(\data_in[1] [2]), .I1(\data_in[2] [2]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n29221));   // verilog/coms.v(128[12] 303[6])
    defparam i15273_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15275_3_lut (.I0(\data_in[1] [1]), .I1(\data_in[2] [1]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n29223));   // verilog/coms.v(128[12] 303[6])
    defparam i15275_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_250_i7_4_lut (.I0(encoder1_position_scaled[6]), .I1(displacement[6]), 
            .I2(n15_adj_5249), .I3(n15_adj_5321), .O(motor_state_23__N_123[6]));   // verilog/TinyFPGA_B.v(285[5] 287[10])
    defparam mux_250_i7_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i15276_3_lut (.I0(\data_in[1] [0]), .I1(\data_in[2] [0]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n29224));   // verilog/coms.v(128[12] 303[6])
    defparam i15276_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i35047_1_lut (.I0(n2940), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n50635));
    defparam i35047_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_1005_i4_3_lut (.I0(duty[3]), .I1(n360), .I2(duty[23]), 
            .I3(GND_net), .O(n4720));   // verilog/TinyFPGA_B.v(118[13] 129[7])
    defparam mux_1005_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15277_3_lut (.I0(\data_in[0] [7]), .I1(\data_in[1] [7]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n29225));   // verilog/coms.v(128[12] 303[6])
    defparam i15277_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2773_23_lut (.I0(n51084), .I1(n2_adj_5411), .I2(n1257), 
            .I3(n39304), .O(encoder0_position_scaled_23__N_51[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2773_23_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2773_23 (.CI(n39304), .I0(n2_adj_5411), .I1(n1257), .CO(n39305));
    SB_LUT4 i16_4_lut (.I0(state_adj_5537[0]), .I1(n49357), .I2(n7210), 
            .I3(n34664), .O(n8));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i16_4_lut.LUT_INIT = 16'h3afa;
    SB_LUT4 add_2773_22_lut (.I0(n51069), .I1(n2_adj_5411), .I2(n1356), 
            .I3(n39303), .O(encoder0_position_scaled_23__N_51[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2773_22_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2773_22 (.CI(n39303), .I0(n2_adj_5411), .I1(n1356), .CO(n39304));
    SB_LUT4 i15289_4_lut (.I0(r_Rx_Data), .I1(rx_data[0]), .I2(n4_adj_5287), 
            .I3(n27131), .O(n29237));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i15289_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i15290_4_lut (.I0(CS_MISO_c), .I1(data_adj_5514[0]), .I2(n11_adj_5367), 
            .I3(state_7__N_4460), .O(n29238));   // verilog/tli4970.v(35[10] 68[6])
    defparam i15290_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 add_2773_21_lut (.I0(n51053), .I1(n2_adj_5411), .I2(n1455), 
            .I3(n39302), .O(encoder0_position_scaled_23__N_51[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2773_21_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 mux_250_i8_4_lut (.I0(encoder1_position_scaled[7]), .I1(displacement[7]), 
            .I2(n15_adj_5249), .I3(n15_adj_5321), .O(motor_state_23__N_123[7]));   // verilog/TinyFPGA_B.v(285[5] 287[10])
    defparam mux_250_i8_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i15291_3_lut (.I0(\data_in[0] [6]), .I1(\data_in[1] [6]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n29239));   // verilog/coms.v(128[12] 303[6])
    defparam i15291_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_250_i9_4_lut (.I0(encoder1_position_scaled[8]), .I1(displacement[8]), 
            .I2(n15_adj_5249), .I3(n15_adj_5321), .O(motor_state_23__N_123[8]));   // verilog/TinyFPGA_B.v(285[5] 287[10])
    defparam mux_250_i9_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_250_i10_4_lut (.I0(encoder1_position_scaled[9]), .I1(displacement[9]), 
            .I2(n15_adj_5249), .I3(n15_adj_5321), .O(motor_state_23__N_123[9]));   // verilog/TinyFPGA_B.v(285[5] 287[10])
    defparam mux_250_i10_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i15292_3_lut (.I0(\data_in[0] [5]), .I1(\data_in[1] [5]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n29240));   // verilog/coms.v(128[12] 303[6])
    defparam i15292_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15293_3_lut (.I0(\data_in[0] [4]), .I1(\data_in[1] [4]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n29241));   // verilog/coms.v(128[12] 303[6])
    defparam i15293_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15294_3_lut (.I0(\data_in[0] [3]), .I1(\data_in[1] [3]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n29242));   // verilog/coms.v(128[12] 303[6])
    defparam i15294_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1005_i5_3_lut (.I0(duty[4]), .I1(n359), .I2(duty[23]), 
            .I3(GND_net), .O(n4719));   // verilog/TinyFPGA_B.v(118[13] 129[7])
    defparam mux_1005_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15295_3_lut (.I0(\data_in[0] [2]), .I1(\data_in[1] [2]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n29243));   // verilog/coms.v(128[12] 303[6])
    defparam i15295_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15296_3_lut (.I0(\data_in[0] [1]), .I1(\data_in[1] [1]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n29244));   // verilog/coms.v(128[12] 303[6])
    defparam i15296_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15598_3_lut (.I0(current[8]), .I1(data_adj_5514[8]), .I2(n28537), 
            .I3(GND_net), .O(n29546));   // verilog/tli4970.v(35[10] 68[6])
    defparam i15598_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15599_3_lut (.I0(current[7]), .I1(data_adj_5514[7]), .I2(n28537), 
            .I3(GND_net), .O(n29547));   // verilog/tli4970.v(35[10] 68[6])
    defparam i15599_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15600_3_lut (.I0(current[6]), .I1(data_adj_5514[6]), .I2(n28537), 
            .I3(GND_net), .O(n29548));   // verilog/tli4970.v(35[10] 68[6])
    defparam i15600_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2_3_lut_adj_1750 (.I0(current_limit[13]), .I1(n26_adj_5384), 
            .I2(current_limit[14]), .I3(GND_net), .O(n46084));
    defparam i2_3_lut_adj_1750.LUT_INIT = 16'hfefe;
    SB_LUT4 i2_3_lut_adj_1751 (.I0(current_limit[13]), .I1(n26_adj_5384), 
            .I2(current_limit[14]), .I3(GND_net), .O(n46081));
    defparam i2_3_lut_adj_1751.LUT_INIT = 16'h8080;
    SB_LUT4 i15601_3_lut (.I0(current[5]), .I1(data_adj_5514[5]), .I2(n28537), 
            .I3(GND_net), .O(n29549));   // verilog/tli4970.v(35[10] 68[6])
    defparam i15601_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15602_3_lut (.I0(current[4]), .I1(data_adj_5514[4]), .I2(n28537), 
            .I3(GND_net), .O(n29550));   // verilog/tli4970.v(35[10] 68[6])
    defparam i15602_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_250_i11_4_lut (.I0(encoder1_position_scaled[10]), .I1(displacement[10]), 
            .I2(n15_adj_5249), .I3(n15_adj_5321), .O(motor_state_23__N_123[10]));   // verilog/TinyFPGA_B.v(285[5] 287[10])
    defparam mux_250_i11_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i1_4_lut_adj_1752 (.I0(current[15]), .I1(current_limit[15]), 
            .I2(n46081), .I3(n46084), .O(n10621));
    defparam i1_4_lut_adj_1752.LUT_INIT = 16'hb3a2;
    SB_LUT4 i15603_3_lut (.I0(current[3]), .I1(data_adj_5514[3]), .I2(n28537), 
            .I3(GND_net), .O(n29551));   // verilog/tli4970.v(35[10] 68[6])
    defparam i15603_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15208_3_lut (.I0(IntegralLimit[3]), .I1(\data_in_frame[13] [3]), 
            .I2(n28521), .I3(GND_net), .O(n29156));   // verilog/coms.v(128[12] 303[6])
    defparam i15208_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15209_3_lut (.I0(IntegralLimit[2]), .I1(\data_in_frame[13] [2]), 
            .I2(n28521), .I3(GND_net), .O(n29157));   // verilog/coms.v(128[12] 303[6])
    defparam i15209_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_250_i12_4_lut (.I0(encoder1_position_scaled[11]), .I1(displacement[11]), 
            .I2(n15_adj_5249), .I3(n15_adj_5321), .O(motor_state_23__N_123[11]));   // verilog/TinyFPGA_B.v(285[5] 287[10])
    defparam mux_250_i12_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i15604_3_lut (.I0(current[2]), .I1(data_adj_5514[2]), .I2(n28537), 
            .I3(GND_net), .O(n29552));   // verilog/tli4970.v(35[10] 68[6])
    defparam i15604_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15605_3_lut (.I0(current[1]), .I1(data_adj_5514[1]), .I2(n28537), 
            .I3(GND_net), .O(n29553));   // verilog/tli4970.v(35[10] 68[6])
    defparam i15605_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15307_3_lut (.I0(\data_in_frame[22] [7]), .I1(rx_data[7]), 
            .I2(n43824), .I3(GND_net), .O(n29255));   // verilog/coms.v(128[12] 303[6])
    defparam i15307_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15308_3_lut (.I0(\data_in_frame[22] [6]), .I1(rx_data[6]), 
            .I2(n43824), .I3(GND_net), .O(n29256));   // verilog/coms.v(128[12] 303[6])
    defparam i15308_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15309_3_lut (.I0(\data_in_frame[22] [5]), .I1(rx_data[5]), 
            .I2(n43824), .I3(GND_net), .O(n29257));   // verilog/coms.v(128[12] 303[6])
    defparam i15309_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15310_3_lut (.I0(\data_in_frame[22] [4]), .I1(rx_data[4]), 
            .I2(n43824), .I3(GND_net), .O(n29258));   // verilog/coms.v(128[12] 303[6])
    defparam i15310_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i35005_1_lut (.I0(n3039), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n50593));
    defparam i35005_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_250_i13_4_lut (.I0(encoder1_position_scaled[12]), .I1(displacement[12]), 
            .I2(n15_adj_5249), .I3(n15_adj_5321), .O(motor_state_23__N_123[12]));   // verilog/TinyFPGA_B.v(285[5] 287[10])
    defparam mux_250_i13_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_250_i14_4_lut (.I0(encoder1_position_scaled[13]), .I1(displacement[13]), 
            .I2(n15_adj_5249), .I3(n15_adj_5321), .O(motor_state_23__N_123[13]));   // verilog/TinyFPGA_B.v(285[5] 287[10])
    defparam mux_250_i14_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i15311_3_lut (.I0(\data_in_frame[22] [3]), .I1(rx_data[3]), 
            .I2(n43824), .I3(GND_net), .O(n29259));   // verilog/coms.v(128[12] 303[6])
    defparam i15311_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15607_3_lut (.I0(PWMLimit[23]), .I1(\data_in_frame[8] [7]), 
            .I2(n28521), .I3(GND_net), .O(n29555));   // verilog/coms.v(128[12] 303[6])
    defparam i15607_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_250_i15_4_lut (.I0(encoder1_position_scaled[14]), .I1(displacement[14]), 
            .I2(n15_adj_5249), .I3(n15_adj_5321), .O(motor_state_23__N_123[14]));   // verilog/TinyFPGA_B.v(285[5] 287[10])
    defparam mux_250_i15_4_lut.LUT_INIT = 16'h0aca;
    SB_CARRY add_2773_21 (.CI(n39302), .I0(n2_adj_5411), .I1(n1455), .CO(n39303));
    SB_LUT4 i15608_3_lut (.I0(PWMLimit[22]), .I1(\data_in_frame[8] [6]), 
            .I2(n28521), .I3(GND_net), .O(n29556));   // verilog/coms.v(128[12] 303[6])
    defparam i15608_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15609_3_lut (.I0(PWMLimit[21]), .I1(\data_in_frame[8] [5]), 
            .I2(n28521), .I3(GND_net), .O(n29557));   // verilog/coms.v(128[12] 303[6])
    defparam i15609_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15312_3_lut (.I0(\data_in_frame[22] [2]), .I1(rx_data[2]), 
            .I2(n43824), .I3(GND_net), .O(n29260));   // verilog/coms.v(128[12] 303[6])
    defparam i15312_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15610_3_lut (.I0(PWMLimit[20]), .I1(\data_in_frame[8] [4]), 
            .I2(n28521), .I3(GND_net), .O(n29558));   // verilog/coms.v(128[12] 303[6])
    defparam i15610_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15611_3_lut (.I0(PWMLimit[19]), .I1(\data_in_frame[8] [3]), 
            .I2(n28521), .I3(GND_net), .O(n29559));   // verilog/coms.v(128[12] 303[6])
    defparam i15611_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15612_3_lut (.I0(PWMLimit[18]), .I1(\data_in_frame[8] [2]), 
            .I2(n28521), .I3(GND_net), .O(n29560));   // verilog/coms.v(128[12] 303[6])
    defparam i15612_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15313_3_lut (.I0(\data_in_frame[22] [1]), .I1(rx_data[1]), 
            .I2(n43824), .I3(GND_net), .O(n29261));   // verilog/coms.v(128[12] 303[6])
    defparam i15313_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15613_3_lut (.I0(PWMLimit[17]), .I1(\data_in_frame[8] [1]), 
            .I2(n28521), .I3(GND_net), .O(n29561));   // verilog/coms.v(128[12] 303[6])
    defparam i15613_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2773_20_lut (.I0(n51036), .I1(n2_adj_5411), .I2(n1554), 
            .I3(n39301), .O(encoder0_position_scaled_23__N_51[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2773_20_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2773_20 (.CI(n39301), .I0(n2_adj_5411), .I1(n1554), .CO(n39302));
    SB_LUT4 i15177_3_lut (.I0(\data_out_frame[4] [6]), .I1(ID[6]), .I2(n24278), 
            .I3(GND_net), .O(n29125));   // verilog/coms.v(128[12] 303[6])
    defparam i15177_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15178_3_lut (.I0(\data_out_frame[4] [5]), .I1(ID[5]), .I2(n24278), 
            .I3(GND_net), .O(n29126));   // verilog/coms.v(128[12] 303[6])
    defparam i15178_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15314_3_lut (.I0(\data_in_frame[22] [0]), .I1(rx_data[0]), 
            .I2(n43824), .I3(GND_net), .O(n29262));   // verilog/coms.v(128[12] 303[6])
    defparam i15314_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_2773_19_lut (.I0(n51018), .I1(n2_adj_5411), .I2(n1653), 
            .I3(n39300), .O(encoder0_position_scaled_23__N_51[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2773_19_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2773_19 (.CI(n39300), .I0(n2_adj_5411), .I1(n1653), .CO(n39301));
    SB_LUT4 i34956_1_lut (.I0(n3138), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n50544));
    defparam i34956_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_250_i16_4_lut (.I0(encoder1_position_scaled[15]), .I1(displacement[15]), 
            .I2(n15_adj_5249), .I3(n15_adj_5321), .O(motor_state_23__N_123[15]));   // verilog/TinyFPGA_B.v(285[5] 287[10])
    defparam mux_250_i16_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i15315_3_lut (.I0(\data_in_frame[21] [7]), .I1(rx_data[7]), 
            .I2(n43822), .I3(GND_net), .O(n29263));   // verilog/coms.v(128[12] 303[6])
    defparam i15315_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15316_3_lut (.I0(\data_in_frame[21] [6]), .I1(rx_data[6]), 
            .I2(n43822), .I3(GND_net), .O(n29264));   // verilog/coms.v(128[12] 303[6])
    defparam i15316_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15614_3_lut (.I0(PWMLimit[16]), .I1(\data_in_frame[8] [0]), 
            .I2(n28521), .I3(GND_net), .O(n29562));   // verilog/coms.v(128[12] 303[6])
    defparam i15614_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15317_3_lut (.I0(\data_in_frame[21] [5]), .I1(rx_data[5]), 
            .I2(n43822), .I3(GND_net), .O(n29265));   // verilog/coms.v(128[12] 303[6])
    defparam i15317_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_2773_18_lut (.I0(n50999), .I1(n2_adj_5411), .I2(n1752), 
            .I3(n39299), .O(encoder0_position_scaled_23__N_51[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2773_18_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 i15615_3_lut (.I0(PWMLimit[15]), .I1(\data_in_frame[9] [7]), 
            .I2(n28521), .I3(GND_net), .O(n29563));   // verilog/coms.v(128[12] 303[6])
    defparam i15615_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15318_3_lut (.I0(\data_in_frame[21] [4]), .I1(rx_data[4]), 
            .I2(n43822), .I3(GND_net), .O(n29266));   // verilog/coms.v(128[12] 303[6])
    defparam i15318_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_2773_18 (.CI(n39299), .I0(n2_adj_5411), .I1(n1752), .CO(n39300));
    SB_LUT4 add_2773_17_lut (.I0(n50979), .I1(n2_adj_5411), .I2(n1851), 
            .I3(n39298), .O(encoder0_position_scaled_23__N_51[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2773_17_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2773_17 (.CI(n39298), .I0(n2_adj_5411), .I1(n1851), .CO(n39299));
    SB_LUT4 add_2773_16_lut (.I0(n50958), .I1(n2_adj_5411), .I2(n1950), 
            .I3(n39297), .O(encoder0_position_scaled_23__N_51[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2773_16_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2773_16 (.CI(n39297), .I0(n2_adj_5411), .I1(n1950), .CO(n39298));
    SB_LUT4 add_157_5_lut (.I0(GND_net), .I1(delay_counter[3]), .I2(GND_net), 
            .I3(n38448), .O(n1325)) /* synthesis syn_instantiated=1 */ ;
    defparam add_157_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_250_i17_4_lut (.I0(encoder1_position_scaled[16]), .I1(displacement[16]), 
            .I2(n15_adj_5249), .I3(n15_adj_5321), .O(motor_state_23__N_123[16]));   // verilog/TinyFPGA_B.v(285[5] 287[10])
    defparam mux_250_i17_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 add_2773_15_lut (.I0(n50937), .I1(n2_adj_5411), .I2(n2049), 
            .I3(n39296), .O(encoder0_position_scaled_23__N_51[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2773_15_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 i15319_3_lut (.I0(\data_in_frame[21] [3]), .I1(rx_data[3]), 
            .I2(n43822), .I3(GND_net), .O(n29267));   // verilog/coms.v(128[12] 303[6])
    defparam i15319_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_2773_15 (.CI(n39296), .I0(n2_adj_5411), .I1(n2049), .CO(n39297));
    SB_LUT4 i15320_3_lut (.I0(\data_in_frame[21] [2]), .I1(rx_data[2]), 
            .I2(n43822), .I3(GND_net), .O(n29268));   // verilog/coms.v(128[12] 303[6])
    defparam i15320_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15616_3_lut (.I0(PWMLimit[14]), .I1(\data_in_frame[9] [6]), 
            .I2(n28521), .I3(GND_net), .O(n29564));   // verilog/coms.v(128[12] 303[6])
    defparam i15616_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15617_3_lut (.I0(PWMLimit[13]), .I1(\data_in_frame[9] [5]), 
            .I2(n28521), .I3(GND_net), .O(n29565));   // verilog/coms.v(128[12] 303[6])
    defparam i15617_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1005_i6_3_lut (.I0(duty[5]), .I1(n358), .I2(duty[23]), 
            .I3(GND_net), .O(n4718));   // verilog/TinyFPGA_B.v(118[13] 129[7])
    defparam mux_1005_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_19_inv_0_i23_1_lut (.I0(duty[22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n3));   // verilog/TinyFPGA_B.v(123[25:30])
    defparam unary_minus_19_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i15321_3_lut (.I0(\data_in_frame[21] [1]), .I1(rx_data[1]), 
            .I2(n43822), .I3(GND_net), .O(n29269));   // verilog/coms.v(128[12] 303[6])
    defparam i15321_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_2773_14_lut (.I0(n50914), .I1(n2_adj_5411), .I2(n2148), 
            .I3(n39295), .O(encoder0_position_scaled_23__N_51[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2773_14_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2773_14 (.CI(n39295), .I0(n2_adj_5411), .I1(n2148), .CO(n39296));
    SB_LUT4 add_2773_13_lut (.I0(n50890), .I1(n2_adj_5411), .I2(n2247), 
            .I3(n39294), .O(encoder0_position_scaled_23__N_51[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2773_13_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 i15322_3_lut (.I0(\data_in_frame[21] [0]), .I1(rx_data[0]), 
            .I2(n43822), .I3(GND_net), .O(n29270));   // verilog/coms.v(128[12] 303[6])
    defparam i15322_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_2773_13 (.CI(n39294), .I0(n2_adj_5411), .I1(n2247), .CO(n39295));
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i27_1_lut (.I0(encoder0_position[26]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n7_adj_5416));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i27_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_2773_12_lut (.I0(n50865), .I1(n2_adj_5411), .I2(n2346), 
            .I3(n39293), .O(encoder0_position_scaled_23__N_51[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2773_12_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2773_12 (.CI(n39293), .I0(n2_adj_5411), .I1(n2346), .CO(n39294));
    SB_LUT4 add_2773_11_lut (.I0(n50784), .I1(n2_adj_5411), .I2(n2445), 
            .I3(n39292), .O(encoder0_position_scaled_23__N_51[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2773_11_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2773_11 (.CI(n39292), .I0(n2_adj_5411), .I1(n2445), .CO(n39293));
    SB_LUT4 add_2773_10_lut (.I0(n50754), .I1(n2_adj_5411), .I2(n2544), 
            .I3(n39291), .O(encoder0_position_scaled_23__N_51[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2773_10_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 i15073_3_lut (.I0(\data_out_frame[12] [6]), .I1(setpoint[22]), 
            .I2(n24278), .I3(GND_net), .O(n29021));   // verilog/coms.v(128[12] 303[6])
    defparam i15073_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2773_10 (.CI(n39291), .I0(n2_adj_5411), .I1(n2544), .CO(n39292));
    SB_LUT4 i15618_3_lut (.I0(PWMLimit[12]), .I1(\data_in_frame[9] [4]), 
            .I2(n28521), .I3(GND_net), .O(n29566));   // verilog/coms.v(128[12] 303[6])
    defparam i15618_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i35481_1_lut (.I0(n1356), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n51069));
    defparam i35481_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_2773_9_lut (.I0(n50702), .I1(n2_adj_5411), .I2(n2643), 
            .I3(n39290), .O(encoder0_position_scaled_23__N_51[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2773_9_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2773_9 (.CI(n39290), .I0(n2_adj_5411), .I1(n2643), .CO(n39291));
    SB_LUT4 add_2773_8_lut (.I0(n50697), .I1(n2_adj_5411), .I2(n2742), 
            .I3(n39289), .O(encoder0_position_scaled_23__N_51[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2773_8_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2773_8 (.CI(n39289), .I0(n2_adj_5411), .I1(n2742), .CO(n39290));
    SB_LUT4 add_2773_7_lut (.I0(n50668), .I1(n2_adj_5411), .I2(n2841), 
            .I3(n39288), .O(encoder0_position_scaled_23__N_51[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2773_7_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2773_7 (.CI(n39288), .I0(n2_adj_5411), .I1(n2841), .CO(n39289));
    SB_LUT4 add_2773_6_lut (.I0(n50635), .I1(n2_adj_5411), .I2(n2940), 
            .I3(n39287), .O(encoder0_position_scaled_23__N_51[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2773_6_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2773_6 (.CI(n39287), .I0(n2_adj_5411), .I1(n2940), .CO(n39288));
    SB_LUT4 add_2773_5_lut (.I0(n50593), .I1(n2_adj_5411), .I2(n3039), 
            .I3(n39286), .O(encoder0_position_scaled_23__N_51[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2773_5_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2773_5 (.CI(n39286), .I0(n2_adj_5411), .I1(n3039), .CO(n39287));
    SB_LUT4 add_2773_4_lut (.I0(n50544), .I1(n2_adj_5411), .I2(n3138), 
            .I3(n39285), .O(encoder0_position_scaled_23__N_51[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2773_4_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2773_4 (.CI(n39285), .I0(n2_adj_5411), .I1(n3138), .CO(n39286));
    SB_LUT4 add_2773_3_lut (.I0(n51192), .I1(n2_adj_5411), .I2(n3237), 
            .I3(n39284), .O(encoder0_position_scaled_23__N_51[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2773_3_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2773_3 (.CI(n39284), .I0(n2_adj_5411), .I1(n3237), .CO(n39285));
    SB_LUT4 add_2773_2_lut (.I0(n51159), .I1(n2_adj_5411), .I2(n35558), 
            .I3(VCC_net), .O(encoder0_position_scaled_23__N_51[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2773_2_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2773_2 (.CI(VCC_net), .I0(n2_adj_5411), .I1(n35558), 
            .CO(n39284));
    SB_LUT4 i15619_3_lut (.I0(PWMLimit[11]), .I1(\data_in_frame[9] [3]), 
            .I2(n28521), .I3(GND_net), .O(n29567));   // verilog/coms.v(128[12] 303[6])
    defparam i15619_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_add_2173_33_lut (.I0(GND_net), .I1(n3204), 
            .I2(VCC_net), .I3(n39283), .O(n3271)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_33_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15340_4_lut (.I0(CS_MISO_c), .I1(data_adj_5514[10]), .I2(n5_adj_5347), 
            .I3(n27174), .O(n29288));   // verilog/tli4970.v(35[10] 68[6])
    defparam i15340_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 encoder0_position_31__I_0_add_2173_32_lut (.I0(GND_net), .I1(n3205), 
            .I2(VCC_net), .I3(n39282), .O(n3272)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_32_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2173_32 (.CI(n39282), .I0(n3205), 
            .I1(VCC_net), .CO(n39283));
    SB_LUT4 i35465_1_lut (.I0(n1455), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n51053));
    defparam i35465_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_add_2173_31_lut (.I0(GND_net), .I1(n3206), 
            .I2(VCC_net), .I3(n39281), .O(n3273)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_31_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15342_4_lut (.I0(CS_MISO_c), .I1(data_adj_5514[11]), .I2(n34690), 
            .I3(n27174), .O(n29290));   // verilog/tli4970.v(35[10] 68[6])
    defparam i15342_4_lut.LUT_INIT = 16'hccac;
    SB_CARRY add_236_8 (.CI(n38482), .I0(encoder1_position[9]), .I1(GND_net), 
            .CO(n38483));
    SB_CARRY encoder0_position_31__I_0_add_2173_31 (.CI(n39281), .I0(n3206), 
            .I1(VCC_net), .CO(n39282));
    SB_LUT4 encoder0_position_31__I_0_add_2173_30_lut (.I0(GND_net), .I1(n3207), 
            .I2(VCC_net), .I3(n39280), .O(n3274)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2173_30 (.CI(n39280), .I0(n3207), 
            .I1(VCC_net), .CO(n39281));
    SB_DFF pwm_setpoint_i1 (.Q(pwm_setpoint[1]), .C(CLK_c), .D(pwm_setpoint_23__N_11[1]));   // verilog/TinyFPGA_B.v(104[9] 130[5])
    SB_LUT4 encoder0_position_31__I_0_add_2173_29_lut (.I0(GND_net), .I1(n3208), 
            .I2(VCC_net), .I3(n39279), .O(n3275)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_29_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15620_3_lut (.I0(PWMLimit[10]), .I1(\data_in_frame[9] [2]), 
            .I2(n28521), .I3(GND_net), .O(n29568));   // verilog/coms.v(128[12] 303[6])
    defparam i15620_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_31__I_0_add_2173_29 (.CI(n39279), .I0(n3208), 
            .I1(VCC_net), .CO(n39280));
    SB_LUT4 i14881_2_lut (.I0(n28482), .I1(dti), .I2(GND_net), .I3(GND_net), 
            .O(n28835));   // verilog/TinyFPGA_B.v(144[9] 223[5])
    defparam i14881_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i34886_4_lut (.I0(commutation_state[1]), .I1(n24462), .I2(dti), 
            .I3(commutation_state[2]), .O(n28482));
    defparam i34886_4_lut.LUT_INIT = 16'hc5cf;
    SB_LUT4 encoder0_position_31__I_0_add_2173_28_lut (.I0(GND_net), .I1(n3209), 
            .I2(VCC_net), .I3(n39278), .O(n3276)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2173_28 (.CI(n39278), .I0(n3209), 
            .I1(VCC_net), .CO(n39279));
    SB_LUT4 encoder0_position_31__I_0_add_2173_27_lut (.I0(GND_net), .I1(n3210), 
            .I2(VCC_net), .I3(n39277), .O(n3277)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_27_lut.LUT_INIT = 16'hC33C;
    SB_IO INLC_pad (.PACKAGE_PIN(INLC), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INLC_c_0));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INLC_pad.PIN_TYPE = 6'b011001;
    defparam INLC_pad.PULLUP = 1'b0;
    defparam INLC_pad.NEG_TRIGGER = 1'b0;
    defparam INLC_pad.IO_STANDARD = "SB_LVCMOS";
    SB_CARRY encoder0_position_31__I_0_add_2173_27 (.CI(n39277), .I0(n3210), 
            .I1(VCC_net), .CO(n39278));
    SB_LUT4 encoder0_position_31__I_0_add_2173_26_lut (.I0(GND_net), .I1(n3211), 
            .I2(VCC_net), .I3(n39276), .O(n3278)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_236_7_lut (.I0(GND_net), .I1(encoder1_position[8]), .I2(GND_net), 
            .I3(n38481), .O(encoder1_position_scaled_23__N_75[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_236_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15621_3_lut (.I0(PWMLimit[9]), .I1(\data_in_frame[9] [1]), 
            .I2(n28521), .I3(GND_net), .O(n29569));   // verilog/coms.v(128[12] 303[6])
    defparam i15621_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15496_3_lut (.I0(neopxl_color[23]), .I1(\data_in_frame[4] [7]), 
            .I2(n28522), .I3(GND_net), .O(n29444));   // verilog/coms.v(128[12] 303[6])
    defparam i15496_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15497_3_lut (.I0(neopxl_color[22]), .I1(\data_in_frame[4] [6]), 
            .I2(n28522), .I3(GND_net), .O(n29445));   // verilog/coms.v(128[12] 303[6])
    defparam i15497_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15498_3_lut (.I0(neopxl_color[21]), .I1(\data_in_frame[4] [5]), 
            .I2(n28522), .I3(GND_net), .O(n29446));   // verilog/coms.v(128[12] 303[6])
    defparam i15498_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_31__I_0_add_2173_26 (.CI(n39276), .I0(n3211), 
            .I1(VCC_net), .CO(n39277));
    SB_LUT4 i15499_3_lut (.I0(neopxl_color[20]), .I1(\data_in_frame[4] [4]), 
            .I2(n28522), .I3(GND_net), .O(n29447));   // verilog/coms.v(128[12] 303[6])
    defparam i15499_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_236_7 (.CI(n38481), .I0(encoder1_position[8]), .I1(GND_net), 
            .CO(n38482));
    SB_LUT4 i15622_3_lut (.I0(PWMLimit[8]), .I1(\data_in_frame[9] [0]), 
            .I2(n28521), .I3(GND_net), .O(n29570));   // verilog/coms.v(128[12] 303[6])
    defparam i15622_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_add_2173_25_lut (.I0(GND_net), .I1(n3212), 
            .I2(VCC_net), .I3(n39275), .O(n3279)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 n51450_bdd_4_lut (.I0(n51450), .I1(n343), .I2(n4488), .I3(n4208), 
            .O(pwm_setpoint_23__N_11[20]));
    defparam n51450_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_CARRY encoder0_position_31__I_0_add_2173_25 (.CI(n39275), .I0(n3212), 
            .I1(VCC_net), .CO(n39276));
    SB_LUT4 i15500_3_lut (.I0(neopxl_color[19]), .I1(\data_in_frame[4] [3]), 
            .I2(n28522), .I3(GND_net), .O(n29448));   // verilog/coms.v(128[12] 303[6])
    defparam i15500_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_add_2173_24_lut (.I0(GND_net), .I1(n3213), 
            .I2(VCC_net), .I3(n39274), .O(n3280)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15501_3_lut (.I0(neopxl_color[18]), .I1(\data_in_frame[4] [2]), 
            .I2(n28522), .I3(GND_net), .O(n29449));   // verilog/coms.v(128[12] 303[6])
    defparam i15501_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_31__I_0_add_2173_24 (.CI(n39274), .I0(n3213), 
            .I1(VCC_net), .CO(n39275));
    SB_LUT4 encoder0_position_31__I_0_add_2173_23_lut (.I0(GND_net), .I1(n3214), 
            .I2(VCC_net), .I3(n39273), .O(n3281)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i35448_1_lut (.I0(n1554), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n51036));
    defparam i35448_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_31__I_0_add_2173_23 (.CI(n39273), .I0(n3214), 
            .I1(VCC_net), .CO(n39274));
    SB_DFFESR delay_counter_i0_i7 (.Q(delay_counter[7]), .C(CLK_c), .E(n7417), 
            .D(n1321), .R(n28933));   // verilog/TinyFPGA_B.v(375[10] 403[6])
    SB_LUT4 encoder0_position_31__I_0_add_2173_22_lut (.I0(GND_net), .I1(n3215), 
            .I2(VCC_net), .I3(n39272), .O(n3282)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2173_22 (.CI(n39272), .I0(n3215), 
            .I1(VCC_net), .CO(n39273));
    SB_LUT4 i15502_3_lut (.I0(neopxl_color[17]), .I1(\data_in_frame[4] [1]), 
            .I2(n28522), .I3(GND_net), .O(n29450));   // verilog/coms.v(128[12] 303[6])
    defparam i15502_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFESR delay_counter_i0_i0 (.Q(delay_counter[0]), .C(CLK_c), .E(n7417), 
            .D(n1328), .R(n28933));   // verilog/TinyFPGA_B.v(375[10] 403[6])
    SB_LUT4 add_157_13_lut (.I0(GND_net), .I1(delay_counter[11]), .I2(GND_net), 
            .I3(n38456), .O(n1317)) /* synthesis syn_instantiated=1 */ ;
    defparam add_157_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_2173_21_lut (.I0(GND_net), .I1(n3216), 
            .I2(VCC_net), .I3(n39271), .O(n3283)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_21_lut.LUT_INIT = 16'hC33C;
    SB_DFFESR delay_counter_i0_i8 (.Q(delay_counter[8]), .C(CLK_c), .E(n7417), 
            .D(n1320), .R(n28933));   // verilog/TinyFPGA_B.v(375[10] 403[6])
    SB_CARRY encoder0_position_31__I_0_add_2173_21 (.CI(n39271), .I0(n3216), 
            .I1(VCC_net), .CO(n39272));
    SB_LUT4 i15503_3_lut (.I0(neopxl_color[16]), .I1(\data_in_frame[4] [0]), 
            .I2(n28522), .I3(GND_net), .O(n29451));   // verilog/coms.v(128[12] 303[6])
    defparam i15503_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_add_2173_20_lut (.I0(GND_net), .I1(n3217), 
            .I2(VCC_net), .I3(n39270), .O(n3284)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_20_lut.LUT_INIT = 16'hC33C;
    SB_DFFESR delay_counter_i0_i9 (.Q(delay_counter[9]), .C(CLK_c), .E(n7417), 
            .D(n1319), .R(n28933));   // verilog/TinyFPGA_B.v(375[10] 403[6])
    SB_CARRY encoder0_position_31__I_0_add_2173_20 (.CI(n39270), .I0(n3217), 
            .I1(VCC_net), .CO(n39271));
    SB_LUT4 encoder0_position_31__I_0_add_2173_19_lut (.I0(GND_net), .I1(n3218), 
            .I2(VCC_net), .I3(n39269), .O(n3285)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2173_19 (.CI(n39269), .I0(n3218), 
            .I1(VCC_net), .CO(n39270));
    SB_LUT4 encoder0_position_31__I_0_add_2173_18_lut (.I0(GND_net), .I1(n3219), 
            .I2(VCC_net), .I3(n39268), .O(n3286)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2173_18 (.CI(n39268), .I0(n3219), 
            .I1(VCC_net), .CO(n39269));
    SB_LUT4 encoder0_position_31__I_0_add_2173_17_lut (.I0(GND_net), .I1(n3220), 
            .I2(VCC_net), .I3(n39267), .O(n3287)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2173_17 (.CI(n39267), .I0(n3220), 
            .I1(VCC_net), .CO(n39268));
    SB_LUT4 encoder0_position_31__I_0_add_2173_16_lut (.I0(GND_net), .I1(n3221), 
            .I2(VCC_net), .I3(n39266), .O(n3288)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2173_16 (.CI(n39266), .I0(n3221), 
            .I1(VCC_net), .CO(n39267));
    SB_LUT4 encoder0_position_31__I_0_add_2173_15_lut (.I0(GND_net), .I1(n3222), 
            .I2(VCC_net), .I3(n39265), .O(n3289)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2173_15 (.CI(n39265), .I0(n3222), 
            .I1(VCC_net), .CO(n39266));
    SB_LUT4 encoder0_position_31__I_0_add_2173_14_lut (.I0(GND_net), .I1(n3223), 
            .I2(VCC_net), .I3(n39264), .O(n3290)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2173_14 (.CI(n39264), .I0(n3223), 
            .I1(VCC_net), .CO(n39265));
    SB_LUT4 encoder0_position_31__I_0_add_2173_13_lut (.I0(GND_net), .I1(n3224), 
            .I2(VCC_net), .I3(n39263), .O(n3291)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2173_13 (.CI(n39263), .I0(n3224), 
            .I1(VCC_net), .CO(n39264));
    SB_LUT4 encoder0_position_31__I_0_add_2173_12_lut (.I0(GND_net), .I1(n3225), 
            .I2(VCC_net), .I3(n39262), .O(n3292)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15504_3_lut (.I0(neopxl_color[15]), .I1(\data_in_frame[5] [7]), 
            .I2(n28522), .I3(GND_net), .O(n29452));   // verilog/coms.v(128[12] 303[6])
    defparam i15504_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15623_3_lut (.I0(PWMLimit[7]), .I1(\data_in_frame[10] [7]), 
            .I2(n28521), .I3(GND_net), .O(n29571));   // verilog/coms.v(128[12] 303[6])
    defparam i15623_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15505_3_lut (.I0(neopxl_color[14]), .I1(\data_in_frame[5] [6]), 
            .I2(n28522), .I3(GND_net), .O(n29453));   // verilog/coms.v(128[12] 303[6])
    defparam i15505_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15624_3_lut (.I0(PWMLimit[6]), .I1(\data_in_frame[10] [6]), 
            .I2(n28521), .I3(GND_net), .O(n29572));   // verilog/coms.v(128[12] 303[6])
    defparam i15624_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i28_1_lut (.I0(encoder0_position[27]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n6_adj_5415));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i28_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i15625_3_lut (.I0(PWMLimit[5]), .I1(\data_in_frame[10] [5]), 
            .I2(n28521), .I3(GND_net), .O(n29573));   // verilog/coms.v(128[12] 303[6])
    defparam i15625_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15506_3_lut (.I0(neopxl_color[13]), .I1(\data_in_frame[5] [5]), 
            .I2(n28522), .I3(GND_net), .O(n29454));   // verilog/coms.v(128[12] 303[6])
    defparam i15506_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15507_3_lut (.I0(neopxl_color[12]), .I1(\data_in_frame[5] [4]), 
            .I2(n28522), .I3(GND_net), .O(n29455));   // verilog/coms.v(128[12] 303[6])
    defparam i15507_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15508_3_lut (.I0(neopxl_color[11]), .I1(\data_in_frame[5] [3]), 
            .I2(n28522), .I3(GND_net), .O(n29456));   // verilog/coms.v(128[12] 303[6])
    defparam i15508_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15509_3_lut (.I0(neopxl_color[10]), .I1(\data_in_frame[5] [2]), 
            .I2(n28522), .I3(GND_net), .O(n29457));   // verilog/coms.v(128[12] 303[6])
    defparam i15509_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15510_3_lut (.I0(neopxl_color[9]), .I1(\data_in_frame[5] [1]), 
            .I2(n28522), .I3(GND_net), .O(n29458));   // verilog/coms.v(128[12] 303[6])
    defparam i15510_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15511_3_lut (.I0(neopxl_color[8]), .I1(\data_in_frame[5] [0]), 
            .I2(n28522), .I3(GND_net), .O(n29459));   // verilog/coms.v(128[12] 303[6])
    defparam i15511_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15373_3_lut (.I0(\data_in_frame[14] [7]), .I1(rx_data[7]), 
            .I2(n43848), .I3(GND_net), .O(n29321));   // verilog/coms.v(128[12] 303[6])
    defparam i15373_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15626_3_lut (.I0(PWMLimit[4]), .I1(\data_in_frame[10] [4]), 
            .I2(n28521), .I3(GND_net), .O(n29574));   // verilog/coms.v(128[12] 303[6])
    defparam i15626_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15374_3_lut (.I0(\data_in_frame[14] [6]), .I1(rx_data[6]), 
            .I2(n43848), .I3(GND_net), .O(n29322));   // verilog/coms.v(128[12] 303[6])
    defparam i15374_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15375_4_lut (.I0(CS_MISO_c), .I1(data_adj_5514[12]), .I2(n34688), 
            .I3(n27143), .O(n29323));   // verilog/tli4970.v(35[10] 68[6])
    defparam i15375_4_lut.LUT_INIT = 16'hccac;
    SB_LUT4 mux_1005_i7_3_lut (.I0(duty[6]), .I1(n357), .I2(duty[23]), 
            .I3(GND_net), .O(n4717));   // verilog/TinyFPGA_B.v(118[13] 129[7])
    defparam mux_1005_i7_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15512_3_lut (.I0(neopxl_color[7]), .I1(\data_in_frame[6] [7]), 
            .I2(n28522), .I3(GND_net), .O(n29460));   // verilog/coms.v(128[12] 303[6])
    defparam i15512_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15513_3_lut (.I0(neopxl_color[6]), .I1(\data_in_frame[6] [6]), 
            .I2(n28522), .I3(GND_net), .O(n29461));   // verilog/coms.v(128[12] 303[6])
    defparam i15513_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15376_4_lut (.I0(CS_MISO_c), .I1(data_adj_5514[15]), .I2(n34688), 
            .I3(n27180), .O(n29324));   // verilog/tli4970.v(35[10] 68[6])
    defparam i15376_4_lut.LUT_INIT = 16'hccac;
    SB_LUT4 i15377_3_lut (.I0(\data_in_frame[14] [5]), .I1(rx_data[5]), 
            .I2(n43848), .I3(GND_net), .O(n29325));   // verilog/coms.v(128[12] 303[6])
    defparam i15377_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15514_3_lut (.I0(neopxl_color[5]), .I1(\data_in_frame[6] [5]), 
            .I2(n28522), .I3(GND_net), .O(n29462));   // verilog/coms.v(128[12] 303[6])
    defparam i15514_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1005_i8_3_lut (.I0(duty[7]), .I1(n356), .I2(duty[23]), 
            .I3(GND_net), .O(n4716));   // verilog/TinyFPGA_B.v(118[13] 129[7])
    defparam mux_1005_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15378_3_lut (.I0(\data_in_frame[14] [4]), .I1(rx_data[4]), 
            .I2(n43848), .I3(GND_net), .O(n29326));   // verilog/coms.v(128[12] 303[6])
    defparam i15378_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15515_3_lut (.I0(neopxl_color[4]), .I1(\data_in_frame[6] [4]), 
            .I2(n28522), .I3(GND_net), .O(n29463));   // verilog/coms.v(128[12] 303[6])
    defparam i15515_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15379_3_lut (.I0(\data_in_frame[14] [3]), .I1(rx_data[3]), 
            .I2(n43848), .I3(GND_net), .O(n29327));   // verilog/coms.v(128[12] 303[6])
    defparam i15379_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_2173_12 (.CI(n39262), .I0(n3225), 
            .I1(VCC_net), .CO(n39263));
    SB_LUT4 encoder0_position_31__I_0_add_2173_11_lut (.I0(GND_net), .I1(n3226), 
            .I2(VCC_net), .I3(n39261), .O(n3293)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2173_11 (.CI(n39261), .I0(n3226), 
            .I1(VCC_net), .CO(n39262));
    SB_LUT4 encoder0_position_31__I_0_add_2173_10_lut (.I0(GND_net), .I1(n3227), 
            .I2(VCC_net), .I3(n39260), .O(n3294)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2173_10 (.CI(n39260), .I0(n3227), 
            .I1(VCC_net), .CO(n39261));
    SB_LUT4 encoder0_position_31__I_0_add_2173_9_lut (.I0(GND_net), .I1(n3228), 
            .I2(VCC_net), .I3(n39259), .O(n3295)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15380_3_lut (.I0(\data_in_frame[14] [2]), .I1(rx_data[2]), 
            .I2(n43848), .I3(GND_net), .O(n29328));   // verilog/coms.v(128[12] 303[6])
    defparam i15380_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_2173_9 (.CI(n39259), .I0(n3228), 
            .I1(VCC_net), .CO(n39260));
    SB_LUT4 i15381_3_lut (.I0(\data_in_frame[14] [1]), .I1(rx_data[1]), 
            .I2(n43848), .I3(GND_net), .O(n29329));   // verilog/coms.v(128[12] 303[6])
    defparam i15381_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15627_3_lut (.I0(PWMLimit[3]), .I1(\data_in_frame[10] [3]), 
            .I2(n28521), .I3(GND_net), .O(n29575));   // verilog/coms.v(128[12] 303[6])
    defparam i15627_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_add_2173_8_lut (.I0(GND_net), .I1(n3229), 
            .I2(GND_net), .I3(n39258), .O(n3296)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15382_3_lut (.I0(\data_in_frame[14] [0]), .I1(rx_data[0]), 
            .I2(n43848), .I3(GND_net), .O(n29330));   // verilog/coms.v(128[12] 303[6])
    defparam i15382_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_2173_8 (.CI(n39258), .I0(n3229), 
            .I1(GND_net), .CO(n39259));
    SB_LUT4 i15383_3_lut (.I0(\data_in_frame[13] [7]), .I1(rx_data[7]), 
            .I2(n43847), .I3(GND_net), .O(n29331));   // verilog/coms.v(128[12] 303[6])
    defparam i15383_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_2173_7_lut (.I0(n3298), .I1(n3230), 
            .I2(GND_net), .I3(n39257), .O(n49339)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_7_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i15516_3_lut (.I0(neopxl_color[3]), .I1(\data_in_frame[6] [3]), 
            .I2(n28522), .I3(GND_net), .O(n29464));   // verilog/coms.v(128[12] 303[6])
    defparam i15516_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15384_3_lut (.I0(\data_in_frame[13] [6]), .I1(rx_data[6]), 
            .I2(n43847), .I3(GND_net), .O(n29332));   // verilog/coms.v(128[12] 303[6])
    defparam i15384_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_2173_7 (.CI(n39257), .I0(n3230), 
            .I1(GND_net), .CO(n39258));
    SB_LUT4 add_236_6_lut (.I0(GND_net), .I1(encoder1_position[7]), .I2(GND_net), 
            .I3(n38480), .O(encoder1_position_scaled_23__N_75[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_236_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_2173_6_lut (.I0(GND_net), .I1(n3231), 
            .I2(VCC_net), .I3(n39256), .O(n3298)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15517_3_lut (.I0(neopxl_color[2]), .I1(\data_in_frame[6] [2]), 
            .I2(n28522), .I3(GND_net), .O(n29465));   // verilog/coms.v(128[12] 303[6])
    defparam i15517_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_31__I_0_add_2173_6 (.CI(n39256), .I0(n3231), 
            .I1(VCC_net), .CO(n39257));
    SB_LUT4 i15385_3_lut (.I0(\data_in_frame[13] [5]), .I1(rx_data[5]), 
            .I2(n43847), .I3(GND_net), .O(n29333));   // verilog/coms.v(128[12] 303[6])
    defparam i15385_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i35430_1_lut (.I0(n1653), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n51018));
    defparam i35430_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_add_2173_5_lut (.I0(GND_net), .I1(n3232), 
            .I2(GND_net), .I3(n39255), .O(n3299)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2173_5 (.CI(n39255), .I0(n3232), 
            .I1(GND_net), .CO(n39256));
    SB_LUT4 i15386_3_lut (.I0(\data_in_frame[13] [4]), .I1(rx_data[4]), 
            .I2(n43847), .I3(GND_net), .O(n29334));   // verilog/coms.v(128[12] 303[6])
    defparam i15386_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_2173_4_lut (.I0(GND_net), .I1(n3233), 
            .I2(VCC_net), .I3(n39254), .O(n3300)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2173_4 (.CI(n39254), .I0(n3233), 
            .I1(VCC_net), .CO(n39255));
    SB_LUT4 encoder0_position_31__I_0_add_2173_3_lut (.I0(GND_net), .I1(n543), 
            .I2(GND_net), .I3(n39253), .O(n3301)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2173_3 (.CI(n39253), .I0(n543), 
            .I1(GND_net), .CO(n39254));
    SB_LUT4 i15387_3_lut (.I0(\data_in_frame[13] [3]), .I1(rx_data[3]), 
            .I2(n43847), .I3(GND_net), .O(n29335));   // verilog/coms.v(128[12] 303[6])
    defparam i15387_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_2173_2 (.CI(VCC_net), .I0(n544), 
            .I1(VCC_net), .CO(n39253));
    SB_LUT4 encoder0_position_31__I_0_add_2106_31_lut (.I0(n50544), .I1(n3105), 
            .I2(VCC_net), .I3(n39252), .O(n3204)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_31_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i15388_3_lut (.I0(\data_in_frame[13] [2]), .I1(rx_data[2]), 
            .I2(n43847), .I3(GND_net), .O(n29336));   // verilog/coms.v(128[12] 303[6])
    defparam i15388_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_2106_30_lut (.I0(GND_net), .I1(n3106), 
            .I2(VCC_net), .I3(n39251), .O(n3173)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_30_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15518_3_lut (.I0(neopxl_color[1]), .I1(\data_in_frame[6] [1]), 
            .I2(n28522), .I3(GND_net), .O(n29466));   // verilog/coms.v(128[12] 303[6])
    defparam i15518_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_31__I_0_add_2106_30 (.CI(n39251), .I0(n3106), 
            .I1(VCC_net), .CO(n39252));
    SB_LUT4 i15390_3_lut (.I0(\data_in_frame[13] [1]), .I1(rx_data[1]), 
            .I2(n43847), .I3(GND_net), .O(n29338));   // verilog/coms.v(128[12] 303[6])
    defparam i15390_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_2106_29_lut (.I0(GND_net), .I1(n3107), 
            .I2(VCC_net), .I3(n39250), .O(n3174)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2106_29 (.CI(n39250), .I0(n3107), 
            .I1(VCC_net), .CO(n39251));
    SB_LUT4 i15519_4_lut (.I0(r_Rx_Data), .I1(rx_data[2]), .I2(n4_adj_5245), 
            .I3(n27131), .O(n29467));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i15519_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i15520_3_lut (.I0(\neo_pixel_transmitter.t0 [31]), .I1(timer[31]), 
            .I2(n42404), .I3(GND_net), .O(n29468));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15520_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_2106_28_lut (.I0(GND_net), .I1(n3108), 
            .I2(VCC_net), .I3(n39249), .O(n3175)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2106_28 (.CI(n39249), .I0(n3108), 
            .I1(VCC_net), .CO(n39250));
    SB_LUT4 encoder0_position_31__I_0_add_2106_27_lut (.I0(GND_net), .I1(n3109), 
            .I2(VCC_net), .I3(n39248), .O(n3176)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2106_27 (.CI(n39248), .I0(n3109), 
            .I1(VCC_net), .CO(n39249));
    SB_LUT4 encoder0_position_31__I_0_add_2106_26_lut (.I0(GND_net), .I1(n3110), 
            .I2(VCC_net), .I3(n39247), .O(n3177)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_26_lut.LUT_INIT = 16'hC33C;
    SB_DFFESR delay_counter_i0_i10 (.Q(delay_counter[10]), .C(CLK_c), .E(n7417), 
            .D(n1318), .R(n28933));   // verilog/TinyFPGA_B.v(375[10] 403[6])
    SB_CARRY encoder0_position_31__I_0_add_2106_26 (.CI(n39247), .I0(n3110), 
            .I1(VCC_net), .CO(n39248));
    SB_LUT4 encoder0_position_31__I_0_add_2106_25_lut (.I0(GND_net), .I1(n3111), 
            .I2(VCC_net), .I3(n39246), .O(n3178)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2106_25 (.CI(n39246), .I0(n3111), 
            .I1(VCC_net), .CO(n39247));
    SB_LUT4 encoder0_position_31__I_0_add_2106_24_lut (.I0(GND_net), .I1(n3112), 
            .I2(VCC_net), .I3(n39245), .O(n3179)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15521_3_lut (.I0(\neo_pixel_transmitter.t0 [30]), .I1(timer[30]), 
            .I2(n42404), .I3(GND_net), .O(n29469));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15521_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15522_3_lut (.I0(\neo_pixel_transmitter.t0 [29]), .I1(timer[29]), 
            .I2(n42404), .I3(GND_net), .O(n29470));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15522_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_2106_24 (.CI(n39245), .I0(n3112), 
            .I1(VCC_net), .CO(n39246));
    SB_LUT4 encoder0_position_31__I_0_add_2106_23_lut (.I0(GND_net), .I1(n3113), 
            .I2(VCC_net), .I3(n39244), .O(n3180)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2106_23 (.CI(n39244), .I0(n3113), 
            .I1(VCC_net), .CO(n39245));
    SB_LUT4 encoder0_position_31__I_0_add_2106_22_lut (.I0(GND_net), .I1(n3114), 
            .I2(VCC_net), .I3(n39243), .O(n3181)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2106_22 (.CI(n39243), .I0(n3114), 
            .I1(VCC_net), .CO(n39244));
    SB_LUT4 encoder0_position_31__I_0_add_2106_21_lut (.I0(GND_net), .I1(n3115), 
            .I2(VCC_net), .I3(n39242), .O(n3182)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15523_3_lut (.I0(\neo_pixel_transmitter.t0 [28]), .I1(timer[28]), 
            .I2(n42404), .I3(GND_net), .O(n29471));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15523_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_2106_21 (.CI(n39242), .I0(n3115), 
            .I1(VCC_net), .CO(n39243));
    SB_LUT4 encoder0_position_31__I_0_add_2106_20_lut (.I0(GND_net), .I1(n3116), 
            .I2(VCC_net), .I3(n39241), .O(n3183)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2106_20 (.CI(n39241), .I0(n3116), 
            .I1(VCC_net), .CO(n39242));
    SB_LUT4 encoder0_position_31__I_0_add_2106_19_lut (.I0(GND_net), .I1(n3117), 
            .I2(VCC_net), .I3(n39240), .O(n3184)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2106_19 (.CI(n39240), .I0(n3117), 
            .I1(VCC_net), .CO(n39241));
    SB_LUT4 encoder0_position_31__I_0_add_2106_18_lut (.I0(GND_net), .I1(n3118), 
            .I2(VCC_net), .I3(n39239), .O(n3185)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2106_18 (.CI(n39239), .I0(n3118), 
            .I1(VCC_net), .CO(n39240));
    SB_LUT4 i15524_3_lut (.I0(\neo_pixel_transmitter.t0 [27]), .I1(timer[27]), 
            .I2(n42404), .I3(GND_net), .O(n29472));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15524_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_2106_17_lut (.I0(GND_net), .I1(n3119), 
            .I2(VCC_net), .I3(n39238), .O(n3186)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_236_6 (.CI(n38480), .I0(encoder1_position[7]), .I1(GND_net), 
            .CO(n38481));
    SB_CARRY encoder0_position_31__I_0_add_2106_17 (.CI(n39238), .I0(n3119), 
            .I1(VCC_net), .CO(n39239));
    SB_LUT4 encoder0_position_31__I_0_add_2106_16_lut (.I0(GND_net), .I1(n3120), 
            .I2(VCC_net), .I3(n39237), .O(n3187)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2106_16 (.CI(n39237), .I0(n3120), 
            .I1(VCC_net), .CO(n39238));
    SB_LUT4 encoder0_position_31__I_0_add_2106_15_lut (.I0(GND_net), .I1(n3121), 
            .I2(VCC_net), .I3(n39236), .O(n3188)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2106_15 (.CI(n39236), .I0(n3121), 
            .I1(VCC_net), .CO(n39237));
    SB_LUT4 encoder0_position_31__I_0_add_2106_14_lut (.I0(GND_net), .I1(n3122), 
            .I2(VCC_net), .I3(n39235), .O(n3189)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2106_14 (.CI(n39235), .I0(n3122), 
            .I1(VCC_net), .CO(n39236));
    SB_LUT4 encoder0_position_31__I_0_add_2106_13_lut (.I0(GND_net), .I1(n3123), 
            .I2(VCC_net), .I3(n39234), .O(n3190)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2106_13 (.CI(n39234), .I0(n3123), 
            .I1(VCC_net), .CO(n39235));
    SB_LUT4 encoder0_position_31__I_0_add_2106_12_lut (.I0(GND_net), .I1(n3124), 
            .I2(VCC_net), .I3(n39233), .O(n3191)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2106_12 (.CI(n39233), .I0(n3124), 
            .I1(VCC_net), .CO(n39234));
    SB_LUT4 encoder0_position_31__I_0_add_2106_11_lut (.I0(GND_net), .I1(n3125), 
            .I2(VCC_net), .I3(n39232), .O(n3192)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2106_11 (.CI(n39232), .I0(n3125), 
            .I1(VCC_net), .CO(n39233));
    SB_LUT4 encoder0_position_31__I_0_add_2106_10_lut (.I0(GND_net), .I1(n3126), 
            .I2(VCC_net), .I3(n39231), .O(n3193)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2106_10 (.CI(n39231), .I0(n3126), 
            .I1(VCC_net), .CO(n39232));
    SB_LUT4 encoder0_position_31__I_0_add_2106_9_lut (.I0(GND_net), .I1(n3127), 
            .I2(VCC_net), .I3(n39230), .O(n3194)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2106_9 (.CI(n39230), .I0(n3127), 
            .I1(VCC_net), .CO(n39231));
    SB_LUT4 encoder0_position_31__I_0_add_2106_8_lut (.I0(GND_net), .I1(n3128), 
            .I2(VCC_net), .I3(n39229), .O(n3195)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2106_8 (.CI(n39229), .I0(n3128), 
            .I1(VCC_net), .CO(n39230));
    SB_LUT4 encoder0_position_31__I_0_add_2106_7_lut (.I0(GND_net), .I1(n3129), 
            .I2(GND_net), .I3(n39228), .O(n3196)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2106_7 (.CI(n39228), .I0(n3129), 
            .I1(GND_net), .CO(n39229));
    SB_LUT4 encoder0_position_31__I_0_add_2106_6_lut (.I0(GND_net), .I1(n3130), 
            .I2(GND_net), .I3(n39227), .O(n3197)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2106_6 (.CI(n39227), .I0(n3130), 
            .I1(GND_net), .CO(n39228));
    SB_LUT4 encoder0_position_31__I_0_add_2106_5_lut (.I0(GND_net), .I1(n3131), 
            .I2(VCC_net), .I3(n39226), .O(n3198)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2106_5 (.CI(n39226), .I0(n3131), 
            .I1(VCC_net), .CO(n39227));
    SB_LUT4 i15525_3_lut (.I0(\neo_pixel_transmitter.t0 [26]), .I1(timer[26]), 
            .I2(n42404), .I3(GND_net), .O(n29473));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15525_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_2106_4_lut (.I0(GND_net), .I1(n3132), 
            .I2(GND_net), .I3(n39225), .O(n3199)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2106_4 (.CI(n39225), .I0(n3132), 
            .I1(GND_net), .CO(n39226));
    SB_LUT4 encoder0_position_31__I_0_add_2106_3_lut (.I0(GND_net), .I1(n3133), 
            .I2(VCC_net), .I3(n39224), .O(n3200)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2106_3 (.CI(n39224), .I0(n3133), 
            .I1(VCC_net), .CO(n39225));
    SB_LUT4 encoder0_position_31__I_0_add_2106_2_lut (.I0(GND_net), .I1(n542), 
            .I2(GND_net), .I3(VCC_net), .O(n3201)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2106_2 (.CI(VCC_net), .I0(n542), 
            .I1(GND_net), .CO(n39224));
    SB_LUT4 encoder0_position_31__I_0_add_2039_30_lut (.I0(n50593), .I1(n3006), 
            .I2(VCC_net), .I3(n39223), .O(n3105)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_30_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_31__I_0_add_2039_29_lut (.I0(GND_net), .I1(n3007), 
            .I2(VCC_net), .I3(n39222), .O(n3074)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_29_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15526_3_lut (.I0(\neo_pixel_transmitter.t0 [25]), .I1(timer[25]), 
            .I2(n42404), .I3(GND_net), .O(n29474));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15526_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_2039_29 (.CI(n39222), .I0(n3007), 
            .I1(VCC_net), .CO(n39223));
    SB_LUT4 encoder0_position_31__I_0_add_2039_28_lut (.I0(GND_net), .I1(n3008), 
            .I2(VCC_net), .I3(n39221), .O(n3075)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2039_28 (.CI(n39221), .I0(n3008), 
            .I1(VCC_net), .CO(n39222));
    SB_LUT4 encoder0_position_31__I_0_add_2039_27_lut (.I0(GND_net), .I1(n3009), 
            .I2(VCC_net), .I3(n39220), .O(n3076)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_27_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15527_3_lut (.I0(\neo_pixel_transmitter.t0 [24]), .I1(timer[24]), 
            .I2(n42404), .I3(GND_net), .O(n29475));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15527_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_2039_27 (.CI(n39220), .I0(n3009), 
            .I1(VCC_net), .CO(n39221));
    SB_LUT4 encoder0_position_31__I_0_add_2039_26_lut (.I0(GND_net), .I1(n3010), 
            .I2(VCC_net), .I3(n39219), .O(n3077)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2039_26 (.CI(n39219), .I0(n3010), 
            .I1(VCC_net), .CO(n39220));
    SB_LUT4 encoder0_position_31__I_0_add_2039_25_lut (.I0(GND_net), .I1(n3011), 
            .I2(VCC_net), .I3(n39218), .O(n3078)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2039_25 (.CI(n39218), .I0(n3011), 
            .I1(VCC_net), .CO(n39219));
    SB_LUT4 encoder0_position_31__I_0_add_2039_24_lut (.I0(GND_net), .I1(n3012), 
            .I2(VCC_net), .I3(n39217), .O(n3079)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2039_24 (.CI(n39217), .I0(n3012), 
            .I1(VCC_net), .CO(n39218));
    SB_LUT4 encoder0_position_31__I_0_add_2039_23_lut (.I0(GND_net), .I1(n3013), 
            .I2(VCC_net), .I3(n39216), .O(n3080)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2039_23 (.CI(n39216), .I0(n3013), 
            .I1(VCC_net), .CO(n39217));
    SB_LUT4 encoder0_position_31__I_0_add_2039_22_lut (.I0(GND_net), .I1(n3014), 
            .I2(VCC_net), .I3(n39215), .O(n3081)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_236_5_lut (.I0(GND_net), .I1(encoder1_position[6]), .I2(GND_net), 
            .I3(n38479), .O(encoder1_position_scaled_23__N_75[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_236_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2039_22 (.CI(n39215), .I0(n3014), 
            .I1(VCC_net), .CO(n39216));
    SB_LUT4 encoder0_position_31__I_0_add_2039_21_lut (.I0(GND_net), .I1(n3015), 
            .I2(VCC_net), .I3(n39214), .O(n3082)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2039_21 (.CI(n39214), .I0(n3015), 
            .I1(VCC_net), .CO(n39215));
    SB_LUT4 encoder0_position_31__I_0_add_2039_20_lut (.I0(GND_net), .I1(n3016), 
            .I2(VCC_net), .I3(n39213), .O(n3083)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2039_20 (.CI(n39213), .I0(n3016), 
            .I1(VCC_net), .CO(n39214));
    SB_LUT4 i15528_3_lut (.I0(\neo_pixel_transmitter.t0 [23]), .I1(timer[23]), 
            .I2(n42404), .I3(GND_net), .O(n29476));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15528_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_2039_19_lut (.I0(GND_net), .I1(n3017), 
            .I2(VCC_net), .I3(n39212), .O(n3084)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2039_19 (.CI(n39212), .I0(n3017), 
            .I1(VCC_net), .CO(n39213));
    SB_LUT4 encoder0_position_31__I_0_add_2039_18_lut (.I0(GND_net), .I1(n3018), 
            .I2(VCC_net), .I3(n39211), .O(n3085)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2039_18 (.CI(n39211), .I0(n3018), 
            .I1(VCC_net), .CO(n39212));
    SB_LUT4 encoder0_position_31__I_0_add_2039_17_lut (.I0(GND_net), .I1(n3019), 
            .I2(VCC_net), .I3(n39210), .O(n3086)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2039_17 (.CI(n39210), .I0(n3019), 
            .I1(VCC_net), .CO(n39211));
    SB_LUT4 encoder0_position_31__I_0_add_2039_16_lut (.I0(GND_net), .I1(n3020), 
            .I2(VCC_net), .I3(n39209), .O(n3087)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2039_16 (.CI(n39209), .I0(n3020), 
            .I1(VCC_net), .CO(n39210));
    SB_LUT4 encoder0_position_31__I_0_add_2039_15_lut (.I0(GND_net), .I1(n3021), 
            .I2(VCC_net), .I3(n39208), .O(n3088)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15529_3_lut (.I0(\neo_pixel_transmitter.t0 [22]), .I1(timer[22]), 
            .I2(n42404), .I3(GND_net), .O(n29477));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15529_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15530_3_lut (.I0(\neo_pixel_transmitter.t0 [21]), .I1(timer[21]), 
            .I2(n42404), .I3(GND_net), .O(n29478));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15530_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_2039_15 (.CI(n39208), .I0(n3021), 
            .I1(VCC_net), .CO(n39209));
    SB_LUT4 encoder0_position_31__I_0_add_2039_14_lut (.I0(GND_net), .I1(n3022), 
            .I2(VCC_net), .I3(n39207), .O(n3089)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2039_14 (.CI(n39207), .I0(n3022), 
            .I1(VCC_net), .CO(n39208));
    SB_LUT4 encoder0_position_31__I_0_add_2039_13_lut (.I0(GND_net), .I1(n3023), 
            .I2(VCC_net), .I3(n39206), .O(n3090)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2039_13 (.CI(n39206), .I0(n3023), 
            .I1(VCC_net), .CO(n39207));
    SB_LUT4 encoder0_position_31__I_0_add_2039_12_lut (.I0(GND_net), .I1(n3024), 
            .I2(VCC_net), .I3(n39205), .O(n3091)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2039_12 (.CI(n39205), .I0(n3024), 
            .I1(VCC_net), .CO(n39206));
    SB_LUT4 encoder0_position_31__I_0_add_2039_11_lut (.I0(GND_net), .I1(n3025), 
            .I2(VCC_net), .I3(n39204), .O(n3092)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_11_lut.LUT_INIT = 16'hC33C;
    SB_IO CS_MISO_pad (.PACKAGE_PIN(CS_MISO), .OUTPUT_ENABLE(VCC_net), .D_IN_0(CS_MISO_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam CS_MISO_pad.PIN_TYPE = 6'b000001;
    defparam CS_MISO_pad.PULLUP = 1'b0;
    defparam CS_MISO_pad.NEG_TRIGGER = 1'b0;
    defparam CS_MISO_pad.IO_STANDARD = "SB_LVCMOS";
    SB_CARRY encoder0_position_31__I_0_add_2039_11 (.CI(n39204), .I0(n3025), 
            .I1(VCC_net), .CO(n39205));
    SB_CARRY add_236_5 (.CI(n38479), .I0(encoder1_position[6]), .I1(GND_net), 
            .CO(n38480));
    SB_LUT4 encoder0_position_31__I_0_add_2039_10_lut (.I0(GND_net), .I1(n3026), 
            .I2(VCC_net), .I3(n39203), .O(n3093)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15531_3_lut (.I0(\neo_pixel_transmitter.t0 [20]), .I1(timer[20]), 
            .I2(n42404), .I3(GND_net), .O(n29479));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15531_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_2039_10 (.CI(n39203), .I0(n3026), 
            .I1(VCC_net), .CO(n39204));
    SB_LUT4 encoder0_position_31__I_0_add_2039_9_lut (.I0(GND_net), .I1(n3027), 
            .I2(VCC_net), .I3(n39202), .O(n3094)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2039_9 (.CI(n39202), .I0(n3027), 
            .I1(VCC_net), .CO(n39203));
    SB_LUT4 encoder0_position_31__I_0_add_2039_8_lut (.I0(GND_net), .I1(n3028), 
            .I2(VCC_net), .I3(n39201), .O(n3095)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2039_8 (.CI(n39201), .I0(n3028), 
            .I1(VCC_net), .CO(n39202));
    SB_LUT4 encoder0_position_31__I_0_add_2039_7_lut (.I0(GND_net), .I1(n3029), 
            .I2(GND_net), .I3(n39200), .O(n3096)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15179_3_lut (.I0(\data_out_frame[4] [4]), .I1(ID[4]), .I2(n24278), 
            .I3(GND_net), .O(n29127));   // verilog/coms.v(128[12] 303[6])
    defparam i15179_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_250_i18_4_lut (.I0(encoder1_position_scaled[17]), .I1(displacement[17]), 
            .I2(n15_adj_5249), .I3(n15_adj_5321), .O(motor_state_23__N_123[17]));   // verilog/TinyFPGA_B.v(285[5] 287[10])
    defparam mux_250_i18_4_lut.LUT_INIT = 16'h0aca;
    SB_CARRY encoder0_position_31__I_0_add_2039_7 (.CI(n39200), .I0(n3029), 
            .I1(GND_net), .CO(n39201));
    SB_LUT4 encoder0_position_31__I_0_add_2039_6_lut (.I0(GND_net), .I1(n3030), 
            .I2(GND_net), .I3(n39199), .O(n3097)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2039_6 (.CI(n39199), .I0(n3030), 
            .I1(GND_net), .CO(n39200));
    SB_LUT4 encoder0_position_31__I_0_add_2039_5_lut (.I0(GND_net), .I1(n3031), 
            .I2(VCC_net), .I3(n39198), .O(n3098)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2039_5 (.CI(n39198), .I0(n3031), 
            .I1(VCC_net), .CO(n39199));
    SB_LUT4 i15180_3_lut (.I0(\data_out_frame[4] [3]), .I1(ID[3]), .I2(n24278), 
            .I3(GND_net), .O(n29128));   // verilog/coms.v(128[12] 303[6])
    defparam i15180_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_add_2039_4_lut (.I0(GND_net), .I1(n3032), 
            .I2(GND_net), .I3(n39197), .O(n3099)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15181_3_lut (.I0(\data_out_frame[4] [2]), .I1(ID[2]), .I2(n24278), 
            .I3(GND_net), .O(n29129));   // verilog/coms.v(128[12] 303[6])
    defparam i15181_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_31__I_0_add_2039_4 (.CI(n39197), .I0(n3032), 
            .I1(GND_net), .CO(n39198));
    SB_LUT4 encoder0_position_31__I_0_add_2039_3_lut (.I0(GND_net), .I1(n3033), 
            .I2(VCC_net), .I3(n39196), .O(n3100)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2039_3 (.CI(n39196), .I0(n3033), 
            .I1(VCC_net), .CO(n39197));
    SB_LUT4 i15532_3_lut (.I0(\neo_pixel_transmitter.t0 [19]), .I1(timer[19]), 
            .I2(n42404), .I3(GND_net), .O(n29480));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15532_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_2039_2_lut (.I0(GND_net), .I1(n541), 
            .I2(GND_net), .I3(VCC_net), .O(n3101)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15533_3_lut (.I0(\neo_pixel_transmitter.t0 [18]), .I1(timer[18]), 
            .I2(n42404), .I3(GND_net), .O(n29481));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15533_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15182_3_lut (.I0(\data_out_frame[4] [1]), .I1(ID[1]), .I2(n24278), 
            .I3(GND_net), .O(n29130));   // verilog/coms.v(128[12] 303[6])
    defparam i15182_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15534_3_lut (.I0(\neo_pixel_transmitter.t0 [17]), .I1(timer[17]), 
            .I2(n42404), .I3(GND_net), .O(n29482));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15534_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15535_3_lut (.I0(\neo_pixel_transmitter.t0 [16]), .I1(timer[16]), 
            .I2(n42404), .I3(GND_net), .O(n29483));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15535_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15183_3_lut (.I0(\data_out_frame[4] [0]), .I1(ID[0]), .I2(n24278), 
            .I3(GND_net), .O(n29131));   // verilog/coms.v(128[12] 303[6])
    defparam i15183_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_31__I_0_add_2039_2 (.CI(VCC_net), .I0(n541), 
            .I1(GND_net), .CO(n39196));
    SB_LUT4 encoder0_position_31__I_0_add_1972_29_lut (.I0(n50635), .I1(n2907), 
            .I2(VCC_net), .I3(n39195), .O(n3006)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_29_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_31__I_0_add_1972_28_lut (.I0(GND_net), .I1(n2908), 
            .I2(VCC_net), .I3(n39194), .O(n2975)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1972_28 (.CI(n39194), .I0(n2908), 
            .I1(VCC_net), .CO(n39195));
    SB_LUT4 encoder0_position_31__I_0_add_1972_27_lut (.I0(GND_net), .I1(n2909), 
            .I2(VCC_net), .I3(n39193), .O(n2976)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_27_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15184_3_lut (.I0(IntegralLimit[23]), .I1(\data_in_frame[11] [7]), 
            .I2(n28521), .I3(GND_net), .O(n29132));   // verilog/coms.v(128[12] 303[6])
    defparam i15184_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15185_3_lut (.I0(IntegralLimit[22]), .I1(\data_in_frame[11] [6]), 
            .I2(n28521), .I3(GND_net), .O(n29133));   // verilog/coms.v(128[12] 303[6])
    defparam i15185_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15186_3_lut (.I0(IntegralLimit[21]), .I1(\data_in_frame[11] [5]), 
            .I2(n28521), .I3(GND_net), .O(n29134));   // verilog/coms.v(128[12] 303[6])
    defparam i15186_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_236_4_lut (.I0(GND_net), .I1(encoder1_position[5]), .I2(GND_net), 
            .I3(n38478), .O(encoder1_position_scaled_23__N_75[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_236_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1972_27 (.CI(n39193), .I0(n2909), 
            .I1(VCC_net), .CO(n39194));
    SB_LUT4 encoder0_position_31__I_0_add_1972_26_lut (.I0(GND_net), .I1(n2910), 
            .I2(VCC_net), .I3(n39192), .O(n2977)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1972_26 (.CI(n39192), .I0(n2910), 
            .I1(VCC_net), .CO(n39193));
    SB_LUT4 encoder0_position_31__I_0_add_1972_25_lut (.I0(GND_net), .I1(n2911), 
            .I2(VCC_net), .I3(n39191), .O(n2978)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1972_25 (.CI(n39191), .I0(n2911), 
            .I1(VCC_net), .CO(n39192));
    SB_LUT4 i15536_3_lut (.I0(\neo_pixel_transmitter.t0 [15]), .I1(timer[15]), 
            .I2(n42404), .I3(GND_net), .O(n29484));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15536_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1972_24_lut (.I0(GND_net), .I1(n2912), 
            .I2(VCC_net), .I3(n39190), .O(n2979)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1972_24 (.CI(n39190), .I0(n2912), 
            .I1(VCC_net), .CO(n39191));
    SB_LUT4 encoder0_position_31__I_0_add_1972_23_lut (.I0(GND_net), .I1(n2913), 
            .I2(VCC_net), .I3(n39189), .O(n2980)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1972_23 (.CI(n39189), .I0(n2913), 
            .I1(VCC_net), .CO(n39190));
    SB_LUT4 encoder0_position_31__I_0_add_1972_22_lut (.I0(GND_net), .I1(n2914), 
            .I2(VCC_net), .I3(n39188), .O(n2981)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15537_3_lut (.I0(\neo_pixel_transmitter.t0 [14]), .I1(timer[14]), 
            .I2(n42404), .I3(GND_net), .O(n29485));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15537_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15538_3_lut (.I0(\neo_pixel_transmitter.t0 [13]), .I1(timer[13]), 
            .I2(n42404), .I3(GND_net), .O(n29486));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15538_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15539_3_lut (.I0(\neo_pixel_transmitter.t0 [12]), .I1(timer[12]), 
            .I2(n42404), .I3(GND_net), .O(n29487));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15539_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_1972_22 (.CI(n39188), .I0(n2914), 
            .I1(VCC_net), .CO(n39189));
    SB_LUT4 i15187_3_lut (.I0(IntegralLimit[20]), .I1(\data_in_frame[11] [4]), 
            .I2(n28521), .I3(GND_net), .O(n29135));   // verilog/coms.v(128[12] 303[6])
    defparam i15187_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_add_1972_21_lut (.I0(GND_net), .I1(n2915), 
            .I2(VCC_net), .I3(n39187), .O(n2982)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1972_21 (.CI(n39187), .I0(n2915), 
            .I1(VCC_net), .CO(n39188));
    SB_LUT4 i15188_3_lut (.I0(IntegralLimit[19]), .I1(\data_in_frame[11] [3]), 
            .I2(n28521), .I3(GND_net), .O(n29136));   // verilog/coms.v(128[12] 303[6])
    defparam i15188_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_add_1972_20_lut (.I0(GND_net), .I1(n2916), 
            .I2(VCC_net), .I3(n39186), .O(n2983)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1972_20 (.CI(n39186), .I0(n2916), 
            .I1(VCC_net), .CO(n39187));
    SB_LUT4 encoder0_position_31__I_0_add_1972_19_lut (.I0(GND_net), .I1(n2917), 
            .I2(VCC_net), .I3(n39185), .O(n2984)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15189_3_lut (.I0(IntegralLimit[18]), .I1(\data_in_frame[11] [2]), 
            .I2(n28521), .I3(GND_net), .O(n29137));   // verilog/coms.v(128[12] 303[6])
    defparam i15189_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_31__I_0_add_1972_19 (.CI(n39185), .I0(n2917), 
            .I1(VCC_net), .CO(n39186));
    SB_LUT4 encoder0_position_31__I_0_add_1972_18_lut (.I0(GND_net), .I1(n2918), 
            .I2(VCC_net), .I3(n39184), .O(n2985)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1972_18 (.CI(n39184), .I0(n2918), 
            .I1(VCC_net), .CO(n39185));
    SB_LUT4 encoder0_position_31__I_0_add_1972_17_lut (.I0(GND_net), .I1(n2919), 
            .I2(VCC_net), .I3(n39183), .O(n2986)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1972_17 (.CI(n39183), .I0(n2919), 
            .I1(VCC_net), .CO(n39184));
    SB_LUT4 encoder0_position_31__I_0_add_1972_16_lut (.I0(GND_net), .I1(n2920), 
            .I2(VCC_net), .I3(n39182), .O(n2987)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1972_16 (.CI(n39182), .I0(n2920), 
            .I1(VCC_net), .CO(n39183));
    SB_LUT4 encoder0_position_31__I_0_add_1972_15_lut (.I0(GND_net), .I1(n2921), 
            .I2(VCC_net), .I3(n39181), .O(n2988)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1972_15 (.CI(n39181), .I0(n2921), 
            .I1(VCC_net), .CO(n39182));
    SB_LUT4 encoder0_position_31__I_0_add_1972_14_lut (.I0(GND_net), .I1(n2922), 
            .I2(VCC_net), .I3(n39180), .O(n2989)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1972_14 (.CI(n39180), .I0(n2922), 
            .I1(VCC_net), .CO(n39181));
    SB_LUT4 encoder0_position_31__I_0_add_1972_13_lut (.I0(GND_net), .I1(n2923), 
            .I2(VCC_net), .I3(n39179), .O(n2990)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1972_13 (.CI(n39179), .I0(n2923), 
            .I1(VCC_net), .CO(n39180));
    SB_LUT4 encoder0_position_31__I_0_add_1972_12_lut (.I0(GND_net), .I1(n2924), 
            .I2(VCC_net), .I3(n39178), .O(n2991)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_236_4 (.CI(n38478), .I0(encoder1_position[5]), .I1(GND_net), 
            .CO(n38479));
    SB_CARRY encoder0_position_31__I_0_add_1972_12 (.CI(n39178), .I0(n2924), 
            .I1(VCC_net), .CO(n39179));
    SB_LUT4 encoder0_position_31__I_0_add_1972_11_lut (.I0(GND_net), .I1(n2925), 
            .I2(VCC_net), .I3(n39177), .O(n2992)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1972_11 (.CI(n39177), .I0(n2925), 
            .I1(VCC_net), .CO(n39178));
    SB_LUT4 encoder0_position_31__I_0_add_1972_10_lut (.I0(GND_net), .I1(n2926), 
            .I2(VCC_net), .I3(n39176), .O(n2993)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1972_10 (.CI(n39176), .I0(n2926), 
            .I1(VCC_net), .CO(n39177));
    SB_LUT4 encoder0_position_31__I_0_add_1972_9_lut (.I0(GND_net), .I1(n2927), 
            .I2(VCC_net), .I3(n39175), .O(n2994)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1972_9 (.CI(n39175), .I0(n2927), 
            .I1(VCC_net), .CO(n39176));
    SB_LUT4 i15540_3_lut (.I0(\neo_pixel_transmitter.t0 [11]), .I1(timer[11]), 
            .I2(n42404), .I3(GND_net), .O(n29488));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15540_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1972_8_lut (.I0(GND_net), .I1(n2928), 
            .I2(VCC_net), .I3(n39174), .O(n2995)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1972_8 (.CI(n39174), .I0(n2928), 
            .I1(VCC_net), .CO(n39175));
    SB_LUT4 encoder0_position_31__I_0_add_1972_7_lut (.I0(GND_net), .I1(n2929), 
            .I2(GND_net), .I3(n39173), .O(n2996)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1972_7 (.CI(n39173), .I0(n2929), 
            .I1(GND_net), .CO(n39174));
    SB_LUT4 encoder0_position_31__I_0_add_1972_6_lut (.I0(GND_net), .I1(n2930), 
            .I2(GND_net), .I3(n39172), .O(n2997)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_250_i19_4_lut (.I0(encoder1_position_scaled[18]), .I1(displacement[18]), 
            .I2(n15_adj_5249), .I3(n15_adj_5321), .O(motor_state_23__N_123[18]));   // verilog/TinyFPGA_B.v(285[5] 287[10])
    defparam mux_250_i19_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 n10621_bdd_4_lut_35819 (.I0(n10621), .I1(current[15]), .I2(duty[19]), 
            .I3(n4208), .O(n51444));
    defparam n10621_bdd_4_lut_35819.LUT_INIT = 16'he4aa;
    SB_CARRY encoder0_position_31__I_0_add_1972_6 (.CI(n39172), .I0(n2930), 
            .I1(GND_net), .CO(n39173));
    SB_LUT4 i15190_4_lut (.I0(CS_MISO_c), .I1(data_adj_5514[4]), .I2(n6_adj_5340), 
            .I3(n27143), .O(n29138));   // verilog/tli4970.v(35[10] 68[6])
    defparam i15190_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i15191_3_lut (.I0(IntegralLimit[17]), .I1(\data_in_frame[11] [1]), 
            .I2(n28521), .I3(GND_net), .O(n29139));   // verilog/coms.v(128[12] 303[6])
    defparam i15191_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_add_1972_5_lut (.I0(GND_net), .I1(n2931), 
            .I2(VCC_net), .I3(n39171), .O(n2998)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1972_5 (.CI(n39171), .I0(n2931), 
            .I1(VCC_net), .CO(n39172));
    SB_LUT4 i15541_3_lut (.I0(\neo_pixel_transmitter.t0 [10]), .I1(timer[10]), 
            .I2(n42404), .I3(GND_net), .O(n29489));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15541_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1972_4_lut (.I0(GND_net), .I1(n2932), 
            .I2(GND_net), .I3(n39170), .O(n2999)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1972_4 (.CI(n39170), .I0(n2932), 
            .I1(GND_net), .CO(n39171));
    SB_LUT4 encoder0_position_31__I_0_add_1972_3_lut (.I0(GND_net), .I1(n2933), 
            .I2(VCC_net), .I3(n39169), .O(n3000)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1972_3 (.CI(n39169), .I0(n2933), 
            .I1(VCC_net), .CO(n39170));
    SB_LUT4 encoder0_position_31__I_0_add_1972_2_lut (.I0(GND_net), .I1(n540), 
            .I2(GND_net), .I3(VCC_net), .O(n3001)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1972_2 (.CI(VCC_net), .I0(n540), 
            .I1(GND_net), .CO(n39169));
    SB_LUT4 encoder0_position_31__I_0_add_1905_28_lut (.I0(n50668), .I1(n2808), 
            .I2(VCC_net), .I3(n39168), .O(n2907)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_28_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_31__I_0_add_1905_27_lut (.I0(GND_net), .I1(n2809), 
            .I2(VCC_net), .I3(n39167), .O(n2876)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1905_27 (.CI(n39167), .I0(n2809), 
            .I1(VCC_net), .CO(n39168));
    SB_LUT4 i15192_3_lut (.I0(IntegralLimit[16]), .I1(\data_in_frame[11] [0]), 
            .I2(n28521), .I3(GND_net), .O(n29140));   // verilog/coms.v(128[12] 303[6])
    defparam i15192_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_add_1905_26_lut (.I0(GND_net), .I1(n2810), 
            .I2(VCC_net), .I3(n39166), .O(n2877)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1905_26 (.CI(n39166), .I0(n2810), 
            .I1(VCC_net), .CO(n39167));
    SB_LUT4 encoder0_position_31__I_0_add_1905_25_lut (.I0(GND_net), .I1(n2811), 
            .I2(VCC_net), .I3(n39165), .O(n2878)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1905_25 (.CI(n39165), .I0(n2811), 
            .I1(VCC_net), .CO(n39166));
    SB_LUT4 encoder0_position_31__I_0_add_1905_24_lut (.I0(GND_net), .I1(n2812), 
            .I2(VCC_net), .I3(n39164), .O(n2879)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_236_3_lut (.I0(GND_net), .I1(encoder1_position[4]), .I2(GND_net), 
            .I3(n38477), .O(encoder1_position_scaled_23__N_75[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_236_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1905_24 (.CI(n39164), .I0(n2812), 
            .I1(VCC_net), .CO(n39165));
    SB_LUT4 encoder0_position_31__I_0_add_1905_23_lut (.I0(GND_net), .I1(n2813), 
            .I2(VCC_net), .I3(n39163), .O(n2880)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1905_23 (.CI(n39163), .I0(n2813), 
            .I1(VCC_net), .CO(n39164));
    SB_LUT4 encoder0_position_31__I_0_add_1905_22_lut (.I0(GND_net), .I1(n2814), 
            .I2(VCC_net), .I3(n39162), .O(n2881)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1905_22 (.CI(n39162), .I0(n2814), 
            .I1(VCC_net), .CO(n39163));
    SB_LUT4 encoder0_position_31__I_0_add_1905_21_lut (.I0(GND_net), .I1(n2815), 
            .I2(VCC_net), .I3(n39161), .O(n2882)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1905_21 (.CI(n39161), .I0(n2815), 
            .I1(VCC_net), .CO(n39162));
    SB_LUT4 encoder0_position_31__I_0_add_1905_20_lut (.I0(GND_net), .I1(n2816), 
            .I2(VCC_net), .I3(n39160), .O(n2883)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1905_20 (.CI(n39160), .I0(n2816), 
            .I1(VCC_net), .CO(n39161));
    SB_LUT4 encoder0_position_31__I_0_add_1905_19_lut (.I0(GND_net), .I1(n2817), 
            .I2(VCC_net), .I3(n39159), .O(n2884)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1905_19 (.CI(n39159), .I0(n2817), 
            .I1(VCC_net), .CO(n39160));
    SB_LUT4 encoder0_position_31__I_0_add_1905_18_lut (.I0(GND_net), .I1(n2818), 
            .I2(VCC_net), .I3(n39158), .O(n2885)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1905_18 (.CI(n39158), .I0(n2818), 
            .I1(VCC_net), .CO(n39159));
    SB_LUT4 encoder0_position_31__I_0_add_1905_17_lut (.I0(GND_net), .I1(n2819), 
            .I2(VCC_net), .I3(n39157), .O(n2886)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_250_i20_4_lut (.I0(encoder1_position_scaled[19]), .I1(displacement[19]), 
            .I2(n15_adj_5249), .I3(n15_adj_5321), .O(motor_state_23__N_123[19]));   // verilog/TinyFPGA_B.v(285[5] 287[10])
    defparam mux_250_i20_4_lut.LUT_INIT = 16'h0aca;
    SB_CARRY encoder0_position_31__I_0_add_1905_17 (.CI(n39157), .I0(n2819), 
            .I1(VCC_net), .CO(n39158));
    SB_LUT4 encoder0_position_31__I_0_add_1905_16_lut (.I0(GND_net), .I1(n2820), 
            .I2(VCC_net), .I3(n39156), .O(n2887)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1905_16 (.CI(n39156), .I0(n2820), 
            .I1(VCC_net), .CO(n39157));
    SB_LUT4 encoder0_position_31__I_0_add_1905_15_lut (.I0(GND_net), .I1(n2821), 
            .I2(VCC_net), .I3(n39155), .O(n2888)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1905_15 (.CI(n39155), .I0(n2821), 
            .I1(VCC_net), .CO(n39156));
    SB_LUT4 encoder0_position_31__I_0_add_1905_14_lut (.I0(GND_net), .I1(n2822), 
            .I2(VCC_net), .I3(n39154), .O(n2889)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1905_14 (.CI(n39154), .I0(n2822), 
            .I1(VCC_net), .CO(n39155));
    SB_LUT4 encoder0_position_31__I_0_add_1905_13_lut (.I0(GND_net), .I1(n2823), 
            .I2(VCC_net), .I3(n39153), .O(n2890)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1905_13 (.CI(n39153), .I0(n2823), 
            .I1(VCC_net), .CO(n39154));
    SB_LUT4 encoder0_position_31__I_0_add_1905_12_lut (.I0(GND_net), .I1(n2824), 
            .I2(VCC_net), .I3(n39152), .O(n2891)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1905_12 (.CI(n39152), .I0(n2824), 
            .I1(VCC_net), .CO(n39153));
    SB_LUT4 encoder0_position_31__I_0_add_1905_11_lut (.I0(GND_net), .I1(n2825), 
            .I2(VCC_net), .I3(n39151), .O(n2892)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1905_11 (.CI(n39151), .I0(n2825), 
            .I1(VCC_net), .CO(n39152));
    SB_LUT4 encoder0_position_31__I_0_add_1905_10_lut (.I0(GND_net), .I1(n2826), 
            .I2(VCC_net), .I3(n39150), .O(n2893)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1905_10 (.CI(n39150), .I0(n2826), 
            .I1(VCC_net), .CO(n39151));
    SB_LUT4 encoder0_position_31__I_0_add_1905_9_lut (.I0(GND_net), .I1(n2827), 
            .I2(VCC_net), .I3(n39149), .O(n2894)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1905_9 (.CI(n39149), .I0(n2827), 
            .I1(VCC_net), .CO(n39150));
    SB_LUT4 encoder0_position_31__I_0_add_1905_8_lut (.I0(GND_net), .I1(n2828), 
            .I2(VCC_net), .I3(n39148), .O(n2895)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1905_8 (.CI(n39148), .I0(n2828), 
            .I1(VCC_net), .CO(n39149));
    SB_CARRY add_157_13 (.CI(n38456), .I0(delay_counter[11]), .I1(GND_net), 
            .CO(n38457));
    SB_LUT4 encoder0_position_31__I_0_add_1905_7_lut (.I0(GND_net), .I1(n2829), 
            .I2(GND_net), .I3(n39147), .O(n2896)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1905_7 (.CI(n39147), .I0(n2829), 
            .I1(GND_net), .CO(n39148));
    SB_LUT4 encoder0_position_31__I_0_add_1905_6_lut (.I0(GND_net), .I1(n2830), 
            .I2(GND_net), .I3(n39146), .O(n2897)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1905_6 (.CI(n39146), .I0(n2830), 
            .I1(GND_net), .CO(n39147));
    SB_LUT4 encoder0_position_31__I_0_add_1905_5_lut (.I0(GND_net), .I1(n2831), 
            .I2(VCC_net), .I3(n39145), .O(n2898)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1905_5 (.CI(n39145), .I0(n2831), 
            .I1(VCC_net), .CO(n39146));
    SB_LUT4 i15193_3_lut (.I0(IntegralLimit[15]), .I1(\data_in_frame[12] [7]), 
            .I2(n28521), .I3(GND_net), .O(n29141));   // verilog/coms.v(128[12] 303[6])
    defparam i15193_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_add_1905_4_lut (.I0(GND_net), .I1(n2832), 
            .I2(GND_net), .I3(n39144), .O(n2899)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1905_4 (.CI(n39144), .I0(n2832), 
            .I1(GND_net), .CO(n39145));
    SB_LUT4 encoder0_position_31__I_0_add_1905_3_lut (.I0(GND_net), .I1(n2833), 
            .I2(VCC_net), .I3(n39143), .O(n2900)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15194_3_lut (.I0(IntegralLimit[14]), .I1(\data_in_frame[12] [6]), 
            .I2(n28521), .I3(GND_net), .O(n29142));   // verilog/coms.v(128[12] 303[6])
    defparam i15194_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_31__I_0_add_1905_3 (.CI(n39143), .I0(n2833), 
            .I1(VCC_net), .CO(n39144));
    SB_LUT4 encoder0_position_31__I_0_add_1905_2_lut (.I0(GND_net), .I1(n539), 
            .I2(GND_net), .I3(VCC_net), .O(n2901)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1905_2 (.CI(VCC_net), .I0(n539), 
            .I1(GND_net), .CO(n39143));
    SB_LUT4 encoder0_position_31__I_0_add_1838_27_lut (.I0(GND_net), .I1(n2709), 
            .I2(VCC_net), .I3(n39142), .O(n2776)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_27_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1838_26_lut (.I0(GND_net), .I1(n2710), 
            .I2(VCC_net), .I3(n39141), .O(n2777)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1838_26 (.CI(n39141), .I0(n2710), 
            .I1(VCC_net), .CO(n39142));
    SB_LUT4 encoder0_position_31__I_0_add_1838_25_lut (.I0(GND_net), .I1(n2711), 
            .I2(VCC_net), .I3(n39140), .O(n2778)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1838_25 (.CI(n39140), .I0(n2711), 
            .I1(VCC_net), .CO(n39141));
    SB_LUT4 i15542_3_lut (.I0(\neo_pixel_transmitter.t0 [9]), .I1(timer[9]), 
            .I2(n42404), .I3(GND_net), .O(n29490));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15542_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1838_24_lut (.I0(GND_net), .I1(n2712), 
            .I2(VCC_net), .I3(n39139), .O(n2779)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i1_3_lut (.I0(encoder0_position[0]), 
            .I1(n33), .I2(encoder0_position[31]), .I3(GND_net), .O(n544));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_mux_3_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15543_3_lut (.I0(\neo_pixel_transmitter.t0 [8]), .I1(timer[8]), 
            .I2(n42404), .I3(GND_net), .O(n29491));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15543_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i35571_1_lut (.I0(n35558), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n51159));
    defparam i35571_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_i2200_3_lut (.I0(n3229), .I1(n3296), 
            .I2(n3237), .I3(GND_net), .O(n13_adj_5447));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i2200_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2191_3_lut (.I0(n3220), .I1(n3287), 
            .I2(n3237), .I3(GND_net), .O(n31_adj_5452));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i2191_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_1838_24 (.CI(n39139), .I0(n2712), 
            .I1(VCC_net), .CO(n39140));
    SB_LUT4 encoder0_position_31__I_0_i2198_3_lut (.I0(n3227), .I1(n3294), 
            .I2(n3237), .I3(GND_net), .O(n17_adj_5448));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i2198_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2197_3_lut (.I0(n3226), .I1(n3293), 
            .I2(n3237), .I3(GND_net), .O(n19_adj_5449));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i2197_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1838_23_lut (.I0(GND_net), .I1(n2713), 
            .I2(VCC_net), .I3(n39138), .O(n2780)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i2196_3_lut (.I0(n3225), .I1(n3292), 
            .I2(n3237), .I3(GND_net), .O(n21_adj_5450));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i2196_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2193_3_lut (.I0(n3222), .I1(n3289), 
            .I2(n3237), .I3(GND_net), .O(n27_adj_5451));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i2193_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1753 (.I0(n3224), .I1(n13_adj_5447), .I2(n3291), 
            .I3(n3237), .O(n46623));
    defparam i1_4_lut_adj_1753.LUT_INIT = 16'heefc;
    SB_LUT4 i1_4_lut_adj_1754 (.I0(n3218), .I1(n31_adj_5452), .I2(n3285), 
            .I3(n3237), .O(n46619));
    defparam i1_4_lut_adj_1754.LUT_INIT = 16'heefc;
    SB_CARRY encoder0_position_31__I_0_add_1838_23 (.CI(n39138), .I0(n2713), 
            .I1(VCC_net), .CO(n39139));
    SB_LUT4 i1_4_lut_adj_1755 (.I0(n3219), .I1(n17_adj_5448), .I2(n3286), 
            .I3(n3237), .O(n46627));
    defparam i1_4_lut_adj_1755.LUT_INIT = 16'heefc;
    SB_LUT4 encoder0_position_31__I_0_add_1838_22_lut (.I0(GND_net), .I1(n2714), 
            .I2(VCC_net), .I3(n39137), .O(n2781)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15628_3_lut (.I0(PWMLimit[2]), .I1(\data_in_frame[10] [2]), 
            .I2(n28521), .I3(GND_net), .O(n29576));   // verilog/coms.v(128[12] 303[6])
    defparam i15628_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1756 (.I0(n3228), .I1(n27_adj_5451), .I2(n3295), 
            .I3(n3237), .O(n46621));
    defparam i1_4_lut_adj_1756.LUT_INIT = 16'heefc;
    SB_CARRY encoder0_position_31__I_0_add_1838_22 (.CI(n39137), .I0(n2714), 
            .I1(VCC_net), .CO(n39138));
    SB_LUT4 i1_4_lut_adj_1757 (.I0(n3223), .I1(n19_adj_5449), .I2(n3290), 
            .I3(n3237), .O(n46617));
    defparam i1_4_lut_adj_1757.LUT_INIT = 16'heefc;
    SB_LUT4 i1_4_lut_adj_1758 (.I0(n3221), .I1(n21_adj_5450), .I2(n3288), 
            .I3(n3237), .O(n46625));
    defparam i1_4_lut_adj_1758.LUT_INIT = 16'heefc;
    SB_LUT4 i15629_3_lut (.I0(PWMLimit[1]), .I1(\data_in_frame[10] [1]), 
            .I2(n28521), .I3(GND_net), .O(n29577));   // verilog/coms.v(128[12] 303[6])
    defparam i15629_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15630_3_lut (.I0(current_limit[15]), .I1(\data_in_frame[20] [7]), 
            .I2(n28521), .I3(GND_net), .O(n29578));   // verilog/coms.v(128[12] 303[6])
    defparam i15630_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1759 (.I0(n46621), .I1(n46627), .I2(n46619), 
            .I3(n46623), .O(n46635));
    defparam i1_4_lut_adj_1759.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_31__I_0_add_1838_21_lut (.I0(GND_net), .I1(n2715), 
            .I2(VCC_net), .I3(n39136), .O(n2782)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i2188_3_lut (.I0(n3217), .I1(n3284), 
            .I2(n3237), .I3(GND_net), .O(n37));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i2188_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1760 (.I0(n37), .I1(n46635), .I2(n46625), .I3(n46617), 
            .O(n46639));
    defparam i1_4_lut_adj_1760.LUT_INIT = 16'hfffe;
    SB_LUT4 i15544_3_lut (.I0(\neo_pixel_transmitter.t0 [7]), .I1(timer[7]), 
            .I2(n42404), .I3(GND_net), .O(n29492));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15544_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1761 (.I0(n3216), .I1(n46639), .I2(n3283), .I3(n3237), 
            .O(n46641));
    defparam i1_4_lut_adj_1761.LUT_INIT = 16'heefc;
    SB_LUT4 i15631_3_lut (.I0(current_limit[14]), .I1(\data_in_frame[20] [6]), 
            .I2(n28521), .I3(GND_net), .O(n29579));   // verilog/coms.v(128[12] 303[6])
    defparam i15631_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i21334_4_lut (.I0(n544), .I1(n543), .I2(n3301), .I3(n3237), 
            .O(n35277));
    defparam i21334_4_lut.LUT_INIT = 16'heefa;
    SB_LUT4 i35411_1_lut (.I0(n1752), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n50999));
    defparam i35411_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i15632_3_lut (.I0(current_limit[13]), .I1(\data_in_frame[20] [5]), 
            .I2(n28521), .I3(GND_net), .O(n29580));   // verilog/coms.v(128[12] 303[6])
    defparam i15632_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_31__I_0_add_1838_21 (.CI(n39136), .I0(n2715), 
            .I1(VCC_net), .CO(n39137));
    SB_LUT4 encoder0_position_31__I_0_i2203_3_lut (.I0(n3232), .I1(n3299), 
            .I2(n3237), .I3(GND_net), .O(n7_adj_5446));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i2203_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16_4_lut_adj_1762 (.I0(n3231), .I1(n49339), .I2(n3237), .I3(n3230), 
            .O(n5_adj_5402));
    defparam i16_4_lut_adj_1762.LUT_INIT = 16'hac0c;
    SB_LUT4 i1_4_lut_adj_1763 (.I0(n3215), .I1(n46641), .I2(n3282), .I3(n3237), 
            .O(n46643));
    defparam i1_4_lut_adj_1763.LUT_INIT = 16'heefc;
    SB_LUT4 i21440_4_lut (.I0(n35277), .I1(n3233), .I2(n3300), .I3(n3237), 
            .O(n35388));
    defparam i21440_4_lut.LUT_INIT = 16'h88a0;
    SB_LUT4 i1_4_lut_adj_1764 (.I0(n35388), .I1(n46643), .I2(n5_adj_5402), 
            .I3(n7_adj_5446), .O(n46645));
    defparam i1_4_lut_adj_1764.LUT_INIT = 16'hfcec;
    SB_LUT4 i1_4_lut_adj_1765 (.I0(n3214), .I1(n46645), .I2(n3281), .I3(n3237), 
            .O(n46647));
    defparam i1_4_lut_adj_1765.LUT_INIT = 16'heefc;
    SB_LUT4 i1_4_lut_adj_1766 (.I0(n3213), .I1(n46647), .I2(n3280), .I3(n3237), 
            .O(n46649));
    defparam i1_4_lut_adj_1766.LUT_INIT = 16'heefc;
    SB_LUT4 i1_4_lut_adj_1767 (.I0(n3212), .I1(n46649), .I2(n3279), .I3(n3237), 
            .O(n46651));
    defparam i1_4_lut_adj_1767.LUT_INIT = 16'heefc;
    SB_LUT4 encoder0_position_31__I_0_add_1838_20_lut (.I0(GND_net), .I1(n2716), 
            .I2(VCC_net), .I3(n39135), .O(n2783)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_20_lut.LUT_INIT = 16'hC33C;
    SB_DFF dti_counter_2244__i7 (.Q(dti_counter[7]), .C(CLK_c), .D(n48));   // verilog/TinyFPGA_B.v(175[23:37])
    SB_DFF dti_counter_2244__i6 (.Q(dti_counter[6]), .C(CLK_c), .D(n49));   // verilog/TinyFPGA_B.v(175[23:37])
    SB_DFF dti_counter_2244__i5 (.Q(dti_counter[5]), .C(CLK_c), .D(n50));   // verilog/TinyFPGA_B.v(175[23:37])
    SB_DFF dti_counter_2244__i4 (.Q(dti_counter[4]), .C(CLK_c), .D(n51));   // verilog/TinyFPGA_B.v(175[23:37])
    SB_DFF dti_counter_2244__i3 (.Q(dti_counter[3]), .C(CLK_c), .D(n52));   // verilog/TinyFPGA_B.v(175[23:37])
    SB_DFF dti_counter_2244__i2 (.Q(dti_counter[2]), .C(CLK_c), .D(n53));   // verilog/TinyFPGA_B.v(175[23:37])
    SB_DFF dti_counter_2244__i1 (.Q(dti_counter[1]), .C(CLK_c), .D(n54));   // verilog/TinyFPGA_B.v(175[23:37])
    SB_LUT4 n51444_bdd_4_lut (.I0(n51444), .I1(n344), .I2(n4489), .I3(n4208), 
            .O(pwm_setpoint_23__N_11[19]));
    defparam n51444_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n10621_bdd_4_lut_35814 (.I0(n10621), .I1(current[15]), .I2(duty[18]), 
            .I3(n4208), .O(n51438));
    defparam n10621_bdd_4_lut_35814.LUT_INIT = 16'he4aa;
    SB_LUT4 n51438_bdd_4_lut (.I0(n51438), .I1(n345), .I2(n4490), .I3(n4208), 
            .O(pwm_setpoint_23__N_11[18]));
    defparam n51438_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_CARRY encoder0_position_31__I_0_add_1838_20 (.CI(n39135), .I0(n2716), 
            .I1(VCC_net), .CO(n39136));
    SB_LUT4 n10621_bdd_4_lut_35809 (.I0(n10621), .I1(current[15]), .I2(duty[17]), 
            .I3(n4208), .O(n51432));
    defparam n10621_bdd_4_lut_35809.LUT_INIT = 16'he4aa;
    SB_LUT4 n51432_bdd_4_lut (.I0(n51432), .I1(n346), .I2(n4491), .I3(n4208), 
            .O(pwm_setpoint_23__N_11[17]));
    defparam n51432_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 encoder0_position_31__I_0_add_1838_19_lut (.I0(GND_net), .I1(n2717), 
            .I2(VCC_net), .I3(n39134), .O(n2784)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1838_19 (.CI(n39134), .I0(n2717), 
            .I1(VCC_net), .CO(n39135));
    SB_LUT4 encoder0_position_31__I_0_add_1838_18_lut (.I0(GND_net), .I1(n2718), 
            .I2(VCC_net), .I3(n39133), .O(n2785)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15545_3_lut (.I0(\neo_pixel_transmitter.t0 [6]), .I1(timer[6]), 
            .I2(n42404), .I3(GND_net), .O(n29493));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15545_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_1838_18 (.CI(n39133), .I0(n2718), 
            .I1(VCC_net), .CO(n39134));
    SB_LUT4 encoder0_position_31__I_0_add_1838_17_lut (.I0(GND_net), .I1(n2719), 
            .I2(VCC_net), .I3(n39132), .O(n2786)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1768 (.I0(n3211), .I1(n46651), .I2(n3278), .I3(n3237), 
            .O(n46653));
    defparam i1_4_lut_adj_1768.LUT_INIT = 16'heefc;
    SB_CARRY encoder0_position_31__I_0_add_1838_17 (.CI(n39132), .I0(n2719), 
            .I1(VCC_net), .CO(n39133));
    SB_LUT4 encoder0_position_31__I_0_add_1838_16_lut (.I0(GND_net), .I1(n2720), 
            .I2(VCC_net), .I3(n39131), .O(n2787)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15633_3_lut (.I0(current_limit[12]), .I1(\data_in_frame[20] [4]), 
            .I2(n28521), .I3(GND_net), .O(n29581));   // verilog/coms.v(128[12] 303[6])
    defparam i15633_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1769 (.I0(n3210), .I1(n46653), .I2(n3277), .I3(n3237), 
            .O(n46655));
    defparam i1_4_lut_adj_1769.LUT_INIT = 16'heefc;
    SB_CARRY encoder0_position_31__I_0_add_1838_16 (.CI(n39131), .I0(n2720), 
            .I1(VCC_net), .CO(n39132));
    SB_LUT4 i1_4_lut_adj_1770 (.I0(n3209), .I1(n46655), .I2(n3276), .I3(n3237), 
            .O(n46657));
    defparam i1_4_lut_adj_1770.LUT_INIT = 16'heefc;
    SB_LUT4 encoder0_position_31__I_0_add_1838_15_lut (.I0(GND_net), .I1(n2721), 
            .I2(VCC_net), .I3(n39130), .O(n2788)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1771 (.I0(n3208), .I1(n46657), .I2(n3275), .I3(n3237), 
            .O(n46659));
    defparam i1_4_lut_adj_1771.LUT_INIT = 16'heefc;
    SB_CARRY encoder0_position_31__I_0_add_1838_15 (.CI(n39130), .I0(n2721), 
            .I1(VCC_net), .CO(n39131));
    SB_LUT4 i1_4_lut_adj_1772 (.I0(n3207), .I1(n46659), .I2(n3274), .I3(n3237), 
            .O(n46661));
    defparam i1_4_lut_adj_1772.LUT_INIT = 16'heefc;
    SB_LUT4 encoder0_position_31__I_0_add_1838_14_lut (.I0(GND_net), .I1(n2722), 
            .I2(VCC_net), .I3(n39129), .O(n2789)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1838_14 (.CI(n39129), .I0(n2722), 
            .I1(VCC_net), .CO(n39130));
    SB_LUT4 i1_4_lut_adj_1773 (.I0(n3206), .I1(n46661), .I2(n3273), .I3(n3237), 
            .O(n46663));
    defparam i1_4_lut_adj_1773.LUT_INIT = 16'heefc;
    SB_LUT4 i1_4_lut_adj_1774 (.I0(n3205), .I1(n46663), .I2(n3272), .I3(n3237), 
            .O(n46665));
    defparam i1_4_lut_adj_1774.LUT_INIT = 16'heefc;
    SB_LUT4 i15546_3_lut (.I0(\neo_pixel_transmitter.t0 [5]), .I1(timer[5]), 
            .I2(n42404), .I3(GND_net), .O(n29494));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15546_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15074_3_lut (.I0(\neo_pixel_transmitter.t0 [0]), .I1(timer[0]), 
            .I2(n42404), .I3(GND_net), .O(n29022));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15074_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i35574_4_lut (.I0(n46665), .I1(n3204), .I2(n3271), .I3(n3237), 
            .O(n35558));
    defparam i35574_4_lut.LUT_INIT = 16'h1105;
    SB_LUT4 encoder0_position_31__I_0_add_1838_13_lut (.I0(GND_net), .I1(n2723), 
            .I2(VCC_net), .I3(n39128), .O(n2790)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1838_13 (.CI(n39128), .I0(n2723), 
            .I1(VCC_net), .CO(n39129));
    SB_LUT4 encoder0_position_31__I_0_i2109_3_lut (.I0(n3106), .I1(n3173), 
            .I2(n3138), .I3(GND_net), .O(n3205));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i2109_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15634_3_lut (.I0(current_limit[11]), .I1(\data_in_frame[20] [3]), 
            .I2(n28521), .I3(GND_net), .O(n29582));   // verilog/coms.v(128[12] 303[6])
    defparam i15634_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_add_1838_12_lut (.I0(GND_net), .I1(n2724), 
            .I2(VCC_net), .I3(n39127), .O(n2791)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i2112_3_lut (.I0(n3109), .I1(n3176), 
            .I2(n3138), .I3(GND_net), .O(n3208));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i2112_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2110_3_lut (.I0(n3107), .I1(n3174), 
            .I2(n3138), .I3(GND_net), .O(n3206));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i2110_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_1838_12 (.CI(n39127), .I0(n2724), 
            .I1(VCC_net), .CO(n39128));
    SB_LUT4 i15635_3_lut (.I0(current_limit[10]), .I1(\data_in_frame[20] [2]), 
            .I2(n28521), .I3(GND_net), .O(n29583));   // verilog/coms.v(128[12] 303[6])
    defparam i15635_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_add_1838_11_lut (.I0(GND_net), .I1(n2725), 
            .I2(VCC_net), .I3(n39126), .O(n2792)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1838_11 (.CI(n39126), .I0(n2725), 
            .I1(VCC_net), .CO(n39127));
    SB_LUT4 i15547_3_lut (.I0(\neo_pixel_transmitter.t0 [4]), .I1(timer[4]), 
            .I2(n42404), .I3(GND_net), .O(n29495));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15547_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1838_10_lut (.I0(GND_net), .I1(n2726), 
            .I2(VCC_net), .I3(n39125), .O(n2793)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1838_10 (.CI(n39125), .I0(n2726), 
            .I1(VCC_net), .CO(n39126));
    SB_LUT4 i15636_3_lut (.I0(current_limit[9]), .I1(\data_in_frame[20] [1]), 
            .I2(n28521), .I3(GND_net), .O(n29584));   // verilog/coms.v(128[12] 303[6])
    defparam i15636_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_add_1838_9_lut (.I0(GND_net), .I1(n2727), 
            .I2(VCC_net), .I3(n39124), .O(n2794)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1838_9 (.CI(n39124), .I0(n2727), 
            .I1(VCC_net), .CO(n39125));
    SB_LUT4 encoder0_position_31__I_0_add_1838_8_lut (.I0(GND_net), .I1(n2728), 
            .I2(VCC_net), .I3(n39123), .O(n2795)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1838_8 (.CI(n39123), .I0(n2728), 
            .I1(VCC_net), .CO(n39124));
    SB_LUT4 encoder0_position_31__I_0_add_1838_7_lut (.I0(GND_net), .I1(n2729), 
            .I2(GND_net), .I3(n39122), .O(n2796)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1838_7 (.CI(n39122), .I0(n2729), 
            .I1(GND_net), .CO(n39123));
    SB_LUT4 encoder0_position_31__I_0_add_1838_6_lut (.I0(GND_net), .I1(n2730), 
            .I2(GND_net), .I3(n39121), .O(n2797)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1838_6 (.CI(n39121), .I0(n2730), 
            .I1(GND_net), .CO(n39122));
    SB_LUT4 encoder0_position_31__I_0_add_1838_5_lut (.I0(GND_net), .I1(n2731), 
            .I2(VCC_net), .I3(n39120), .O(n2798)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1838_5 (.CI(n39120), .I0(n2731), 
            .I1(VCC_net), .CO(n39121));
    SB_LUT4 encoder0_position_31__I_0_add_1838_4_lut (.I0(GND_net), .I1(n2732), 
            .I2(GND_net), .I3(n39119), .O(n2799)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1838_4 (.CI(n39119), .I0(n2732), 
            .I1(GND_net), .CO(n39120));
    SB_LUT4 encoder0_position_31__I_0_add_1838_3_lut (.I0(GND_net), .I1(n2733), 
            .I2(VCC_net), .I3(n39118), .O(n2800)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1838_3 (.CI(n39118), .I0(n2733), 
            .I1(VCC_net), .CO(n39119));
    SB_LUT4 encoder0_position_31__I_0_add_1838_2_lut (.I0(GND_net), .I1(n538), 
            .I2(GND_net), .I3(VCC_net), .O(n2801)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1838_2 (.CI(VCC_net), .I0(n538), 
            .I1(GND_net), .CO(n39118));
    SB_LUT4 encoder0_position_31__I_0_add_1771_26_lut (.I0(n50702), .I1(n2610), 
            .I2(VCC_net), .I3(n39117), .O(n2709)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_26_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_31__I_0_add_1771_25_lut (.I0(GND_net), .I1(n2611), 
            .I2(VCC_net), .I3(n39116), .O(n2678)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1771_25 (.CI(n39116), .I0(n2611), 
            .I1(VCC_net), .CO(n39117));
    SB_LUT4 encoder0_position_31__I_0_add_1771_24_lut (.I0(GND_net), .I1(n2612), 
            .I2(VCC_net), .I3(n39115), .O(n2679)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1771_24 (.CI(n39115), .I0(n2612), 
            .I1(VCC_net), .CO(n39116));
    SB_LUT4 encoder0_position_31__I_0_add_1771_23_lut (.I0(GND_net), .I1(n2613), 
            .I2(VCC_net), .I3(n39114), .O(n2680)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1771_23 (.CI(n39114), .I0(n2613), 
            .I1(VCC_net), .CO(n39115));
    SB_LUT4 encoder0_position_31__I_0_i2111_3_lut (.I0(n3108), .I1(n3175), 
            .I2(n3138), .I3(GND_net), .O(n3207));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i2111_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1771_22_lut (.I0(GND_net), .I1(n2614), 
            .I2(VCC_net), .I3(n39113), .O(n2681)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i2116_3_lut (.I0(n3113), .I1(n3180), 
            .I2(n3138), .I3(GND_net), .O(n3212));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i2116_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_1771_22 (.CI(n39113), .I0(n2614), 
            .I1(VCC_net), .CO(n39114));
    SB_LUT4 encoder0_position_31__I_0_add_1771_21_lut (.I0(GND_net), .I1(n2615), 
            .I2(VCC_net), .I3(n39112), .O(n2682)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1771_21 (.CI(n39112), .I0(n2615), 
            .I1(VCC_net), .CO(n39113));
    SB_LUT4 encoder0_position_31__I_0_add_1771_20_lut (.I0(GND_net), .I1(n2616), 
            .I2(VCC_net), .I3(n39111), .O(n2683)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1771_20 (.CI(n39111), .I0(n2616), 
            .I1(VCC_net), .CO(n39112));
    SB_LUT4 encoder0_position_31__I_0_add_1771_19_lut (.I0(GND_net), .I1(n2617), 
            .I2(VCC_net), .I3(n39110), .O(n2684)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1771_19 (.CI(n39110), .I0(n2617), 
            .I1(VCC_net), .CO(n39111));
    SB_LUT4 encoder0_position_31__I_0_add_1771_18_lut (.I0(GND_net), .I1(n2618), 
            .I2(VCC_net), .I3(n39109), .O(n2685)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1771_18 (.CI(n39109), .I0(n2618), 
            .I1(VCC_net), .CO(n39110));
    SB_LUT4 encoder0_position_31__I_0_add_1771_17_lut (.I0(GND_net), .I1(n2619), 
            .I2(VCC_net), .I3(n39108), .O(n2686)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1771_17 (.CI(n39108), .I0(n2619), 
            .I1(VCC_net), .CO(n39109));
    SB_LUT4 encoder0_position_31__I_0_i2120_3_lut (.I0(n3117), .I1(n3184), 
            .I2(n3138), .I3(GND_net), .O(n3216));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i2120_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1771_16_lut (.I0(GND_net), .I1(n2620), 
            .I2(VCC_net), .I3(n39107), .O(n2687)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1771_16 (.CI(n39107), .I0(n2620), 
            .I1(VCC_net), .CO(n39108));
    SB_LUT4 encoder0_position_31__I_0_add_1771_15_lut (.I0(GND_net), .I1(n2621), 
            .I2(VCC_net), .I3(n39106), .O(n2688)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1771_15 (.CI(n39106), .I0(n2621), 
            .I1(VCC_net), .CO(n39107));
    SB_LUT4 encoder0_position_31__I_0_add_1771_14_lut (.I0(GND_net), .I1(n2622), 
            .I2(VCC_net), .I3(n39105), .O(n2689)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1771_14 (.CI(n39105), .I0(n2622), 
            .I1(VCC_net), .CO(n39106));
    SB_LUT4 encoder0_position_31__I_0_add_1771_13_lut (.I0(GND_net), .I1(n2623), 
            .I2(VCC_net), .I3(n39104), .O(n2690)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1771_13 (.CI(n39104), .I0(n2623), 
            .I1(VCC_net), .CO(n39105));
    SB_LUT4 encoder0_position_31__I_0_add_1771_12_lut (.I0(GND_net), .I1(n2624), 
            .I2(VCC_net), .I3(n39103), .O(n2691)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1771_12 (.CI(n39103), .I0(n2624), 
            .I1(VCC_net), .CO(n39104));
    SB_LUT4 encoder0_position_31__I_0_add_1771_11_lut (.I0(GND_net), .I1(n2625), 
            .I2(VCC_net), .I3(n39102), .O(n2692)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1771_11 (.CI(n39102), .I0(n2625), 
            .I1(VCC_net), .CO(n39103));
    SB_LUT4 encoder0_position_31__I_0_add_1771_10_lut (.I0(GND_net), .I1(n2626), 
            .I2(VCC_net), .I3(n39101), .O(n2693)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1771_10 (.CI(n39101), .I0(n2626), 
            .I1(VCC_net), .CO(n39102));
    SB_LUT4 encoder0_position_31__I_0_add_1771_9_lut (.I0(GND_net), .I1(n2627), 
            .I2(VCC_net), .I3(n39100), .O(n2694)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1771_9 (.CI(n39100), .I0(n2627), 
            .I1(VCC_net), .CO(n39101));
    SB_LUT4 encoder0_position_31__I_0_add_1771_8_lut (.I0(GND_net), .I1(n2628), 
            .I2(VCC_net), .I3(n39099), .O(n2695)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1771_8 (.CI(n39099), .I0(n2628), 
            .I1(VCC_net), .CO(n39100));
    SB_LUT4 encoder0_position_31__I_0_add_1771_7_lut (.I0(GND_net), .I1(n2629), 
            .I2(GND_net), .I3(n39098), .O(n2696)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1771_7 (.CI(n39098), .I0(n2629), 
            .I1(GND_net), .CO(n39099));
    SB_LUT4 encoder0_position_31__I_0_add_1771_6_lut (.I0(GND_net), .I1(n2630), 
            .I2(GND_net), .I3(n39097), .O(n2697)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1771_6 (.CI(n39097), .I0(n2630), 
            .I1(GND_net), .CO(n39098));
    SB_LUT4 encoder0_position_31__I_0_add_1771_5_lut (.I0(GND_net), .I1(n2631), 
            .I2(VCC_net), .I3(n39096), .O(n2698)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1771_5 (.CI(n39096), .I0(n2631), 
            .I1(VCC_net), .CO(n39097));
    SB_LUT4 encoder0_position_31__I_0_add_1771_4_lut (.I0(GND_net), .I1(n2632), 
            .I2(GND_net), .I3(n39095), .O(n2699)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1771_4 (.CI(n39095), .I0(n2632), 
            .I1(GND_net), .CO(n39096));
    SB_LUT4 encoder0_position_31__I_0_add_1771_3_lut (.I0(GND_net), .I1(n2633), 
            .I2(VCC_net), .I3(n39094), .O(n2700)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1771_3 (.CI(n39094), .I0(n2633), 
            .I1(VCC_net), .CO(n39095));
    SB_LUT4 encoder0_position_31__I_0_add_1771_2_lut (.I0(GND_net), .I1(n537), 
            .I2(GND_net), .I3(VCC_net), .O(n2701)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1771_2 (.CI(VCC_net), .I0(n537), 
            .I1(GND_net), .CO(n39094));
    SB_LUT4 encoder0_position_31__I_0_add_1704_25_lut (.I0(n50754), .I1(n2511), 
            .I2(VCC_net), .I3(n39093), .O(n2610)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_25_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_31__I_0_add_1704_24_lut (.I0(GND_net), .I1(n2512), 
            .I2(VCC_net), .I3(n39092), .O(n2579)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1704_24 (.CI(n39092), .I0(n2512), 
            .I1(VCC_net), .CO(n39093));
    SB_LUT4 i15548_3_lut (.I0(\neo_pixel_transmitter.t0 [3]), .I1(timer[3]), 
            .I2(n42404), .I3(GND_net), .O(n29496));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15548_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1704_23_lut (.I0(GND_net), .I1(n2513), 
            .I2(VCC_net), .I3(n39091), .O(n2580)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1704_23 (.CI(n39091), .I0(n2513), 
            .I1(VCC_net), .CO(n39092));
    SB_LUT4 encoder0_position_31__I_0_add_1704_22_lut (.I0(GND_net), .I1(n2514), 
            .I2(VCC_net), .I3(n39090), .O(n2581)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1704_22 (.CI(n39090), .I0(n2514), 
            .I1(VCC_net), .CO(n39091));
    SB_LUT4 encoder0_position_31__I_0_add_1704_21_lut (.I0(GND_net), .I1(n2515), 
            .I2(VCC_net), .I3(n39089), .O(n2582)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1704_21 (.CI(n39089), .I0(n2515), 
            .I1(VCC_net), .CO(n39090));
    SB_LUT4 encoder0_position_31__I_0_add_1704_20_lut (.I0(GND_net), .I1(n2516), 
            .I2(VCC_net), .I3(n39088), .O(n2583)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1704_20 (.CI(n39088), .I0(n2516), 
            .I1(VCC_net), .CO(n39089));
    SB_LUT4 encoder0_position_31__I_0_add_1704_19_lut (.I0(GND_net), .I1(n2517), 
            .I2(VCC_net), .I3(n39087), .O(n2584)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1704_19 (.CI(n39087), .I0(n2517), 
            .I1(VCC_net), .CO(n39088));
    SB_LUT4 encoder0_position_31__I_0_add_1704_18_lut (.I0(GND_net), .I1(n2518), 
            .I2(VCC_net), .I3(n39086), .O(n2585)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1704_18 (.CI(n39086), .I0(n2518), 
            .I1(VCC_net), .CO(n39087));
    SB_LUT4 encoder0_position_31__I_0_add_1704_17_lut (.I0(GND_net), .I1(n2519), 
            .I2(VCC_net), .I3(n39085), .O(n2586)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1704_17 (.CI(n39085), .I0(n2519), 
            .I1(VCC_net), .CO(n39086));
    SB_LUT4 encoder0_position_31__I_0_add_1704_16_lut (.I0(GND_net), .I1(n2520), 
            .I2(VCC_net), .I3(n39084), .O(n2587)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1704_16 (.CI(n39084), .I0(n2520), 
            .I1(VCC_net), .CO(n39085));
    SB_LUT4 encoder0_position_31__I_0_add_1704_15_lut (.I0(GND_net), .I1(n2521), 
            .I2(VCC_net), .I3(n39083), .O(n2588)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1704_15 (.CI(n39083), .I0(n2521), 
            .I1(VCC_net), .CO(n39084));
    SB_LUT4 encoder0_position_31__I_0_add_1704_14_lut (.I0(GND_net), .I1(n2522), 
            .I2(VCC_net), .I3(n39082), .O(n2589)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1704_14 (.CI(n39082), .I0(n2522), 
            .I1(VCC_net), .CO(n39083));
    SB_LUT4 encoder0_position_31__I_0_add_1704_13_lut (.I0(GND_net), .I1(n2523), 
            .I2(VCC_net), .I3(n39081), .O(n2590)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1704_13 (.CI(n39081), .I0(n2523), 
            .I1(VCC_net), .CO(n39082));
    SB_LUT4 encoder0_position_31__I_0_add_1704_12_lut (.I0(GND_net), .I1(n2524), 
            .I2(VCC_net), .I3(n39080), .O(n2591)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1704_12 (.CI(n39080), .I0(n2524), 
            .I1(VCC_net), .CO(n39081));
    SB_LUT4 encoder0_position_31__I_0_add_1704_11_lut (.I0(GND_net), .I1(n2525), 
            .I2(VCC_net), .I3(n39079), .O(n2592)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1704_11 (.CI(n39079), .I0(n2525), 
            .I1(VCC_net), .CO(n39080));
    SB_LUT4 encoder0_position_31__I_0_add_1704_10_lut (.I0(GND_net), .I1(n2526), 
            .I2(VCC_net), .I3(n39078), .O(n2593)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1704_10 (.CI(n39078), .I0(n2526), 
            .I1(VCC_net), .CO(n39079));
    SB_LUT4 encoder0_position_31__I_0_add_1704_9_lut (.I0(GND_net), .I1(n2527), 
            .I2(VCC_net), .I3(n39077), .O(n2594)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1704_9 (.CI(n39077), .I0(n2527), 
            .I1(VCC_net), .CO(n39078));
    SB_LUT4 encoder0_position_31__I_0_add_1704_8_lut (.I0(GND_net), .I1(n2528), 
            .I2(VCC_net), .I3(n39076), .O(n2595)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1704_8 (.CI(n39076), .I0(n2528), 
            .I1(VCC_net), .CO(n39077));
    SB_LUT4 encoder0_position_31__I_0_i2128_3_lut (.I0(n3125), .I1(n3192), 
            .I2(n3138), .I3(GND_net), .O(n3224));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i2128_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2126_3_lut (.I0(n3123), .I1(n3190), 
            .I2(n3138), .I3(GND_net), .O(n3222));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i2126_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1704_7_lut (.I0(GND_net), .I1(n2529), 
            .I2(GND_net), .I3(n39075), .O(n2596)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15549_3_lut (.I0(\neo_pixel_transmitter.t0 [2]), .I1(timer[2]), 
            .I2(n42404), .I3(GND_net), .O(n29497));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15549_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2121_3_lut (.I0(n3118), .I1(n3185), 
            .I2(n3138), .I3(GND_net), .O(n3217));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i2121_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2134_3_lut (.I0(n3131), .I1(n3198), 
            .I2(n3138), .I3(GND_net), .O(n3230));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i2134_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2133_3_lut (.I0(n3130), .I1(n3197), 
            .I2(n3138), .I3(GND_net), .O(n3229));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i2133_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2123_3_lut (.I0(n3120), .I1(n3187), 
            .I2(n3138), .I3(GND_net), .O(n3219));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i2123_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2122_3_lut (.I0(n3119), .I1(n3186), 
            .I2(n3138), .I3(GND_net), .O(n3218));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i2122_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15550_3_lut (.I0(\neo_pixel_transmitter.t0 [1]), .I1(timer[1]), 
            .I2(n42404), .I3(GND_net), .O(n29498));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15550_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2124_3_lut (.I0(n3121), .I1(n3188), 
            .I2(n3138), .I3(GND_net), .O(n3220));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i2124_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2125_3_lut (.I0(n3122), .I1(n3189), 
            .I2(n3138), .I3(GND_net), .O(n3221));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i2125_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2129_3_lut (.I0(n3126), .I1(n3193), 
            .I2(n3138), .I3(GND_net), .O(n3225));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i2129_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2115_3_lut (.I0(n3112), .I1(n3179), 
            .I2(n3138), .I3(GND_net), .O(n3211));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i2115_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_1704_7 (.CI(n39075), .I0(n2529), 
            .I1(GND_net), .CO(n39076));
    SB_LUT4 encoder0_position_31__I_0_add_1704_6_lut (.I0(GND_net), .I1(n2530), 
            .I2(GND_net), .I3(n39074), .O(n2597)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_6_lut.LUT_INIT = 16'hC33C;
    SB_IO RX_pad (.PACKAGE_PIN(RX), .OUTPUT_ENABLE(VCC_net), .D_IN_0(RX_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam RX_pad.PIN_TYPE = 6'b000001;
    defparam RX_pad.PULLUP = 1'b0;
    defparam RX_pad.NEG_TRIGGER = 1'b0;
    defparam RX_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO ENCODER1_B_pad (.PACKAGE_PIN(ENCODER1_B), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(ENCODER1_B_N));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ENCODER1_B_pad.PIN_TYPE = 6'b000001;
    defparam ENCODER1_B_pad.PULLUP = 1'b0;
    defparam ENCODER1_B_pad.NEG_TRIGGER = 1'b0;
    defparam ENCODER1_B_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO ENCODER1_A_pad (.PACKAGE_PIN(ENCODER1_A), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(ENCODER1_A_N));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ENCODER1_A_pad.PIN_TYPE = 6'b000001;
    defparam ENCODER1_A_pad.PULLUP = 1'b0;
    defparam ENCODER1_A_pad.NEG_TRIGGER = 1'b0;
    defparam ENCODER1_A_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO ENCODER0_B_pad (.PACKAGE_PIN(ENCODER0_B), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(ENCODER0_B_N));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ENCODER0_B_pad.PIN_TYPE = 6'b000001;
    defparam ENCODER0_B_pad.PULLUP = 1'b0;
    defparam ENCODER0_B_pad.NEG_TRIGGER = 1'b0;
    defparam ENCODER0_B_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO ENCODER0_A_pad (.PACKAGE_PIN(ENCODER0_A), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(ENCODER0_A_N));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ENCODER0_A_pad.PIN_TYPE = 6'b000001;
    defparam ENCODER0_A_pad.PULLUP = 1'b0;
    defparam ENCODER0_A_pad.NEG_TRIGGER = 1'b0;
    defparam ENCODER0_A_pad.IO_STANDARD = "SB_LVCMOS";
    SB_GB_IO CLK_pad (.PACKAGE_PIN(CLK), .OUTPUT_ENABLE(VCC_net), .GLOBAL_BUFFER_OUTPUT(CLK_c));   // verilog/TinyFPGA_B.v(3[9:12])
    defparam CLK_pad.PIN_TYPE = 6'b000001;
    defparam CLK_pad.PULLUP = 1'b0;
    defparam CLK_pad.NEG_TRIGGER = 1'b0;
    defparam CLK_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO INHA_pad (.PACKAGE_PIN(INHA), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INHA_c_0));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INHA_pad.PIN_TYPE = 6'b011001;
    defparam INHA_pad.PULLUP = 1'b0;
    defparam INHA_pad.NEG_TRIGGER = 1'b0;
    defparam INHA_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO INLA_pad (.PACKAGE_PIN(INLA), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INLA_c_0));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INLA_pad.PIN_TYPE = 6'b011001;
    defparam INLA_pad.PULLUP = 1'b0;
    defparam INLA_pad.NEG_TRIGGER = 1'b0;
    defparam INLA_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO INHB_pad (.PACKAGE_PIN(INHB), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INHB_c_0));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INHB_pad.PIN_TYPE = 6'b011001;
    defparam INHB_pad.PULLUP = 1'b0;
    defparam INHB_pad.NEG_TRIGGER = 1'b0;
    defparam INHB_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO INLB_pad (.PACKAGE_PIN(INLB), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INLB_c_0));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INLB_pad.PIN_TYPE = 6'b011001;
    defparam INLB_pad.PULLUP = 1'b0;
    defparam INLB_pad.NEG_TRIGGER = 1'b0;
    defparam INLB_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO INHC_pad (.PACKAGE_PIN(INHC), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INHC_c_0));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INHC_pad.PIN_TYPE = 6'b011001;
    defparam INHC_pad.PULLUP = 1'b0;
    defparam INHC_pad.NEG_TRIGGER = 1'b0;
    defparam INHC_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO CS_CLK_pad (.PACKAGE_PIN(CS_CLK), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(CS_CLK_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam CS_CLK_pad.PIN_TYPE = 6'b011001;
    defparam CS_CLK_pad.PULLUP = 1'b0;
    defparam CS_CLK_pad.NEG_TRIGGER = 1'b0;
    defparam CS_CLK_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 encoder0_position_31__I_0_i2114_3_lut (.I0(n3111), .I1(n3178), 
            .I2(n3138), .I3(GND_net), .O(n3210));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i2114_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2113_3_lut (.I0(n3110), .I1(n3177), 
            .I2(n3138), .I3(GND_net), .O(n3209));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i2113_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2119_3_lut (.I0(n3116), .I1(n3183), 
            .I2(n3138), .I3(GND_net), .O(n3215));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i2119_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15637_3_lut (.I0(current_limit[8]), .I1(\data_in_frame[20] [0]), 
            .I2(n28521), .I3(GND_net), .O(n29585));   // verilog/coms.v(128[12] 303[6])
    defparam i15637_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15638_3_lut (.I0(current_limit[7]), .I1(\data_in_frame[21] [7]), 
            .I2(n28521), .I3(GND_net), .O(n29586));   // verilog/coms.v(128[12] 303[6])
    defparam i15638_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15639_3_lut (.I0(current_limit[6]), .I1(\data_in_frame[21] [6]), 
            .I2(n28521), .I3(GND_net), .O(n29587));   // verilog/coms.v(128[12] 303[6])
    defparam i15639_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i2118_3_lut (.I0(n3115), .I1(n3182), 
            .I2(n3138), .I3(GND_net), .O(n3214));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i2118_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2117_3_lut (.I0(n3114), .I1(n3181), 
            .I2(n3138), .I3(GND_net), .O(n3213));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i2117_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2130_3_lut (.I0(n3127), .I1(n3194), 
            .I2(n3138), .I3(GND_net), .O(n3226));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i2130_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15551_3_lut (.I0(\data_out_frame[25] [7]), .I1(neopxl_color[7]), 
            .I2(n24278), .I3(GND_net), .O(n29499));   // verilog/coms.v(128[12] 303[6])
    defparam i15551_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i2132_3_lut (.I0(n3129), .I1(n3196), 
            .I2(n3138), .I3(GND_net), .O(n3228));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i2132_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2131_3_lut (.I0(n3128), .I1(n3195), 
            .I2(n3138), .I3(GND_net), .O(n3227));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i2131_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2127_3_lut (.I0(n3124), .I1(n3191), 
            .I2(n3138), .I3(GND_net), .O(n3223));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i2127_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2137_3_lut (.I0(n542), .I1(n3201), 
            .I2(n3138), .I3(GND_net), .O(n3233));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i2137_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15640_3_lut (.I0(current_limit[5]), .I1(\data_in_frame[21] [5]), 
            .I2(n28521), .I3(GND_net), .O(n29588));   // verilog/coms.v(128[12] 303[6])
    defparam i15640_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15075_3_lut (.I0(\data_out_frame[12] [5]), .I1(setpoint[21]), 
            .I2(n24278), .I3(GND_net), .O(n29023));   // verilog/coms.v(128[12] 303[6])
    defparam i15075_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i2136_3_lut (.I0(n3133), .I1(n3200), 
            .I2(n3138), .I3(GND_net), .O(n3232));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i2136_3_lut.LUT_INIT = 16'hacac;
    SB_IO DE_pad (.PACKAGE_PIN(DE), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DE_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DE_pad.PIN_TYPE = 6'b011001;
    defparam DE_pad.PULLUP = 1'b0;
    defparam DE_pad.NEG_TRIGGER = 1'b0;
    defparam DE_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 encoder0_position_31__I_0_i2135_3_lut (.I0(n3132), .I1(n3199), 
            .I2(n3138), .I3(GND_net), .O(n3231));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i2135_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i2_3_lut (.I0(encoder0_position[1]), 
            .I1(n32), .I2(encoder0_position[31]), .I3(GND_net), .O(n543));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_mux_3_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15552_3_lut (.I0(\data_out_frame[25] [6]), .I1(neopxl_color[6]), 
            .I2(n24278), .I3(GND_net), .O(n29500));   // verilog/coms.v(128[12] 303[6])
    defparam i15552_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15641_3_lut (.I0(current_limit[4]), .I1(\data_in_frame[21] [4]), 
            .I2(n28521), .I3(GND_net), .O(n29589));   // verilog/coms.v(128[12] 303[6])
    defparam i15641_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_236_8_lut (.I0(GND_net), .I1(encoder1_position[9]), .I2(GND_net), 
            .I3(n38482), .O(encoder1_position_scaled_23__N_75[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_236_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 n10621_bdd_4_lut_35804 (.I0(n10621), .I1(current[15]), .I2(duty[16]), 
            .I3(n4208), .O(n51426));
    defparam n10621_bdd_4_lut_35804.LUT_INIT = 16'he4aa;
    SB_LUT4 n51426_bdd_4_lut (.I0(n51426), .I1(n347), .I2(n4492), .I3(n4208), 
            .O(pwm_setpoint_23__N_11[16]));
    defparam n51426_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n10621_bdd_4_lut_35799 (.I0(n10621), .I1(current[15]), .I2(duty[15]), 
            .I3(n4208), .O(n51420));
    defparam n10621_bdd_4_lut_35799.LUT_INIT = 16'he4aa;
    SB_LUT4 n51420_bdd_4_lut (.I0(n51420), .I1(n348), .I2(n4493), .I3(n4208), 
            .O(pwm_setpoint_23__N_11[15]));
    defparam n51420_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n10621_bdd_4_lut_35794 (.I0(n10621), .I1(current[15]), .I2(duty[14]), 
            .I3(n4208), .O(n51414));
    defparam n10621_bdd_4_lut_35794.LUT_INIT = 16'he4aa;
    SB_LUT4 n51414_bdd_4_lut (.I0(n51414), .I1(n349), .I2(n4494), .I3(n4208), 
            .O(pwm_setpoint_23__N_11[14]));
    defparam n51414_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n10621_bdd_4_lut_35789 (.I0(n10621), .I1(current[15]), .I2(duty[13]), 
            .I3(n4208), .O(n51408));
    defparam n10621_bdd_4_lut_35789.LUT_INIT = 16'he4aa;
    SB_LUT4 n51408_bdd_4_lut (.I0(n51408), .I1(n350), .I2(n4495), .I3(n4208), 
            .O(pwm_setpoint_23__N_11[13]));
    defparam n51408_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n10621_bdd_4_lut_35784 (.I0(n10621), .I1(current[15]), .I2(duty[12]), 
            .I3(n4208), .O(n51402));
    defparam n10621_bdd_4_lut_35784.LUT_INIT = 16'he4aa;
    SB_LUT4 n51402_bdd_4_lut (.I0(n51402), .I1(n351), .I2(n4496), .I3(n4208), 
            .O(pwm_setpoint_23__N_11[12]));
    defparam n51402_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n10621_bdd_4_lut_35779 (.I0(n10621), .I1(current[11]), .I2(duty[11]), 
            .I3(n4208), .O(n51396));
    defparam n10621_bdd_4_lut_35779.LUT_INIT = 16'he4aa;
    SB_LUT4 n51396_bdd_4_lut (.I0(n51396), .I1(n352), .I2(n4497), .I3(n4208), 
            .O(pwm_setpoint_23__N_11[11]));
    defparam n51396_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n10621_bdd_4_lut_35774 (.I0(n10621), .I1(current[10]), .I2(duty[10]), 
            .I3(n4208), .O(n51390));
    defparam n10621_bdd_4_lut_35774.LUT_INIT = 16'he4aa;
    SB_LUT4 n51390_bdd_4_lut (.I0(n51390), .I1(n353), .I2(n4498), .I3(n4208), 
            .O(pwm_setpoint_23__N_11[10]));
    defparam n51390_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n10621_bdd_4_lut_35769 (.I0(n10621), .I1(current[9]), .I2(duty[9]), 
            .I3(n4208), .O(n51384));
    defparam n10621_bdd_4_lut_35769.LUT_INIT = 16'he4aa;
    SB_LUT4 n51384_bdd_4_lut (.I0(n51384), .I1(n354), .I2(n4499), .I3(n4208), 
            .O(pwm_setpoint_23__N_11[9]));
    defparam n51384_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_CARRY encoder0_position_31__I_0_add_1704_6 (.CI(n39074), .I0(n2530), 
            .I1(GND_net), .CO(n39075));
    SB_LUT4 encoder0_position_31__I_0_add_1704_5_lut (.I0(GND_net), .I1(n2531), 
            .I2(VCC_net), .I3(n39073), .O(n2598)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15076_3_lut (.I0(\data_out_frame[12] [4]), .I1(setpoint[20]), 
            .I2(n24278), .I3(GND_net), .O(n29024));   // verilog/coms.v(128[12] 303[6])
    defparam i15076_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_31__I_0_add_1704_5 (.CI(n39073), .I0(n2531), 
            .I1(VCC_net), .CO(n39074));
    SB_LUT4 encoder0_position_31__I_0_add_1704_4_lut (.I0(GND_net), .I1(n2532), 
            .I2(GND_net), .I3(n39072), .O(n2599)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1704_4 (.CI(n39072), .I0(n2532), 
            .I1(GND_net), .CO(n39073));
    SB_LUT4 encoder0_position_31__I_0_add_1704_3_lut (.I0(GND_net), .I1(n2533), 
            .I2(VCC_net), .I3(n39071), .O(n2600)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1704_3 (.CI(n39071), .I0(n2533), 
            .I1(VCC_net), .CO(n39072));
    SB_LUT4 encoder0_position_31__I_0_add_1704_2_lut (.I0(GND_net), .I1(n950), 
            .I2(GND_net), .I3(VCC_net), .O(n2601)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1704_2 (.CI(VCC_net), .I0(n950), 
            .I1(GND_net), .CO(n39071));
    SB_LUT4 mux_1005_i12_3_lut (.I0(duty[11]), .I1(n352), .I2(duty[23]), 
            .I3(GND_net), .O(n4712));   // verilog/TinyFPGA_B.v(118[13] 129[7])
    defparam mux_1005_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i35604_1_lut (.I0(n3237), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n51192));
    defparam i35604_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_add_1637_24_lut (.I0(n50784), .I1(n2412), 
            .I2(VCC_net), .I3(n39070), .O(n2511)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1637_24_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_31__I_0_add_1637_23_lut (.I0(GND_net), .I1(n2413), 
            .I2(VCC_net), .I3(n39069), .O(n2480)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1637_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1637_23 (.CI(n39069), .I0(n2413), 
            .I1(VCC_net), .CO(n39070));
    SB_LUT4 encoder0_position_31__I_0_add_1637_22_lut (.I0(GND_net), .I1(n2414), 
            .I2(VCC_net), .I3(n39068), .O(n2481)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1637_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1637_22 (.CI(n39068), .I0(n2414), 
            .I1(VCC_net), .CO(n39069));
    SB_LUT4 encoder0_position_31__I_0_add_1637_21_lut (.I0(GND_net), .I1(n2415), 
            .I2(VCC_net), .I3(n39067), .O(n2482)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1637_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1637_21 (.CI(n39067), .I0(n2415), 
            .I1(VCC_net), .CO(n39068));
    SB_LUT4 i15553_3_lut (.I0(\data_out_frame[25] [5]), .I1(neopxl_color[5]), 
            .I2(n24278), .I3(GND_net), .O(n29501));   // verilog/coms.v(128[12] 303[6])
    defparam i15553_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15642_3_lut (.I0(current_limit[3]), .I1(\data_in_frame[21] [3]), 
            .I2(n28521), .I3(GND_net), .O(n29590));   // verilog/coms.v(128[12] 303[6])
    defparam i15642_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15643_3_lut (.I0(current_limit[2]), .I1(\data_in_frame[21] [2]), 
            .I2(n28521), .I3(GND_net), .O(n29591));   // verilog/coms.v(128[12] 303[6])
    defparam i15643_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_add_1637_20_lut (.I0(GND_net), .I1(n2416), 
            .I2(VCC_net), .I3(n39066), .O(n2483)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1637_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1637_20 (.CI(n39066), .I0(n2416), 
            .I1(VCC_net), .CO(n39067));
    SB_LUT4 i15644_3_lut (.I0(current_limit[1]), .I1(\data_in_frame[21] [1]), 
            .I2(n28521), .I3(GND_net), .O(n29592));   // verilog/coms.v(128[12] 303[6])
    defparam i15644_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15645_3_lut (.I0(control_mode[7]), .I1(\data_in_frame[1] [7]), 
            .I2(n28521), .I3(GND_net), .O(n29593));   // verilog/coms.v(128[12] 303[6])
    defparam i15645_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_add_1637_19_lut (.I0(GND_net), .I1(n2417), 
            .I2(VCC_net), .I3(n39065), .O(n2484)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1637_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i21501_4_lut (.I0(n543), .I1(n3231), .I2(n3232), .I3(n3233), 
            .O(n35450));
    defparam i21501_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 i15646_3_lut (.I0(control_mode[6]), .I1(\data_in_frame[1] [6]), 
            .I2(n28521), .I3(GND_net), .O(n29594));   // verilog/coms.v(128[12] 303[6])
    defparam i15646_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_31__I_0_add_1637_19 (.CI(n39065), .I0(n2417), 
            .I1(VCC_net), .CO(n39066));
    SB_LUT4 encoder0_position_31__I_0_add_1637_18_lut (.I0(GND_net), .I1(n2418), 
            .I2(VCC_net), .I3(n39064), .O(n2485)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1637_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1637_18 (.CI(n39064), .I0(n2418), 
            .I1(VCC_net), .CO(n39065));
    SB_LUT4 i1_3_lut_adj_1775 (.I0(n3225), .I1(n3221), .I2(n3220), .I3(GND_net), 
            .O(n47157));
    defparam i1_3_lut_adj_1775.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_2_lut_adj_1776 (.I0(n3218), .I1(n3219), .I2(GND_net), .I3(GND_net), 
            .O(n47201));
    defparam i1_2_lut_adj_1776.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_1777 (.I0(n3229), .I1(n47157), .I2(n35450), .I3(n3230), 
            .O(n47159));
    defparam i1_4_lut_adj_1777.LUT_INIT = 16'heccc;
    SB_LUT4 encoder0_position_31__I_0_add_1637_17_lut (.I0(GND_net), .I1(n2419), 
            .I2(VCC_net), .I3(n39063), .O(n2486)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1637_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15554_4_lut (.I0(r_Rx_Data), .I1(rx_data[3]), .I2(n4_adj_5245), 
            .I3(n27126), .O(n29502));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i15554_4_lut.LUT_INIT = 16'hccca;
    SB_CARRY encoder0_position_31__I_0_add_1637_17 (.CI(n39063), .I0(n2419), 
            .I1(VCC_net), .CO(n39064));
    SB_LUT4 encoder0_position_31__I_0_add_1637_16_lut (.I0(GND_net), .I1(n2420), 
            .I2(VCC_net), .I3(n39062), .O(n2487)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1637_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1778 (.I0(n3223), .I1(n3227), .I2(n3228), .I3(n3226), 
            .O(n47173));
    defparam i1_4_lut_adj_1778.LUT_INIT = 16'hfffe;
    SB_LUT4 i15210_3_lut (.I0(IntegralLimit[1]), .I1(\data_in_frame[13] [1]), 
            .I2(n28521), .I3(GND_net), .O(n29158));   // verilog/coms.v(128[12] 303[6])
    defparam i15210_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15555_3_lut (.I0(\data_out_frame[25] [4]), .I1(neopxl_color[4]), 
            .I2(n24278), .I3(GND_net), .O(n29503));   // verilog/coms.v(128[12] 303[6])
    defparam i15555_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_31__I_0_add_1637_16 (.CI(n39062), .I0(n2420), 
            .I1(VCC_net), .CO(n39063));
    SB_LUT4 encoder0_position_31__I_0_add_1637_15_lut (.I0(GND_net), .I1(n2421), 
            .I2(VCC_net), .I3(n39061), .O(n2488)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1637_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1637_15 (.CI(n39061), .I0(n2421), 
            .I1(VCC_net), .CO(n39062));
    SB_LUT4 encoder0_position_31__I_0_add_1637_14_lut (.I0(GND_net), .I1(n2422), 
            .I2(VCC_net), .I3(n39060), .O(n2489)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1637_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1637_14 (.CI(n39060), .I0(n2422), 
            .I1(VCC_net), .CO(n39061));
    SB_LUT4 i15556_3_lut (.I0(\data_out_frame[25] [3]), .I1(neopxl_color[3]), 
            .I2(n24278), .I3(GND_net), .O(n29504));   // verilog/coms.v(128[12] 303[6])
    defparam i15556_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1779 (.I0(n3217), .I1(n47173), .I2(n3222), .I3(n3224), 
            .O(n47177));
    defparam i1_4_lut_adj_1779.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_31__I_0_add_1637_13_lut (.I0(GND_net), .I1(n2423), 
            .I2(VCC_net), .I3(n39059), .O(n2490)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1637_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1637_13 (.CI(n39059), .I0(n2423), 
            .I1(VCC_net), .CO(n39060));
    SB_LUT4 encoder0_position_31__I_0_add_1637_12_lut (.I0(GND_net), .I1(n2424), 
            .I2(VCC_net), .I3(n39058), .O(n2491)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1637_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1637_12 (.CI(n39058), .I0(n2424), 
            .I1(VCC_net), .CO(n39059));
    SB_LUT4 i20718_2_lut (.I0(n24462), .I1(dti), .I2(GND_net), .I3(GND_net), 
            .O(n34648));
    defparam i20718_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 encoder0_position_31__I_0_add_1637_11_lut (.I0(GND_net), .I1(n2425), 
            .I2(VCC_net), .I3(n39057), .O(n2492)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1637_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1637_11 (.CI(n39057), .I0(n2425), 
            .I1(VCC_net), .CO(n39058));
    SB_LUT4 encoder0_position_31__I_0_add_1637_10_lut (.I0(GND_net), .I1(n2426), 
            .I2(VCC_net), .I3(n39056), .O(n2493)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1637_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1637_10 (.CI(n39056), .I0(n2426), 
            .I1(VCC_net), .CO(n39057));
    SB_LUT4 encoder0_position_31__I_0_add_1637_9_lut (.I0(GND_net), .I1(n2427), 
            .I2(VCC_net), .I3(n39055), .O(n2494)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1637_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1637_9 (.CI(n39055), .I0(n2427), 
            .I1(VCC_net), .CO(n39056));
    SB_LUT4 encoder0_position_31__I_0_add_1637_8_lut (.I0(GND_net), .I1(n2428), 
            .I2(VCC_net), .I3(n39054), .O(n2495)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1637_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1637_8 (.CI(n39054), .I0(n2428), 
            .I1(VCC_net), .CO(n39055));
    SB_LUT4 encoder0_position_31__I_0_add_1637_7_lut (.I0(GND_net), .I1(n2429), 
            .I2(GND_net), .I3(n39053), .O(n2496)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1637_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1780 (.I0(n3213), .I1(n3214), .I2(n3215), .I3(n47177), 
            .O(n47183));
    defparam i1_4_lut_adj_1780.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1781 (.I0(n3209), .I1(n3210), .I2(n3211), .I3(n47183), 
            .O(n47189));
    defparam i1_4_lut_adj_1781.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1782 (.I0(n3216), .I1(n47159), .I2(n3212), .I3(n47201), 
            .O(n47161));
    defparam i1_4_lut_adj_1782.LUT_INIT = 16'hfffe;
    SB_CARRY encoder0_position_31__I_0_add_1637_7 (.CI(n39053), .I0(n2429), 
            .I1(GND_net), .CO(n39054));
    SB_LUT4 encoder0_position_31__I_0_add_1637_6_lut (.I0(GND_net), .I1(n2430), 
            .I2(GND_net), .I3(n39052), .O(n2497)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1637_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1637_6 (.CI(n39052), .I0(n2430), 
            .I1(GND_net), .CO(n39053));
    SB_LUT4 encoder0_position_31__I_0_add_1637_5_lut (.I0(GND_net), .I1(n2431), 
            .I2(VCC_net), .I3(n39051), .O(n2498)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1637_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1637_5 (.CI(n39051), .I0(n2431), 
            .I1(VCC_net), .CO(n39052));
    SB_LUT4 encoder0_position_31__I_0_add_1637_4_lut (.I0(GND_net), .I1(n2432), 
            .I2(GND_net), .I3(n39050), .O(n2499)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1637_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1637_4 (.CI(n39050), .I0(n2432), 
            .I1(GND_net), .CO(n39051));
    SB_LUT4 encoder0_position_31__I_0_add_1637_3_lut (.I0(GND_net), .I1(n2433), 
            .I2(VCC_net), .I3(n39049), .O(n2500)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1637_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1637_3 (.CI(n39049), .I0(n2433), 
            .I1(VCC_net), .CO(n39050));
    SB_LUT4 encoder0_position_31__I_0_add_1637_2_lut (.I0(GND_net), .I1(n535), 
            .I2(GND_net), .I3(VCC_net), .O(n2501)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1637_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1637_2 (.CI(VCC_net), .I0(n535), 
            .I1(GND_net), .CO(n39049));
    SB_LUT4 encoder0_position_31__I_0_add_1570_23_lut (.I0(n50865), .I1(n2313), 
            .I2(VCC_net), .I3(n39048), .O(n2412)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1570_23_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_4_lut_adj_1783 (.I0(n3207), .I1(n3206), .I2(n3208), .I3(n47189), 
            .O(n46128));
    defparam i1_4_lut_adj_1783.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_31__I_0_add_1570_22_lut (.I0(GND_net), .I1(n2314), 
            .I2(VCC_net), .I3(n39047), .O(n2381)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1570_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 n10621_bdd_4_lut_35764 (.I0(n10621), .I1(current[8]), .I2(duty[8]), 
            .I3(n4208), .O(n51378));
    defparam n10621_bdd_4_lut_35764.LUT_INIT = 16'he4aa;
    SB_CARRY encoder0_position_31__I_0_add_1570_22 (.CI(n39047), .I0(n2314), 
            .I1(VCC_net), .CO(n39048));
    SB_LUT4 encoder0_position_31__I_0_add_1570_21_lut (.I0(GND_net), .I1(n2315), 
            .I2(VCC_net), .I3(n39046), .O(n2382)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1570_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 n51378_bdd_4_lut (.I0(n51378), .I1(n355), .I2(n4500), .I3(n4208), 
            .O(pwm_setpoint_23__N_11[8]));
    defparam n51378_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_CARRY encoder0_position_31__I_0_add_1570_21 (.CI(n39046), .I0(n2315), 
            .I1(VCC_net), .CO(n39047));
    SB_LUT4 encoder0_position_31__I_0_add_1570_20_lut (.I0(GND_net), .I1(n2316), 
            .I2(VCC_net), .I3(n39045), .O(n2383)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1570_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1570_20 (.CI(n39045), .I0(n2316), 
            .I1(VCC_net), .CO(n39046));
    SB_LUT4 encoder0_position_31__I_0_add_1570_19_lut (.I0(GND_net), .I1(n2317), 
            .I2(VCC_net), .I3(n39044), .O(n2384)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1570_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1570_19 (.CI(n39044), .I0(n2317), 
            .I1(VCC_net), .CO(n39045));
    SB_LUT4 encoder0_position_31__I_0_add_1570_18_lut (.I0(GND_net), .I1(n2318), 
            .I2(VCC_net), .I3(n39043), .O(n2385)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1570_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1570_18 (.CI(n39043), .I0(n2318), 
            .I1(VCC_net), .CO(n39044));
    SB_LUT4 add_157_12_lut (.I0(GND_net), .I1(delay_counter[10]), .I2(GND_net), 
            .I3(n38455), .O(n1318)) /* synthesis syn_instantiated=1 */ ;
    defparam add_157_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1570_17_lut (.I0(GND_net), .I1(n2319), 
            .I2(VCC_net), .I3(n39042), .O(n2386)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1570_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1570_17 (.CI(n39042), .I0(n2319), 
            .I1(VCC_net), .CO(n39043));
    SB_LUT4 i35608_4_lut (.I0(n3205), .I1(n46128), .I2(n3204), .I3(n47161), 
            .O(n3237));
    defparam i35608_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_31__I_0_i2043_3_lut (.I0(n3008), .I1(n3075), 
            .I2(n3039), .I3(GND_net), .O(n3107));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i2043_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15557_3_lut (.I0(\data_out_frame[25] [2]), .I1(neopxl_color[2]), 
            .I2(n24278), .I3(GND_net), .O(n29505));   // verilog/coms.v(128[12] 303[6])
    defparam i15557_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_add_1570_16_lut (.I0(GND_net), .I1(n2320), 
            .I2(VCC_net), .I3(n39041), .O(n2387)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1570_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1570_16 (.CI(n39041), .I0(n2320), 
            .I1(VCC_net), .CO(n39042));
    SB_LUT4 encoder0_position_31__I_0_add_1570_15_lut (.I0(GND_net), .I1(n2321), 
            .I2(VCC_net), .I3(n39040), .O(n2388)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1570_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1570_15 (.CI(n39040), .I0(n2321), 
            .I1(VCC_net), .CO(n39041));
    SB_LUT4 encoder0_position_31__I_0_add_1570_14_lut (.I0(GND_net), .I1(n2322), 
            .I2(VCC_net), .I3(n39039), .O(n2389)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1570_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1570_14 (.CI(n39039), .I0(n2322), 
            .I1(VCC_net), .CO(n39040));
    SB_LUT4 encoder0_position_31__I_0_add_1570_13_lut (.I0(GND_net), .I1(n2323), 
            .I2(VCC_net), .I3(n39038), .O(n2390)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1570_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1570_13 (.CI(n39038), .I0(n2323), 
            .I1(VCC_net), .CO(n39039));
    SB_LUT4 encoder0_position_31__I_0_add_1570_12_lut (.I0(GND_net), .I1(n2324), 
            .I2(VCC_net), .I3(n39037), .O(n2391)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1570_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1570_12 (.CI(n39037), .I0(n2324), 
            .I1(VCC_net), .CO(n39038));
    SB_LUT4 encoder0_position_31__I_0_add_1570_11_lut (.I0(GND_net), .I1(n2325), 
            .I2(VCC_net), .I3(n39036), .O(n2392)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1570_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_19_inv_0_i3_1_lut (.I0(duty[2]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_5268));   // verilog/TinyFPGA_B.v(123[25:30])
    defparam unary_minus_19_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_31__I_0_add_1570_11 (.CI(n39036), .I0(n2325), 
            .I1(VCC_net), .CO(n39037));
    SB_LUT4 encoder0_position_31__I_0_add_1570_10_lut (.I0(GND_net), .I1(n2326), 
            .I2(VCC_net), .I3(n39035), .O(n2393)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1570_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1570_10 (.CI(n39035), .I0(n2326), 
            .I1(VCC_net), .CO(n39036));
    SB_LUT4 encoder0_position_31__I_0_add_1570_9_lut (.I0(GND_net), .I1(n2327), 
            .I2(VCC_net), .I3(n39034), .O(n2394)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1570_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_236_3 (.CI(n38477), .I0(encoder1_position[4]), .I1(GND_net), 
            .CO(n38478));
    SB_CARRY encoder0_position_31__I_0_add_1570_9 (.CI(n39034), .I0(n2327), 
            .I1(VCC_net), .CO(n39035));
    SB_CARRY add_157_12 (.CI(n38455), .I0(delay_counter[10]), .I1(GND_net), 
            .CO(n38456));
    SB_LUT4 encoder0_position_31__I_0_add_1570_8_lut (.I0(GND_net), .I1(n2328), 
            .I2(VCC_net), .I3(n39033), .O(n2395)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1570_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_236_2_lut (.I0(GND_net), .I1(encoder1_position[3]), .I2(encoder1_position_scaled_23__N_303), 
            .I3(GND_net), .O(encoder1_position_scaled_23__N_75[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_236_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1570_8 (.CI(n39033), .I0(n2328), 
            .I1(VCC_net), .CO(n39034));
    SB_LUT4 encoder0_position_31__I_0_i2042_3_lut (.I0(n3007), .I1(n3074), 
            .I2(n3039), .I3(GND_net), .O(n3106));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i2042_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2046_3_lut (.I0(n3011), .I1(n3078), 
            .I2(n3039), .I3(GND_net), .O(n3110));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i2046_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2045_3_lut (.I0(n3010), .I1(n3077), 
            .I2(n3039), .I3(GND_net), .O(n3109));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i2045_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1570_7_lut (.I0(GND_net), .I1(n2329), 
            .I2(GND_net), .I3(n39032), .O(n2396)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1570_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1570_7 (.CI(n39032), .I0(n2329), 
            .I1(GND_net), .CO(n39033));
    SB_LUT4 encoder0_position_31__I_0_add_1570_6_lut (.I0(GND_net), .I1(n2330), 
            .I2(GND_net), .I3(n39031), .O(n2397)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1570_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1570_6 (.CI(n39031), .I0(n2330), 
            .I1(GND_net), .CO(n39032));
    SB_LUT4 encoder0_position_31__I_0_add_1570_5_lut (.I0(GND_net), .I1(n2331), 
            .I2(VCC_net), .I3(n39030), .O(n2398)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1570_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i2044_3_lut (.I0(n3009), .I1(n3076), 
            .I2(n3039), .I3(GND_net), .O(n3108));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i2044_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_1570_5 (.CI(n39030), .I0(n2331), 
            .I1(VCC_net), .CO(n39031));
    SB_LUT4 encoder0_position_31__I_0_add_1570_4_lut (.I0(GND_net), .I1(n2332), 
            .I2(GND_net), .I3(n39029), .O(n2399)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1570_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1570_4 (.CI(n39029), .I0(n2332), 
            .I1(GND_net), .CO(n39030));
    SB_LUT4 encoder0_position_31__I_0_add_1570_3_lut (.I0(GND_net), .I1(n2333), 
            .I2(VCC_net), .I3(n39028), .O(n2400)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1570_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1570_3 (.CI(n39028), .I0(n2333), 
            .I1(VCC_net), .CO(n39029));
    SB_LUT4 encoder0_position_31__I_0_add_1570_2_lut (.I0(GND_net), .I1(n534), 
            .I2(GND_net), .I3(VCC_net), .O(n2401)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1570_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1570_2 (.CI(VCC_net), .I0(n534), 
            .I1(GND_net), .CO(n39028));
    SB_LUT4 encoder0_position_31__I_0_add_1503_22_lut (.I0(GND_net), .I1(n2214), 
            .I2(VCC_net), .I3(n39027), .O(n2281)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1503_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15558_3_lut (.I0(\data_out_frame[25] [1]), .I1(neopxl_color[1]), 
            .I2(n24278), .I3(GND_net), .O(n29506));   // verilog/coms.v(128[12] 303[6])
    defparam i15558_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_add_1503_21_lut (.I0(GND_net), .I1(n2215), 
            .I2(VCC_net), .I3(n39026), .O(n2282)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1503_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1503_21 (.CI(n39026), .I0(n2215), 
            .I1(VCC_net), .CO(n39027));
    SB_LUT4 encoder0_position_31__I_0_add_1503_20_lut (.I0(GND_net), .I1(n2216), 
            .I2(VCC_net), .I3(n39025), .O(n2283)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1503_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1503_20 (.CI(n39025), .I0(n2216), 
            .I1(VCC_net), .CO(n39026));
    SB_LUT4 encoder0_position_31__I_0_add_1503_19_lut (.I0(GND_net), .I1(n2217), 
            .I2(VCC_net), .I3(n39024), .O(n2284)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1503_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1503_19 (.CI(n39024), .I0(n2217), 
            .I1(VCC_net), .CO(n39025));
    SB_LUT4 encoder0_position_31__I_0_add_1503_18_lut (.I0(GND_net), .I1(n2218), 
            .I2(VCC_net), .I3(n39023), .O(n2285)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1503_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1503_18 (.CI(n39023), .I0(n2218), 
            .I1(VCC_net), .CO(n39024));
    SB_LUT4 encoder0_position_31__I_0_add_1503_17_lut (.I0(GND_net), .I1(n2219), 
            .I2(VCC_net), .I3(n39022), .O(n2286)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1503_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15077_3_lut (.I0(h3), .I1(reg_B[0]), .I2(n46440), .I3(GND_net), 
            .O(n29025));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    defparam i15077_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_1503_17 (.CI(n39022), .I0(n2219), 
            .I1(VCC_net), .CO(n39023));
    SB_LUT4 encoder0_position_31__I_0_add_1503_16_lut (.I0(GND_net), .I1(n2220), 
            .I2(VCC_net), .I3(n39021), .O(n2287)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1503_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1503_16 (.CI(n39021), .I0(n2220), 
            .I1(VCC_net), .CO(n39022));
    SB_LUT4 encoder0_position_31__I_0_add_1503_15_lut (.I0(GND_net), .I1(n2221), 
            .I2(VCC_net), .I3(n39020), .O(n2288)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1503_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1503_15 (.CI(n39020), .I0(n2221), 
            .I1(VCC_net), .CO(n39021));
    SB_LUT4 encoder0_position_31__I_0_add_1503_14_lut (.I0(GND_net), .I1(n2222), 
            .I2(VCC_net), .I3(n39019), .O(n2289)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1503_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1503_14 (.CI(n39019), .I0(n2222), 
            .I1(VCC_net), .CO(n39020));
    SB_LUT4 encoder0_position_31__I_0_add_1503_13_lut (.I0(GND_net), .I1(n2223), 
            .I2(VCC_net), .I3(n39018), .O(n2290)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1503_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1503_13 (.CI(n39018), .I0(n2223), 
            .I1(VCC_net), .CO(n39019));
    SB_CARRY add_236_2 (.CI(GND_net), .I0(encoder1_position[3]), .I1(encoder1_position_scaled_23__N_303), 
            .CO(n38477));
    SB_LUT4 encoder0_position_31__I_0_i2067_3_lut (.I0(n3032), .I1(n3099), 
            .I2(n3039), .I3(GND_net), .O(n3131));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i2067_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1503_12_lut (.I0(GND_net), .I1(n2224), 
            .I2(VCC_net), .I3(n39017), .O(n2291)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1503_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1503_12 (.CI(n39017), .I0(n2224), 
            .I1(VCC_net), .CO(n39018));
    SB_LUT4 encoder0_position_31__I_0_add_1503_11_lut (.I0(GND_net), .I1(n2225), 
            .I2(VCC_net), .I3(n39016), .O(n2292)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1503_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1503_11 (.CI(n39016), .I0(n2225), 
            .I1(VCC_net), .CO(n39017));
    SB_LUT4 encoder0_position_31__I_0_add_1503_10_lut (.I0(GND_net), .I1(n2226), 
            .I2(VCC_net), .I3(n39015), .O(n2293)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1503_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1503_10 (.CI(n39015), .I0(n2226), 
            .I1(VCC_net), .CO(n39016));
    SB_LUT4 encoder0_position_31__I_0_add_1503_9_lut (.I0(GND_net), .I1(n2227), 
            .I2(VCC_net), .I3(n39014), .O(n2294)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1503_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1503_9 (.CI(n39014), .I0(n2227), 
            .I1(VCC_net), .CO(n39015));
    SB_LUT4 encoder0_position_31__I_0_add_1503_8_lut (.I0(GND_net), .I1(n2228), 
            .I2(VCC_net), .I3(n39013), .O(n2295)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1503_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1503_8 (.CI(n39013), .I0(n2228), 
            .I1(VCC_net), .CO(n39014));
    SB_LUT4 encoder0_position_31__I_0_add_1503_7_lut (.I0(GND_net), .I1(n2229), 
            .I2(GND_net), .I3(n39012), .O(n2296)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1503_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1503_7 (.CI(n39012), .I0(n2229), 
            .I1(GND_net), .CO(n39013));
    SB_LUT4 encoder0_position_31__I_0_add_1503_6_lut (.I0(GND_net), .I1(n2230), 
            .I2(GND_net), .I3(n39011), .O(n2297)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1503_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1503_6 (.CI(n39011), .I0(n2230), 
            .I1(GND_net), .CO(n39012));
    SB_LUT4 encoder0_position_31__I_0_add_1503_5_lut (.I0(GND_net), .I1(n2231), 
            .I2(VCC_net), .I3(n39010), .O(n2298)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1503_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1503_5 (.CI(n39010), .I0(n2231), 
            .I1(VCC_net), .CO(n39011));
    SB_LUT4 encoder0_position_31__I_0_add_1503_4_lut (.I0(GND_net), .I1(n2232), 
            .I2(GND_net), .I3(n39009), .O(n2299)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1503_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1503_4 (.CI(n39009), .I0(n2232), 
            .I1(GND_net), .CO(n39010));
    SB_LUT4 encoder0_position_31__I_0_add_1503_3_lut (.I0(GND_net), .I1(n2233), 
            .I2(VCC_net), .I3(n39008), .O(n2300)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1503_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_157_5 (.CI(n38448), .I0(delay_counter[3]), .I1(GND_net), 
            .CO(n38449));
    SB_CARRY encoder0_position_31__I_0_add_1503_3 (.CI(n39008), .I0(n2233), 
            .I1(VCC_net), .CO(n39009));
    SB_LUT4 encoder0_position_31__I_0_add_1503_2_lut (.I0(GND_net), .I1(n533), 
            .I2(GND_net), .I3(VCC_net), .O(n2301)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1503_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1503_2 (.CI(VCC_net), .I0(n533), 
            .I1(GND_net), .CO(n39008));
    SB_LUT4 encoder0_position_31__I_0_add_1436_21_lut (.I0(n50914), .I1(n2115), 
            .I2(VCC_net), .I3(n39007), .O(n2214)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1436_21_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_31__I_0_add_1436_20_lut (.I0(GND_net), .I1(n2116), 
            .I2(VCC_net), .I3(n39006), .O(n2183)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1436_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1436_20 (.CI(n39006), .I0(n2116), 
            .I1(VCC_net), .CO(n39007));
    SB_LUT4 encoder0_position_31__I_0_add_1436_19_lut (.I0(GND_net), .I1(n2117), 
            .I2(VCC_net), .I3(n39005), .O(n2184)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1436_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1436_19 (.CI(n39005), .I0(n2117), 
            .I1(VCC_net), .CO(n39006));
    SB_LUT4 encoder0_position_31__I_0_add_1436_18_lut (.I0(GND_net), .I1(n2118), 
            .I2(VCC_net), .I3(n39004), .O(n2185)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1436_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1436_18 (.CI(n39004), .I0(n2118), 
            .I1(VCC_net), .CO(n39005));
    SB_LUT4 encoder0_position_31__I_0_add_1436_17_lut (.I0(GND_net), .I1(n2119), 
            .I2(VCC_net), .I3(n39003), .O(n2186)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1436_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1436_17 (.CI(n39003), .I0(n2119), 
            .I1(VCC_net), .CO(n39004));
    SB_LUT4 encoder0_position_31__I_0_add_1436_16_lut (.I0(GND_net), .I1(n2120), 
            .I2(VCC_net), .I3(n39002), .O(n2187)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1436_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1436_16 (.CI(n39002), .I0(n2120), 
            .I1(VCC_net), .CO(n39003));
    SB_LUT4 encoder0_position_31__I_0_add_1436_15_lut (.I0(GND_net), .I1(n2121), 
            .I2(VCC_net), .I3(n39001), .O(n2188)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1436_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1436_15 (.CI(n39001), .I0(n2121), 
            .I1(VCC_net), .CO(n39002));
    SB_LUT4 encoder0_position_31__I_0_add_1436_14_lut (.I0(GND_net), .I1(n2122), 
            .I2(VCC_net), .I3(n39000), .O(n2189)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1436_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1436_14 (.CI(n39000), .I0(n2122), 
            .I1(VCC_net), .CO(n39001));
    SB_LUT4 encoder0_position_31__I_0_add_1436_13_lut (.I0(GND_net), .I1(n2123), 
            .I2(VCC_net), .I3(n38999), .O(n2190)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1436_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1436_13 (.CI(n38999), .I0(n2123), 
            .I1(VCC_net), .CO(n39000));
    SB_LUT4 encoder0_position_31__I_0_add_1436_12_lut (.I0(GND_net), .I1(n2124), 
            .I2(VCC_net), .I3(n38998), .O(n2191)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1436_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i2066_3_lut (.I0(n3031), .I1(n3098), 
            .I2(n3039), .I3(GND_net), .O(n3130));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i2066_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_1436_12 (.CI(n38998), .I0(n2124), 
            .I1(VCC_net), .CO(n38999));
    SB_LUT4 encoder0_position_31__I_0_add_1436_11_lut (.I0(GND_net), .I1(n2125), 
            .I2(VCC_net), .I3(n38997), .O(n2192)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1436_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1436_11 (.CI(n38997), .I0(n2125), 
            .I1(VCC_net), .CO(n38998));
    SB_LUT4 encoder0_position_31__I_0_add_1436_10_lut (.I0(GND_net), .I1(n2126), 
            .I2(VCC_net), .I3(n38996), .O(n2193)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1436_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1436_10 (.CI(n38996), .I0(n2126), 
            .I1(VCC_net), .CO(n38997));
    SB_LUT4 encoder0_position_31__I_0_add_1436_9_lut (.I0(GND_net), .I1(n2127), 
            .I2(VCC_net), .I3(n38995), .O(n2194)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1436_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1436_9 (.CI(n38995), .I0(n2127), 
            .I1(VCC_net), .CO(n38996));
    SB_LUT4 encoder0_position_31__I_0_add_1436_8_lut (.I0(GND_net), .I1(n2128), 
            .I2(VCC_net), .I3(n38994), .O(n2195_adj_5401)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1436_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1436_8 (.CI(n38994), .I0(n2128), 
            .I1(VCC_net), .CO(n38995));
    SB_LUT4 encoder0_position_31__I_0_add_1436_7_lut (.I0(GND_net), .I1(n2129), 
            .I2(GND_net), .I3(n38993), .O(n2196)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1436_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1436_7 (.CI(n38993), .I0(n2129), 
            .I1(GND_net), .CO(n38994));
    SB_LUT4 encoder0_position_31__I_0_add_1436_6_lut (.I0(GND_net), .I1(n2130), 
            .I2(GND_net), .I3(n38992), .O(n2197)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1436_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1436_6 (.CI(n38992), .I0(n2130), 
            .I1(GND_net), .CO(n38993));
    SB_LUT4 encoder0_position_31__I_0_add_1436_5_lut (.I0(GND_net), .I1(n2131), 
            .I2(VCC_net), .I3(n38991), .O(n2198)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1436_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1436_5 (.CI(n38991), .I0(n2131), 
            .I1(VCC_net), .CO(n38992));
    SB_LUT4 encoder0_position_31__I_0_add_1436_4_lut (.I0(GND_net), .I1(n2132), 
            .I2(GND_net), .I3(n38990), .O(n2199)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1436_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1436_4 (.CI(n38990), .I0(n2132), 
            .I1(GND_net), .CO(n38991));
    SB_LUT4 encoder0_position_31__I_0_add_1436_3_lut (.I0(GND_net), .I1(n2133), 
            .I2(VCC_net), .I3(n38989), .O(n2200)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1436_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1436_3 (.CI(n38989), .I0(n2133), 
            .I1(VCC_net), .CO(n38990));
    SB_LUT4 encoder0_position_31__I_0_add_1436_2_lut (.I0(GND_net), .I1(n532), 
            .I2(GND_net), .I3(VCC_net), .O(n2201)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1436_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1436_2 (.CI(VCC_net), .I0(n532), 
            .I1(GND_net), .CO(n38989));
    SB_LUT4 encoder0_position_31__I_0_i2065_3_lut (.I0(n3030), .I1(n3097), 
            .I2(n3039), .I3(GND_net), .O(n3129));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i2065_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1369_20_lut (.I0(n50937), .I1(n2016), 
            .I2(VCC_net), .I3(n38988), .O(n2115)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1369_20_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_31__I_0_i2069_3_lut (.I0(n541), .I1(n3101), 
            .I2(n3039), .I3(GND_net), .O(n3133));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i2069_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1369_19_lut (.I0(GND_net), .I1(n2017), 
            .I2(VCC_net), .I3(n38987), .O(n2084)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1369_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1369_19 (.CI(n38987), .I0(n2017), 
            .I1(VCC_net), .CO(n38988));
    SB_LUT4 encoder0_position_31__I_0_add_1369_18_lut (.I0(GND_net), .I1(n2018), 
            .I2(VCC_net), .I3(n38986), .O(n2085)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1369_18_lut.LUT_INIT = 16'hC33C;
    SB_DFF displacement_i23 (.Q(displacement[23]), .C(CLK_c), .D(displacement_23__N_99[23]));   // verilog/TinyFPGA_B.v(337[10] 341[6])
    SB_LUT4 i15078_3_lut (.I0(IntegralLimit[0]), .I1(\data_in_frame[13] [0]), 
            .I2(n28521), .I3(GND_net), .O(n29026));   // verilog/coms.v(128[12] 303[6])
    defparam i15078_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i2068_3_lut (.I0(n3033), .I1(n3100), 
            .I2(n3039), .I3(GND_net), .O(n3132));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i2068_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15079_4_lut (.I0(state_7__N_4267[3]), .I1(data[1]), .I2(n10_adj_5410), 
            .I3(n27152), .O(n29027));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i15079_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i3_3_lut (.I0(encoder0_position[2]), 
            .I1(n31), .I2(encoder0_position[31]), .I3(GND_net), .O(n542));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_mux_3_i3_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i2059_3_lut (.I0(n3024), .I1(n3091), 
            .I2(n3039), .I3(GND_net), .O(n3123));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i2059_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_1369_18 (.CI(n38986), .I0(n2018), 
            .I1(VCC_net), .CO(n38987));
    SB_LUT4 encoder0_position_31__I_0_add_1369_17_lut (.I0(GND_net), .I1(n2019), 
            .I2(VCC_net), .I3(n38985), .O(n2086)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1369_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1369_17 (.CI(n38985), .I0(n2019), 
            .I1(VCC_net), .CO(n38986));
    SB_LUT4 add_157_33_lut (.I0(GND_net), .I1(delay_counter[31]), .I2(GND_net), 
            .I3(n38476), .O(n1297)) /* synthesis syn_instantiated=1 */ ;
    defparam add_157_33_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15560_4_lut (.I0(r_Rx_Data), .I1(rx_data[4]), .I2(n4_adj_5362), 
            .I3(n27131), .O(n29508));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i15560_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 encoder0_position_31__I_0_add_1369_16_lut (.I0(GND_net), .I1(n2020), 
            .I2(VCC_net), .I3(n38984), .O(n2087)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1369_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i2062_3_lut (.I0(n3027), .I1(n3094), 
            .I2(n3039), .I3(GND_net), .O(n3126));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i2062_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2052_3_lut (.I0(n3017), .I1(n3084), 
            .I2(n3039), .I3(GND_net), .O(n3116));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i2052_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15080_4_lut (.I0(state_7__N_4267[3]), .I1(data[2]), .I2(n4_adj_5346), 
            .I3(n27147), .O(n29028));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i15080_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i15081_4_lut (.I0(state_7__N_4267[3]), .I1(data[3]), .I2(n4_adj_5346), 
            .I3(n27152), .O(n29029));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i15081_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 encoder0_position_31__I_0_i2061_3_lut (.I0(n3026), .I1(n3093), 
            .I2(n3039), .I3(GND_net), .O(n3125));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i2061_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2063_3_lut (.I0(n3028), .I1(n3095), 
            .I2(n3039), .I3(GND_net), .O(n3127));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i2063_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2055_3_lut (.I0(n3020), .I1(n3087), 
            .I2(n3039), .I3(GND_net), .O(n3119));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i2055_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15082_4_lut (.I0(state_7__N_4267[3]), .I1(data[4]), .I2(n4_adj_5248), 
            .I3(n27147), .O(n29030));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i15082_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 encoder0_position_31__I_0_i2056_3_lut (.I0(n3021), .I1(n3088), 
            .I2(n3039), .I3(GND_net), .O(n3120));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i2056_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2054_3_lut (.I0(n3019), .I1(n3086), 
            .I2(n3039), .I3(GND_net), .O(n3118));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i2054_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2049_3_lut (.I0(n3014), .I1(n3081), 
            .I2(n3039), .I3(GND_net), .O(n3113));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i2049_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_3_lut_adj_1784 (.I0(state_adj_5510[1]), .I1(read), .I2(n44835), 
            .I3(GND_net), .O(n12_adj_5286));   // verilog/eeprom.v(26[8] 58[4])
    defparam i1_3_lut_adj_1784.LUT_INIT = 16'ha2a2;
    SB_LUT4 i1_4_lut_adj_1785 (.I0(n34717), .I1(n12_adj_5286), .I2(state_adj_5510[0]), 
            .I3(n44835), .O(n43380));   // verilog/eeprom.v(26[8] 58[4])
    defparam i1_4_lut_adj_1785.LUT_INIT = 16'h88a8;
    SB_LUT4 i15083_4_lut (.I0(state_7__N_4267[3]), .I1(data[5]), .I2(n4_adj_5248), 
            .I3(n27152), .O(n29031));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i15083_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 encoder0_position_31__I_0_i2048_3_lut (.I0(n3013), .I1(n3080), 
            .I2(n3039), .I3(GND_net), .O(n3112));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i2048_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15084_4_lut (.I0(state_7__N_4267[3]), .I1(data[6]), .I2(n34660), 
            .I3(n27147), .O(n29032));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i15084_4_lut.LUT_INIT = 16'hccac;
    SB_CARRY encoder0_position_31__I_0_add_1369_16 (.CI(n38984), .I0(n2020), 
            .I1(VCC_net), .CO(n38985));
    SB_LUT4 add_157_11_lut (.I0(GND_net), .I1(delay_counter[9]), .I2(GND_net), 
            .I3(n38454), .O(n1319)) /* synthesis syn_instantiated=1 */ ;
    defparam add_157_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i2047_3_lut (.I0(n3012), .I1(n3079), 
            .I2(n3039), .I3(GND_net), .O(n3111));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i2047_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15085_4_lut (.I0(state_7__N_4267[3]), .I1(data[7]), .I2(n34660), 
            .I3(n27152), .O(n29033));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i15085_4_lut.LUT_INIT = 16'hccac;
    SB_LUT4 i15562_4_lut (.I0(r_Rx_Data), .I1(rx_data[5]), .I2(n4_adj_5362), 
            .I3(n27126), .O(n29510));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i15562_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 encoder0_position_31__I_0_i2051_3_lut (.I0(n3016), .I1(n3083), 
            .I2(n3039), .I3(GND_net), .O(n3115));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i2051_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2050_3_lut (.I0(n3015), .I1(n3082), 
            .I2(n3039), .I3(GND_net), .O(n3114));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i2050_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1786 (.I0(h3), .I1(commutation_state[1]), .I2(h2), 
            .I3(h1), .O(n43630));   // verilog/TinyFPGA_B.v(144[9] 223[5])
    defparam i1_4_lut_adj_1786.LUT_INIT = 16'hd054;
    SB_LUT4 encoder0_position_31__I_0_i2053_3_lut (.I0(n3018), .I1(n3085), 
            .I2(n3039), .I3(GND_net), .O(n3117));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i2053_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15092_3_lut (.I0(\data_in[0] [0]), .I1(\data_in[1] [0]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n29040));   // verilog/coms.v(128[12] 303[6])
    defparam i15092_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i2064_3_lut (.I0(n3029), .I1(n3096), 
            .I2(n3039), .I3(GND_net), .O(n3128));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i2064_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2057_3_lut (.I0(n3022), .I1(n3089), 
            .I2(n3039), .I3(GND_net), .O(n3121));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i2057_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1369_15_lut (.I0(GND_net), .I1(n2021), 
            .I2(VCC_net), .I3(n38983), .O(n2088)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1369_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1369_15 (.CI(n38983), .I0(n2021), 
            .I1(VCC_net), .CO(n38984));
    SB_LUT4 encoder0_position_31__I_0_add_1369_14_lut (.I0(GND_net), .I1(n2022), 
            .I2(VCC_net), .I3(n38982), .O(n2089)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1369_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i2058_3_lut (.I0(n3023), .I1(n3090), 
            .I2(n3039), .I3(GND_net), .O(n3122));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i2058_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2060_3_lut (.I0(n3025), .I1(n3092), 
            .I2(n3039), .I3(GND_net), .O(n3124));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i2060_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_1369_14 (.CI(n38982), .I0(n2022), 
            .I1(VCC_net), .CO(n38983));
    SB_LUT4 i15093_3_lut (.I0(Kp[0]), .I1(\data_in_frame[3] [0]), .I2(n28521), 
            .I3(GND_net), .O(n29041));   // verilog/coms.v(128[12] 303[6])
    defparam i15093_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_add_1369_13_lut (.I0(GND_net), .I1(n2023), 
            .I2(VCC_net), .I3(n38981), .O(n2090)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1369_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1369_13 (.CI(n38981), .I0(n2023), 
            .I1(VCC_net), .CO(n38982));
    SB_LUT4 n51462_bdd_4_lut (.I0(n51462), .I1(n341), .I2(n4486), .I3(n4208), 
            .O(pwm_setpoint_23__N_11[22]));
    defparam n51462_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n10621_bdd_4_lut_35834 (.I0(n10621), .I1(current[15]), .I2(duty[22]), 
            .I3(n4208), .O(n51462));
    defparam n10621_bdd_4_lut_35834.LUT_INIT = 16'he4aa;
    SB_LUT4 n51468_bdd_4_lut (.I0(n51468), .I1(n340), .I2(n4485), .I3(n4208), 
            .O(pwm_setpoint_23__N_11[23]));
    defparam n51468_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n10621_bdd_4_lut_35759 (.I0(n10621), .I1(current[7]), .I2(duty[7]), 
            .I3(n4208), .O(n51372));
    defparam n10621_bdd_4_lut_35759.LUT_INIT = 16'he4aa;
    SB_LUT4 n51372_bdd_4_lut (.I0(n51372), .I1(n356), .I2(n4501), .I3(n4208), 
            .O(pwm_setpoint_23__N_11[7]));
    defparam n51372_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n10621_bdd_4_lut_35754 (.I0(n10621), .I1(current[6]), .I2(duty[6]), 
            .I3(n4208), .O(n51366));
    defparam n10621_bdd_4_lut_35754.LUT_INIT = 16'he4aa;
    SB_LUT4 n51366_bdd_4_lut (.I0(n51366), .I1(n357), .I2(n4502), .I3(n4208), 
            .O(pwm_setpoint_23__N_11[6]));
    defparam n51366_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n10621_bdd_4_lut_35749 (.I0(n10621), .I1(current[5]), .I2(duty[5]), 
            .I3(n4208), .O(n51360));
    defparam n10621_bdd_4_lut_35749.LUT_INIT = 16'he4aa;
    SB_LUT4 n51360_bdd_4_lut (.I0(n51360), .I1(n358), .I2(n4503), .I3(n4208), 
            .O(pwm_setpoint_23__N_11[5]));
    defparam n51360_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n10621_bdd_4_lut_35744 (.I0(n10621), .I1(current[4]), .I2(duty[4]), 
            .I3(n4208), .O(n51354));
    defparam n10621_bdd_4_lut_35744.LUT_INIT = 16'he4aa;
    SB_LUT4 n51354_bdd_4_lut (.I0(n51354), .I1(n359), .I2(n4504), .I3(n4208), 
            .O(pwm_setpoint_23__N_11[4]));
    defparam n51354_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n10621_bdd_4_lut_35739 (.I0(n10621), .I1(current[3]), .I2(duty[3]), 
            .I3(n4208), .O(n51348));
    defparam n10621_bdd_4_lut_35739.LUT_INIT = 16'he4aa;
    SB_LUT4 n51348_bdd_4_lut (.I0(n51348), .I1(n360), .I2(n4505), .I3(n4208), 
            .O(pwm_setpoint_23__N_11[3]));
    defparam n51348_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n10621_bdd_4_lut_35734 (.I0(n10621), .I1(current[2]), .I2(duty[2]), 
            .I3(n4208), .O(n51342));
    defparam n10621_bdd_4_lut_35734.LUT_INIT = 16'he4aa;
    SB_LUT4 n51342_bdd_4_lut (.I0(n51342), .I1(n361), .I2(n4506), .I3(n4208), 
            .O(pwm_setpoint_23__N_11[2]));
    defparam n51342_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n10621_bdd_4_lut_35729 (.I0(n10621), .I1(current[1]), .I2(duty[1]), 
            .I3(n4208), .O(n51336));
    defparam n10621_bdd_4_lut_35729.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_4_lut_adj_1787 (.I0(n5_adj_5368), .I1(\ID_READOUT_FSM.state [0]), 
            .I2(n2204), .I3(read_N_445), .O(n25_adj_5270));   // verilog/TinyFPGA_B.v(375[10] 403[6])
    defparam i1_4_lut_adj_1787.LUT_INIT = 16'h7350;
    SB_LUT4 i32450_2_lut (.I0(data_ready), .I1(\ID_READOUT_FSM.state [0]), 
            .I2(GND_net), .I3(GND_net), .O(n47975));
    defparam i32450_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i15094_3_lut (.I0(Ki[0]), .I1(\data_in_frame[5] [0]), .I2(n28521), 
            .I3(GND_net), .O(n29042));   // verilog/coms.v(128[12] 303[6])
    defparam i15094_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1788 (.I0(n3124), .I1(n3122), .I2(n3121), .I3(n3128), 
            .O(n46717));
    defparam i1_4_lut_adj_1788.LUT_INIT = 16'hfffe;
    SB_LUT4 i35530_4_lut (.I0(\ID_READOUT_FSM.state [1]), .I1(n7494), .I2(n47975), 
            .I3(n25_adj_5270), .O(n17_adj_5271));   // verilog/TinyFPGA_B.v(375[10] 403[6])
    defparam i35530_4_lut.LUT_INIT = 16'h88ba;
    SB_LUT4 i1_4_lut_adj_1789 (.I0(n3118), .I1(n3120), .I2(n3119), .I3(n3127), 
            .O(n46719));
    defparam i1_4_lut_adj_1789.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1790 (.I0(n3125), .I1(n3116), .I2(n3126), .I3(n3123), 
            .O(n45800));
    defparam i1_4_lut_adj_1790.LUT_INIT = 16'hfffe;
    SB_LUT4 i15095_3_lut (.I0(neopxl_color[0]), .I1(\data_in_frame[6] [0]), 
            .I2(n28522), .I3(GND_net), .O(n29043));   // verilog/coms.v(128[12] 303[6])
    defparam i15095_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i21444_3_lut (.I0(n542), .I1(n3132), .I2(n3133), .I3(GND_net), 
            .O(n35392));
    defparam i21444_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i1_4_lut_adj_1791 (.I0(n45800), .I1(n3117), .I2(n46719), .I3(n46717), 
            .O(n46725));
    defparam i1_4_lut_adj_1791.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1792 (.I0(n3129), .I1(n35392), .I2(n3130), .I3(n3131), 
            .O(n45016));
    defparam i1_4_lut_adj_1792.LUT_INIT = 16'ha080;
    SB_LUT4 i15568_4_lut (.I0(r_Rx_Data), .I1(rx_data[6]), .I2(n34695), 
            .I3(n27131), .O(n29516));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i15568_4_lut.LUT_INIT = 16'hccac;
    SB_LUT4 i1_4_lut_adj_1793 (.I0(n3114), .I1(n45016), .I2(n46725), .I3(n3115), 
            .O(n46731));
    defparam i1_4_lut_adj_1793.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1794 (.I0(n3111), .I1(n3112), .I2(n3113), .I3(n46731), 
            .O(n46737));
    defparam i1_4_lut_adj_1794.LUT_INIT = 16'hfffe;
    SB_LUT4 i15569_3_lut (.I0(\data_out_frame[25] [0]), .I1(neopxl_color[0]), 
            .I2(n24278), .I3(GND_net), .O(n29517));   // verilog/coms.v(128[12] 303[6])
    defparam i15569_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_add_1369_12_lut (.I0(GND_net), .I1(n2024), 
            .I2(VCC_net), .I3(n38980), .O(n2091)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1369_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1369_12 (.CI(n38980), .I0(n2024), 
            .I1(VCC_net), .CO(n38981));
    SB_LUT4 encoder0_position_31__I_0_add_1369_11_lut (.I0(GND_net), .I1(n2025), 
            .I2(VCC_net), .I3(n38979), .O(n2092)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1369_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1369_11 (.CI(n38979), .I0(n2025), 
            .I1(VCC_net), .CO(n38980));
    SB_LUT4 i15570_3_lut (.I0(\data_out_frame[24] [7]), .I1(neopxl_color[15]), 
            .I2(n24278), .I3(GND_net), .O(n29518));   // verilog/coms.v(128[12] 303[6])
    defparam i15570_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15571_3_lut (.I0(\data_out_frame[24] [6]), .I1(neopxl_color[14]), 
            .I2(n24278), .I3(GND_net), .O(n29519));   // verilog/coms.v(128[12] 303[6])
    defparam i15571_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF displacement_i22 (.Q(displacement[22]), .C(CLK_c), .D(displacement_23__N_99[22]));   // verilog/TinyFPGA_B.v(337[10] 341[6])
    SB_LUT4 encoder0_position_31__I_0_add_1369_10_lut (.I0(GND_net), .I1(n2026), 
            .I2(VCC_net), .I3(n38978), .O(n2093)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1369_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1795 (.I0(n3108), .I1(n3109), .I2(n3110), .I3(n46737), 
            .O(n46743));
    defparam i1_4_lut_adj_1795.LUT_INIT = 16'hfffe;
    SB_LUT4 i15572_3_lut (.I0(\data_out_frame[24] [5]), .I1(neopxl_color[13]), 
            .I2(n24278), .I3(GND_net), .O(n29520));   // verilog/coms.v(128[12] 303[6])
    defparam i15572_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15573_3_lut (.I0(\data_out_frame[24] [4]), .I1(neopxl_color[12]), 
            .I2(n24278), .I3(GND_net), .O(n29521));   // verilog/coms.v(128[12] 303[6])
    defparam i15573_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF displacement_i21 (.Q(displacement[21]), .C(CLK_c), .D(displacement_23__N_99[21]));   // verilog/TinyFPGA_B.v(337[10] 341[6])
    SB_DFF displacement_i20 (.Q(displacement[20]), .C(CLK_c), .D(displacement_23__N_99[20]));   // verilog/TinyFPGA_B.v(337[10] 341[6])
    SB_DFF displacement_i19 (.Q(displacement[19]), .C(CLK_c), .D(displacement_23__N_99[19]));   // verilog/TinyFPGA_B.v(337[10] 341[6])
    SB_DFF displacement_i18 (.Q(displacement[18]), .C(CLK_c), .D(displacement_23__N_99[18]));   // verilog/TinyFPGA_B.v(337[10] 341[6])
    SB_DFF displacement_i17 (.Q(displacement[17]), .C(CLK_c), .D(displacement_23__N_99[17]));   // verilog/TinyFPGA_B.v(337[10] 341[6])
    SB_DFF displacement_i16 (.Q(displacement[16]), .C(CLK_c), .D(displacement_23__N_99[16]));   // verilog/TinyFPGA_B.v(337[10] 341[6])
    SB_DFF displacement_i15 (.Q(displacement[15]), .C(CLK_c), .D(displacement_23__N_99[15]));   // verilog/TinyFPGA_B.v(337[10] 341[6])
    SB_DFF displacement_i14 (.Q(displacement[14]), .C(CLK_c), .D(displacement_23__N_99[14]));   // verilog/TinyFPGA_B.v(337[10] 341[6])
    SB_DFF displacement_i13 (.Q(displacement[13]), .C(CLK_c), .D(displacement_23__N_99[13]));   // verilog/TinyFPGA_B.v(337[10] 341[6])
    SB_DFF displacement_i12 (.Q(displacement[12]), .C(CLK_c), .D(displacement_23__N_99[12]));   // verilog/TinyFPGA_B.v(337[10] 341[6])
    SB_DFF displacement_i11 (.Q(displacement[11]), .C(CLK_c), .D(displacement_23__N_99[11]));   // verilog/TinyFPGA_B.v(337[10] 341[6])
    SB_DFF displacement_i10 (.Q(displacement[10]), .C(CLK_c), .D(displacement_23__N_99[10]));   // verilog/TinyFPGA_B.v(337[10] 341[6])
    SB_DFF displacement_i9 (.Q(displacement[9]), .C(CLK_c), .D(displacement_23__N_99[9]));   // verilog/TinyFPGA_B.v(337[10] 341[6])
    SB_DFF displacement_i8 (.Q(displacement[8]), .C(CLK_c), .D(displacement_23__N_99[8]));   // verilog/TinyFPGA_B.v(337[10] 341[6])
    SB_DFF displacement_i7 (.Q(displacement[7]), .C(CLK_c), .D(displacement_23__N_99[7]));   // verilog/TinyFPGA_B.v(337[10] 341[6])
    SB_DFF displacement_i6 (.Q(displacement[6]), .C(CLK_c), .D(displacement_23__N_99[6]));   // verilog/TinyFPGA_B.v(337[10] 341[6])
    SB_DFF displacement_i5 (.Q(displacement[5]), .C(CLK_c), .D(displacement_23__N_99[5]));   // verilog/TinyFPGA_B.v(337[10] 341[6])
    SB_DFF displacement_i4 (.Q(displacement[4]), .C(CLK_c), .D(displacement_23__N_99[4]));   // verilog/TinyFPGA_B.v(337[10] 341[6])
    SB_DFF displacement_i3 (.Q(displacement[3]), .C(CLK_c), .D(displacement_23__N_99[3]));   // verilog/TinyFPGA_B.v(337[10] 341[6])
    SB_DFF displacement_i2 (.Q(displacement[2]), .C(CLK_c), .D(displacement_23__N_99[2]));   // verilog/TinyFPGA_B.v(337[10] 341[6])
    SB_DFF displacement_i1 (.Q(displacement[1]), .C(CLK_c), .D(displacement_23__N_99[1]));   // verilog/TinyFPGA_B.v(337[10] 341[6])
    SB_DFF encoder1_position_scaled_i23 (.Q(encoder1_position_scaled[23]), 
           .C(CLK_c), .D(encoder1_position_scaled_23__N_75[23]));   // verilog/TinyFPGA_B.v(337[10] 341[6])
    SB_DFF encoder1_position_scaled_i22 (.Q(encoder1_position_scaled[22]), 
           .C(CLK_c), .D(encoder1_position_scaled_23__N_75[22]));   // verilog/TinyFPGA_B.v(337[10] 341[6])
    SB_DFF encoder1_position_scaled_i21 (.Q(encoder1_position_scaled[21]), 
           .C(CLK_c), .D(encoder1_position_scaled_23__N_75[21]));   // verilog/TinyFPGA_B.v(337[10] 341[6])
    SB_DFF encoder1_position_scaled_i20 (.Q(encoder1_position_scaled[20]), 
           .C(CLK_c), .D(encoder1_position_scaled_23__N_75[20]));   // verilog/TinyFPGA_B.v(337[10] 341[6])
    SB_DFF encoder1_position_scaled_i19 (.Q(encoder1_position_scaled[19]), 
           .C(CLK_c), .D(encoder1_position_scaled_23__N_75[19]));   // verilog/TinyFPGA_B.v(337[10] 341[6])
    SB_DFF encoder1_position_scaled_i18 (.Q(encoder1_position_scaled[18]), 
           .C(CLK_c), .D(encoder1_position_scaled_23__N_75[18]));   // verilog/TinyFPGA_B.v(337[10] 341[6])
    SB_DFF encoder1_position_scaled_i17 (.Q(encoder1_position_scaled[17]), 
           .C(CLK_c), .D(encoder1_position_scaled_23__N_75[17]));   // verilog/TinyFPGA_B.v(337[10] 341[6])
    SB_DFF encoder1_position_scaled_i16 (.Q(encoder1_position_scaled[16]), 
           .C(CLK_c), .D(encoder1_position_scaled_23__N_75[16]));   // verilog/TinyFPGA_B.v(337[10] 341[6])
    SB_DFF encoder1_position_scaled_i15 (.Q(encoder1_position_scaled[15]), 
           .C(CLK_c), .D(encoder1_position_scaled_23__N_75[15]));   // verilog/TinyFPGA_B.v(337[10] 341[6])
    SB_DFF encoder1_position_scaled_i14 (.Q(encoder1_position_scaled[14]), 
           .C(CLK_c), .D(encoder1_position_scaled_23__N_75[14]));   // verilog/TinyFPGA_B.v(337[10] 341[6])
    SB_DFF encoder1_position_scaled_i13 (.Q(encoder1_position_scaled[13]), 
           .C(CLK_c), .D(encoder1_position_scaled_23__N_75[13]));   // verilog/TinyFPGA_B.v(337[10] 341[6])
    SB_DFF encoder1_position_scaled_i12 (.Q(encoder1_position_scaled[12]), 
           .C(CLK_c), .D(encoder1_position_scaled_23__N_75[12]));   // verilog/TinyFPGA_B.v(337[10] 341[6])
    SB_DFF encoder1_position_scaled_i11 (.Q(encoder1_position_scaled[11]), 
           .C(CLK_c), .D(encoder1_position_scaled_23__N_75[11]));   // verilog/TinyFPGA_B.v(337[10] 341[6])
    SB_DFF encoder1_position_scaled_i10 (.Q(encoder1_position_scaled[10]), 
           .C(CLK_c), .D(encoder1_position_scaled_23__N_75[10]));   // verilog/TinyFPGA_B.v(337[10] 341[6])
    SB_DFF encoder1_position_scaled_i9 (.Q(encoder1_position_scaled[9]), .C(CLK_c), 
           .D(encoder1_position_scaled_23__N_75[9]));   // verilog/TinyFPGA_B.v(337[10] 341[6])
    SB_DFF encoder1_position_scaled_i8 (.Q(encoder1_position_scaled[8]), .C(CLK_c), 
           .D(encoder1_position_scaled_23__N_75[8]));   // verilog/TinyFPGA_B.v(337[10] 341[6])
    SB_DFF encoder1_position_scaled_i7 (.Q(encoder1_position_scaled[7]), .C(CLK_c), 
           .D(encoder1_position_scaled_23__N_75[7]));   // verilog/TinyFPGA_B.v(337[10] 341[6])
    SB_DFF encoder1_position_scaled_i6 (.Q(encoder1_position_scaled[6]), .C(CLK_c), 
           .D(encoder1_position_scaled_23__N_75[6]));   // verilog/TinyFPGA_B.v(337[10] 341[6])
    SB_DFF encoder1_position_scaled_i5 (.Q(encoder1_position_scaled[5]), .C(CLK_c), 
           .D(encoder1_position_scaled_23__N_75[5]));   // verilog/TinyFPGA_B.v(337[10] 341[6])
    SB_DFF encoder1_position_scaled_i4 (.Q(encoder1_position_scaled[4]), .C(CLK_c), 
           .D(encoder1_position_scaled_23__N_75[4]));   // verilog/TinyFPGA_B.v(337[10] 341[6])
    SB_DFF encoder1_position_scaled_i3 (.Q(encoder1_position_scaled[3]), .C(CLK_c), 
           .D(encoder1_position_scaled_23__N_75[3]));   // verilog/TinyFPGA_B.v(337[10] 341[6])
    SB_DFF encoder1_position_scaled_i2 (.Q(encoder1_position_scaled[2]), .C(CLK_c), 
           .D(encoder1_position_scaled_23__N_75[2]));   // verilog/TinyFPGA_B.v(337[10] 341[6])
    SB_DFF encoder1_position_scaled_i1 (.Q(encoder1_position_scaled[1]), .C(CLK_c), 
           .D(encoder1_position_scaled_23__N_75[1]));   // verilog/TinyFPGA_B.v(337[10] 341[6])
    SB_CARRY encoder0_position_31__I_0_add_1369_10 (.CI(n38978), .I0(n2026), 
            .I1(VCC_net), .CO(n38979));
    SB_LUT4 encoder0_position_31__I_0_add_1369_9_lut (.I0(GND_net), .I1(n2027), 
            .I2(VCC_net), .I3(n38977), .O(n2094)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1369_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1369_9 (.CI(n38977), .I0(n2027), 
            .I1(VCC_net), .CO(n38978));
    SB_LUT4 encoder0_position_31__I_0_add_1369_8_lut (.I0(GND_net), .I1(n2028), 
            .I2(VCC_net), .I3(n38976), .O(n2095)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1369_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1369_8 (.CI(n38976), .I0(n2028), 
            .I1(VCC_net), .CO(n38977));
    SB_LUT4 encoder0_position_31__I_0_add_1369_7_lut (.I0(GND_net), .I1(n2029), 
            .I2(GND_net), .I3(n38975), .O(n2096)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1369_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1369_7 (.CI(n38975), .I0(n2029), 
            .I1(GND_net), .CO(n38976));
    SB_LUT4 encoder0_position_31__I_0_add_1369_6_lut (.I0(GND_net), .I1(n2030), 
            .I2(GND_net), .I3(n38974), .O(n2097)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1369_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1369_6 (.CI(n38974), .I0(n2030), 
            .I1(GND_net), .CO(n38975));
    SB_LUT4 encoder0_position_31__I_0_add_1369_5_lut (.I0(GND_net), .I1(n2031), 
            .I2(VCC_net), .I3(n38973), .O(n2098)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1369_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1369_5 (.CI(n38973), .I0(n2031), 
            .I1(VCC_net), .CO(n38974));
    SB_LUT4 encoder0_position_31__I_0_add_1369_4_lut (.I0(GND_net), .I1(n2032), 
            .I2(GND_net), .I3(n38972), .O(n2099)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1369_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1369_4 (.CI(n38972), .I0(n2032), 
            .I1(GND_net), .CO(n38973));
    SB_LUT4 encoder0_position_31__I_0_add_1369_3_lut (.I0(GND_net), .I1(n2033), 
            .I2(VCC_net), .I3(n38971), .O(n2100)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1369_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1369_3 (.CI(n38971), .I0(n2033), 
            .I1(VCC_net), .CO(n38972));
    SB_LUT4 encoder0_position_31__I_0_add_1369_2_lut (.I0(GND_net), .I1(n531), 
            .I2(GND_net), .I3(VCC_net), .O(n2101)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1369_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1369_2 (.CI(VCC_net), .I0(n531), 
            .I1(GND_net), .CO(n38971));
    SB_LUT4 encoder0_position_31__I_0_add_1302_19_lut (.I0(n50958), .I1(n1917), 
            .I2(VCC_net), .I3(n38970), .O(n2016)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1302_19_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_31__I_0_add_1302_18_lut (.I0(GND_net), .I1(n1918), 
            .I2(VCC_net), .I3(n38969), .O(n1985)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1302_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1302_18 (.CI(n38969), .I0(n1918), 
            .I1(VCC_net), .CO(n38970));
    SB_LUT4 encoder0_position_31__I_0_add_1302_17_lut (.I0(GND_net), .I1(n1919), 
            .I2(VCC_net), .I3(n38968), .O(n1986)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1302_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1302_17 (.CI(n38968), .I0(n1919), 
            .I1(VCC_net), .CO(n38969));
    SB_LUT4 encoder0_position_31__I_0_add_1302_16_lut (.I0(GND_net), .I1(n1920), 
            .I2(VCC_net), .I3(n38967), .O(n1987)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1302_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1302_16 (.CI(n38967), .I0(n1920), 
            .I1(VCC_net), .CO(n38968));
    SB_LUT4 encoder0_position_31__I_0_add_1302_15_lut (.I0(GND_net), .I1(n1921), 
            .I2(VCC_net), .I3(n38966), .O(n1988)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1302_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1302_15 (.CI(n38966), .I0(n1921), 
            .I1(VCC_net), .CO(n38967));
    SB_LUT4 encoder0_position_31__I_0_add_1302_14_lut (.I0(GND_net), .I1(n1922), 
            .I2(VCC_net), .I3(n38965), .O(n1989)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1302_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1302_14 (.CI(n38965), .I0(n1922), 
            .I1(VCC_net), .CO(n38966));
    SB_LUT4 encoder0_position_31__I_0_add_1302_13_lut (.I0(GND_net), .I1(n1923), 
            .I2(VCC_net), .I3(n38964), .O(n1990)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1302_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15574_3_lut (.I0(\data_out_frame[24] [3]), .I1(neopxl_color[11]), 
            .I2(n24278), .I3(GND_net), .O(n29522));   // verilog/coms.v(128[12] 303[6])
    defparam i15574_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1005_i13_3_lut (.I0(duty[12]), .I1(n351), .I2(duty[23]), 
            .I3(GND_net), .O(n4711));   // verilog/TinyFPGA_B.v(118[13] 129[7])
    defparam mux_1005_i13_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_31__I_0_add_1302_13 (.CI(n38964), .I0(n1923), 
            .I1(VCC_net), .CO(n38965));
    SB_LUT4 i15575_3_lut (.I0(\data_out_frame[24] [2]), .I1(neopxl_color[10]), 
            .I2(n24278), .I3(GND_net), .O(n29523));   // verilog/coms.v(128[12] 303[6])
    defparam i15575_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34959_4_lut (.I0(n3106), .I1(n3105), .I2(n3107), .I3(n46743), 
            .O(n3138));
    defparam i34959_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_31__I_0_i1976_3_lut (.I0(n2909), .I1(n2976), 
            .I2(n2940), .I3(GND_net), .O(n3008));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1976_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15097_3_lut (.I0(control_mode[0]), .I1(\data_in_frame[1] [0]), 
            .I2(n28521), .I3(GND_net), .O(n29045));   // verilog/coms.v(128[12] 303[6])
    defparam i15097_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15098_3_lut (.I0(current_limit[0]), .I1(\data_in_frame[21] [0]), 
            .I2(n28521), .I3(GND_net), .O(n29046));   // verilog/coms.v(128[12] 303[6])
    defparam i15098_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i1975_3_lut (.I0(n2908), .I1(n2975), 
            .I2(n2940), .I3(GND_net), .O(n3007));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1975_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15099_3_lut (.I0(PWMLimit[0]), .I1(\data_in_frame[10] [0]), 
            .I2(n28521), .I3(GND_net), .O(n29047));   // verilog/coms.v(128[12] 303[6])
    defparam i15099_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i1979_3_lut (.I0(n2912), .I1(n2979), 
            .I2(n2940), .I3(GND_net), .O(n3011));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1979_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1978_3_lut (.I0(n2911), .I1(n2978), 
            .I2(n2940), .I3(GND_net), .O(n3010));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1978_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1977_3_lut (.I0(n2910), .I1(n2977), 
            .I2(n2940), .I3(GND_net), .O(n3009));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1977_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1999_3_lut (.I0(n2932), .I1(n2999), 
            .I2(n2940), .I3(GND_net), .O(n3031));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1999_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1998_3_lut (.I0(n2931), .I1(n2998), 
            .I2(n2940), .I3(GND_net), .O(n3030));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1998_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15576_4_lut (.I0(r_Rx_Data), .I1(rx_data[7]), .I2(n34695), 
            .I3(n27126), .O(n29524));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i15576_4_lut.LUT_INIT = 16'hccac;
    SB_DFF encoder0_position_scaled_i23 (.Q(encoder0_position_scaled[23]), 
           .C(CLK_c), .D(encoder0_position_scaled_23__N_51[23]));   // verilog/TinyFPGA_B.v(337[10] 341[6])
    SB_LUT4 i15577_3_lut (.I0(\data_out_frame[24] [1]), .I1(neopxl_color[9]), 
            .I2(n24278), .I3(GND_net), .O(n29525));   // verilog/coms.v(128[12] 303[6])
    defparam i15577_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i1997_3_lut (.I0(n2930), .I1(n2997), 
            .I2(n2940), .I3(GND_net), .O(n3029));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1997_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1302_12_lut (.I0(GND_net), .I1(n1924), 
            .I2(VCC_net), .I3(n38963), .O(n1991)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1302_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15578_3_lut (.I0(\data_out_frame[24] [0]), .I1(neopxl_color[8]), 
            .I2(n24278), .I3(GND_net), .O(n29526));   // verilog/coms.v(128[12] 303[6])
    defparam i15578_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i2001_3_lut (.I0(n540), .I1(n3001), 
            .I2(n2940), .I3(GND_net), .O(n3033));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i2001_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2000_3_lut (.I0(n2933), .I1(n3000), 
            .I2(n2940), .I3(GND_net), .O(n3032));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i2000_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i4_3_lut (.I0(encoder0_position[3]), 
            .I1(n30), .I2(encoder0_position[31]), .I3(GND_net), .O(n541));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_mux_3_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i1994_3_lut (.I0(n2927), .I1(n2994), 
            .I2(n2940), .I3(GND_net), .O(n3026));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1994_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1996_3_lut (.I0(n2929), .I1(n2996), 
            .I2(n2940), .I3(GND_net), .O(n3028));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1996_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1990_3_lut (.I0(n2923), .I1(n2990), 
            .I2(n2940), .I3(GND_net), .O(n3022));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1990_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1995_3_lut (.I0(n2928), .I1(n2995), 
            .I2(n2940), .I3(GND_net), .O(n3027));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1995_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1982_3_lut (.I0(n2915), .I1(n2982), 
            .I2(n2940), .I3(GND_net), .O(n3014));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1982_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 unary_minus_19_inv_0_i4_1_lut (.I0(duty[3]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n22_adj_5267));   // verilog/TinyFPGA_B.v(123[25:30])
    defparam unary_minus_19_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_31__I_0_add_1302_12 (.CI(n38963), .I0(n1924), 
            .I1(VCC_net), .CO(n38964));
    SB_DFF encoder0_position_scaled_i22 (.Q(encoder0_position_scaled[22]), 
           .C(CLK_c), .D(encoder0_position_scaled_23__N_51[22]));   // verilog/TinyFPGA_B.v(337[10] 341[6])
    SB_DFF encoder0_position_scaled_i21 (.Q(encoder0_position_scaled[21]), 
           .C(CLK_c), .D(encoder0_position_scaled_23__N_51[21]));   // verilog/TinyFPGA_B.v(337[10] 341[6])
    SB_LUT4 encoder0_position_31__I_0_add_1302_11_lut (.I0(GND_net), .I1(n1925), 
            .I2(VCC_net), .I3(n38962), .O(n1992)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1302_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1302_11 (.CI(n38962), .I0(n1925), 
            .I1(VCC_net), .CO(n38963));
    SB_LUT4 encoder0_position_31__I_0_add_1302_10_lut (.I0(GND_net), .I1(n1926), 
            .I2(VCC_net), .I3(n38961), .O(n1993)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1302_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_157_11 (.CI(n38454), .I0(delay_counter[9]), .I1(GND_net), 
            .CO(n38455));
    SB_LUT4 add_157_4_lut (.I0(GND_net), .I1(delay_counter[2]), .I2(GND_net), 
            .I3(n38447), .O(n1326)) /* synthesis syn_instantiated=1 */ ;
    defparam add_157_4_lut.LUT_INIT = 16'hC33C;
    SB_DFF \ID_READOUT_FSM.state__i0  (.Q(\ID_READOUT_FSM.state [0]), .C(CLK_c), 
           .D(n42724));   // verilog/TinyFPGA_B.v(375[10] 403[6])
    SB_CARRY encoder0_position_31__I_0_add_1302_10 (.CI(n38961), .I0(n1926), 
            .I1(VCC_net), .CO(n38962));
    SB_LUT4 add_157_32_lut (.I0(GND_net), .I1(delay_counter[30]), .I2(GND_net), 
            .I3(n38475), .O(n1298)) /* synthesis syn_instantiated=1 */ ;
    defparam add_157_32_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1302_9_lut (.I0(GND_net), .I1(n1927), 
            .I2(VCC_net), .I3(n38960), .O(n1994)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1302_9_lut.LUT_INIT = 16'hC33C;
    SB_DFF encoder0_position_scaled_i20 (.Q(encoder0_position_scaled[20]), 
           .C(CLK_c), .D(encoder0_position_scaled_23__N_51[20]));   // verilog/TinyFPGA_B.v(337[10] 341[6])
    SB_CARRY add_157_32 (.CI(n38475), .I0(delay_counter[30]), .I1(GND_net), 
            .CO(n38476));
    SB_CARRY encoder0_position_31__I_0_add_1302_9 (.CI(n38960), .I0(n1927), 
            .I1(VCC_net), .CO(n38961));
    SB_DFF encoder0_position_scaled_i19 (.Q(encoder0_position_scaled[19]), 
           .C(CLK_c), .D(encoder0_position_scaled_23__N_51[19]));   // verilog/TinyFPGA_B.v(337[10] 341[6])
    SB_LUT4 n51336_bdd_4_lut (.I0(n51336), .I1(n362), .I2(n4507), .I3(n4208), 
            .O(pwm_setpoint_23__N_11[1]));
    defparam n51336_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF encoder0_position_scaled_i18 (.Q(encoder0_position_scaled[18]), 
           .C(CLK_c), .D(encoder0_position_scaled_23__N_51[18]));   // verilog/TinyFPGA_B.v(337[10] 341[6])
    SB_DFF encoder0_position_scaled_i17 (.Q(encoder0_position_scaled[17]), 
           .C(CLK_c), .D(encoder0_position_scaled_23__N_51[17]));   // verilog/TinyFPGA_B.v(337[10] 341[6])
    SB_LUT4 encoder0_position_31__I_0_add_1302_8_lut (.I0(GND_net), .I1(n1928), 
            .I2(VCC_net), .I3(n38959), .O(n1995)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1302_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1302_8 (.CI(n38959), .I0(n1928), 
            .I1(VCC_net), .CO(n38960));
    SB_DFF encoder0_position_scaled_i16 (.Q(encoder0_position_scaled[16]), 
           .C(CLK_c), .D(encoder0_position_scaled_23__N_51[16]));   // verilog/TinyFPGA_B.v(337[10] 341[6])
    SB_DFF encoder0_position_scaled_i15 (.Q(encoder0_position_scaled[15]), 
           .C(CLK_c), .D(encoder0_position_scaled_23__N_51[15]));   // verilog/TinyFPGA_B.v(337[10] 341[6])
    SB_DFF encoder0_position_scaled_i14 (.Q(encoder0_position_scaled[14]), 
           .C(CLK_c), .D(encoder0_position_scaled_23__N_51[14]));   // verilog/TinyFPGA_B.v(337[10] 341[6])
    SB_DFF encoder0_position_scaled_i13 (.Q(encoder0_position_scaled[13]), 
           .C(CLK_c), .D(encoder0_position_scaled_23__N_51[13]));   // verilog/TinyFPGA_B.v(337[10] 341[6])
    SB_DFF encoder0_position_scaled_i12 (.Q(encoder0_position_scaled[12]), 
           .C(CLK_c), .D(encoder0_position_scaled_23__N_51[12]));   // verilog/TinyFPGA_B.v(337[10] 341[6])
    SB_DFF encoder0_position_scaled_i11 (.Q(encoder0_position_scaled[11]), 
           .C(CLK_c), .D(encoder0_position_scaled_23__N_51[11]));   // verilog/TinyFPGA_B.v(337[10] 341[6])
    SB_DFF encoder0_position_scaled_i10 (.Q(encoder0_position_scaled[10]), 
           .C(CLK_c), .D(encoder0_position_scaled_23__N_51[10]));   // verilog/TinyFPGA_B.v(337[10] 341[6])
    SB_DFF encoder0_position_scaled_i9 (.Q(encoder0_position_scaled[9]), .C(CLK_c), 
           .D(encoder0_position_scaled_23__N_51[9]));   // verilog/TinyFPGA_B.v(337[10] 341[6])
    SB_DFF encoder0_position_scaled_i8 (.Q(encoder0_position_scaled[8]), .C(CLK_c), 
           .D(encoder0_position_scaled_23__N_51[8]));   // verilog/TinyFPGA_B.v(337[10] 341[6])
    SB_DFF encoder0_position_scaled_i7 (.Q(encoder0_position_scaled[7]), .C(CLK_c), 
           .D(encoder0_position_scaled_23__N_51[7]));   // verilog/TinyFPGA_B.v(337[10] 341[6])
    SB_DFF encoder0_position_scaled_i6 (.Q(encoder0_position_scaled[6]), .C(CLK_c), 
           .D(encoder0_position_scaled_23__N_51[6]));   // verilog/TinyFPGA_B.v(337[10] 341[6])
    SB_DFF encoder0_position_scaled_i5 (.Q(encoder0_position_scaled[5]), .C(CLK_c), 
           .D(encoder0_position_scaled_23__N_51[5]));   // verilog/TinyFPGA_B.v(337[10] 341[6])
    SB_DFF encoder0_position_scaled_i4 (.Q(encoder0_position_scaled[4]), .C(CLK_c), 
           .D(encoder0_position_scaled_23__N_51[4]));   // verilog/TinyFPGA_B.v(337[10] 341[6])
    SB_DFF encoder0_position_scaled_i3 (.Q(encoder0_position_scaled[3]), .C(CLK_c), 
           .D(encoder0_position_scaled_23__N_51[3]));   // verilog/TinyFPGA_B.v(337[10] 341[6])
    SB_DFF encoder0_position_scaled_i2 (.Q(encoder0_position_scaled[2]), .C(CLK_c), 
           .D(encoder0_position_scaled_23__N_51[2]));   // verilog/TinyFPGA_B.v(337[10] 341[6])
    SB_DFF encoder0_position_scaled_i1 (.Q(encoder0_position_scaled[1]), .C(CLK_c), 
           .D(encoder0_position_scaled_23__N_51[1]));   // verilog/TinyFPGA_B.v(337[10] 341[6])
    SB_LUT4 encoder0_position_31__I_0_i1981_3_lut (.I0(n2914), .I1(n2981), 
            .I2(n2940), .I3(GND_net), .O(n3013));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1981_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1302_7_lut (.I0(GND_net), .I1(n1929), 
            .I2(GND_net), .I3(n38958), .O(n1996)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1302_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1980_3_lut (.I0(n2913), .I1(n2980), 
            .I2(n2940), .I3(GND_net), .O(n3012));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1980_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1984_3_lut (.I0(n2917), .I1(n2984), 
            .I2(n2940), .I3(GND_net), .O(n3016));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1984_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1983_3_lut (.I0(n2916), .I1(n2983), 
            .I2(n2940), .I3(GND_net), .O(n3015));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1983_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1986_3_lut (.I0(n2919), .I1(n2986), 
            .I2(n2940), .I3(GND_net), .O(n3018));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1986_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1985_3_lut (.I0(n2918), .I1(n2985), 
            .I2(n2940), .I3(GND_net), .O(n3017));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1985_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1988_3_lut (.I0(n2921), .I1(n2988), 
            .I2(n2940), .I3(GND_net), .O(n3020));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1988_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1987_3_lut (.I0(n2920), .I1(n2987), 
            .I2(n2940), .I3(GND_net), .O(n3019));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1987_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1993_3_lut (.I0(n2926), .I1(n2993), 
            .I2(n2940), .I3(GND_net), .O(n3025));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1993_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i34640_3_lut (.I0(n2826), .I1(n2893), .I2(n2841), .I3(GND_net), 
            .O(n2925));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam i34640_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i34641_3_lut (.I0(n2925), .I1(n2992), .I2(n2940), .I3(GND_net), 
            .O(n3024));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam i34641_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1989_3_lut (.I0(n2922), .I1(n2989), 
            .I2(n2940), .I3(GND_net), .O(n3021));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1989_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1991_3_lut (.I0(n2924), .I1(n2991), 
            .I2(n2940), .I3(GND_net), .O(n3023));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1991_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1796 (.I0(n3023), .I1(n3021), .I2(n3024), .I3(n3025), 
            .O(n47119));
    defparam i1_4_lut_adj_1796.LUT_INIT = 16'hfffe;
    SB_CARRY encoder0_position_31__I_0_add_1302_7 (.CI(n38958), .I0(n1929), 
            .I1(GND_net), .CO(n38959));
    SB_LUT4 encoder0_position_31__I_0_add_1302_6_lut (.I0(GND_net), .I1(n1930), 
            .I2(GND_net), .I3(n38957), .O(n1997)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1302_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1302_6 (.CI(n38957), .I0(n1930), 
            .I1(GND_net), .CO(n38958));
    SB_LUT4 encoder0_position_31__I_0_add_1302_5_lut (.I0(GND_net), .I1(n1931), 
            .I2(VCC_net), .I3(n38956), .O(n1998)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1302_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1302_5 (.CI(n38956), .I0(n1931), 
            .I1(VCC_net), .CO(n38957));
    SB_LUT4 add_157_31_lut (.I0(GND_net), .I1(delay_counter[29]), .I2(GND_net), 
            .I3(n38474), .O(n1299)) /* synthesis syn_instantiated=1 */ ;
    defparam add_157_31_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1302_4_lut (.I0(GND_net), .I1(n1932), 
            .I2(GND_net), .I3(n38955), .O(n1999)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1302_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1302_4 (.CI(n38955), .I0(n1932), 
            .I1(GND_net), .CO(n38956));
    SB_DFF dti_counter_2244__i0 (.Q(dti_counter[0]), .C(CLK_c), .D(n55));   // verilog/TinyFPGA_B.v(175[23:37])
    SB_LUT4 add_157_10_lut (.I0(GND_net), .I1(delay_counter[8]), .I2(GND_net), 
            .I3(n38453), .O(n1320)) /* synthesis syn_instantiated=1 */ ;
    defparam add_157_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1302_3_lut (.I0(GND_net), .I1(n1933), 
            .I2(VCC_net), .I3(n38954), .O(n2000)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1302_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1302_3 (.CI(n38954), .I0(n1933), 
            .I1(VCC_net), .CO(n38955));
    SB_LUT4 encoder0_position_31__I_0_add_1302_2_lut (.I0(GND_net), .I1(n530), 
            .I2(GND_net), .I3(VCC_net), .O(n2001)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1302_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1302_2 (.CI(VCC_net), .I0(n530), 
            .I1(GND_net), .CO(n38954));
    SB_LUT4 encoder0_position_31__I_0_add_1235_18_lut (.I0(n50979), .I1(n1818), 
            .I2(VCC_net), .I3(n38953), .O(n1917)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1235_18_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_31__I_0_add_1235_17_lut (.I0(GND_net), .I1(n1819), 
            .I2(VCC_net), .I3(n38952), .O(n1886)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1235_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_33_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n2_adj_5411), .I3(n39523), .O(n2_adj_5313)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_33_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1235_17 (.CI(n38952), .I0(n1819), 
            .I1(VCC_net), .CO(n38953));
    SB_LUT4 i1_4_lut_adj_1797 (.I0(n3027), .I1(n3022), .I2(n3028), .I3(n3026), 
            .O(n47117));
    defparam i1_4_lut_adj_1797.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_31__I_0_add_1235_16_lut (.I0(GND_net), .I1(n1820), 
            .I2(VCC_net), .I3(n38951), .O(n1887)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1235_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1235_16 (.CI(n38951), .I0(n1820), 
            .I1(VCC_net), .CO(n38952));
    SB_LUT4 encoder0_position_31__I_0_add_1235_15_lut (.I0(GND_net), .I1(n1821), 
            .I2(VCC_net), .I3(n38950), .O(n1888)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1235_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1235_15 (.CI(n38950), .I0(n1821), 
            .I1(VCC_net), .CO(n38951));
    SB_LUT4 encoder0_position_31__I_0_add_1235_14_lut (.I0(GND_net), .I1(n1822), 
            .I2(VCC_net), .I3(n38949), .O(n1889)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1235_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1235_14 (.CI(n38949), .I0(n1822), 
            .I1(VCC_net), .CO(n38950));
    SB_LUT4 i1_3_lut_adj_1798 (.I0(n47119), .I1(n3019), .I2(n3020), .I3(GND_net), 
            .O(n47121));
    defparam i1_3_lut_adj_1798.LUT_INIT = 16'hfefe;
    SB_LUT4 i21446_3_lut (.I0(n541), .I1(n3032), .I2(n3033), .I3(GND_net), 
            .O(n35394));
    defparam i21446_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i1_4_lut_adj_1799 (.I0(n3017), .I1(n47121), .I2(n3018), .I3(n47117), 
            .O(n47127));
    defparam i1_4_lut_adj_1799.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1800 (.I0(n3029), .I1(n35394), .I2(n3030), .I3(n3031), 
            .O(n45056));
    defparam i1_4_lut_adj_1800.LUT_INIT = 16'ha080;
    SB_LUT4 i1_4_lut_adj_1801 (.I0(n3015), .I1(n3016), .I2(n45056), .I3(n47127), 
            .O(n47133));
    defparam i1_4_lut_adj_1801.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1802 (.I0(n3012), .I1(n3013), .I2(n3014), .I3(n47133), 
            .O(n47139));
    defparam i1_4_lut_adj_1802.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1803 (.I0(n3009), .I1(n3010), .I2(n3011), .I3(n47139), 
            .O(n47145));
    defparam i1_4_lut_adj_1803.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_31__I_0_add_1235_13_lut (.I0(GND_net), .I1(n1823), 
            .I2(VCC_net), .I3(n38948), .O(n1890)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1235_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1235_13 (.CI(n38948), .I0(n1823), 
            .I1(VCC_net), .CO(n38949));
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_32_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n3_adj_5412), .I3(n39522), .O(n3_adj_5312)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_32_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_32 (.CI(n39522), 
            .I0(GND_net), .I1(n3_adj_5412), .CO(n39523));
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_31_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n4_adj_5413), .I3(n39521), .O(n4_adj_5311)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_31_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_31 (.CI(n39521), 
            .I0(GND_net), .I1(n4_adj_5413), .CO(n39522));
    SB_LUT4 encoder0_position_31__I_0_add_1235_12_lut (.I0(GND_net), .I1(n1824), 
            .I2(VCC_net), .I3(n38947), .O(n1891_adj_5399)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1235_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1235_12 (.CI(n38947), .I0(n1824), 
            .I1(VCC_net), .CO(n38948));
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_30_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n5_adj_5414), .I3(n39520), .O(n5_adj_5310)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_30_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1235_11_lut (.I0(GND_net), .I1(n1825), 
            .I2(VCC_net), .I3(n38946), .O(n1892)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1235_11_lut.LUT_INIT = 16'hC33C;
    SB_DFF ID_i0_i0 (.Q(ID[0]), .C(CLK_c), .D(n29059));   // verilog/TinyFPGA_B.v(375[10] 403[6])
    SB_DFF commutation_state_prev_i2 (.Q(commutation_state_prev[2]), .C(CLK_c), 
           .D(commutation_state[2]));   // verilog/TinyFPGA_B.v(144[9] 223[5])
    SB_DFF commutation_state_prev_i1 (.Q(commutation_state_prev[1]), .C(CLK_c), 
           .D(commutation_state[1]));   // verilog/TinyFPGA_B.v(144[9] 223[5])
    SB_CARRY encoder0_position_31__I_0_add_1235_11 (.CI(n38946), .I0(n1825), 
            .I1(VCC_net), .CO(n38947));
    SB_DFF pwm_setpoint_i23 (.Q(pwm_setpoint[23]), .C(CLK_c), .D(pwm_setpoint_23__N_11[23]));   // verilog/TinyFPGA_B.v(104[9] 130[5])
    SB_DFF pwm_setpoint_i22 (.Q(pwm_setpoint[22]), .C(CLK_c), .D(pwm_setpoint_23__N_11[22]));   // verilog/TinyFPGA_B.v(104[9] 130[5])
    SB_DFF pwm_setpoint_i21 (.Q(pwm_setpoint[21]), .C(CLK_c), .D(pwm_setpoint_23__N_11[21]));   // verilog/TinyFPGA_B.v(104[9] 130[5])
    SB_DFF pwm_setpoint_i20 (.Q(pwm_setpoint[20]), .C(CLK_c), .D(pwm_setpoint_23__N_11[20]));   // verilog/TinyFPGA_B.v(104[9] 130[5])
    SB_DFF pwm_setpoint_i19 (.Q(pwm_setpoint[19]), .C(CLK_c), .D(pwm_setpoint_23__N_11[19]));   // verilog/TinyFPGA_B.v(104[9] 130[5])
    SB_DFF pwm_setpoint_i18 (.Q(pwm_setpoint[18]), .C(CLK_c), .D(pwm_setpoint_23__N_11[18]));   // verilog/TinyFPGA_B.v(104[9] 130[5])
    SB_DFF pwm_setpoint_i17 (.Q(pwm_setpoint[17]), .C(CLK_c), .D(pwm_setpoint_23__N_11[17]));   // verilog/TinyFPGA_B.v(104[9] 130[5])
    SB_DFF pwm_setpoint_i16 (.Q(pwm_setpoint[16]), .C(CLK_c), .D(pwm_setpoint_23__N_11[16]));   // verilog/TinyFPGA_B.v(104[9] 130[5])
    SB_DFF pwm_setpoint_i15 (.Q(pwm_setpoint[15]), .C(CLK_c), .D(pwm_setpoint_23__N_11[15]));   // verilog/TinyFPGA_B.v(104[9] 130[5])
    SB_DFF pwm_setpoint_i14 (.Q(pwm_setpoint[14]), .C(CLK_c), .D(pwm_setpoint_23__N_11[14]));   // verilog/TinyFPGA_B.v(104[9] 130[5])
    SB_DFF pwm_setpoint_i13 (.Q(pwm_setpoint[13]), .C(CLK_c), .D(pwm_setpoint_23__N_11[13]));   // verilog/TinyFPGA_B.v(104[9] 130[5])
    SB_DFF pwm_setpoint_i12 (.Q(pwm_setpoint[12]), .C(CLK_c), .D(pwm_setpoint_23__N_11[12]));   // verilog/TinyFPGA_B.v(104[9] 130[5])
    SB_DFF pwm_setpoint_i11 (.Q(pwm_setpoint[11]), .C(CLK_c), .D(pwm_setpoint_23__N_11[11]));   // verilog/TinyFPGA_B.v(104[9] 130[5])
    SB_DFF pwm_setpoint_i10 (.Q(pwm_setpoint[10]), .C(CLK_c), .D(pwm_setpoint_23__N_11[10]));   // verilog/TinyFPGA_B.v(104[9] 130[5])
    SB_DFF pwm_setpoint_i9 (.Q(pwm_setpoint[9]), .C(CLK_c), .D(pwm_setpoint_23__N_11[9]));   // verilog/TinyFPGA_B.v(104[9] 130[5])
    SB_DFF pwm_setpoint_i8 (.Q(pwm_setpoint[8]), .C(CLK_c), .D(pwm_setpoint_23__N_11[8]));   // verilog/TinyFPGA_B.v(104[9] 130[5])
    SB_DFF pwm_setpoint_i7 (.Q(pwm_setpoint[7]), .C(CLK_c), .D(pwm_setpoint_23__N_11[7]));   // verilog/TinyFPGA_B.v(104[9] 130[5])
    SB_DFF pwm_setpoint_i6 (.Q(pwm_setpoint[6]), .C(CLK_c), .D(pwm_setpoint_23__N_11[6]));   // verilog/TinyFPGA_B.v(104[9] 130[5])
    SB_DFF pwm_setpoint_i5 (.Q(pwm_setpoint[5]), .C(CLK_c), .D(pwm_setpoint_23__N_11[5]));   // verilog/TinyFPGA_B.v(104[9] 130[5])
    SB_DFF pwm_setpoint_i4 (.Q(pwm_setpoint[4]), .C(CLK_c), .D(pwm_setpoint_23__N_11[4]));   // verilog/TinyFPGA_B.v(104[9] 130[5])
    SB_DFF pwm_setpoint_i3 (.Q(pwm_setpoint[3]), .C(CLK_c), .D(pwm_setpoint_23__N_11[3]));   // verilog/TinyFPGA_B.v(104[9] 130[5])
    SB_DFF pwm_setpoint_i2 (.Q(pwm_setpoint[2]), .C(CLK_c), .D(pwm_setpoint_23__N_11[2]));   // verilog/TinyFPGA_B.v(104[9] 130[5])
    GND i1 (.Y(GND_net));
    SB_LUT4 n10621_bdd_4_lut_35724 (.I0(n10621), .I1(current[0]), .I2(duty[0]), 
            .I3(n4208), .O(n51330));
    defparam n10621_bdd_4_lut_35724.LUT_INIT = 16'he4aa;
    SB_LUT4 n51330_bdd_4_lut (.I0(n51330), .I1(n363), .I2(n4508), .I3(n4208), 
            .O(pwm_setpoint_23__N_11[0]));
    defparam n51330_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i35009_4_lut (.I0(n3007), .I1(n3006), .I2(n3008), .I3(n47145), 
            .O(n3039));
    defparam i35009_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 n51456_bdd_4_lut (.I0(n51456), .I1(n342), .I2(n4487), .I3(n4208), 
            .O(pwm_setpoint_23__N_11[21]));
    defparam n51456_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n10621_bdd_4_lut_35829 (.I0(n10621), .I1(current[15]), .I2(duty[21]), 
            .I3(n4208), .O(n51456));
    defparam n10621_bdd_4_lut_35829.LUT_INIT = 16'he4aa;
    SB_LUT4 encoder0_position_31__I_0_i1909_3_lut (.I0(n2810), .I1(n2877), 
            .I2(n2841), .I3(GND_net), .O(n2909));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1909_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1908_3_lut (.I0(n2809), .I1(n2876), 
            .I2(n2841), .I3(GND_net), .O(n2908));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1908_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1235_10_lut (.I0(GND_net), .I1(n1826), 
            .I2(VCC_net), .I3(n38945), .O(n1893)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1235_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1912_3_lut (.I0(n2813), .I1(n2880), 
            .I2(n2841), .I3(GND_net), .O(n2912));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1912_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1911_3_lut (.I0(n2812), .I1(n2879), 
            .I2(n2841), .I3(GND_net), .O(n2911));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1911_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1910_3_lut (.I0(n2811), .I1(n2878), 
            .I2(n2841), .I3(GND_net), .O(n2910));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1910_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1933_3_lut (.I0(n539), .I1(n2901), 
            .I2(n2841), .I3(GND_net), .O(n2933));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1933_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_1235_10 (.CI(n38945), .I0(n1826), 
            .I1(VCC_net), .CO(n38946));
    SB_LUT4 encoder0_position_31__I_0_i1932_3_lut (.I0(n2833), .I1(n2900), 
            .I2(n2841), .I3(GND_net), .O(n2932));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1932_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1931_3_lut (.I0(n2832), .I1(n2899), 
            .I2(n2841), .I3(GND_net), .O(n2931));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1931_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i5_3_lut (.I0(encoder0_position[4]), 
            .I1(n29), .I2(encoder0_position[31]), .I3(GND_net), .O(n540));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_mux_3_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i1923_3_lut (.I0(n2824), .I1(n2891), 
            .I2(n2841), .I3(GND_net), .O(n2923));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1923_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1919_3_lut (.I0(n2820), .I1(n2887), 
            .I2(n2841), .I3(GND_net), .O(n2919));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1919_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1928_3_lut (.I0(n2829), .I1(n2896), 
            .I2(n2841), .I3(GND_net), .O(n2928));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1928_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1921_3_lut (.I0(n2822), .I1(n2889), 
            .I2(n2841), .I3(GND_net), .O(n2921));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1921_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1922_3_lut (.I0(n2823), .I1(n2890), 
            .I2(n2841), .I3(GND_net), .O(n2922));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1922_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1915_3_lut (.I0(n2816), .I1(n2883), 
            .I2(n2841), .I3(GND_net), .O(n2915));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1915_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1914_3_lut (.I0(n2815), .I1(n2882), 
            .I2(n2841), .I3(GND_net), .O(n2914));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1914_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1913_3_lut (.I0(n2814), .I1(n2881), 
            .I2(n2841), .I3(GND_net), .O(n2913));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1913_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1930_3_lut (.I0(n2831), .I1(n2898), 
            .I2(n2841), .I3(GND_net), .O(n2930));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1930_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1929_3_lut (.I0(n2830), .I1(n2897), 
            .I2(n2841), .I3(GND_net), .O(n2929));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1929_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1918_3_lut (.I0(n2819), .I1(n2886), 
            .I2(n2841), .I3(GND_net), .O(n2918));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1918_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1917_3_lut (.I0(n2818), .I1(n2885), 
            .I2(n2841), .I3(GND_net), .O(n2917));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1917_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1916_3_lut (.I0(n2817), .I1(n2884), 
            .I2(n2841), .I3(GND_net), .O(n2916));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1916_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1926_3_lut (.I0(n2827), .I1(n2894), 
            .I2(n2841), .I3(GND_net), .O(n2926));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1926_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1920_3_lut (.I0(n2821), .I1(n2888), 
            .I2(n2841), .I3(GND_net), .O(n2920));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1920_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1927_3_lut (.I0(n2828), .I1(n2895), 
            .I2(n2841), .I3(GND_net), .O(n2927));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1927_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1924_3_lut (.I0(n2825), .I1(n2892), 
            .I2(n2841), .I3(GND_net), .O(n2924));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1924_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1804 (.I0(n2924), .I1(n2927), .I2(n2920), .I3(n2926), 
            .O(n46677));
    defparam i1_4_lut_adj_1804.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1805 (.I0(n2925), .I1(n2922), .I2(n2921), .I3(n2928), 
            .O(n46679));
    defparam i1_4_lut_adj_1805.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1806 (.I0(n46679), .I1(n46677), .I2(n2919), .I3(n2923), 
            .O(n46683));
    defparam i1_4_lut_adj_1806.LUT_INIT = 16'hfffe;
    SB_LUT4 i21507_4_lut (.I0(n540), .I1(n2931), .I2(n2932), .I3(n2933), 
            .O(n35456));
    defparam i21507_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 i1_4_lut_adj_1807 (.I0(n2916), .I1(n2917), .I2(n46683), .I3(n2918), 
            .O(n46689));
    defparam i1_4_lut_adj_1807.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1808 (.I0(n46689), .I1(n2929), .I2(n35456), .I3(n2930), 
            .O(n46691));
    defparam i1_4_lut_adj_1808.LUT_INIT = 16'heaaa;
    SB_LUT4 i1_4_lut_adj_1809 (.I0(n2913), .I1(n2914), .I2(n2915), .I3(n46691), 
            .O(n46697));
    defparam i1_4_lut_adj_1809.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1810 (.I0(n2910), .I1(n2911), .I2(n2912), .I3(n46697), 
            .O(n46703));
    defparam i1_4_lut_adj_1810.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_31__I_0_add_1235_9_lut (.I0(GND_net), .I1(n1827), 
            .I2(VCC_net), .I3(n38944), .O(n1894)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1235_9_lut.LUT_INIT = 16'hC33C;
    SB_DFFESR delay_counter_i0_i1 (.Q(delay_counter[1]), .C(CLK_c), .E(n7417), 
            .D(n1327), .R(n28933));   // verilog/TinyFPGA_B.v(375[10] 403[6])
    SB_DFFESR delay_counter_i0_i2 (.Q(delay_counter[2]), .C(CLK_c), .E(n7417), 
            .D(n1326), .R(n28933));   // verilog/TinyFPGA_B.v(375[10] 403[6])
    SB_CARRY encoder0_position_31__I_0_add_1235_9 (.CI(n38944), .I0(n1827), 
            .I1(VCC_net), .CO(n38945));
    SB_LUT4 encoder0_position_31__I_0_add_1235_8_lut (.I0(GND_net), .I1(n1828), 
            .I2(VCC_net), .I3(n38943), .O(n1895)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1235_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1235_8 (.CI(n38943), .I0(n1828), 
            .I1(VCC_net), .CO(n38944));
    SB_LUT4 encoder0_position_31__I_0_add_1235_7_lut (.I0(GND_net), .I1(n1829), 
            .I2(GND_net), .I3(n38942), .O(n1896_adj_5400)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1235_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1235_7 (.CI(n38942), .I0(n1829), 
            .I1(GND_net), .CO(n38943));
    SB_LUT4 encoder0_position_31__I_0_add_1235_6_lut (.I0(GND_net), .I1(n1830), 
            .I2(GND_net), .I3(n38941), .O(n1897)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1235_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1235_6 (.CI(n38941), .I0(n1830), 
            .I1(GND_net), .CO(n38942));
    SB_LUT4 encoder0_position_31__I_0_add_1235_5_lut (.I0(GND_net), .I1(n1831), 
            .I2(VCC_net), .I3(n38940), .O(n1898)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1235_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1235_5 (.CI(n38940), .I0(n1831), 
            .I1(VCC_net), .CO(n38941));
    SB_LUT4 encoder0_position_31__I_0_add_1235_4_lut (.I0(GND_net), .I1(n1832), 
            .I2(GND_net), .I3(n38939), .O(n1899)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1235_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1235_4 (.CI(n38939), .I0(n1832), 
            .I1(GND_net), .CO(n38940));
    SB_LUT4 encoder0_position_31__I_0_add_1235_3_lut (.I0(GND_net), .I1(n1833), 
            .I2(VCC_net), .I3(n38938), .O(n1900)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1235_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i35051_4_lut (.I0(n2908), .I1(n2907), .I2(n2909), .I3(n46703), 
            .O(n2940));
    defparam i35051_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_31__I_0_i1842_3_lut (.I0(n2711), .I1(n2778), 
            .I2(n2742), .I3(GND_net), .O(n2810));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1842_3_lut.LUT_INIT = 16'hacac;
    SB_DFFESR delay_counter_i0_i3 (.Q(delay_counter[3]), .C(CLK_c), .E(n7417), 
            .D(n1325), .R(n28933));   // verilog/TinyFPGA_B.v(375[10] 403[6])
    SB_LUT4 i15101_3_lut (.I0(\data_out_frame[12] [3]), .I1(setpoint[19]), 
            .I2(n24278), .I3(GND_net), .O(n29049));   // verilog/coms.v(128[12] 303[6])
    defparam i15101_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i1840_3_lut (.I0(n2709), .I1(n2776), 
            .I2(n2742), .I3(GND_net), .O(n2808));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1840_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1841_3_lut (.I0(n2710), .I1(n2777), 
            .I2(n2742), .I3(GND_net), .O(n2809));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1841_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1845_3_lut (.I0(n2714), .I1(n2781), 
            .I2(n2742), .I3(GND_net), .O(n2813));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1845_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1844_3_lut (.I0(n2713), .I1(n2780), 
            .I2(n2742), .I3(GND_net), .O(n2812));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1844_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15102_3_lut (.I0(\data_out_frame[12] [2]), .I1(setpoint[18]), 
            .I2(n24278), .I3(GND_net), .O(n29050));   // verilog/coms.v(128[12] 303[6])
    defparam i15102_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i1843_3_lut (.I0(n2712), .I1(n2779), 
            .I2(n2742), .I3(GND_net), .O(n2811));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1843_3_lut.LUT_INIT = 16'hacac;
    SB_DFFESR delay_counter_i0_i4 (.Q(delay_counter[4]), .C(CLK_c), .E(n7417), 
            .D(n1324), .R(n28933));   // verilog/TinyFPGA_B.v(375[10] 403[6])
    SB_CARRY encoder0_position_31__I_0_add_1235_3 (.CI(n38938), .I0(n1833), 
            .I1(VCC_net), .CO(n38939));
    SB_LUT4 encoder0_position_31__I_0_add_1235_2_lut (.I0(GND_net), .I1(n529), 
            .I2(GND_net), .I3(VCC_net), .O(n1901)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1235_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1235_2 (.CI(VCC_net), .I0(n529), 
            .I1(GND_net), .CO(n38938));
    SB_LUT4 encoder0_position_31__I_0_add_1168_17_lut (.I0(n50999), .I1(n1719), 
            .I2(VCC_net), .I3(n38937), .O(n1818)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1168_17_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_31__I_0_add_1168_16_lut (.I0(GND_net), .I1(n1720), 
            .I2(VCC_net), .I3(n38936), .O(n1787)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1168_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1168_16 (.CI(n38936), .I0(n1720), 
            .I1(VCC_net), .CO(n38937));
    SB_LUT4 encoder0_position_31__I_0_add_1168_15_lut (.I0(GND_net), .I1(n1721), 
            .I2(VCC_net), .I3(n38935), .O(n1788)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1168_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1168_15 (.CI(n38935), .I0(n1721), 
            .I1(VCC_net), .CO(n38936));
    SB_LUT4 encoder0_position_31__I_0_add_1168_14_lut (.I0(GND_net), .I1(n1722), 
            .I2(VCC_net), .I3(n38934), .O(n1789)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1168_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1168_14 (.CI(n38934), .I0(n1722), 
            .I1(VCC_net), .CO(n38935));
    SB_LUT4 encoder0_position_31__I_0_add_1168_13_lut (.I0(GND_net), .I1(n1723), 
            .I2(VCC_net), .I3(n38933), .O(n1790)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1168_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1168_13 (.CI(n38933), .I0(n1723), 
            .I1(VCC_net), .CO(n38934));
    SB_IO NEOPXL_pad (.PACKAGE_PIN(NEOPXL), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(NEOPXL_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam NEOPXL_pad.PIN_TYPE = 6'b011001;
    defparam NEOPXL_pad.PULLUP = 1'b0;
    defparam NEOPXL_pad.NEG_TRIGGER = 1'b0;
    defparam NEOPXL_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO USBPU_pad (.PACKAGE_PIN(USBPU), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(GND_net));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam USBPU_pad.PIN_TYPE = 6'b011001;
    defparam USBPU_pad.PULLUP = 1'b0;
    defparam USBPU_pad.NEG_TRIGGER = 1'b0;
    defparam USBPU_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 encoder0_position_31__I_0_add_1168_12_lut (.I0(GND_net), .I1(n1724), 
            .I2(VCC_net), .I3(n38932), .O(n1791)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1168_12_lut.LUT_INIT = 16'hC33C;
    SB_IO LED_pad (.PACKAGE_PIN(LED), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(LED_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam LED_pad.PIN_TYPE = 6'b011001;
    defparam LED_pad.PULLUP = 1'b0;
    defparam LED_pad.NEG_TRIGGER = 1'b0;
    defparam LED_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 encoder0_position_31__I_0_i1848_3_lut (.I0(n2717), .I1(n2784), 
            .I2(n2742), .I3(GND_net), .O(n2816));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1848_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1847_3_lut (.I0(n2716), .I1(n2783), 
            .I2(n2742), .I3(GND_net), .O(n2815));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1847_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1846_3_lut (.I0(n2715), .I1(n2782), 
            .I2(n2742), .I3(GND_net), .O(n2814));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1846_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_1168_12 (.CI(n38932), .I0(n1724), 
            .I1(VCC_net), .CO(n38933));
    SB_LUT4 encoder0_position_31__I_0_add_1168_11_lut (.I0(GND_net), .I1(n1725), 
            .I2(VCC_net), .I3(n38931), .O(n1792)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1168_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1168_11 (.CI(n38931), .I0(n1725), 
            .I1(VCC_net), .CO(n38932));
    SB_LUT4 encoder0_position_31__I_0_add_1168_10_lut (.I0(GND_net), .I1(n1726), 
            .I2(VCC_net), .I3(n38930), .O(n1793)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1168_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1168_10 (.CI(n38930), .I0(n1726), 
            .I1(VCC_net), .CO(n38931));
    SB_LUT4 encoder0_position_31__I_0_add_1168_9_lut (.I0(GND_net), .I1(n1727), 
            .I2(VCC_net), .I3(n38929), .O(n1794)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1168_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1168_9 (.CI(n38929), .I0(n1727), 
            .I1(VCC_net), .CO(n38930));
    SB_LUT4 encoder0_position_31__I_0_add_1168_8_lut (.I0(GND_net), .I1(n1728), 
            .I2(VCC_net), .I3(n38928), .O(n1795)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1168_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1168_8 (.CI(n38928), .I0(n1728), 
            .I1(VCC_net), .CO(n38929));
    SB_LUT4 i15103_3_lut (.I0(current[0]), .I1(data_adj_5514[0]), .I2(n28537), 
            .I3(GND_net), .O(n29051));   // verilog/tli4970.v(35[10] 68[6])
    defparam i15103_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_add_1168_7_lut (.I0(GND_net), .I1(n1729), 
            .I2(GND_net), .I3(n38927), .O(n1796)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1168_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1168_7 (.CI(n38927), .I0(n1729), 
            .I1(GND_net), .CO(n38928));
    SB_LUT4 encoder0_position_31__I_0_add_1168_6_lut (.I0(GND_net), .I1(n1730), 
            .I2(GND_net), .I3(n38926), .O(n1797)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1168_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1862_3_lut (.I0(n2731), .I1(n2798), 
            .I2(n2742), .I3(GND_net), .O(n2830));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1862_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1861_3_lut (.I0(n2730), .I1(n2797), 
            .I2(n2742), .I3(GND_net), .O(n2829));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1861_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1851_3_lut (.I0(n2720), .I1(n2787), 
            .I2(n2742), .I3(GND_net), .O(n2819));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1851_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_30 (.CI(n39520), 
            .I0(GND_net), .I1(n5_adj_5414), .CO(n39521));
    SB_LUT4 encoder0_position_31__I_0_i1850_3_lut (.I0(n2719), .I1(n2786), 
            .I2(n2742), .I3(GND_net), .O(n2818));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1850_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_1168_6 (.CI(n38926), .I0(n1730), 
            .I1(GND_net), .CO(n38927));
    SB_LUT4 i15104_4_lut (.I0(CS_MISO_c), .I1(data_adj_5514[1]), .I2(n10_adj_5341), 
            .I3(n27167), .O(n29052));   // verilog/tli4970.v(35[10] 68[6])
    defparam i15104_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i1_4_lut_adj_1811 (.I0(enable_slow_N_4354), .I1(data_ready), 
            .I2(state_adj_5510[1]), .I3(state_adj_5510[0]), .O(n43506));   // verilog/eeprom.v(26[8] 58[4])
    defparam i1_4_lut_adj_1811.LUT_INIT = 16'hccd0;
    SB_LUT4 i15106_4_lut (.I0(rw), .I1(state_adj_5510[0]), .I2(state_adj_5510[1]), 
            .I3(n6130), .O(n29054));   // verilog/eeprom.v(26[8] 58[4])
    defparam i15106_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 encoder0_position_31__I_0_add_1168_5_lut (.I0(GND_net), .I1(n1731), 
            .I2(VCC_net), .I3(n38925), .O(n1798)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1168_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1849_3_lut (.I0(n2718), .I1(n2785), 
            .I2(n2742), .I3(GND_net), .O(n2817));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1849_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_1168_5 (.CI(n38925), .I0(n1731), 
            .I1(VCC_net), .CO(n38926));
    SB_LUT4 encoder0_position_31__I_0_add_1168_4_lut (.I0(GND_net), .I1(n1732), 
            .I2(GND_net), .I3(n38924), .O(n1799)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1168_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15107_3_lut (.I0(\data_out_frame[12] [1]), .I1(setpoint[17]), 
            .I2(n24278), .I3(GND_net), .O(n29055));   // verilog/coms.v(128[12] 303[6])
    defparam i15107_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i1854_3_lut (.I0(n2723), .I1(n2790), 
            .I2(n2742), .I3(GND_net), .O(n2822));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1854_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1855_3_lut (.I0(n2724), .I1(n2791), 
            .I2(n2742), .I3(GND_net), .O(n2823));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1855_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15647_3_lut (.I0(control_mode[5]), .I1(\data_in_frame[1] [5]), 
            .I2(n28521), .I3(GND_net), .O(n29595));   // verilog/coms.v(128[12] 303[6])
    defparam i15647_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_31__I_0_add_1168_4 (.CI(n38924), .I0(n1732), 
            .I1(GND_net), .CO(n38925));
    SB_LUT4 encoder0_position_31__I_0_i1865_3_lut (.I0(n538), .I1(n2801), 
            .I2(n2742), .I3(GND_net), .O(n2833));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1865_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1864_3_lut (.I0(n2733), .I1(n2800), 
            .I2(n2742), .I3(GND_net), .O(n2832));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1864_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1863_3_lut (.I0(n2732), .I1(n2799), 
            .I2(n2742), .I3(GND_net), .O(n2831));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1863_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i6_3_lut (.I0(encoder0_position[5]), 
            .I1(n28), .I2(encoder0_position[31]), .I3(GND_net), .O(n539));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_mux_3_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i1856_rep_15_3_lut (.I0(n2725), .I1(n2792), 
            .I2(n2742), .I3(GND_net), .O(n2824));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1856_rep_15_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15648_3_lut (.I0(control_mode[4]), .I1(\data_in_frame[1] [4]), 
            .I2(n28521), .I3(GND_net), .O(n29596));   // verilog/coms.v(128[12] 303[6])
    defparam i15648_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i1853_rep_14_3_lut (.I0(n2722), .I1(n2789), 
            .I2(n2742), .I3(GND_net), .O(n2821));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1853_rep_14_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1168_3_lut (.I0(GND_net), .I1(n1733), 
            .I2(VCC_net), .I3(n38923), .O(n1800)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1168_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1168_3 (.CI(n38923), .I0(n1733), 
            .I1(VCC_net), .CO(n38924));
    SB_LUT4 encoder0_position_31__I_0_add_1168_2_lut (.I0(GND_net), .I1(n528), 
            .I2(GND_net), .I3(VCC_net), .O(n1801)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1168_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1168_2 (.CI(VCC_net), .I0(n528), 
            .I1(GND_net), .CO(n38923));
    SB_LUT4 encoder0_position_31__I_0_i1859_3_lut (.I0(n2728), .I1(n2795), 
            .I2(n2742), .I3(GND_net), .O(n2827));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1859_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1858_rep_12_3_lut (.I0(n2727), .I1(n2794), 
            .I2(n2742), .I3(GND_net), .O(n2826));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1858_rep_12_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1857_3_lut (.I0(n2726), .I1(n2793), 
            .I2(n2742), .I3(GND_net), .O(n2825));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1857_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1852_3_lut (.I0(n2721), .I1(n2788), 
            .I2(n2742), .I3(GND_net), .O(n2820));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1852_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15649_3_lut (.I0(control_mode[3]), .I1(\data_in_frame[1] [3]), 
            .I2(n28521), .I3(GND_net), .O(n29597));   // verilog/coms.v(128[12] 303[6])
    defparam i15649_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i1860_3_lut (.I0(n2729), .I1(n2796), 
            .I2(n2742), .I3(GND_net), .O(n2828));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1860_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1101_16_lut (.I0(n51018), .I1(n1620), 
            .I2(VCC_net), .I3(n38922), .O(n1719)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1101_16_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i15650_3_lut (.I0(control_mode[2]), .I1(\data_in_frame[1] [2]), 
            .I2(n28521), .I3(GND_net), .O(n29598));   // verilog/coms.v(128[12] 303[6])
    defparam i15650_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut_adj_1812 (.I0(n2828), .I1(n2820), .I2(n2825), .I3(GND_net), 
            .O(n47069));
    defparam i1_3_lut_adj_1812.LUT_INIT = 16'hfefe;
    SB_LUT4 encoder0_position_31__I_0_add_1101_15_lut (.I0(GND_net), .I1(n1621), 
            .I2(VCC_net), .I3(n38921), .O(n1688)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1101_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1101_15 (.CI(n38921), .I0(n1621), 
            .I1(VCC_net), .CO(n38922));
    SB_LUT4 encoder0_position_31__I_0_add_1101_14_lut (.I0(GND_net), .I1(n1622), 
            .I2(VCC_net), .I3(n38920), .O(n1689)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1101_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1101_14 (.CI(n38920), .I0(n1622), 
            .I1(VCC_net), .CO(n38921));
    SB_LUT4 i1_4_lut_adj_1813 (.I0(n2826), .I1(n2827), .I2(n2821), .I3(n2824), 
            .O(n47071));
    defparam i1_4_lut_adj_1813.LUT_INIT = 16'hfffe;
    SB_LUT4 i15651_3_lut (.I0(control_mode[1]), .I1(\data_in_frame[1] [1]), 
            .I2(n28521), .I3(GND_net), .O(n29599));   // verilog/coms.v(128[12] 303[6])
    defparam i15651_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1814 (.I0(n47071), .I1(n47069), .I2(n2823), .I3(n2822), 
            .O(n47075));
    defparam i1_4_lut_adj_1814.LUT_INIT = 16'hfffe;
    SB_LUT4 i21509_4_lut (.I0(n539), .I1(n2831), .I2(n2832), .I3(n2833), 
            .O(n35458));
    defparam i21509_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 encoder0_position_31__I_0_add_1101_13_lut (.I0(GND_net), .I1(n1623), 
            .I2(VCC_net), .I3(n38919), .O(n1690)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1101_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1101_13 (.CI(n38919), .I0(n1623), 
            .I1(VCC_net), .CO(n38920));
    SB_LUT4 encoder0_position_31__I_0_add_1101_12_lut (.I0(GND_net), .I1(n1624), 
            .I2(VCC_net), .I3(n38918), .O(n1691)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1101_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1101_12 (.CI(n38918), .I0(n1624), 
            .I1(VCC_net), .CO(n38919));
    SB_LUT4 i1_4_lut_adj_1815 (.I0(n2817), .I1(n2818), .I2(n47075), .I3(n2819), 
            .O(n47081));
    defparam i1_4_lut_adj_1815.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1816 (.I0(n47081), .I1(n2829), .I2(n35458), .I3(n2830), 
            .O(n47083));
    defparam i1_4_lut_adj_1816.LUT_INIT = 16'heaaa;
    SB_LUT4 i1_4_lut_adj_1817 (.I0(n2814), .I1(n2815), .I2(n2816), .I3(n47083), 
            .O(n47089));
    defparam i1_4_lut_adj_1817.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1818 (.I0(n2811), .I1(n2812), .I2(n2813), .I3(n47089), 
            .O(n47095));
    defparam i1_4_lut_adj_1818.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_31__I_0_add_1101_11_lut (.I0(GND_net), .I1(n1625), 
            .I2(VCC_net), .I3(n38917), .O(n1692)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1101_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i35083_4_lut (.I0(n2809), .I1(n2808), .I2(n2810), .I3(n47095), 
            .O(n2841));
    defparam i35083_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_31__I_0_i1775_3_lut (.I0(n2612), .I1(n2679), 
            .I2(n2643), .I3(GND_net), .O(n2711));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1775_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1785_3_lut (.I0(n2622), .I1(n2689), 
            .I2(n2643), .I3(GND_net), .O(n2721));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1785_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_1101_11 (.CI(n38917), .I0(n1625), 
            .I1(VCC_net), .CO(n38918));
    SB_LUT4 encoder0_position_31__I_0_add_1101_10_lut (.I0(GND_net), .I1(n1626), 
            .I2(VCC_net), .I3(n38916), .O(n1693)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1101_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1101_10 (.CI(n38916), .I0(n1626), 
            .I1(VCC_net), .CO(n38917));
    SB_LUT4 encoder0_position_31__I_0_add_1101_9_lut (.I0(GND_net), .I1(n1627), 
            .I2(VCC_net), .I3(n38915), .O(n1694)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1101_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1101_9 (.CI(n38915), .I0(n1627), 
            .I1(VCC_net), .CO(n38916));
    SB_LUT4 encoder0_position_31__I_0_add_1101_8_lut (.I0(GND_net), .I1(n1628), 
            .I2(VCC_net), .I3(n38914), .O(n1695)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1101_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15654_3_lut (.I0(\data_out_frame[22] [6]), .I1(current[6]), 
            .I2(n24278), .I3(GND_net), .O(n29602));   // verilog/coms.v(128[12] 303[6])
    defparam i15654_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i1783_3_lut (.I0(n2620), .I1(n2687), 
            .I2(n2643), .I3(GND_net), .O(n2719));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1783_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_1005_i14_3_lut (.I0(duty[13]), .I1(n350), .I2(duty[23]), 
            .I3(GND_net), .O(n4710));   // verilog/TinyFPGA_B.v(118[13] 129[7])
    defparam mux_1005_i14_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i1774_3_lut (.I0(n2611), .I1(n2678), 
            .I2(n2643), .I3(GND_net), .O(n2710));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1774_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_1101_8 (.CI(n38914), .I0(n1628), 
            .I1(VCC_net), .CO(n38915));
    SB_LUT4 encoder0_position_31__I_0_add_1101_7_lut (.I0(GND_net), .I1(n1629), 
            .I2(GND_net), .I3(n38913), .O(n1696)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1101_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1101_7 (.CI(n38913), .I0(n1629), 
            .I1(GND_net), .CO(n38914));
    SB_LUT4 encoder0_position_31__I_0_add_1101_6_lut (.I0(GND_net), .I1(n1630), 
            .I2(GND_net), .I3(n38912), .O(n1697)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1101_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1776_3_lut (.I0(n2613), .I1(n2680), 
            .I2(n2643), .I3(GND_net), .O(n2712));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1776_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1779_3_lut (.I0(n2616), .I1(n2683), 
            .I2(n2643), .I3(GND_net), .O(n2715));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1779_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1778_3_lut (.I0(n2615), .I1(n2682), 
            .I2(n2643), .I3(GND_net), .O(n2714));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1778_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_1101_6 (.CI(n38912), .I0(n1630), 
            .I1(GND_net), .CO(n38913));
    SB_LUT4 encoder0_position_31__I_0_i1777_3_lut (.I0(n2614), .I1(n2681), 
            .I2(n2643), .I3(GND_net), .O(n2713));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1777_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1101_5_lut (.I0(GND_net), .I1(n1631), 
            .I2(VCC_net), .I3(n38911), .O(n1698)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1101_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1101_5 (.CI(n38911), .I0(n1631), 
            .I1(VCC_net), .CO(n38912));
    SB_LUT4 encoder0_position_31__I_0_add_1101_4_lut (.I0(GND_net), .I1(n1632), 
            .I2(GND_net), .I3(n38910), .O(n1699)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1101_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_29_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n6_adj_5415), .I3(n39519), .O(n6_adj_5309)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_29_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1787_3_lut (.I0(n2624), .I1(n2691), 
            .I2(n2643), .I3(GND_net), .O(n2723));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1787_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1791_3_lut (.I0(n2628), .I1(n2695), 
            .I2(n2643), .I3(GND_net), .O(n2727));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1791_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_1101_4 (.CI(n38910), .I0(n1632), 
            .I1(GND_net), .CO(n38911));
    SB_LUT4 encoder0_position_31__I_0_add_1101_3_lut (.I0(GND_net), .I1(n1633), 
            .I2(VCC_net), .I3(n38909), .O(n1700)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1101_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1101_3 (.CI(n38909), .I0(n1633), 
            .I1(VCC_net), .CO(n38910));
    SB_LUT4 encoder0_position_31__I_0_add_1101_2_lut (.I0(GND_net), .I1(n527), 
            .I2(GND_net), .I3(VCC_net), .O(n1701)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1101_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15656_3_lut (.I0(\data_out_frame[22] [5]), .I1(current[5]), 
            .I2(n24278), .I3(GND_net), .O(n29604));   // verilog/coms.v(128[12] 303[6])
    defparam i15656_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i1780_3_lut (.I0(n2617), .I1(n2684), 
            .I2(n2643), .I3(GND_net), .O(n2716));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1780_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_1101_2 (.CI(VCC_net), .I0(n527), 
            .I1(GND_net), .CO(n38909));
    SB_LUT4 encoder0_position_31__I_0_add_1034_15_lut (.I0(n51036), .I1(n1521), 
            .I2(VCC_net), .I3(n38908), .O(n1620)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1034_15_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_31__I_0_add_1034_14_lut (.I0(GND_net), .I1(n1522), 
            .I2(VCC_net), .I3(n38907), .O(n1589)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1034_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1034_14 (.CI(n38907), .I0(n1522), 
            .I1(VCC_net), .CO(n38908));
    SB_LUT4 i15657_3_lut (.I0(\data_out_frame[22] [4]), .I1(current[4]), 
            .I2(n24278), .I3(GND_net), .O(n29605));   // verilog/coms.v(128[12] 303[6])
    defparam i15657_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15658_3_lut (.I0(\data_out_frame[22] [3]), .I1(current[3]), 
            .I2(n24278), .I3(GND_net), .O(n29606));   // verilog/coms.v(128[12] 303[6])
    defparam i15658_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_add_1034_13_lut (.I0(GND_net), .I1(n1523), 
            .I2(VCC_net), .I3(n38906), .O(n1590)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1034_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1034_13 (.CI(n38906), .I0(n1523), 
            .I1(VCC_net), .CO(n38907));
    SB_LUT4 encoder0_position_31__I_0_add_1034_12_lut (.I0(GND_net), .I1(n1524), 
            .I2(VCC_net), .I3(n38905), .O(n1591)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1034_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1034_12 (.CI(n38905), .I0(n1524), 
            .I1(VCC_net), .CO(n38906));
    SB_LUT4 i15659_3_lut (.I0(\data_out_frame[22] [2]), .I1(current[2]), 
            .I2(n24278), .I3(GND_net), .O(n29607));   // verilog/coms.v(128[12] 303[6])
    defparam i15659_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15660_3_lut (.I0(\data_out_frame[22] [1]), .I1(current[1]), 
            .I2(n24278), .I3(GND_net), .O(n29608));   // verilog/coms.v(128[12] 303[6])
    defparam i15660_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i1781_3_lut (.I0(n2618), .I1(n2685), 
            .I2(n2643), .I3(GND_net), .O(n2717));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1781_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1782_3_lut (.I0(n2619), .I1(n2686), 
            .I2(n2643), .I3(GND_net), .O(n2718));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1782_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1034_11_lut (.I0(GND_net), .I1(n1525), 
            .I2(VCC_net), .I3(n38904), .O(n1592)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1034_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1034_11 (.CI(n38904), .I0(n1525), 
            .I1(VCC_net), .CO(n38905));
    SB_LUT4 encoder0_position_31__I_0_add_1034_10_lut (.I0(GND_net), .I1(n1526), 
            .I2(VCC_net), .I3(n38903), .O(n1593)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1034_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1034_10 (.CI(n38903), .I0(n1526), 
            .I1(VCC_net), .CO(n38904));
    SB_LUT4 encoder0_position_31__I_0_i1788_3_lut (.I0(n2625), .I1(n2692), 
            .I2(n2643), .I3(GND_net), .O(n2724));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1788_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1786_3_lut (.I0(n2623), .I1(n2690), 
            .I2(n2643), .I3(GND_net), .O(n2722));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1786_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1792_3_lut (.I0(n2629), .I1(n2696), 
            .I2(n2643), .I3(GND_net), .O(n2728));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1792_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15661_3_lut (.I0(\data_out_frame[22] [0]), .I1(current[0]), 
            .I2(n24278), .I3(GND_net), .O(n29609));   // verilog/coms.v(128[12] 303[6])
    defparam i15661_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i1790_3_lut (.I0(n2627), .I1(n2694), 
            .I2(n2643), .I3(GND_net), .O(n2726));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1790_3_lut.LUT_INIT = 16'hacac;
    SB_DFFESR GHC_196 (.Q(GHC), .C(CLK_c), .E(n28482), .D(GHC_N_427), 
            .R(n28835));   // verilog/TinyFPGA_B.v(144[9] 223[5])
    SB_LUT4 encoder0_position_31__I_0_i1789_3_lut (.I0(n2626), .I1(n2693), 
            .I2(n2643), .I3(GND_net), .O(n2725));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1789_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1034_9_lut (.I0(GND_net), .I1(n1527), 
            .I2(VCC_net), .I3(n38902), .O(n1594)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1034_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1034_9 (.CI(n38902), .I0(n1527), 
            .I1(VCC_net), .CO(n38903));
    SB_LUT4 encoder0_position_31__I_0_add_1034_8_lut (.I0(GND_net), .I1(n1528), 
            .I2(VCC_net), .I3(n38901), .O(n1595)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1034_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1034_8 (.CI(n38901), .I0(n1528), 
            .I1(VCC_net), .CO(n38902));
    SB_LUT4 encoder0_position_31__I_0_i1784_3_lut (.I0(n2621), .I1(n2688), 
            .I2(n2643), .I3(GND_net), .O(n2720));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1784_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1795_3_lut (.I0(n2632), .I1(n2699), 
            .I2(n2643), .I3(GND_net), .O(n2731));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1795_3_lut.LUT_INIT = 16'hacac;
    SB_DFFESR GHB_194 (.Q(GHB), .C(CLK_c), .E(n28482), .D(GHB_N_413), 
            .R(n28835));   // verilog/TinyFPGA_B.v(144[9] 223[5])
    SB_LUT4 encoder0_position_31__I_0_i1794_3_lut (.I0(n2631), .I1(n2698), 
            .I2(n2643), .I3(GND_net), .O(n2730));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1794_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1034_7_lut (.I0(GND_net), .I1(n1529), 
            .I2(GND_net), .I3(n38900), .O(n1596)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1034_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1034_7 (.CI(n38900), .I0(n1529), 
            .I1(GND_net), .CO(n38901));
    SB_LUT4 encoder0_position_31__I_0_add_1034_6_lut (.I0(GND_net), .I1(n1530), 
            .I2(GND_net), .I3(n38899), .O(n1597)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1034_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1034_6 (.CI(n38899), .I0(n1530), 
            .I1(GND_net), .CO(n38900));
    SB_LUT4 encoder0_position_31__I_0_i1793_3_lut (.I0(n2630), .I1(n2697), 
            .I2(n2643), .I3(GND_net), .O(n2729));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1793_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1797_3_lut (.I0(n537), .I1(n2701), 
            .I2(n2643), .I3(GND_net), .O(n2733));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1797_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 unary_minus_19_inv_0_i5_1_lut (.I0(duty[4]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_5266));   // verilog/TinyFPGA_B.v(123[25:30])
    defparam unary_minus_19_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_add_1034_5_lut (.I0(GND_net), .I1(n1531), 
            .I2(VCC_net), .I3(n38898), .O(n1598)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1034_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1034_5 (.CI(n38898), .I0(n1531), 
            .I1(VCC_net), .CO(n38899));
    SB_LUT4 encoder0_position_31__I_0_add_1034_4_lut (.I0(GND_net), .I1(n1532), 
            .I2(GND_net), .I3(n38897), .O(n1599)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1034_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1034_4 (.CI(n38897), .I0(n1532), 
            .I1(GND_net), .CO(n38898));
    SB_LUT4 i15662_3_lut (.I0(\data_out_frame[21] [7]), .I1(current[15]), 
            .I2(n24278), .I3(GND_net), .O(n29610));   // verilog/coms.v(128[12] 303[6])
    defparam i15662_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i1796_3_lut (.I0(n2633), .I1(n2700), 
            .I2(n2643), .I3(GND_net), .O(n2732));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1796_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i7_3_lut (.I0(encoder0_position[6]), 
            .I1(n27), .I2(encoder0_position[31]), .I3(GND_net), .O(n538));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_mux_3_i7_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_add_1034_3_lut (.I0(GND_net), .I1(n1533), 
            .I2(VCC_net), .I3(n38896), .O(n1600)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1034_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15663_3_lut (.I0(\data_out_frame[21] [6]), .I1(current[15]), 
            .I2(n24278), .I3(GND_net), .O(n29611));   // verilog/coms.v(128[12] 303[6])
    defparam i15663_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_31__I_0_add_1034_3 (.CI(n38896), .I0(n1533), 
            .I1(VCC_net), .CO(n38897));
    SB_LUT4 encoder0_position_31__I_0_add_1034_2_lut (.I0(GND_net), .I1(n526), 
            .I2(GND_net), .I3(VCC_net), .O(n1601)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1034_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1034_2 (.CI(VCC_net), .I0(n526), 
            .I1(GND_net), .CO(n38896));
    SB_LUT4 i35109_1_lut (.I0(n2742), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n50697));
    defparam i35109_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i21450_3_lut (.I0(n538), .I1(n2732), .I2(n2733), .I3(GND_net), 
            .O(n35398));
    defparam i21450_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 encoder0_position_31__I_0_add_967_14_lut (.I0(n51053), .I1(n1422), 
            .I2(VCC_net), .I3(n38895), .O(n1521)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_967_14_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_31__I_0_add_967_13_lut (.I0(GND_net), .I1(n1423), 
            .I2(VCC_net), .I3(n38894), .O(n1490)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_967_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15664_3_lut (.I0(\data_out_frame[21] [5]), .I1(current[15]), 
            .I2(n24278), .I3(GND_net), .O(n29612));   // verilog/coms.v(128[12] 303[6])
    defparam i15664_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_31__I_0_add_967_13 (.CI(n38894), .I0(n1423), 
            .I1(VCC_net), .CO(n38895));
    SB_LUT4 encoder0_position_31__I_0_add_967_12_lut (.I0(GND_net), .I1(n1424), 
            .I2(VCC_net), .I3(n38893), .O(n1491)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_967_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_967_12 (.CI(n38893), .I0(n1424), 
            .I1(VCC_net), .CO(n38894));
    SB_LUT4 i1_4_lut_adj_1819 (.I0(n2729), .I1(n35398), .I2(n2730), .I3(n2731), 
            .O(n44993));
    defparam i1_4_lut_adj_1819.LUT_INIT = 16'ha080;
    SB_LUT4 i1_3_lut_adj_1820 (.I0(n2728), .I1(n2722), .I2(n2724), .I3(GND_net), 
            .O(n46975));
    defparam i1_3_lut_adj_1820.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_4_lut_adj_1821 (.I0(n2720), .I1(n46975), .I2(n2725), .I3(n2726), 
            .O(n46979));
    defparam i1_4_lut_adj_1821.LUT_INIT = 16'hfffe;
    SB_LUT4 i15665_3_lut (.I0(\data_out_frame[21] [4]), .I1(current[15]), 
            .I2(n24278), .I3(GND_net), .O(n29613));   // verilog/coms.v(128[12] 303[6])
    defparam i15665_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1822 (.I0(n2716), .I1(n44993), .I2(n2727), .I3(n2723), 
            .O(n46561));
    defparam i1_4_lut_adj_1822.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1823 (.I0(n46561), .I1(n2718), .I2(n2717), .I3(n46979), 
            .O(n46563));
    defparam i1_4_lut_adj_1823.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1824 (.I0(n2713), .I1(n2714), .I2(n2715), .I3(n46563), 
            .O(n46569));
    defparam i1_4_lut_adj_1824.LUT_INIT = 16'hfffe;
    SB_LUT4 i15666_3_lut (.I0(\data_out_frame[21] [3]), .I1(current[11]), 
            .I2(n24278), .I3(GND_net), .O(n29614));   // verilog/coms.v(128[12] 303[6])
    defparam i15666_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1825 (.I0(n2712), .I1(n2710), .I2(n2719), .I3(n2721), 
            .O(n45290));
    defparam i1_4_lut_adj_1825.LUT_INIT = 16'hfffe;
    SB_LUT4 i35113_4_lut (.I0(n2709), .I1(n45290), .I2(n2711), .I3(n46569), 
            .O(n2742));
    defparam i35113_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_31__I_0_add_967_11_lut (.I0(GND_net), .I1(n1425), 
            .I2(VCC_net), .I3(n38892), .O(n1492)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_967_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_967_11 (.CI(n38892), .I0(n1425), 
            .I1(VCC_net), .CO(n38893));
    SB_LUT4 encoder0_position_31__I_0_add_967_10_lut (.I0(GND_net), .I1(n1426), 
            .I2(VCC_net), .I3(n38891), .O(n1493)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_967_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_967_10 (.CI(n38891), .I0(n1426), 
            .I1(VCC_net), .CO(n38892));
    SB_LUT4 i15667_3_lut (.I0(\data_out_frame[21] [2]), .I1(current[10]), 
            .I2(n24278), .I3(GND_net), .O(n29615));   // verilog/coms.v(128[12] 303[6])
    defparam i15667_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i1708_3_lut (.I0(n2513), .I1(n2580), 
            .I2(n2544), .I3(GND_net), .O(n2612));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1708_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1707_3_lut (.I0(n2512), .I1(n2579), 
            .I2(n2544), .I3(GND_net), .O(n2611));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1707_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_967_9_lut (.I0(GND_net), .I1(n1427), 
            .I2(VCC_net), .I3(n38890), .O(n1494)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_967_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1711_3_lut (.I0(n2516), .I1(n2583), 
            .I2(n2544), .I3(GND_net), .O(n2615));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1711_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_967_9 (.CI(n38890), .I0(n1427), 
            .I1(VCC_net), .CO(n38891));
    SB_LUT4 encoder0_position_31__I_0_add_967_8_lut (.I0(GND_net), .I1(n1428), 
            .I2(VCC_net), .I3(n38889), .O(n1495)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_967_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_967_8 (.CI(n38889), .I0(n1428), 
            .I1(VCC_net), .CO(n38890));
    SB_LUT4 i15668_3_lut (.I0(\data_out_frame[21] [1]), .I1(current[9]), 
            .I2(n24278), .I3(GND_net), .O(n29616));   // verilog/coms.v(128[12] 303[6])
    defparam i15668_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_add_967_7_lut (.I0(GND_net), .I1(n1429), 
            .I2(GND_net), .I3(n38888), .O(n1496)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_967_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15669_3_lut (.I0(\data_out_frame[21] [0]), .I1(current[8]), 
            .I2(n24278), .I3(GND_net), .O(n29617));   // verilog/coms.v(128[12] 303[6])
    defparam i15669_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i1710_3_lut (.I0(n2515), .I1(n2582), 
            .I2(n2544), .I3(GND_net), .O(n2614));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1710_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15670_3_lut (.I0(\data_out_frame[20] [7]), .I1(displacement[7]), 
            .I2(n24278), .I3(GND_net), .O(n29618));   // verilog/coms.v(128[12] 303[6])
    defparam i15670_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i1709_3_lut (.I0(n2514), .I1(n2581), 
            .I2(n2544), .I3(GND_net), .O(n2613));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1709_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1727_3_lut (.I0(n2532), .I1(n2599), 
            .I2(n2544), .I3(GND_net), .O(n2631));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1727_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_967_7 (.CI(n38888), .I0(n1429), 
            .I1(GND_net), .CO(n38889));
    SB_LUT4 encoder0_position_31__I_0_i1726_3_lut (.I0(n2531), .I1(n2598), 
            .I2(n2544), .I3(GND_net), .O(n2630));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1726_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15671_3_lut (.I0(\data_out_frame[20] [6]), .I1(displacement[6]), 
            .I2(n24278), .I3(GND_net), .O(n29619));   // verilog/coms.v(128[12] 303[6])
    defparam i15671_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i1725_3_lut (.I0(n2530), .I1(n2597), 
            .I2(n2544), .I3(GND_net), .O(n2629));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1725_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1716_3_lut (.I0(n2521), .I1(n2588), 
            .I2(n2544), .I3(GND_net), .O(n2620));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1716_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1715_3_lut (.I0(n2520), .I1(n2587), 
            .I2(n2544), .I3(GND_net), .O(n2619));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1715_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15672_3_lut (.I0(\data_out_frame[20] [5]), .I1(displacement[5]), 
            .I2(n24278), .I3(GND_net), .O(n29620));   // verilog/coms.v(128[12] 303[6])
    defparam i15672_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15673_3_lut (.I0(\data_out_frame[20] [4]), .I1(displacement[4]), 
            .I2(n24278), .I3(GND_net), .O(n29621));   // verilog/coms.v(128[12] 303[6])
    defparam i15673_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_add_967_6_lut (.I0(GND_net), .I1(n1430), 
            .I2(GND_net), .I3(n38887), .O(n1497)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_967_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_967_6 (.CI(n38887), .I0(n1430), 
            .I1(GND_net), .CO(n38888));
    SB_LUT4 encoder0_position_31__I_0_i1714_3_lut (.I0(n2519), .I1(n2586), 
            .I2(n2544), .I3(GND_net), .O(n2618));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1714_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_967_5_lut (.I0(GND_net), .I1(n1431), 
            .I2(VCC_net), .I3(n38886), .O(n1498)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_967_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15674_3_lut (.I0(\data_out_frame[20] [3]), .I1(displacement[3]), 
            .I2(n24278), .I3(GND_net), .O(n29622));   // verilog/coms.v(128[12] 303[6])
    defparam i15674_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i1729_rep_16_3_lut (.I0(n950), .I1(n2601), 
            .I2(n2544), .I3(GND_net), .O(n2633));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1729_rep_16_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15675_3_lut (.I0(\data_out_frame[20] [2]), .I1(displacement[2]), 
            .I2(n24278), .I3(GND_net), .O(n29623));   // verilog/coms.v(128[12] 303[6])
    defparam i15675_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i1728_3_lut (.I0(n2533), .I1(n2600), 
            .I2(n2544), .I3(GND_net), .O(n2632));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1728_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i8_3_lut (.I0(encoder0_position[7]), 
            .I1(n26), .I2(encoder0_position[31]), .I3(GND_net), .O(n537));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_mux_3_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i1724_3_lut (.I0(n2529), .I1(n2596), 
            .I2(n2544), .I3(GND_net), .O(n2628));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1724_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1718_3_lut (.I0(n2523), .I1(n2590), 
            .I2(n2544), .I3(GND_net), .O(n2622));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1718_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_967_5 (.CI(n38886), .I0(n1431), 
            .I1(VCC_net), .CO(n38887));
    SB_LUT4 i15676_3_lut (.I0(\data_out_frame[20] [1]), .I1(displacement[1]), 
            .I2(n24278), .I3(GND_net), .O(n29624));   // verilog/coms.v(128[12] 303[6])
    defparam i15676_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_add_967_4_lut (.I0(GND_net), .I1(n1432), 
            .I2(GND_net), .I3(n38885), .O(n1499)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_967_4_lut.LUT_INIT = 16'hC33C;
    SB_DFFESR GHA_192 (.Q(GHA), .C(CLK_c), .E(n28482), .D(GHA_N_391), 
            .R(n28835));   // verilog/TinyFPGA_B.v(144[9] 223[5])
    SB_CARRY encoder0_position_31__I_0_add_967_4 (.CI(n38885), .I0(n1432), 
            .I1(GND_net), .CO(n38886));
    SB_LUT4 i15677_3_lut (.I0(\data_out_frame[20] [0]), .I1(displacement[0]), 
            .I2(n24278), .I3(GND_net), .O(n29625));   // verilog/coms.v(128[12] 303[6])
    defparam i15677_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_add_967_3_lut (.I0(GND_net), .I1(n1433), 
            .I2(VCC_net), .I3(n38884), .O(n1500)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_967_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15678_3_lut (.I0(\data_out_frame[19] [7]), .I1(displacement[15]), 
            .I2(n24278), .I3(GND_net), .O(n29626));   // verilog/coms.v(128[12] 303[6])
    defparam i15678_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34647_3_lut (.I0(n2425), .I1(n2492), .I2(n2445), .I3(GND_net), 
            .O(n2524));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam i34647_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i34639_3_lut (.I0(n2524), .I1(n2591), .I2(n2544), .I3(GND_net), 
            .O(n2623));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam i34639_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1722_3_lut (.I0(n2527), .I1(n2594), 
            .I2(n2544), .I3(GND_net), .O(n2626));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1722_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i34649_3_lut (.I0(n2423), .I1(n2490), .I2(n2445), .I3(GND_net), 
            .O(n2522));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam i34649_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i34637_3_lut (.I0(n2522), .I1(n2589), .I2(n2544), .I3(GND_net), 
            .O(n2621));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam i34637_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_967_3 (.CI(n38884), .I0(n1433), 
            .I1(VCC_net), .CO(n38885));
    SB_LUT4 encoder0_position_31__I_0_add_967_2_lut (.I0(GND_net), .I1(n525), 
            .I2(GND_net), .I3(VCC_net), .O(n1501)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_967_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_967_2 (.CI(VCC_net), .I0(n525), 
            .I1(GND_net), .CO(n38884));
    SB_LUT4 encoder0_position_31__I_0_add_900_13_lut (.I0(n51069), .I1(n1323_adj_5393), 
            .I2(VCC_net), .I3(n38883), .O(n1422)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_900_13_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_31__I_0_add_900_12_lut (.I0(GND_net), .I1(n1324_adj_5394), 
            .I2(VCC_net), .I3(n38882), .O(n1391)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_900_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_900_12 (.CI(n38882), .I0(n1324_adj_5394), 
            .I1(VCC_net), .CO(n38883));
    SB_LUT4 encoder0_position_31__I_0_add_900_11_lut (.I0(GND_net), .I1(n1325_adj_5395), 
            .I2(VCC_net), .I3(n38881), .O(n1392)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_900_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_900_11 (.CI(n38881), .I0(n1325_adj_5395), 
            .I1(VCC_net), .CO(n38882));
    SB_LUT4 encoder0_position_31__I_0_i1720_3_lut (.I0(n2525), .I1(n2592), 
            .I2(n2544), .I3(GND_net), .O(n2624));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1720_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1721_3_lut (.I0(n2526), .I1(n2593), 
            .I2(n2544), .I3(GND_net), .O(n2625));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1721_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1723_3_lut (.I0(n2528), .I1(n2595), 
            .I2(n2544), .I3(GND_net), .O(n2627));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1723_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1713_3_lut (.I0(n2518), .I1(n2585), 
            .I2(n2544), .I3(GND_net), .O(n2617));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1713_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1712_3_lut (.I0(n2517), .I1(n2584), 
            .I2(n2544), .I3(GND_net), .O(n2616));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1712_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_adj_1826 (.I0(n2627), .I1(n2625), .I2(GND_net), .I3(GND_net), 
            .O(n47023));
    defparam i1_2_lut_adj_1826.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_1827 (.I0(n2624), .I1(n2621), .I2(n2626), .I3(n2623), 
            .O(n47031));
    defparam i1_4_lut_adj_1827.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_31__I_0_add_900_10_lut (.I0(GND_net), .I1(n1326_adj_5396), 
            .I2(VCC_net), .I3(n38880), .O(n1393)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_900_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1828 (.I0(n2622), .I1(n47031), .I2(n47023), .I3(n2628), 
            .O(n47033));
    defparam i1_4_lut_adj_1828.LUT_INIT = 16'hfffe;
    SB_LUT4 i21452_3_lut (.I0(n537), .I1(n2632), .I2(n2633), .I3(GND_net), 
            .O(n35400));
    defparam i21452_3_lut.LUT_INIT = 16'hc8c8;
    SB_CARRY encoder0_position_31__I_0_add_900_10 (.CI(n38880), .I0(n1326_adj_5396), 
            .I1(VCC_net), .CO(n38881));
    SB_LUT4 encoder0_position_31__I_0_add_900_9_lut (.I0(GND_net), .I1(n1327_adj_5397), 
            .I2(VCC_net), .I3(n38879), .O(n1394)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_900_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_900_9 (.CI(n38879), .I0(n1327_adj_5397), 
            .I1(VCC_net), .CO(n38880));
    SB_LUT4 encoder0_position_31__I_0_add_900_8_lut (.I0(GND_net), .I1(n1328_adj_5398), 
            .I2(VCC_net), .I3(n38878), .O(n1395)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_900_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15679_3_lut (.I0(\data_out_frame[19] [6]), .I1(displacement[14]), 
            .I2(n24278), .I3(GND_net), .O(n29627));   // verilog/coms.v(128[12] 303[6])
    defparam i15679_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15108_3_lut (.I0(\data_out_frame[12] [0]), .I1(setpoint[16]), 
            .I2(n24278), .I3(GND_net), .O(n29056));   // verilog/coms.v(128[12] 303[6])
    defparam i15108_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15109_3_lut (.I0(CS_c), .I1(state_adj_5516[0]), .I2(state_adj_5516[1]), 
            .I3(GND_net), .O(n29057));   // verilog/tli4970.v(35[10] 68[6])
    defparam i15109_3_lut.LUT_INIT = 16'ha3a3;
    SB_LUT4 i35614_4_lut (.I0(n15_adj_5339), .I1(clk_out), .I2(state_adj_5516[0]), 
            .I3(state_adj_5516[1]), .O(n9_adj_5289));   // verilog/tli4970.v(35[10] 68[6])
    defparam i35614_4_lut.LUT_INIT = 16'hc8fc;
    SB_LUT4 i1_4_lut_adj_1829 (.I0(n2618), .I1(n2619), .I2(n47033), .I3(n2620), 
            .O(n47039));
    defparam i1_4_lut_adj_1829.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_3_lut_adj_1830 (.I0(data_ready), .I1(\ID_READOUT_FSM.state [1]), 
            .I2(\ID_READOUT_FSM.state [0]), .I3(GND_net), .O(n46410));
    defparam i2_3_lut_adj_1830.LUT_INIT = 16'hdfdf;
    SB_LUT4 i15111_3_lut (.I0(ID[0]), .I1(data[0]), .I2(n46410), .I3(GND_net), 
            .O(n29059));   // verilog/TinyFPGA_B.v(375[10] 403[6])
    defparam i15111_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1831 (.I0(n2629), .I1(n35400), .I2(n2630), .I3(n2631), 
            .O(n45028));
    defparam i1_4_lut_adj_1831.LUT_INIT = 16'ha080;
    SB_LUT4 i1_4_lut_adj_1832 (.I0(n2616), .I1(n2617), .I2(n45028), .I3(n47039), 
            .O(n47045));
    defparam i1_4_lut_adj_1832.LUT_INIT = 16'hfffe;
    SB_LUT4 i15112_3_lut (.I0(\data_out_frame[11] [7]), .I1(encoder1_position_scaled[7]), 
            .I2(n24278), .I3(GND_net), .O(n29060));   // verilog/coms.v(128[12] 303[6])
    defparam i15112_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15113_3_lut (.I0(\data_out_frame[11] [6]), .I1(encoder1_position_scaled[6]), 
            .I2(n24278), .I3(GND_net), .O(n29061));   // verilog/coms.v(128[12] 303[6])
    defparam i15113_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_31__I_0_add_900_8 (.CI(n38878), .I0(n1328_adj_5398), 
            .I1(VCC_net), .CO(n38879));
    SB_LUT4 encoder0_position_31__I_0_add_900_7_lut (.I0(GND_net), .I1(n1329), 
            .I2(GND_net), .I3(n38877), .O(n1396)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_900_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_900_7 (.CI(n38877), .I0(n1329), 
            .I1(GND_net), .CO(n38878));
    SB_LUT4 encoder0_position_31__I_0_add_900_6_lut (.I0(GND_net), .I1(n1330), 
            .I2(GND_net), .I3(n38876), .O(n1397)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_900_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_19_add_3_25_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_setpoint_23__N_239), 
            .I3(n38553), .O(n340)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_19_add_3_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1833 (.I0(n2613), .I1(n2614), .I2(n2615), .I3(n47045), 
            .O(n47051));
    defparam i1_4_lut_adj_1833.LUT_INIT = 16'hfffe;
    SB_LUT4 i35142_4_lut (.I0(n2611), .I1(n2610), .I2(n2612), .I3(n47051), 
            .O(n2643));
    defparam i35142_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i15114_3_lut (.I0(\data_out_frame[11] [5]), .I1(encoder1_position_scaled[5]), 
            .I2(n24278), .I3(GND_net), .O(n29062));   // verilog/coms.v(128[12] 303[6])
    defparam i15114_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_29 (.CI(n39519), 
            .I0(GND_net), .I1(n6_adj_5415), .CO(n39520));
    SB_LUT4 i15115_3_lut (.I0(\data_out_frame[11] [4]), .I1(encoder1_position_scaled[4]), 
            .I2(n24278), .I3(GND_net), .O(n29063));   // verilog/coms.v(128[12] 303[6])
    defparam i15115_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15116_3_lut (.I0(\data_out_frame[11] [3]), .I1(encoder1_position_scaled[3]), 
            .I2(n24278), .I3(GND_net), .O(n29064));   // verilog/coms.v(128[12] 303[6])
    defparam i15116_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4598_4_lut (.I0(n27028), .I1(delay_counter[11]), .I2(delay_counter[10]), 
            .I3(delay_counter[9]), .O(n24_adj_5403));
    defparam i4598_4_lut.LUT_INIT = 16'hc8c0;
    SB_LUT4 i15195_3_lut (.I0(IntegralLimit[13]), .I1(\data_in_frame[12] [5]), 
            .I2(n28521), .I3(GND_net), .O(n29143));   // verilog/coms.v(128[12] 303[6])
    defparam i15195_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_31__I_0_add_900_6 (.CI(n38876), .I0(n1330), 
            .I1(GND_net), .CO(n38877));
    SB_LUT4 encoder0_position_31__I_0_add_900_5_lut (.I0(GND_net), .I1(n1331), 
            .I2(VCC_net), .I3(n38875), .O(n1398)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_900_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15196_3_lut (.I0(IntegralLimit[12]), .I1(\data_in_frame[12] [4]), 
            .I2(n28521), .I3(GND_net), .O(n29144));   // verilog/coms.v(128[12] 303[6])
    defparam i15196_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_157_31 (.CI(n38474), .I0(delay_counter[29]), .I1(GND_net), 
            .CO(n38475));
    SB_CARRY add_157_4 (.CI(n38447), .I0(delay_counter[2]), .I1(GND_net), 
            .CO(n38448));
    SB_LUT4 i15117_3_lut (.I0(\data_out_frame[11] [2]), .I1(encoder1_position_scaled[2]), 
            .I2(n24278), .I3(GND_net), .O(n29065));   // verilog/coms.v(128[12] 303[6])
    defparam i15117_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15197_3_lut (.I0(IntegralLimit[11]), .I1(\data_in_frame[12] [3]), 
            .I2(n28521), .I3(GND_net), .O(n29145));   // verilog/coms.v(128[12] 303[6])
    defparam i15197_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2_4_lut (.I0(n24_adj_5403), .I1(delay_counter[14]), .I2(delay_counter[12]), 
            .I3(delay_counter[13]), .O(n45933));
    defparam i2_4_lut.LUT_INIT = 16'hc800;
    SB_LUT4 i15198_4_lut (.I0(saved_addr[0]), .I1(rw), .I2(state_7__N_4251[0]), 
            .I3(enable_slow_N_4354), .O(n29146));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i15198_4_lut.LUT_INIT = 16'haaca;
    SB_LUT4 i2_3_lut_adj_1834 (.I0(n45933), .I1(delay_counter[18]), .I2(n27034), 
            .I3(GND_net), .O(n46347));
    defparam i2_3_lut_adj_1834.LUT_INIT = 16'hfefe;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_28_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n7_adj_5416), .I3(n39518), .O(n7_adj_5308)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_28_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15199_3_lut (.I0(IntegralLimit[10]), .I1(\data_in_frame[12] [2]), 
            .I2(n28521), .I3(GND_net), .O(n29147));   // verilog/coms.v(128[12] 303[6])
    defparam i15199_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15200_3_lut (.I0(IntegralLimit[9]), .I1(\data_in_frame[12] [1]), 
            .I2(n28521), .I3(GND_net), .O(n29148));   // verilog/coms.v(128[12] 303[6])
    defparam i15200_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2_4_lut_adj_1835 (.I0(delay_counter[23]), .I1(n46347), .I2(delay_counter[20]), 
            .I3(delay_counter[19]), .O(n7_adj_5273));
    defparam i2_4_lut_adj_1835.LUT_INIT = 16'heaaa;
    SB_LUT4 i15201_3_lut (.I0(IntegralLimit[8]), .I1(\data_in_frame[12] [0]), 
            .I2(n28521), .I3(GND_net), .O(n29149));   // verilog/coms.v(128[12] 303[6])
    defparam i15201_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_19_add_3_24_lut (.I0(GND_net), .I1(GND_net), .I2(n3), 
            .I3(n38552), .O(n341)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_19_add_3_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_19_inv_0_i1_1_lut (.I0(duty[0]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n25));   // verilog/TinyFPGA_B.v(123[25:30])
    defparam unary_minus_19_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i15118_4_lut (.I0(tx_active), .I1(r_SM_Main_adj_5525[1]), .I2(n19541), 
            .I3(n4_adj_5272), .O(n29066));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i15118_4_lut.LUT_INIT = 16'h32aa;
    SB_CARRY unary_minus_19_add_3_24 (.CI(n38552), .I0(GND_net), .I1(n3), 
            .CO(n38553));
    SB_LUT4 i4_4_lut (.I0(n7_adj_5273), .I1(delay_counter[21]), .I2(delay_counter[22]), 
            .I3(n27037), .O(n62));
    defparam i4_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_4_lut (.I0(control_mode[0]), .I1(control_mode[6]), 
            .I2(n10_adj_5453), .I3(control_mode[2]), .O(n27015));   // verilog/TinyFPGA_B.v(286[5:22])
    defparam i1_2_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_2_lut (.I0(ID[2]), .I1(ID[4]), .I2(GND_net), .I3(GND_net), 
            .O(n10_adj_5283));   // verilog/TinyFPGA_B.v(393[7:11])
    defparam i2_2_lut.LUT_INIT = 16'heeee;
    SB_CARRY encoder0_position_31__I_0_add_900_5 (.CI(n38875), .I0(n1331), 
            .I1(VCC_net), .CO(n38876));
    SB_LUT4 i6_4_lut_adj_1836 (.I0(ID[7]), .I1(ID[5]), .I2(ID[1]), .I3(ID[0]), 
            .O(n14_adj_5282));   // verilog/TinyFPGA_B.v(393[7:11])
    defparam i6_4_lut_adj_1836.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_4_lut (.I0(ID[3]), .I1(n14_adj_5282), .I2(n10_adj_5283), 
            .I3(ID[6]), .O(n27013));   // verilog/TinyFPGA_B.v(393[7:11])
    defparam i7_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i15119_3_lut (.I0(\data_out_frame[11] [1]), .I1(encoder1_position_scaled[1]), 
            .I2(n24278), .I3(GND_net), .O(n29067));   // verilog/coms.v(128[12] 303[6])
    defparam i15119_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 \ID_READOUT_FSM.state_2__I_0_i5_2_lut  (.I0(\ID_READOUT_FSM.state [0]), 
            .I1(\ID_READOUT_FSM.state [1]), .I2(GND_net), .I3(GND_net), 
            .O(n5_adj_5368));   // verilog/TinyFPGA_B.v(393[7:11])
    defparam \ID_READOUT_FSM.state_2__I_0_i5_2_lut .LUT_INIT = 16'hbbbb;
    SB_LUT4 i5_4_lut (.I0(delay_counter[27]), .I1(delay_counter[29]), .I2(delay_counter[24]), 
            .I3(delay_counter[26]), .O(n12_adj_5276));
    defparam i5_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i29_1_lut (.I0(encoder0_position[28]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n5_adj_5414));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i29_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i6_4_lut_adj_1837 (.I0(delay_counter[28]), .I1(n12_adj_5276), 
            .I2(delay_counter[25]), .I3(delay_counter[30]), .O(n27037));
    defparam i6_4_lut_adj_1837.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_3_lut_adj_1838 (.I0(delay_counter[17]), .I1(delay_counter[16]), 
            .I2(delay_counter[15]), .I3(GND_net), .O(n27034));
    defparam i2_3_lut_adj_1838.LUT_INIT = 16'hfefe;
    SB_LUT4 inv_1004_i1_1_lut (.I0(current[0]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n4698));   // verilog/TinyFPGA_B.v(118[13] 129[7])
    defparam inv_1004_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i5_3_lut_adj_1839 (.I0(delay_counter[3]), .I1(delay_counter[5]), 
            .I2(delay_counter[4]), .I3(GND_net), .O(n14));
    defparam i5_3_lut_adj_1839.LUT_INIT = 16'hfefe;
    SB_LUT4 i15213_3_lut (.I0(h1), .I1(reg_B[2]), .I2(n46440), .I3(GND_net), 
            .O(n29161));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    defparam i15213_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i6_4_lut_adj_1840 (.I0(delay_counter[8]), .I1(delay_counter[7]), 
            .I2(delay_counter[1]), .I3(delay_counter[0]), .O(n15_adj_5244));
    defparam i6_4_lut_adj_1840.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i30_1_lut (.I0(encoder0_position[29]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n4_adj_5413));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i30_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i31_1_lut (.I0(encoder0_position[30]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n3_adj_5412));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i31_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i8_4_lut (.I0(n15_adj_5244), .I1(delay_counter[2]), .I2(n14), 
            .I3(delay_counter[6]), .O(n27028));
    defparam i8_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i15579_3_lut (.I0(\data_out_frame[23] [7]), .I1(neopxl_color[23]), 
            .I2(n24278), .I3(GND_net), .O(n29527));   // verilog/coms.v(128[12] 303[6])
    defparam i15579_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15202_3_lut (.I0(IntegralLimit[7]), .I1(\data_in_frame[13] [7]), 
            .I2(n28521), .I3(GND_net), .O(n29150));   // verilog/coms.v(128[12] 303[6])
    defparam i15202_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_1841 (.I0(delay_counter[12]), .I1(delay_counter[11]), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_5243));
    defparam i1_2_lut_adj_1841.LUT_INIT = 16'heeee;
    SB_LUT4 unary_minus_17_inv_0_i2_1_lut (.I0(current[1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n24));   // verilog/TinyFPGA_B.v(122[16:24])
    defparam unary_minus_17_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i2_4_lut_adj_1842 (.I0(delay_counter[9]), .I1(n4_adj_5243), 
            .I2(delay_counter[10]), .I3(n27028), .O(n45355));
    defparam i2_4_lut_adj_1842.LUT_INIT = 16'hfcec;
    SB_LUT4 i2_2_lut_adj_1843 (.I0(dti_counter[1]), .I1(dti_counter[2]), 
            .I2(GND_net), .I3(GND_net), .O(n10_adj_5444));   // verilog/TinyFPGA_B.v(172[9:23])
    defparam i2_2_lut_adj_1843.LUT_INIT = 16'heeee;
    SB_LUT4 i2_4_lut_adj_1844 (.I0(n45355), .I1(n27034), .I2(delay_counter[13]), 
            .I3(delay_counter[14]), .O(n46354));
    defparam i2_4_lut_adj_1844.LUT_INIT = 16'hffec;
    SB_LUT4 i6_4_lut_adj_1845 (.I0(dti_counter[7]), .I1(dti_counter[4]), 
            .I2(dti_counter[5]), .I3(dti_counter[6]), .O(n14_adj_5443));   // verilog/TinyFPGA_B.v(172[9:23])
    defparam i6_4_lut_adj_1845.LUT_INIT = 16'hfffe;
    SB_LUT4 i15121_4_lut (.I0(n44637), .I1(state[1]), .I2(state_3__N_552[1]), 
            .I3(n28592), .O(n29069));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15121_4_lut.LUT_INIT = 16'hfaee;
    SB_LUT4 i3_3_lut_adj_1846 (.I0(delay_counter[20]), .I1(delay_counter[21]), 
            .I2(delay_counter[23]), .I3(GND_net), .O(n8_adj_5280));
    defparam i3_3_lut_adj_1846.LUT_INIT = 16'h8080;
    SB_LUT4 i7_4_lut_adj_1847 (.I0(dti_counter[0]), .I1(n14_adj_5443), .I2(n10_adj_5444), 
            .I3(dti_counter[3]), .O(n24462));   // verilog/TinyFPGA_B.v(172[9:23])
    defparam i7_4_lut_adj_1847.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_4_lut_adj_1848 (.I0(delay_counter[22]), .I1(n46354), .I2(delay_counter[19]), 
            .I3(delay_counter[18]), .O(n7_adj_5281));
    defparam i2_4_lut_adj_1848.LUT_INIT = 16'ha8a0;
    SB_LUT4 i1_4_lut_adj_1849 (.I0(commutation_state[2]), .I1(commutation_state[1]), 
            .I2(commutation_state_prev[2]), .I3(commutation_state_prev[1]), 
            .O(n4));   // verilog/TinyFPGA_B.v(147[7:48])
    defparam i1_4_lut_adj_1849.LUT_INIT = 16'h7bde;
    SB_LUT4 i20854_4_lut (.I0(n7_adj_5281), .I1(delay_counter[31]), .I2(n27037), 
            .I3(n8_adj_5280), .O(n1415));   // verilog/TinyFPGA_B.v(396[14:38])
    defparam i20854_4_lut.LUT_INIT = 16'h3230;
    SB_LUT4 i20849_2_lut (.I0(n62), .I1(delay_counter[31]), .I2(GND_net), 
            .I3(GND_net), .O(read_N_445));   // verilog/TinyFPGA_B.v(381[12:35])
    defparam i20849_2_lut.LUT_INIT = 16'h2222;
    SB_DFFESS commutation_state_i0 (.Q(commutation_state[0]), .C(CLK_c), 
            .E(n6_adj_5454), .D(commutation_state_7__N_240[0]), .S(commutation_state_7__N_248));   // verilog/TinyFPGA_B.v(144[9] 223[5])
    SB_LUT4 i35391_1_lut (.I0(n1851), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n50979));
    defparam i35391_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i15125_4_lut (.I0(CS_MISO_c), .I1(data_adj_5514[2]), .I2(n10_adj_5341), 
            .I3(n27177), .O(n29073));   // verilog/tli4970.v(35[10] 68[6])
    defparam i15125_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i2_2_lut_3_lut (.I0(h1), .I1(h3), .I2(h2), .I3(GND_net), 
            .O(commutation_state_7__N_248));   // verilog/TinyFPGA_B.v(167[7:23])
    defparam i2_2_lut_3_lut.LUT_INIT = 16'h0404;
    SB_LUT4 i2_3_lut_4_lut (.I0(data_ready), .I1(n62), .I2(delay_counter[31]), 
            .I3(\ID_READOUT_FSM.state [0]), .O(n6_adj_5445));   // verilog/TinyFPGA_B.v(375[10] 403[6])
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h080c;
    SB_LUT4 i2050_4_lut_4_lut (.I0(\ID_READOUT_FSM.state [0]), .I1(\ID_READOUT_FSM.state [1]), 
            .I2(n1415), .I3(n27013), .O(n7494));   // verilog/TinyFPGA_B.v(378[5] 402[12])
    defparam i2050_4_lut_4_lut.LUT_INIT = 16'hcc8c;
    SB_LUT4 i35555_2_lut (.I0(n24462), .I1(dti), .I2(GND_net), .I3(GND_net), 
            .O(dti_N_440));
    defparam i35555_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 encoder0_position_31__I_0_add_900_4_lut (.I0(GND_net), .I1(n1332), 
            .I2(GND_net), .I3(n38874), .O(n1399)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_900_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i3_4_lut_4_lut (.I0(r_SM_Main_adj_5525[2]), .I1(r_SM_Main_adj_5525[0]), 
            .I2(r_SM_Main_2__N_3777[1]), .I3(r_SM_Main_adj_5525[1]), .O(n51602));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i3_4_lut_4_lut.LUT_INIT = 16'h4000;
    SB_LUT4 i15014_4_lut (.I0(n7417), .I1(n1415), .I2(n49335), .I3(n27014), 
            .O(n28933));   // verilog/TinyFPGA_B.v(375[10] 403[6])
    defparam i15014_4_lut.LUT_INIT = 16'ha088;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_28 (.CI(n39518), 
            .I0(GND_net), .I1(n7_adj_5416), .CO(n39519));
    SB_LUT4 i15126_3_lut (.I0(\data_out_frame[11] [0]), .I1(encoder1_position_scaled[0]), 
            .I2(n24278), .I3(GND_net), .O(n29074));   // verilog/coms.v(128[12] 303[6])
    defparam i15126_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_31__I_0_add_900_4 (.CI(n38874), .I0(n1332), 
            .I1(GND_net), .CO(n38875));
    SB_LUT4 encoder0_position_31__I_0_add_900_3_lut (.I0(GND_net), .I1(n1333), 
            .I2(VCC_net), .I3(n38873), .O(n1400)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_900_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_900_3 (.CI(n38873), .I0(n1333), 
            .I1(VCC_net), .CO(n38874));
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_27_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n8_adj_5417), .I3(n39517), .O(n8_adj_5307)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_27_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_900_2_lut (.I0(GND_net), .I1(n938), 
            .I2(GND_net), .I3(VCC_net), .O(n1401)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_900_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_19_add_3_23_lut (.I0(GND_net), .I1(GND_net), .I2(n4_adj_5255), 
            .I3(n38551), .O(n342)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_19_add_3_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_900_2 (.CI(VCC_net), .I0(n938), 
            .I1(GND_net), .CO(n38873));
    SB_LUT4 encoder0_position_31__I_0_add_833_12_lut (.I0(n51084), .I1(n1224), 
            .I2(VCC_net), .I3(n38872), .O(n1323_adj_5393)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_833_12_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_31__I_0_add_833_11_lut (.I0(GND_net), .I1(n1225), 
            .I2(VCC_net), .I3(n38871), .O(n1292)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_833_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_27 (.CI(n39517), 
            .I0(GND_net), .I1(n8_adj_5417), .CO(n39518));
    SB_CARRY encoder0_position_31__I_0_add_833_11 (.CI(n38871), .I0(n1225), 
            .I1(VCC_net), .CO(n38872));
    SB_LUT4 encoder0_position_31__I_0_add_833_10_lut (.I0(GND_net), .I1(n1226), 
            .I2(VCC_net), .I3(n38870), .O(n1293)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_833_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_833_10 (.CI(n38870), .I0(n1226), 
            .I1(VCC_net), .CO(n38871));
    SB_LUT4 encoder0_position_31__I_0_add_833_9_lut (.I0(GND_net), .I1(n1227), 
            .I2(VCC_net), .I3(n38869), .O(n1294)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_833_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_26_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n9_adj_5418), .I3(n39516), .O(n9_adj_5306)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_833_9 (.CI(n38869), .I0(n1227), 
            .I1(VCC_net), .CO(n38870));
    SB_LUT4 encoder0_position_31__I_0_add_833_8_lut (.I0(GND_net), .I1(n1228), 
            .I2(VCC_net), .I3(n38868), .O(n1295)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_833_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_26 (.CI(n39516), 
            .I0(GND_net), .I1(n9_adj_5418), .CO(n39517));
    SB_CARRY encoder0_position_31__I_0_add_833_8 (.CI(n38868), .I0(n1228), 
            .I1(VCC_net), .CO(n38869));
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_25_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n10_adj_5419), .I3(n39515), .O(n10_adj_5305)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_833_7_lut (.I0(GND_net), .I1(n1229), 
            .I2(GND_net), .I3(n38867), .O(n1296)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_833_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_25 (.CI(n39515), 
            .I0(GND_net), .I1(n10_adj_5419), .CO(n39516));
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_24_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n11_adj_5420), .I3(n39514), .O(n11_adj_5304)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_833_7 (.CI(n38867), .I0(n1229), 
            .I1(GND_net), .CO(n38868));
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_24 (.CI(n39514), 
            .I0(GND_net), .I1(n11_adj_5420), .CO(n39515));
    SB_LUT4 encoder0_position_31__I_0_add_833_6_lut (.I0(GND_net), .I1(n1230), 
            .I2(GND_net), .I3(n38866), .O(n1297_adj_5388)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_833_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_23_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n12_adj_5421), .I3(n39513), .O(n12_adj_5303)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_833_6 (.CI(n38866), .I0(n1230), 
            .I1(GND_net), .CO(n38867));
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_23 (.CI(n39513), 
            .I0(GND_net), .I1(n12_adj_5421), .CO(n39514));
    SB_LUT4 encoder0_position_31__I_0_add_833_5_lut (.I0(GND_net), .I1(n1231), 
            .I2(VCC_net), .I3(n38865), .O(n1298_adj_5389)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_833_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_22_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n13_adj_5422), .I3(n39512), .O(n13_adj_5302)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_833_5 (.CI(n38865), .I0(n1231), 
            .I1(VCC_net), .CO(n38866));
    SB_LUT4 encoder0_position_31__I_0_add_833_4_lut (.I0(GND_net), .I1(n1232), 
            .I2(GND_net), .I3(n38864), .O(n1299_adj_5390)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_833_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_22 (.CI(n39512), 
            .I0(GND_net), .I1(n13_adj_5422), .CO(n39513));
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_21_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n14_adj_5423), .I3(n39511), .O(n14_adj_5301)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_21 (.CI(n39511), 
            .I0(GND_net), .I1(n14_adj_5423), .CO(n39512));
    SB_CARRY encoder0_position_31__I_0_add_833_4 (.CI(n38864), .I0(n1232), 
            .I1(GND_net), .CO(n38865));
    SB_LUT4 encoder0_position_31__I_0_add_833_3_lut (.I0(GND_net), .I1(n1233), 
            .I2(VCC_net), .I3(n38863), .O(n1300_adj_5391)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_833_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_833_3 (.CI(n38863), .I0(n1233), 
            .I1(VCC_net), .CO(n38864));
    SB_CARRY unary_minus_19_add_3_23 (.CI(n38551), .I0(GND_net), .I1(n4_adj_5255), 
            .CO(n38552));
    SB_LUT4 encoder0_position_31__I_0_add_833_2_lut (.I0(GND_net), .I1(n937), 
            .I2(GND_net), .I3(VCC_net), .O(n1301_adj_5392)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_833_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_833_2 (.CI(VCC_net), .I0(n937), 
            .I1(GND_net), .CO(n38863));
    SB_LUT4 encoder0_position_31__I_0_add_766_11_lut (.I0(n51099), .I1(n1125), 
            .I2(VCC_net), .I3(n38862), .O(n1224)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_766_11_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_20_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n15_adj_5424), .I3(n39510), .O(n15_adj_5300)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_20 (.CI(n39510), 
            .I0(GND_net), .I1(n15_adj_5424), .CO(n39511));
    SB_LUT4 encoder0_position_31__I_0_add_766_10_lut (.I0(GND_net), .I1(n1126), 
            .I2(VCC_net), .I3(n38861), .O(n1193)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_766_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_19_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n16_adj_5425), .I3(n39509), .O(n16_adj_5299)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_19_add_3_22_lut (.I0(GND_net), .I1(GND_net), .I2(n5), 
            .I3(n38550), .O(n343)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_19_add_3_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_157_30_lut (.I0(GND_net), .I1(delay_counter[28]), .I2(GND_net), 
            .I3(n38473), .O(n1300)) /* synthesis syn_instantiated=1 */ ;
    defparam add_157_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_766_10 (.CI(n38861), .I0(n1126), 
            .I1(VCC_net), .CO(n38862));
    SB_LUT4 encoder0_position_31__I_0_add_766_9_lut (.I0(GND_net), .I1(n1127), 
            .I2(VCC_net), .I3(n38860), .O(n1194)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_766_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_766_9 (.CI(n38860), .I0(n1127), 
            .I1(VCC_net), .CO(n38861));
    SB_LUT4 encoder0_position_31__I_0_add_766_8_lut (.I0(GND_net), .I1(n1128), 
            .I2(VCC_net), .I3(n38859), .O(n1195)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_766_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_19 (.CI(n39509), 
            .I0(GND_net), .I1(n16_adj_5425), .CO(n39510));
    SB_CARRY add_157_10 (.CI(n38453), .I0(delay_counter[8]), .I1(GND_net), 
            .CO(n38454));
    SB_LUT4 add_157_9_lut (.I0(GND_net), .I1(delay_counter[7]), .I2(GND_net), 
            .I3(n38452), .O(n1321)) /* synthesis syn_instantiated=1 */ ;
    defparam add_157_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_766_8 (.CI(n38859), .I0(n1128), 
            .I1(VCC_net), .CO(n38860));
    SB_LUT4 encoder0_position_31__I_0_add_766_7_lut (.I0(GND_net), .I1(n1129), 
            .I2(GND_net), .I3(n38858), .O(n1196)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_766_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_766_7 (.CI(n38858), .I0(n1129), 
            .I1(GND_net), .CO(n38859));
    SB_LUT4 encoder0_position_31__I_0_add_766_6_lut (.I0(GND_net), .I1(n1130), 
            .I2(GND_net), .I3(n38857), .O(n1197)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_766_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_766_6 (.CI(n38857), .I0(n1130), 
            .I1(GND_net), .CO(n38858));
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_18_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n17_adj_5426), .I3(n39508), .O(n17_adj_5298)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_157_30 (.CI(n38473), .I0(delay_counter[28]), .I1(GND_net), 
            .CO(n38474));
    SB_LUT4 encoder0_position_31__I_0_add_766_5_lut (.I0(GND_net), .I1(n1131), 
            .I2(VCC_net), .I3(n38856), .O(n1198)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_766_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_766_5 (.CI(n38856), .I0(n1131), 
            .I1(VCC_net), .CO(n38857));
    SB_LUT4 encoder0_position_31__I_0_add_766_4_lut (.I0(GND_net), .I1(n1132), 
            .I2(GND_net), .I3(n38855), .O(n1199)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_766_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_18 (.CI(n39508), 
            .I0(GND_net), .I1(n17_adj_5426), .CO(n39509));
    SB_CARRY encoder0_position_31__I_0_add_766_4 (.CI(n38855), .I0(n1132), 
            .I1(GND_net), .CO(n38856));
    SB_LUT4 add_157_3_lut (.I0(GND_net), .I1(delay_counter[1]), .I2(GND_net), 
            .I3(n38446), .O(n1327)) /* synthesis syn_instantiated=1 */ ;
    defparam add_157_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_17_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n18_adj_5427), .I3(n39507), .O(n18_adj_5297)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_766_3_lut (.I0(GND_net), .I1(n1133), 
            .I2(VCC_net), .I3(n38854), .O(n1200)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_766_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_17 (.CI(n39507), 
            .I0(GND_net), .I1(n18_adj_5427), .CO(n39508));
    SB_CARRY encoder0_position_31__I_0_add_766_3 (.CI(n38854), .I0(n1133), 
            .I1(VCC_net), .CO(n38855));
    SB_LUT4 i15214_3_lut (.I0(h2), .I1(reg_B[1]), .I2(n46440), .I3(GND_net), 
            .O(n29162));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    defparam i15214_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_16_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n19_adj_5428), .I3(n39506), .O(n19_adj_5296)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_16 (.CI(n39506), 
            .I0(GND_net), .I1(n19_adj_5428), .CO(n39507));
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_15_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n20_adj_5429), .I3(n39505), .O(n20_adj_5295)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_15 (.CI(n39505), 
            .I0(GND_net), .I1(n20_adj_5429), .CO(n39506));
    SB_LUT4 add_157_29_lut (.I0(GND_net), .I1(delay_counter[27]), .I2(GND_net), 
            .I3(n38472), .O(n1301)) /* synthesis syn_instantiated=1 */ ;
    defparam add_157_29_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_766_2_lut (.I0(GND_net), .I1(n522), 
            .I2(GND_net), .I3(VCC_net), .O(n1201)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_766_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_766_2 (.CI(VCC_net), .I0(n522), 
            .I1(GND_net), .CO(n38854));
    SB_LUT4 encoder0_position_31__I_0_add_699_10_lut (.I0(GND_net), .I1(n1026), 
            .I2(VCC_net), .I3(n38853), .O(n1093)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_699_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_699_9_lut (.I0(GND_net), .I1(n1027), 
            .I2(VCC_net), .I3(n38852), .O(n1094)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_699_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_14_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n21_adj_5430), .I3(n39504), .O(n21_adj_5294)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_699_9 (.CI(n38852), .I0(n1027), 
            .I1(VCC_net), .CO(n38853));
    SB_LUT4 encoder0_position_31__I_0_add_699_8_lut (.I0(GND_net), .I1(n1028), 
            .I2(VCC_net), .I3(n38851), .O(n1095)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_699_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15127_3_lut (.I0(\data_out_frame[10] [7]), .I1(encoder1_position_scaled[15]), 
            .I2(n24278), .I3(GND_net), .O(n29075));   // verilog/coms.v(128[12] 303[6])
    defparam i15127_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_157_29 (.CI(n38472), .I0(delay_counter[27]), .I1(GND_net), 
            .CO(n38473));
    SB_CARRY encoder0_position_31__I_0_add_699_8 (.CI(n38851), .I0(n1028), 
            .I1(VCC_net), .CO(n38852));
    SB_LUT4 encoder0_position_31__I_0_add_699_7_lut (.I0(GND_net), .I1(n1029), 
            .I2(GND_net), .I3(n38850), .O(n1096)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_699_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15128_3_lut (.I0(\data_out_frame[10] [6]), .I1(encoder1_position_scaled[14]), 
            .I2(n24278), .I3(GND_net), .O(n29076));   // verilog/coms.v(128[12] 303[6])
    defparam i15128_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY unary_minus_19_add_3_22 (.CI(n38550), .I0(GND_net), .I1(n5), 
            .CO(n38551));
    SB_CARRY encoder0_position_31__I_0_add_699_7 (.CI(n38850), .I0(n1029), 
            .I1(GND_net), .CO(n38851));
    SB_LUT4 encoder0_position_31__I_0_add_699_6_lut (.I0(GND_net), .I1(n1030), 
            .I2(GND_net), .I3(n38849), .O(n1097)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_699_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_14 (.CI(n39504), 
            .I0(GND_net), .I1(n21_adj_5430), .CO(n39505));
    SB_CARRY encoder0_position_31__I_0_add_699_6 (.CI(n38849), .I0(n1030), 
            .I1(GND_net), .CO(n38850));
    SB_CARRY add_157_9 (.CI(n38452), .I0(delay_counter[7]), .I1(GND_net), 
            .CO(n38453));
    SB_LUT4 encoder0_position_31__I_0_add_699_5_lut (.I0(GND_net), .I1(n1031), 
            .I2(VCC_net), .I3(n38848), .O(n1098)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_699_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_699_5 (.CI(n38848), .I0(n1031), 
            .I1(VCC_net), .CO(n38849));
    SB_LUT4 encoder0_position_31__I_0_add_699_4_lut (.I0(GND_net), .I1(n1032), 
            .I2(GND_net), .I3(n38847), .O(n1099)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_699_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_699_4 (.CI(n38847), .I0(n1032), 
            .I1(GND_net), .CO(n38848));
    SB_LUT4 encoder0_position_31__I_0_add_699_3_lut (.I0(GND_net), .I1(n1033), 
            .I2(VCC_net), .I3(n38846), .O(n1100)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_699_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_13_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n22_adj_5431), .I3(n39503), .O(n22_adj_5293)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_699_3 (.CI(n38846), .I0(n1033), 
            .I1(VCC_net), .CO(n38847));
    SB_LUT4 unary_minus_19_add_3_21_lut (.I0(GND_net), .I1(GND_net), .I2(n6_adj_5256), 
            .I3(n38549), .O(n344)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_19_add_3_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_699_2_lut (.I0(GND_net), .I1(n521), 
            .I2(GND_net), .I3(VCC_net), .O(n1101)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_699_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_19_add_3_21 (.CI(n38549), .I0(GND_net), .I1(n6_adj_5256), 
            .CO(n38550));
    SB_CARRY encoder0_position_31__I_0_add_699_2 (.CI(VCC_net), .I0(n521), 
            .I1(GND_net), .CO(n38846));
    SB_LUT4 encoder0_position_31__I_0_add_632_9_lut (.I0(n960), .I1(n927), 
            .I2(VCC_net), .I3(n38845), .O(n1026)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_632_9_lut.LUT_INIT = 16'h8228;
    SB_LUT4 add_236_25_lut (.I0(GND_net), .I1(encoder1_position[26]), .I2(GND_net), 
            .I3(n38499), .O(encoder1_position_scaled_23__N_75[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_236_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_157_28_lut (.I0(GND_net), .I1(delay_counter[26]), .I2(GND_net), 
            .I3(n38471), .O(n1302)) /* synthesis syn_instantiated=1 */ ;
    defparam add_157_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_157_28 (.CI(n38471), .I0(delay_counter[26]), .I1(GND_net), 
            .CO(n38472));
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_13 (.CI(n39503), 
            .I0(GND_net), .I1(n22_adj_5431), .CO(n39504));
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_12_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n23_adj_5432), .I3(n39502), .O(n23_adj_5292)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_12 (.CI(n39502), 
            .I0(GND_net), .I1(n23_adj_5432), .CO(n39503));
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_11_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n24_adj_5433), .I3(n39501), .O(n24_adj_5291)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_11 (.CI(n39501), 
            .I0(GND_net), .I1(n24_adj_5433), .CO(n39502));
    SB_LUT4 unary_minus_19_add_3_20_lut (.I0(GND_net), .I1(GND_net), .I2(n7), 
            .I3(n38548), .O(n345)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_19_add_3_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_236_24_lut (.I0(GND_net), .I1(encoder1_position[25]), .I2(GND_net), 
            .I3(n38498), .O(encoder1_position_scaled_23__N_75[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_236_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_632_8_lut (.I0(GND_net), .I1(n928), 
            .I2(VCC_net), .I3(n38844), .O(n995)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_632_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_632_8 (.CI(n38844), .I0(n928), 
            .I1(VCC_net), .CO(n38845));
    SB_LUT4 encoder0_position_31__I_0_add_632_7_lut (.I0(GND_net), .I1(n929), 
            .I2(GND_net), .I3(n38843), .O(n996)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_632_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_10_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n25_adj_5434), .I3(n39500), .O(n25_adj_5290)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_10 (.CI(n39500), 
            .I0(GND_net), .I1(n25_adj_5434), .CO(n39501));
    SB_CARRY unary_minus_19_add_3_20 (.CI(n38548), .I0(GND_net), .I1(n7), 
            .CO(n38549));
    SB_LUT4 add_157_27_lut (.I0(GND_net), .I1(delay_counter[25]), .I2(GND_net), 
            .I3(n38470), .O(n1303)) /* synthesis syn_instantiated=1 */ ;
    defparam add_157_27_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_9_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n26_adj_5435), .I3(n39499), .O(n26)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_157_27 (.CI(n38470), .I0(delay_counter[25]), .I1(GND_net), 
            .CO(n38471));
    SB_LUT4 unary_minus_19_add_3_19_lut (.I0(GND_net), .I1(GND_net), .I2(n8_adj_5257), 
            .I3(n38547), .O(n346)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_19_add_3_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_632_7 (.CI(n38843), .I0(n929), 
            .I1(GND_net), .CO(n38844));
    SB_LUT4 encoder0_position_31__I_0_add_632_6_lut (.I0(GND_net), .I1(n930), 
            .I2(GND_net), .I3(n38842), .O(n997)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_632_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_9 (.CI(n39499), 
            .I0(GND_net), .I1(n26_adj_5435), .CO(n39500));
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_8_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n27_adj_5436), .I3(n39498), .O(n27)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_8 (.CI(n39498), 
            .I0(GND_net), .I1(n27_adj_5436), .CO(n39499));
    SB_CARRY unary_minus_19_add_3_19 (.CI(n38547), .I0(GND_net), .I1(n8_adj_5257), 
            .CO(n38548));
    SB_CARRY add_236_24 (.CI(n38498), .I0(encoder1_position[25]), .I1(GND_net), 
            .CO(n38499));
    SB_CARRY encoder0_position_31__I_0_add_632_6 (.CI(n38842), .I0(n930), 
            .I1(GND_net), .CO(n38843));
    SB_LUT4 encoder0_position_31__I_0_add_632_5_lut (.I0(GND_net), .I1(n931), 
            .I2(VCC_net), .I3(n38841), .O(n998)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_632_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15070_3_lut (.I0(\data_out_frame[13] [1]), .I1(setpoint[9]), 
            .I2(n24278), .I3(GND_net), .O(n29018));   // verilog/coms.v(128[12] 303[6])
    defparam i15070_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15129_3_lut (.I0(\data_out_frame[10] [5]), .I1(encoder1_position_scaled[13]), 
            .I2(n24278), .I3(GND_net), .O(n29077));   // verilog/coms.v(128[12] 303[6])
    defparam i15129_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15130_3_lut (.I0(\data_out_frame[10] [4]), .I1(encoder1_position_scaled[12]), 
            .I2(n24278), .I3(GND_net), .O(n29078));   // verilog/coms.v(128[12] 303[6])
    defparam i15130_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15131_3_lut (.I0(\data_out_frame[10] [3]), .I1(encoder1_position_scaled[11]), 
            .I2(n24278), .I3(GND_net), .O(n29079));   // verilog/coms.v(128[12] 303[6])
    defparam i15131_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15132_3_lut (.I0(\data_out_frame[10] [2]), .I1(encoder1_position_scaled[10]), 
            .I2(n24278), .I3(GND_net), .O(n29080));   // verilog/coms.v(128[12] 303[6])
    defparam i15132_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 RX_I_0_1_lut (.I0(RX_c), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(RX_N_10));   // verilog/TinyFPGA_B.v(261[10:13])
    defparam RX_I_0_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_i1641_3_lut (.I0(n2414), .I1(n2481), 
            .I2(n2445), .I3(GND_net), .O(n2513));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1641_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1640_3_lut (.I0(n2413), .I1(n2480), 
            .I2(n2445), .I3(GND_net), .O(n2512));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1640_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1644_3_lut (.I0(n2417), .I1(n2484), 
            .I2(n2445), .I3(GND_net), .O(n2516));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1644_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_632_5 (.CI(n38841), .I0(n931), 
            .I1(VCC_net), .CO(n38842));
    SB_LUT4 i15133_3_lut (.I0(\data_out_frame[10] [1]), .I1(encoder1_position_scaled[9]), 
            .I2(n24278), .I3(GND_net), .O(n29081));   // verilog/coms.v(128[12] 303[6])
    defparam i15133_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFESR GLA_193 (.Q(INLA_c_0), .C(CLK_c), .E(n28482), .D(GLA_N_408), 
            .R(n28835));   // verilog/TinyFPGA_B.v(144[9] 223[5])
    SB_LUT4 i15134_3_lut (.I0(\data_out_frame[10] [0]), .I1(encoder1_position_scaled[8]), 
            .I2(n24278), .I3(GND_net), .O(n29082));   // verilog/coms.v(128[12] 303[6])
    defparam i15134_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_add_632_4_lut (.I0(GND_net), .I1(n932), 
            .I2(GND_net), .I3(n38840), .O(n999)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_632_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15135_3_lut (.I0(\data_out_frame[9] [7]), .I1(encoder1_position_scaled[23]), 
            .I2(n24278), .I3(GND_net), .O(n29083));   // verilog/coms.v(128[12] 303[6])
    defparam i15135_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i1643_3_lut (.I0(n2416), .I1(n2483), 
            .I2(n2445), .I3(GND_net), .O(n2515));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1643_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15136_3_lut (.I0(\data_out_frame[9] [6]), .I1(encoder1_position_scaled[22]), 
            .I2(n24278), .I3(GND_net), .O(n29084));   // verilog/coms.v(128[12] 303[6])
    defparam i15136_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i1642_3_lut (.I0(n2415), .I1(n2482), 
            .I2(n2445), .I3(GND_net), .O(n2514));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1642_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_7_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n28_adj_5437), .I3(n39497), .O(n28)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1659_3_lut (.I0(n2432), .I1(n2499), 
            .I2(n2445), .I3(GND_net), .O(n2531));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1659_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_7 (.CI(n39497), 
            .I0(GND_net), .I1(n28_adj_5437), .CO(n39498));
    SB_LUT4 add_236_23_lut (.I0(GND_net), .I1(encoder1_position[24]), .I2(GND_net), 
            .I3(n38497), .O(encoder1_position_scaled_23__N_75[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_236_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_6_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n29_adj_5438), .I3(n39496), .O(n29)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_19_add_3_18_lut (.I0(GND_net), .I1(GND_net), .I2(n9), 
            .I3(n38546), .O(n347)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_19_add_3_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_19_add_3_18 (.CI(n38546), .I0(GND_net), .I1(n9), 
            .CO(n38547));
    SB_CARRY add_236_23 (.CI(n38497), .I0(encoder1_position[24]), .I1(GND_net), 
            .CO(n38498));
    SB_CARRY encoder0_position_31__I_0_add_632_4 (.CI(n38840), .I0(n932), 
            .I1(GND_net), .CO(n38841));
    SB_LUT4 encoder0_position_31__I_0_add_632_3_lut (.I0(GND_net), .I1(n933), 
            .I2(VCC_net), .I3(n38839), .O(n1000)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_632_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_632_3 (.CI(n38839), .I0(n933), 
            .I1(VCC_net), .CO(n38840));
    SB_LUT4 encoder0_position_31__I_0_add_632_2_lut (.I0(GND_net), .I1(n520), 
            .I2(GND_net), .I3(VCC_net), .O(n1001)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_632_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_6 (.CI(n39496), 
            .I0(GND_net), .I1(n29_adj_5438), .CO(n39497));
    SB_LUT4 add_157_26_lut (.I0(GND_net), .I1(delay_counter[24]), .I2(GND_net), 
            .I3(n38469), .O(n1304)) /* synthesis syn_instantiated=1 */ ;
    defparam add_157_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_632_2 (.CI(VCC_net), .I0(n520), 
            .I1(GND_net), .CO(n38839));
    SB_LUT4 i15137_3_lut (.I0(\data_out_frame[9] [5]), .I1(encoder1_position_scaled[21]), 
            .I2(n24278), .I3(GND_net), .O(n29085));   // verilog/coms.v(128[12] 303[6])
    defparam i15137_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_add_565_8_lut (.I0(n861), .I1(n828), 
            .I2(VCC_net), .I3(n38838), .O(n927)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_565_8_lut.LUT_INIT = 16'h8228;
    SB_LUT4 unary_minus_19_add_3_17_lut (.I0(GND_net), .I1(GND_net), .I2(n10), 
            .I3(n38545), .O(n348)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_19_add_3_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_565_7_lut (.I0(GND_net), .I1(n829), 
            .I2(GND_net), .I3(n38837), .O(n896)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_565_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_19_add_3_17 (.CI(n38545), .I0(GND_net), .I1(n10), 
            .CO(n38546));
    SB_CARRY encoder0_position_31__I_0_add_565_7 (.CI(n38837), .I0(n829), 
            .I1(GND_net), .CO(n38838));
    SB_LUT4 encoder0_position_31__I_0_add_565_6_lut (.I0(GND_net), .I1(n830), 
            .I2(GND_net), .I3(n38836), .O(n897)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_565_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_565_6 (.CI(n38836), .I0(n830), 
            .I1(GND_net), .CO(n38837));
    SB_LUT4 encoder0_position_31__I_0_add_565_5_lut (.I0(GND_net), .I1(n831), 
            .I2(VCC_net), .I3(n38835), .O(n898)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_565_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1658_3_lut (.I0(n2431), .I1(n2498), 
            .I2(n2445), .I3(GND_net), .O(n2530));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1658_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_565_5 (.CI(n38835), .I0(n831), 
            .I1(VCC_net), .CO(n38836));
    SB_LUT4 i15138_3_lut (.I0(\data_out_frame[9] [4]), .I1(encoder1_position_scaled[20]), 
            .I2(n24278), .I3(GND_net), .O(n29086));   // verilog/coms.v(128[12] 303[6])
    defparam i15138_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_add_565_4_lut (.I0(GND_net), .I1(n832), 
            .I2(GND_net), .I3(n38834), .O(n899)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_565_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_19_add_3_16_lut (.I0(GND_net), .I1(GND_net), .I2(n11_adj_5258), 
            .I3(n38544), .O(n349)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_19_add_3_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_565_4 (.CI(n38834), .I0(n832), 
            .I1(GND_net), .CO(n38835));
    SB_LUT4 encoder0_position_31__I_0_add_565_3_lut (.I0(GND_net), .I1(n833), 
            .I2(VCC_net), .I3(n38833), .O(n900)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_565_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_5_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n30_adj_5439), .I3(n39495), .O(n30)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_236_22_lut (.I0(GND_net), .I1(encoder1_position[23]), .I2(GND_net), 
            .I3(n38496), .O(encoder1_position_scaled_23__N_75[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_236_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_565_3 (.CI(n38833), .I0(n833), 
            .I1(VCC_net), .CO(n38834));
    SB_LUT4 encoder0_position_31__I_0_i1657_3_lut (.I0(n2430), .I1(n2497), 
            .I2(n2445), .I3(GND_net), .O(n2529));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1657_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15139_3_lut (.I0(\data_out_frame[9] [3]), .I1(encoder1_position_scaled[19]), 
            .I2(n24278), .I3(GND_net), .O(n29087));   // verilog/coms.v(128[12] 303[6])
    defparam i15139_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_add_565_2_lut (.I0(GND_net), .I1(n519), 
            .I2(GND_net), .I3(VCC_net), .O(n901)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_565_2_lut.LUT_INIT = 16'hC33C;
    SB_DFFESR GLB_195 (.Q(INLB_c_0), .C(CLK_c), .E(n28482), .D(GLB_N_422), 
            .R(n28835));   // verilog/TinyFPGA_B.v(144[9] 223[5])
    SB_CARRY encoder0_position_31__I_0_add_565_2 (.CI(VCC_net), .I0(n519), 
            .I1(GND_net), .CO(n38833));
    SB_LUT4 add_2723_7_lut (.I0(GND_net), .I1(n621), .I2(GND_net), .I3(n38832), 
            .O(n8408)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2723_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_5 (.CI(n39495), 
            .I0(GND_net), .I1(n30_adj_5439), .CO(n39496));
    SB_CARRY add_236_22 (.CI(n38496), .I0(encoder1_position[23]), .I1(GND_net), 
            .CO(n38497));
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_4_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n31_adj_5440), .I3(n39494), .O(n31)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_4 (.CI(n39494), 
            .I0(GND_net), .I1(n31_adj_5440), .CO(n39495));
    SB_LUT4 add_2723_6_lut (.I0(GND_net), .I1(n622), .I2(GND_net), .I3(n38831), 
            .O(n8409)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2723_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_236_21_lut (.I0(GND_net), .I1(encoder1_position[22]), .I2(GND_net), 
            .I3(n38495), .O(encoder1_position_scaled_23__N_75[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_236_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_236_21 (.CI(n38495), .I0(encoder1_position[22]), .I1(GND_net), 
            .CO(n38496));
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_3_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n32_adj_5441), .I3(n39493), .O(n32)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2723_6 (.CI(n38831), .I0(n622), .I1(GND_net), .CO(n38832));
    SB_LUT4 add_2723_5_lut (.I0(GND_net), .I1(n623), .I2(VCC_net), .I3(n38830), 
            .O(n8410)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2723_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_157_26 (.CI(n38469), .I0(delay_counter[24]), .I1(GND_net), 
            .CO(n38470));
    SB_CARRY add_2723_5 (.CI(n38830), .I0(n623), .I1(VCC_net), .CO(n38831));
    SB_CARRY unary_minus_19_add_3_16 (.CI(n38544), .I0(GND_net), .I1(n11_adj_5258), 
            .CO(n38545));
    SB_LUT4 add_2723_4_lut (.I0(GND_net), .I1(n516), .I2(GND_net), .I3(n38829), 
            .O(n8411)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2723_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2723_4 (.CI(n38829), .I0(n516), .I1(GND_net), .CO(n38830));
    SB_LUT4 i15140_3_lut (.I0(\data_out_frame[9] [2]), .I1(encoder1_position_scaled[18]), 
            .I2(n24278), .I3(GND_net), .O(n29088));   // verilog/coms.v(128[12] 303[6])
    defparam i15140_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_3 (.CI(n39493), 
            .I0(GND_net), .I1(n32_adj_5441), .CO(n39494));
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_2_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n33_adj_5442), .I3(VCC_net), .O(n33)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_2 (.CI(VCC_net), 
            .I0(GND_net), .I1(n33_adj_5442), .CO(n39493));
    SB_LUT4 add_2723_3_lut (.I0(GND_net), .I1(n517), .I2(VCC_net), .I3(n38828), 
            .O(n8412)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2723_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2723_3 (.CI(n38828), .I0(n517), .I1(VCC_net), .CO(n38829));
    SB_LUT4 i15141_3_lut (.I0(\data_out_frame[9] [1]), .I1(encoder1_position_scaled[17]), 
            .I2(n24278), .I3(GND_net), .O(n29089));   // verilog/coms.v(128[12] 303[6])
    defparam i15141_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_236_20_lut (.I0(GND_net), .I1(encoder1_position[21]), .I2(GND_net), 
            .I3(n38494), .O(encoder1_position_scaled_23__N_75[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_236_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_19_add_3_15_lut (.I0(GND_net), .I1(GND_net), .I2(n12), 
            .I3(n38543), .O(n350)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_19_add_3_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_19_add_3_15 (.CI(n38543), .I0(GND_net), .I1(n12), 
            .CO(n38544));
    SB_LUT4 add_2723_2_lut (.I0(GND_net), .I1(n731), .I2(GND_net), .I3(VCC_net), 
            .O(n8413)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2723_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2723_2 (.CI(VCC_net), .I0(n731), .I1(GND_net), .CO(n38828));
    SB_LUT4 encoder0_position_31__I_0_i1646_3_lut (.I0(n2419), .I1(n2486), 
            .I2(n2445), .I3(GND_net), .O(n2518));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1646_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_1006_25_lut (.I0(GND_net), .I1(n4700), .I2(n2), .I3(n38675), 
            .O(n4485)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1006_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_236_20 (.CI(n38494), .I0(encoder1_position[21]), .I1(GND_net), 
            .CO(n38495));
    SB_LUT4 encoder0_position_31__I_0_i1645_3_lut (.I0(n2418), .I1(n2485), 
            .I2(n2445), .I3(GND_net), .O(n2517));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1645_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_1006_24_lut (.I0(GND_net), .I1(n4701), .I2(n2), .I3(n38674), 
            .O(n4486)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1006_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_157_25_lut (.I0(GND_net), .I1(delay_counter[23]), .I2(GND_net), 
            .I3(n38468), .O(n1305)) /* synthesis syn_instantiated=1 */ ;
    defparam add_157_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_236_19_lut (.I0(GND_net), .I1(encoder1_position[20]), .I2(GND_net), 
            .I3(n38493), .O(encoder1_position_scaled_23__N_75[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_236_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1006_24 (.CI(n38674), .I0(n4701), .I1(n2), .CO(n38675));
    SB_LUT4 unary_minus_19_add_3_14_lut (.I0(GND_net), .I1(GND_net), .I2(n13), 
            .I3(n38542), .O(n351)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_19_add_3_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_19_add_3_14 (.CI(n38542), .I0(GND_net), .I1(n13), 
            .CO(n38543));
    SB_LUT4 unary_minus_19_add_3_13_lut (.I0(GND_net), .I1(GND_net), .I2(n14_adj_5259), 
            .I3(n38541), .O(n352)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_19_add_3_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_157_25 (.CI(n38468), .I0(delay_counter[23]), .I1(GND_net), 
            .CO(n38469));
    SB_LUT4 add_1006_23_lut (.I0(GND_net), .I1(n4702), .I2(n2), .I3(n38673), 
            .O(n4487)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1006_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1006_23 (.CI(n38673), .I0(n4702), .I1(n2), .CO(n38674));
    SB_LUT4 add_1006_22_lut (.I0(GND_net), .I1(n4703), .I2(n2), .I3(n38672), 
            .O(n4488)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1006_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_157_24_lut (.I0(GND_net), .I1(delay_counter[22]), .I2(GND_net), 
            .I3(n38467), .O(n1306)) /* synthesis syn_instantiated=1 */ ;
    defparam add_157_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_19_add_3_13 (.CI(n38541), .I0(GND_net), .I1(n14_adj_5259), 
            .CO(n38542));
    SB_CARRY add_236_19 (.CI(n38493), .I0(encoder1_position[20]), .I1(GND_net), 
            .CO(n38494));
    SB_LUT4 add_236_18_lut (.I0(GND_net), .I1(encoder1_position[19]), .I2(GND_net), 
            .I3(n38492), .O(encoder1_position_scaled_23__N_75[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_236_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1006_22 (.CI(n38672), .I0(n4703), .I1(n2), .CO(n38673));
    SB_LUT4 unary_minus_19_add_3_12_lut (.I0(GND_net), .I1(GND_net), .I2(n15_adj_5260), 
            .I3(n38540), .O(n353)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_19_add_3_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15142_3_lut (.I0(\data_out_frame[9] [0]), .I1(encoder1_position_scaled[16]), 
            .I2(n24278), .I3(GND_net), .O(n29090));   // verilog/coms.v(128[12] 303[6])
    defparam i15142_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_157_24 (.CI(n38467), .I0(delay_counter[22]), .I1(GND_net), 
            .CO(n38468));
    SB_CARRY unary_minus_19_add_3_12 (.CI(n38540), .I0(GND_net), .I1(n15_adj_5260), 
            .CO(n38541));
    SB_LUT4 unary_minus_19_add_3_11_lut (.I0(GND_net), .I1(GND_net), .I2(n16_adj_5261), 
            .I3(n38539), .O(n354)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_19_add_3_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_17_inv_0_i3_1_lut (.I0(current[2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_5254));   // verilog/TinyFPGA_B.v(122[16:24])
    defparam unary_minus_17_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i15143_3_lut (.I0(\data_out_frame[8] [7]), .I1(encoder0_position_scaled[7]), 
            .I2(n24278), .I3(GND_net), .O(n29091));   // verilog/coms.v(128[12] 303[6])
    defparam i15143_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_1006_21_lut (.I0(GND_net), .I1(n4704), .I2(n2), .I3(n38671), 
            .O(n4489)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1006_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1655_3_lut (.I0(n2428), .I1(n2495), 
            .I2(n2445), .I3(GND_net), .O(n2527));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1655_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_1006_21 (.CI(n38671), .I0(n4704), .I1(n2), .CO(n38672));
    SB_LUT4 add_1006_20_lut (.I0(GND_net), .I1(n4705), .I2(n2), .I3(n38670), 
            .O(n4490)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1006_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1006_20 (.CI(n38670), .I0(n4705), .I1(n2), .CO(n38671));
    SB_LUT4 add_157_23_lut (.I0(GND_net), .I1(delay_counter[21]), .I2(GND_net), 
            .I3(n38466), .O(n1307)) /* synthesis syn_instantiated=1 */ ;
    defparam add_157_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_19_add_3_11 (.CI(n38539), .I0(GND_net), .I1(n16_adj_5261), 
            .CO(n38540));
    SB_LUT4 i15144_3_lut (.I0(\data_out_frame[8] [6]), .I1(encoder0_position_scaled[6]), 
            .I2(n24278), .I3(GND_net), .O(n29092));   // verilog/coms.v(128[12] 303[6])
    defparam i15144_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_1006_19_lut (.I0(GND_net), .I1(n4706), .I2(n2), .I3(n38669), 
            .O(n4491)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1006_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_19_add_3_10_lut (.I0(GND_net), .I1(GND_net), .I2(n17_adj_5262), 
            .I3(n38538), .O(n355)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_19_add_3_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_19_add_3_10 (.CI(n38538), .I0(GND_net), .I1(n17_adj_5262), 
            .CO(n38539));
    SB_CARRY add_1006_19 (.CI(n38669), .I0(n4706), .I1(n2), .CO(n38670));
    SB_CARRY add_236_18 (.CI(n38492), .I0(encoder1_position[19]), .I1(GND_net), 
            .CO(n38493));
    SB_LUT4 add_1006_18_lut (.I0(GND_net), .I1(n4707), .I2(n2), .I3(n38668), 
            .O(n4492)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1006_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_236_17_lut (.I0(GND_net), .I1(encoder1_position[18]), .I2(GND_net), 
            .I3(n38491), .O(encoder1_position_scaled_23__N_75[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_236_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_236_17 (.CI(n38491), .I0(encoder1_position[18]), .I1(GND_net), 
            .CO(n38492));
    SB_LUT4 i15145_3_lut (.I0(\data_out_frame[8] [5]), .I1(encoder0_position_scaled[5]), 
            .I2(n24278), .I3(GND_net), .O(n29093));   // verilog/coms.v(128[12] 303[6])
    defparam i15145_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_157_23 (.CI(n38466), .I0(delay_counter[21]), .I1(GND_net), 
            .CO(n38467));
    SB_CARRY add_1006_18 (.CI(n38668), .I0(n4707), .I1(n2), .CO(n38669));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_25_lut (.I0(GND_net), .I1(encoder0_position_scaled[23]), 
            .I2(n2_adj_5278), .I3(n38811), .O(displacement_23__N_99[23])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1649_3_lut (.I0(n2422), .I1(n2489), 
            .I2(n2445), .I3(GND_net), .O(n2521));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1649_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_24_lut (.I0(GND_net), .I1(encoder0_position_scaled[22]), 
            .I2(n3_adj_5338), .I3(n38810), .O(displacement_23__N_99[22])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_24 (.CI(n38810), .I0(encoder0_position_scaled[22]), 
            .I1(n3_adj_5338), .CO(n38811));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_23_lut (.I0(GND_net), .I1(encoder0_position_scaled[21]), 
            .I2(n4_adj_5337), .I3(n38809), .O(displacement_23__N_99[21])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_19_add_3_9_lut (.I0(GND_net), .I1(GND_net), .I2(n18_adj_5263), 
            .I3(n38537), .O(n356)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_19_add_3_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_23 (.CI(n38809), .I0(encoder0_position_scaled[21]), 
            .I1(n4_adj_5337), .CO(n38810));
    SB_LUT4 add_157_22_lut (.I0(GND_net), .I1(delay_counter[20]), .I2(GND_net), 
            .I3(n38465), .O(n1308)) /* synthesis syn_instantiated=1 */ ;
    defparam add_157_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_22_lut (.I0(GND_net), .I1(encoder0_position_scaled[20]), 
            .I2(n5_adj_5336), .I3(n38808), .O(displacement_23__N_99[20])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_157_8_lut (.I0(GND_net), .I1(delay_counter[6]), .I2(GND_net), 
            .I3(n38451), .O(n1322)) /* synthesis syn_instantiated=1 */ ;
    defparam add_157_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_1006_17_lut (.I0(GND_net), .I1(n4708), .I2(n2), .I3(n38667), 
            .O(n4493)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1006_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_22 (.CI(n38808), .I0(encoder0_position_scaled[20]), 
            .I1(n5_adj_5336), .CO(n38809));
    SB_CARRY add_157_22 (.CI(n38465), .I0(delay_counter[20]), .I1(GND_net), 
            .CO(n38466));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_21_lut (.I0(GND_net), .I1(encoder0_position_scaled[19]), 
            .I2(n6_adj_5335), .I3(n38807), .O(displacement_23__N_99[19])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1006_17 (.CI(n38667), .I0(n4708), .I1(n2), .CO(n38668));
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_21 (.CI(n38807), .I0(encoder0_position_scaled[19]), 
            .I1(n6_adj_5335), .CO(n38808));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_20_lut (.I0(GND_net), .I1(encoder0_position_scaled[18]), 
            .I2(n7_adj_5334), .I3(n38806), .O(displacement_23__N_99[18])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_236_16_lut (.I0(GND_net), .I1(encoder1_position[17]), .I2(GND_net), 
            .I3(n38490), .O(encoder1_position_scaled_23__N_75[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_236_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_236_16 (.CI(n38490), .I0(encoder1_position[17]), .I1(GND_net), 
            .CO(n38491));
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_20 (.CI(n38806), .I0(encoder0_position_scaled[18]), 
            .I1(n7_adj_5334), .CO(n38807));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_19_lut (.I0(GND_net), .I1(encoder0_position_scaled[17]), 
            .I2(n8_adj_5333), .I3(n38805), .O(displacement_23__N_99[17])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_19 (.CI(n38805), .I0(encoder0_position_scaled[17]), 
            .I1(n8_adj_5333), .CO(n38806));
    SB_CARRY unary_minus_19_add_3_9 (.CI(n38537), .I0(GND_net), .I1(n18_adj_5263), 
            .CO(n38538));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_18_lut (.I0(GND_net), .I1(encoder0_position_scaled[16]), 
            .I2(n9_adj_5332), .I3(n38804), .O(displacement_23__N_99[16])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_236_15_lut (.I0(GND_net), .I1(encoder1_position[16]), .I2(GND_net), 
            .I3(n38489), .O(encoder1_position_scaled_23__N_75[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_236_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_18 (.CI(n38804), .I0(encoder0_position_scaled[16]), 
            .I1(n9_adj_5332), .CO(n38805));
    SB_LUT4 add_1006_16_lut (.I0(GND_net), .I1(n4709), .I2(n2), .I3(n38666), 
            .O(n4494)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1006_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_17_lut (.I0(GND_net), .I1(encoder0_position_scaled[15]), 
            .I2(n10_adj_5331), .I3(n38803), .O(displacement_23__N_99[15])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_17 (.CI(n38803), .I0(encoder0_position_scaled[15]), 
            .I1(n10_adj_5331), .CO(n38804));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_16_lut (.I0(GND_net), .I1(encoder0_position_scaled[14]), 
            .I2(n11_adj_5330), .I3(n38802), .O(displacement_23__N_99[14])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_16 (.CI(n38802), .I0(encoder0_position_scaled[14]), 
            .I1(n11_adj_5330), .CO(n38803));
    SB_LUT4 unary_minus_19_add_3_8_lut (.I0(GND_net), .I1(GND_net), .I2(n19_adj_5264), 
            .I3(n38536), .O(n357)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_19_add_3_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_15_lut (.I0(GND_net), .I1(encoder0_position_scaled[13]), 
            .I2(n12_adj_5329), .I3(n38801), .O(displacement_23__N_99[13])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_15 (.CI(n38801), .I0(encoder0_position_scaled[13]), 
            .I1(n12_adj_5329), .CO(n38802));
    SB_CARRY unary_minus_19_add_3_8 (.CI(n38536), .I0(GND_net), .I1(n19_adj_5264), 
            .CO(n38537));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_14_lut (.I0(GND_net), .I1(encoder0_position_scaled[12]), 
            .I2(n13_adj_5328), .I3(n38800), .O(displacement_23__N_99[12])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_236_15 (.CI(n38489), .I0(encoder1_position[16]), .I1(GND_net), 
            .CO(n38490));
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_14 (.CI(n38800), .I0(encoder0_position_scaled[12]), 
            .I1(n13_adj_5328), .CO(n38801));
    SB_LUT4 i15146_3_lut (.I0(\data_out_frame[8] [4]), .I1(encoder0_position_scaled[4]), 
            .I2(n24278), .I3(GND_net), .O(n29094));   // verilog/coms.v(128[12] 303[6])
    defparam i15146_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15147_3_lut (.I0(\data_out_frame[8] [3]), .I1(encoder0_position_scaled[3]), 
            .I2(n24278), .I3(GND_net), .O(n29095));   // verilog/coms.v(128[12] 303[6])
    defparam i15147_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_13_lut (.I0(GND_net), .I1(encoder0_position_scaled[11]), 
            .I2(n14_adj_5327), .I3(n38799), .O(displacement_23__N_99[11])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_19_add_3_7_lut (.I0(GND_net), .I1(GND_net), .I2(n20_adj_5265), 
            .I3(n38535), .O(n358)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_19_add_3_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_13 (.CI(n38799), .I0(encoder0_position_scaled[11]), 
            .I1(n14_adj_5327), .CO(n38800));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_12_lut (.I0(GND_net), .I1(encoder0_position_scaled[10]), 
            .I2(n15_adj_5326), .I3(n38798), .O(displacement_23__N_99[10])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_12 (.CI(n38798), .I0(encoder0_position_scaled[10]), 
            .I1(n15_adj_5326), .CO(n38799));
    SB_LUT4 i15148_3_lut (.I0(\data_out_frame[8] [2]), .I1(encoder0_position_scaled[2]), 
            .I2(n24278), .I3(GND_net), .O(n29096));   // verilog/coms.v(128[12] 303[6])
    defparam i15148_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_11_lut (.I0(GND_net), .I1(encoder0_position_scaled[9]), 
            .I2(n16_adj_5325), .I3(n38797), .O(displacement_23__N_99[9])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_11 (.CI(n38797), .I0(encoder0_position_scaled[9]), 
            .I1(n16_adj_5325), .CO(n38798));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_10_lut (.I0(GND_net), .I1(encoder0_position_scaled[8]), 
            .I2(n17_adj_5324), .I3(n38796), .O(displacement_23__N_99[8])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_10 (.CI(n38796), .I0(encoder0_position_scaled[8]), 
            .I1(n17_adj_5324), .CO(n38797));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_9_lut (.I0(GND_net), .I1(encoder0_position_scaled[7]), 
            .I2(n18_adj_5323), .I3(n38795), .O(displacement_23__N_99[7])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_9 (.CI(n38795), .I0(encoder0_position_scaled[7]), 
            .I1(n18_adj_5323), .CO(n38796));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_8_lut (.I0(GND_net), .I1(encoder0_position_scaled[6]), 
            .I2(n19_adj_5322), .I3(n38794), .O(displacement_23__N_99[6])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_8 (.CI(n38794), .I0(encoder0_position_scaled[6]), 
            .I1(n19_adj_5322), .CO(n38795));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_7_lut (.I0(GND_net), .I1(encoder0_position_scaled[5]), 
            .I2(n20_adj_5320), .I3(n38793), .O(displacement_23__N_99[5])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_7 (.CI(n38793), .I0(encoder0_position_scaled[5]), 
            .I1(n20_adj_5320), .CO(n38794));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_6_lut (.I0(GND_net), .I1(encoder0_position_scaled[4]), 
            .I2(n21_adj_5319), .I3(n38792), .O(displacement_23__N_99[4])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_6 (.CI(n38792), .I0(encoder0_position_scaled[4]), 
            .I1(n21_adj_5319), .CO(n38793));
    SB_DFF ID_i0_i1 (.Q(ID[1]), .C(CLK_c), .D(n29536));   // verilog/TinyFPGA_B.v(375[10] 403[6])
    SB_DFF ID_i0_i2 (.Q(ID[2]), .C(CLK_c), .D(n29535));   // verilog/TinyFPGA_B.v(375[10] 403[6])
    SB_DFF ID_i0_i3 (.Q(ID[3]), .C(CLK_c), .D(n29534));   // verilog/TinyFPGA_B.v(375[10] 403[6])
    SB_LUT4 encoder0_position_31__I_0_i1648_3_lut (.I0(n2421), .I1(n2488), 
            .I2(n2445), .I3(GND_net), .O(n2520));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1648_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1647_3_lut (.I0(n2420), .I1(n2487), 
            .I2(n2445), .I3(GND_net), .O(n2519));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1647_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_5_lut (.I0(GND_net), .I1(encoder0_position_scaled[3]), 
            .I2(n22_adj_5317), .I3(n38791), .O(displacement_23__N_99[3])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_5 (.CI(n38791), .I0(encoder0_position_scaled[3]), 
            .I1(n22_adj_5317), .CO(n38792));
    SB_LUT4 encoder0_position_31__I_0_i1661_3_lut (.I0(n535), .I1(n2501), 
            .I2(n2445), .I3(GND_net), .O(n2533));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1661_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1660_3_lut (.I0(n2433), .I1(n2500), 
            .I2(n2445), .I3(GND_net), .O(n2532));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1660_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_4_lut (.I0(GND_net), .I1(encoder0_position_scaled[2]), 
            .I2(n23_adj_5316), .I3(n38790), .O(displacement_23__N_99[2])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_4 (.CI(n38790), .I0(encoder0_position_scaled[2]), 
            .I1(n23_adj_5316), .CO(n38791));
    SB_LUT4 encoder0_position_31__I_0_mux_3_i9_3_lut (.I0(encoder0_position[8]), 
            .I1(n25_adj_5290), .I2(encoder0_position[31]), .I3(GND_net), 
            .O(n950));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_mux_3_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_3_lut (.I0(GND_net), .I1(encoder0_position_scaled[1]), 
            .I2(n24_adj_5315), .I3(n38789), .O(displacement_23__N_99[1])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1656_3_lut (.I0(n2429), .I1(n2496), 
            .I2(n2445), .I3(GND_net), .O(n2528));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1656_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY unary_minus_19_add_3_7 (.CI(n38535), .I0(GND_net), .I1(n20_adj_5265), 
            .CO(n38536));
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_3 (.CI(n38789), .I0(encoder0_position_scaled[1]), 
            .I1(n24_adj_5315), .CO(n38790));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_2_lut (.I0(GND_net), .I1(encoder0_position_scaled[0]), 
            .I2(n25_adj_5314), .I3(VCC_net), .O(displacement_23__N_99[0])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_2 (.CI(VCC_net), .I0(encoder0_position_scaled[0]), 
            .I1(n25_adj_5314), .CO(n38789));
    SB_LUT4 unary_minus_17_add_3_15_lut (.I0(GND_net), .I1(GND_net), .I2(n2), 
            .I3(n38788), .O(n321)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_17_add_3_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_17_add_3_14_lut (.I0(GND_net), .I1(GND_net), .I2(n2), 
            .I3(n38787), .O(n325)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_17_add_3_14_lut.LUT_INIT = 16'hC33C;
    SB_DFF ID_i0_i4 (.Q(ID[4]), .C(CLK_c), .D(n29533));   // verilog/TinyFPGA_B.v(375[10] 403[6])
    SB_DFF ID_i0_i5 (.Q(ID[5]), .C(CLK_c), .D(n29532));   // verilog/TinyFPGA_B.v(375[10] 403[6])
    SB_DFF ID_i0_i6 (.Q(ID[6]), .C(CLK_c), .D(n29531));   // verilog/TinyFPGA_B.v(375[10] 403[6])
    SB_CARRY unary_minus_17_add_3_14 (.CI(n38787), .I0(GND_net), .I1(n2), 
            .CO(n38788));
    SB_LUT4 unary_minus_17_add_3_13_lut (.I0(GND_net), .I1(GND_net), .I2(n14_adj_5250), 
            .I3(n38786), .O(n326)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_17_add_3_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_17_add_3_13 (.CI(n38786), .I0(GND_net), .I1(n14_adj_5250), 
            .CO(n38787));
    SB_LUT4 add_236_14_lut (.I0(GND_net), .I1(encoder1_position[15]), .I2(GND_net), 
            .I3(n38488), .O(encoder1_position_scaled_23__N_75[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_236_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_17_add_3_12_lut (.I0(GND_net), .I1(GND_net), .I2(n15_adj_5251), 
            .I3(n38785), .O(n327)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_17_add_3_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_17_add_3_12 (.CI(n38785), .I0(GND_net), .I1(n15_adj_5251), 
            .CO(n38786));
    SB_LUT4 unary_minus_17_add_3_11_lut (.I0(GND_net), .I1(GND_net), .I2(n16_adj_5252), 
            .I3(n38784), .O(n328)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_17_add_3_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15149_3_lut (.I0(\data_out_frame[8] [1]), .I1(encoder0_position_scaled[1]), 
            .I2(n24278), .I3(GND_net), .O(n29097));   // verilog/coms.v(128[12] 303[6])
    defparam i15149_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15150_3_lut (.I0(\data_out_frame[8] [0]), .I1(encoder0_position_scaled[0]), 
            .I2(n24278), .I3(GND_net), .O(n29098));   // verilog/coms.v(128[12] 303[6])
    defparam i15150_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15151_3_lut (.I0(\data_out_frame[7] [7]), .I1(encoder0_position_scaled[15]), 
            .I2(n24278), .I3(GND_net), .O(n29099));   // verilog/coms.v(128[12] 303[6])
    defparam i15151_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15152_3_lut (.I0(\data_out_frame[7] [6]), .I1(encoder0_position_scaled[14]), 
            .I2(n24278), .I3(GND_net), .O(n29100));   // verilog/coms.v(128[12] 303[6])
    defparam i15152_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY unary_minus_17_add_3_11 (.CI(n38784), .I0(GND_net), .I1(n16_adj_5252), 
            .CO(n38785));
    SB_LUT4 unary_minus_17_add_3_10_lut (.I0(GND_net), .I1(GND_net), .I2(n17_adj_5253), 
            .I3(n38783), .O(n329)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_17_add_3_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_17_add_3_10 (.CI(n38783), .I0(GND_net), .I1(n17_adj_5253), 
            .CO(n38784));
    SB_LUT4 i15153_3_lut (.I0(\data_out_frame[7] [5]), .I1(encoder0_position_scaled[13]), 
            .I2(n24278), .I3(GND_net), .O(n29101));   // verilog/coms.v(128[12] 303[6])
    defparam i15153_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_17_add_3_9_lut (.I0(GND_net), .I1(GND_net), .I2(n18), 
            .I3(n38782), .O(n330)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_17_add_3_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15154_3_lut (.I0(\data_out_frame[7] [4]), .I1(encoder0_position_scaled[12]), 
            .I2(n24278), .I3(GND_net), .O(n29102));   // verilog/coms.v(128[12] 303[6])
    defparam i15154_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF ID_i0_i7 (.Q(ID[7]), .C(CLK_c), .D(n29530));   // verilog/TinyFPGA_B.v(375[10] 403[6])
    SB_CARRY unary_minus_17_add_3_9 (.CI(n38782), .I0(GND_net), .I1(n18), 
            .CO(n38783));
    SB_LUT4 i34446_3_lut (.I0(n2325), .I1(n2392), .I2(n2346), .I3(GND_net), 
            .O(n2424));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam i34446_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i34447_3_lut (.I0(n2424), .I1(n2491), .I2(n2445), .I3(GND_net), 
            .O(n2523));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam i34447_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i34450_3_lut (.I0(n2327), .I1(n2394), .I2(n2346), .I3(GND_net), 
            .O(n2426));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam i34450_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 unary_minus_17_add_3_8_lut (.I0(GND_net), .I1(GND_net), .I2(n19), 
            .I3(n38781), .O(n331)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_17_add_3_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_17_add_3_8 (.CI(n38781), .I0(GND_net), .I1(n19), 
            .CO(n38782));
    SB_LUT4 unary_minus_17_add_3_7_lut (.I0(GND_net), .I1(GND_net), .I2(n20), 
            .I3(n38780), .O(n332)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_17_add_3_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_17_add_3_7 (.CI(n38780), .I0(GND_net), .I1(n20), 
            .CO(n38781));
    SB_LUT4 unary_minus_17_add_3_6_lut (.I0(GND_net), .I1(GND_net), .I2(n21), 
            .I3(n38779), .O(n333)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_17_add_3_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_17_add_3_6 (.CI(n38779), .I0(GND_net), .I1(n21), 
            .CO(n38780));
    SB_LUT4 unary_minus_17_add_3_5_lut (.I0(GND_net), .I1(GND_net), .I2(n22), 
            .I3(n38778), .O(n334)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_17_add_3_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_17_add_3_5 (.CI(n38778), .I0(GND_net), .I1(n22), 
            .CO(n38779));
    SB_LUT4 unary_minus_17_add_3_4_lut (.I0(GND_net), .I1(GND_net), .I2(n23_adj_5254), 
            .I3(n38777), .O(n335)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_17_add_3_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_17_add_3_4 (.CI(n38777), .I0(GND_net), .I1(n23_adj_5254), 
            .CO(n38778));
    SB_LUT4 i34451_3_lut (.I0(n2426), .I1(n2493), .I2(n2445), .I3(GND_net), 
            .O(n2525));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam i34451_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 unary_minus_17_add_3_3_lut (.I0(GND_net), .I1(GND_net), .I2(n24), 
            .I3(n38776), .O(n336)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_17_add_3_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i34452_3_lut (.I0(n2328), .I1(n2395), .I2(n2346), .I3(GND_net), 
            .O(n2427));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam i34452_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY unary_minus_17_add_3_3 (.CI(n38776), .I0(GND_net), .I1(n24), 
            .CO(n38777));
    SB_LUT4 unary_minus_17_add_3_2_lut (.I0(n25), .I1(GND_net), .I2(n4698), 
            .I3(VCC_net), .O(n49289)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_17_add_3_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY unary_minus_17_add_3_2 (.CI(VCC_net), .I0(GND_net), .I1(n4698), 
            .CO(n38776));
    SB_CARRY add_1006_16 (.CI(n38666), .I0(n4709), .I1(n2), .CO(n38667));
    SB_CARRY add_236_14 (.CI(n38488), .I0(encoder1_position[15]), .I1(GND_net), 
            .CO(n38489));
    SB_LUT4 unary_minus_19_add_3_6_lut (.I0(GND_net), .I1(GND_net), .I2(n21_adj_5266), 
            .I3(n38534), .O(n359)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_19_add_3_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_236_13_lut (.I0(GND_net), .I1(encoder1_position[14]), .I2(GND_net), 
            .I3(n38487), .O(encoder1_position_scaled_23__N_75[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_236_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_157_21_lut (.I0(GND_net), .I1(delay_counter[19]), .I2(GND_net), 
            .I3(n38464), .O(n1309)) /* synthesis syn_instantiated=1 */ ;
    defparam add_157_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_1006_15_lut (.I0(GND_net), .I1(n4710), .I2(n2), .I3(n38665), 
            .O(n4495)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1006_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_19_add_3_6 (.CI(n38534), .I0(GND_net), .I1(n21_adj_5266), 
            .CO(n38535));
    SB_CARRY add_1006_15 (.CI(n38665), .I0(n4710), .I1(n2), .CO(n38666));
    SB_CARRY add_157_21 (.CI(n38464), .I0(delay_counter[19]), .I1(GND_net), 
            .CO(n38465));
    SB_CARRY add_236_13 (.CI(n38487), .I0(encoder1_position[14]), .I1(GND_net), 
            .CO(n38488));
    SB_LUT4 add_236_12_lut (.I0(GND_net), .I1(encoder1_position[13]), .I2(GND_net), 
            .I3(n38486), .O(encoder1_position_scaled_23__N_75[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_236_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_19_add_3_5_lut (.I0(GND_net), .I1(GND_net), .I2(n22_adj_5267), 
            .I3(n38533), .O(n360)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_19_add_3_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_157_20_lut (.I0(GND_net), .I1(delay_counter[18]), .I2(GND_net), 
            .I3(n38463), .O(n1310)) /* synthesis syn_instantiated=1 */ ;
    defparam add_157_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_1006_14_lut (.I0(GND_net), .I1(n4711), .I2(n2), .I3(n38664), 
            .O(n4496)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1006_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_157_20 (.CI(n38463), .I0(delay_counter[18]), .I1(GND_net), 
            .CO(n38464));
    SB_LUT4 add_157_19_lut (.I0(GND_net), .I1(delay_counter[17]), .I2(GND_net), 
            .I3(n38462), .O(n1311)) /* synthesis syn_instantiated=1 */ ;
    defparam add_157_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_157_19 (.CI(n38462), .I0(delay_counter[17]), .I1(GND_net), 
            .CO(n38463));
    SB_CARRY unary_minus_19_add_3_5 (.CI(n38533), .I0(GND_net), .I1(n22_adj_5267), 
            .CO(n38534));
    SB_DFF \ID_READOUT_FSM.state__i1  (.Q(\ID_READOUT_FSM.state [1]), .C(CLK_c), 
           .D(n17_adj_5271));   // verilog/TinyFPGA_B.v(375[10] 403[6])
    SB_DFF commutation_state_i1 (.Q(commutation_state[1]), .C(CLK_c), .D(n43630));   // verilog/TinyFPGA_B.v(144[9] 223[5])
    SB_CARRY add_1006_14 (.CI(n38664), .I0(n4711), .I1(n2), .CO(n38665));
    SB_DFF commutation_state_i2 (.Q(commutation_state[2]), .C(CLK_c), .D(n44694));   // verilog/TinyFPGA_B.v(144[9] 223[5])
    SB_LUT4 unary_minus_19_add_3_4_lut (.I0(GND_net), .I1(GND_net), .I2(n23_adj_5268), 
            .I3(n38532), .O(n361)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_19_add_3_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_1006_13_lut (.I0(GND_net), .I1(n4712), .I2(n14_adj_5250), 
            .I3(n38663), .O(n4497)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1006_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_19_add_3_4 (.CI(n38532), .I0(GND_net), .I1(n23_adj_5268), 
            .CO(n38533));
    SB_CARRY add_1006_13 (.CI(n38663), .I0(n4712), .I1(n14_adj_5250), 
            .CO(n38664));
    SB_LUT4 i15155_4_lut (.I0(CS_MISO_c), .I1(data_adj_5514[3]), .I2(n10_adj_5341), 
            .I3(n27180), .O(n29103));   // verilog/tli4970.v(35[10] 68[6])
    defparam i15155_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i34453_3_lut (.I0(n2427), .I1(n2494), .I2(n2445), .I3(GND_net), 
            .O(n2526));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam i34453_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_248_i1_3_lut_4_lut (.I0(n27015), .I1(control_mode[1]), .I2(motor_state_23__N_123[0]), 
            .I3(encoder0_position_scaled[0]), .O(motor_state[0]));   // verilog/TinyFPGA_B.v(284[5:22])
    defparam mux_248_i1_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 add_1006_12_lut (.I0(GND_net), .I1(n4713), .I2(n15_adj_5251), 
            .I3(n38662), .O(n4498)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1006_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15211_4_lut (.I0(state_7__N_4267[3]), .I1(data[0]), .I2(n10_adj_5410), 
            .I3(n27147), .O(n29159));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i15211_4_lut.LUT_INIT = 16'hccca;
    SB_CARRY add_1006_12 (.CI(n38662), .I0(n4713), .I1(n15_adj_5251), 
            .CO(n38663));
    SB_LUT4 i1_4_lut_adj_1850 (.I0(n2526), .I1(n2525), .I2(n2523), .I3(n2528), 
            .O(n46531));
    defparam i1_4_lut_adj_1850.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1851 (.I0(n2524), .I1(n2521), .I2(n2527), .I3(n2522), 
            .O(n46533));
    defparam i1_4_lut_adj_1851.LUT_INIT = 16'hfffe;
    SB_LUT4 i21454_3_lut (.I0(n950), .I1(n2532), .I2(n2533), .I3(GND_net), 
            .O(n35402));
    defparam i21454_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 add_1006_11_lut (.I0(GND_net), .I1(n4714), .I2(n16_adj_5252), 
            .I3(n38661), .O(n4499)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1006_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1006_11 (.CI(n38661), .I0(n4714), .I1(n16_adj_5252), 
            .CO(n38662));
    SB_LUT4 unary_minus_19_add_3_3_lut (.I0(GND_net), .I1(GND_net), .I2(n24_adj_5269), 
            .I3(n38531), .O(n362)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_19_add_3_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_19_add_3_3 (.CI(n38531), .I0(GND_net), .I1(n24_adj_5269), 
            .CO(n38532));
    SB_CARRY add_236_12 (.CI(n38486), .I0(encoder1_position[13]), .I1(GND_net), 
            .CO(n38487));
    SB_LUT4 add_1006_10_lut (.I0(GND_net), .I1(n4715), .I2(n17_adj_5253), 
            .I3(n38660), .O(n4500)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1006_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1852 (.I0(n2519), .I1(n2520), .I2(n46533), .I3(n46531), 
            .O(n46539));
    defparam i1_4_lut_adj_1852.LUT_INIT = 16'hfffe;
    SB_LUT4 mux_248_i2_3_lut_4_lut (.I0(n27015), .I1(control_mode[1]), .I2(motor_state_23__N_123[1]), 
            .I3(encoder0_position_scaled[1]), .O(motor_state[1]));   // verilog/TinyFPGA_B.v(284[5:22])
    defparam mux_248_i2_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 mux_248_i3_3_lut_4_lut (.I0(n27015), .I1(control_mode[1]), .I2(motor_state_23__N_123[2]), 
            .I3(encoder0_position_scaled[2]), .O(motor_state[2]));   // verilog/TinyFPGA_B.v(284[5:22])
    defparam mux_248_i3_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 i1_4_lut_adj_1853 (.I0(n2529), .I1(n35402), .I2(n2530), .I3(n2531), 
            .O(n44987));
    defparam i1_4_lut_adj_1853.LUT_INIT = 16'ha080;
    SB_LUT4 i15156_3_lut (.I0(\data_out_frame[7] [3]), .I1(encoder0_position_scaled[11]), 
            .I2(n24278), .I3(GND_net), .O(n29104));   // verilog/coms.v(128[12] 303[6])
    defparam i15156_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_248_i4_3_lut_4_lut (.I0(n27015), .I1(control_mode[1]), .I2(motor_state_23__N_123[3]), 
            .I3(encoder0_position_scaled[3]), .O(motor_state[3]));   // verilog/TinyFPGA_B.v(284[5:22])
    defparam mux_248_i4_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 i15680_3_lut (.I0(\data_out_frame[19] [5]), .I1(displacement[13]), 
            .I2(n24278), .I3(GND_net), .O(n29628));   // verilog/coms.v(128[12] 303[6])
    defparam i15680_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15681_3_lut (.I0(\data_out_frame[19] [4]), .I1(displacement[12]), 
            .I2(n24278), .I3(GND_net), .O(n29629));   // verilog/coms.v(128[12] 303[6])
    defparam i15681_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1854 (.I0(n2517), .I1(n44987), .I2(n2518), .I3(n46539), 
            .O(n46545));
    defparam i1_4_lut_adj_1854.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1855 (.I0(n2514), .I1(n2515), .I2(n2516), .I3(n46545), 
            .O(n46551));
    defparam i1_4_lut_adj_1855.LUT_INIT = 16'hfffe;
    SB_CARRY add_157_3 (.CI(n38446), .I0(delay_counter[1]), .I1(GND_net), 
            .CO(n38447));
    SB_LUT4 i35170_4_lut (.I0(n2512), .I1(n2511), .I2(n2513), .I3(n46551), 
            .O(n2544));
    defparam i35170_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 add_157_18_lut (.I0(GND_net), .I1(delay_counter[16]), .I2(GND_net), 
            .I3(n38461), .O(n1312)) /* synthesis syn_instantiated=1 */ ;
    defparam add_157_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1006_10 (.CI(n38660), .I0(n4715), .I1(n17_adj_5253), 
            .CO(n38661));
    SB_LUT4 unary_minus_17_inv_0_i4_1_lut (.I0(current[3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n22));   // verilog/TinyFPGA_B.v(122[16:24])
    defparam unary_minus_17_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_19_add_3_2_lut (.I0(GND_net), .I1(GND_net), .I2(n25), 
            .I3(VCC_net), .O(n363)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_19_add_3_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_1006_9_lut (.I0(GND_net), .I1(n4716), .I2(n18), .I3(n38659), 
            .O(n4501)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1006_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_157_8 (.CI(n38451), .I0(delay_counter[6]), .I1(GND_net), 
            .CO(n38452));
    SB_CARRY unary_minus_19_add_3_2 (.CI(VCC_net), .I0(GND_net), .I1(n25), 
            .CO(n38531));
    SB_CARRY add_1006_9 (.CI(n38659), .I0(n4716), .I1(n18), .CO(n38660));
    SB_LUT4 add_1006_8_lut (.I0(GND_net), .I1(n4717), .I2(n19), .I3(n38658), 
            .O(n4502)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1006_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_248_i5_3_lut_4_lut (.I0(n27015), .I1(control_mode[1]), .I2(motor_state_23__N_123[4]), 
            .I3(encoder0_position_scaled[4]), .O(motor_state[4]));   // verilog/TinyFPGA_B.v(284[5:22])
    defparam mux_248_i5_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 add_236_11_lut (.I0(GND_net), .I1(encoder1_position[12]), .I2(GND_net), 
            .I3(n38485), .O(encoder1_position_scaled_23__N_75[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_236_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_248_i6_3_lut_4_lut (.I0(n27015), .I1(control_mode[1]), .I2(motor_state_23__N_123[5]), 
            .I3(encoder0_position_scaled[5]), .O(motor_state[5]));   // verilog/TinyFPGA_B.v(284[5:22])
    defparam mux_248_i6_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_CARRY add_236_11 (.CI(n38485), .I0(encoder1_position[12]), .I1(GND_net), 
            .CO(n38486));
    SB_CARRY add_1006_8 (.CI(n38658), .I0(n4717), .I1(n19), .CO(n38659));
    SB_LUT4 mux_248_i7_3_lut_4_lut (.I0(n27015), .I1(control_mode[1]), .I2(motor_state_23__N_123[6]), 
            .I3(encoder0_position_scaled[6]), .O(motor_state[6]));   // verilog/TinyFPGA_B.v(284[5:22])
    defparam mux_248_i7_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 add_236_10_lut (.I0(GND_net), .I1(encoder1_position[11]), .I2(GND_net), 
            .I3(n38484), .O(encoder1_position_scaled_23__N_75[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_236_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_236_10 (.CI(n38484), .I0(encoder1_position[11]), .I1(GND_net), 
            .CO(n38485));
    SB_CARRY add_157_18 (.CI(n38461), .I0(delay_counter[16]), .I1(GND_net), 
            .CO(n38462));
    SB_LUT4 add_1006_7_lut (.I0(GND_net), .I1(n4718), .I2(n20), .I3(n38657), 
            .O(n4503)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1006_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_157_2_lut (.I0(GND_net), .I1(delay_counter[0]), .I2(GND_net), 
            .I3(VCC_net), .O(n1328)) /* synthesis syn_instantiated=1 */ ;
    defparam add_157_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_157_7_lut (.I0(GND_net), .I1(delay_counter[5]), .I2(GND_net), 
            .I3(n38450), .O(n1323)) /* synthesis syn_instantiated=1 */ ;
    defparam add_157_7_lut.LUT_INIT = 16'hC33C;
    SB_DFFESR GLC_197 (.Q(INLC_c_0), .C(CLK_c), .E(n28482), .D(GLC_N_436), 
            .R(n28835));   // verilog/TinyFPGA_B.v(144[9] 223[5])
    SB_LUT4 i15682_3_lut (.I0(\data_out_frame[19] [3]), .I1(displacement[11]), 
            .I2(n24278), .I3(GND_net), .O(n29630));   // verilog/coms.v(128[12] 303[6])
    defparam i15682_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15216_4_lut (.I0(CS_MISO_c), .I1(data_adj_5514[8]), .I2(n6), 
            .I3(n27143), .O(n29164));   // verilog/tli4970.v(35[10] 68[6])
    defparam i15216_4_lut.LUT_INIT = 16'hccca;
    SB_CARRY add_1006_7 (.CI(n38657), .I0(n4718), .I1(n20), .CO(n38658));
    SB_CARRY add_157_7 (.CI(n38450), .I0(delay_counter[5]), .I1(GND_net), 
            .CO(n38451));
    SB_LUT4 add_157_17_lut (.I0(GND_net), .I1(delay_counter[15]), .I2(GND_net), 
            .I3(n38460), .O(n1313)) /* synthesis syn_instantiated=1 */ ;
    defparam add_157_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_157_17 (.CI(n38460), .I0(delay_counter[15]), .I1(GND_net), 
            .CO(n38461));
    SB_LUT4 add_1006_6_lut (.I0(GND_net), .I1(n4719), .I2(n21), .I3(n38656), 
            .O(n4504)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1006_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_236_9_lut (.I0(GND_net), .I1(encoder1_position[10]), .I2(GND_net), 
            .I3(n38483), .O(encoder1_position_scaled_23__N_75[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_236_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1006_6 (.CI(n38656), .I0(n4719), .I1(n21), .CO(n38657));
    SB_LUT4 i15683_3_lut (.I0(\data_out_frame[19] [2]), .I1(displacement[10]), 
            .I2(n24278), .I3(GND_net), .O(n29631));   // verilog/coms.v(128[12] 303[6])
    defparam i15683_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF pwm_setpoint_i0 (.Q(pwm_setpoint[0]), .C(CLK_c), .D(pwm_setpoint_23__N_11[0]));   // verilog/TinyFPGA_B.v(104[9] 130[5])
    SB_LUT4 add_157_16_lut (.I0(GND_net), .I1(delay_counter[14]), .I2(GND_net), 
            .I3(n38459), .O(n1314)) /* synthesis syn_instantiated=1 */ ;
    defparam add_157_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_157_16 (.CI(n38459), .I0(delay_counter[14]), .I1(GND_net), 
            .CO(n38460));
    SB_LUT4 add_1006_5_lut (.I0(GND_net), .I1(n4720), .I2(n22), .I3(n38655), 
            .O(n4505)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1006_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1006_5 (.CI(n38655), .I0(n4720), .I1(n22), .CO(n38656));
    SB_CARRY add_236_9 (.CI(n38483), .I0(encoder1_position[10]), .I1(GND_net), 
            .CO(n38484));
    SB_LUT4 add_1006_4_lut (.I0(GND_net), .I1(n4721), .I2(n23_adj_5254), 
            .I3(n38654), .O(n4506)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1006_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1006_4 (.CI(n38654), .I0(n4721), .I1(n23_adj_5254), .CO(n38655));
    SB_LUT4 add_1006_3_lut (.I0(GND_net), .I1(n4722), .I2(n24), .I3(n38653), 
            .O(n4507)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1006_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_157_15_lut (.I0(GND_net), .I1(delay_counter[13]), .I2(GND_net), 
            .I3(n38458), .O(n1315)) /* synthesis syn_instantiated=1 */ ;
    defparam add_157_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_157_6_lut (.I0(GND_net), .I1(delay_counter[4]), .I2(GND_net), 
            .I3(n38449), .O(n1324)) /* synthesis syn_instantiated=1 */ ;
    defparam add_157_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_157_15 (.CI(n38458), .I0(delay_counter[13]), .I1(GND_net), 
            .CO(n38459));
    SB_DFF read_201 (.Q(read), .C(CLK_c), .D(n46412));   // verilog/TinyFPGA_B.v(375[10] 403[6])
    SB_LUT4 mux_248_i8_3_lut_4_lut (.I0(n27015), .I1(control_mode[1]), .I2(motor_state_23__N_123[7]), 
            .I3(encoder0_position_scaled[7]), .O(motor_state[7]));   // verilog/TinyFPGA_B.v(284[5:22])
    defparam mux_248_i8_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_CARRY add_157_2 (.CI(VCC_net), .I0(delay_counter[0]), .I1(GND_net), 
            .CO(n38446));
    motorControl control (.\Kp[13] (Kp[13]), .GND_net(GND_net), .\Kp[14] (Kp[14]), 
            .\Kp[1] (Kp[1]), .\Kp[0] (Kp[0]), .\Kp[15] (Kp[15]), .\Ki[6] (Ki[6]), 
            .\Ki[3] (Ki[3]), .\Ki[4] (Ki[4]), .\Kp[2] (Kp[2]), .\Kp[3] (Kp[3]), 
            .\Ki[5] (Ki[5]), .\Kp[4] (Kp[4]), .PWMLimit({PWMLimit}), .\Kp[5] (Kp[5]), 
            .\Ki[7] (Ki[7]), .\Kp[9] (Kp[9]), .\Ki[8] (Ki[8]), .\Kp[6] (Kp[6]), 
            .\Ki[2] (Ki[2]), .\Ki[9] (Ki[9]), .\Ki[10] (Ki[10]), .\Ki[1] (Ki[1]), 
            .\Ki[0] (Ki[0]), .\Ki[11] (Ki[11]), .\Kp[10] (Kp[10]), .\Kp[7] (Kp[7]), 
            .\Kp[8] (Kp[8]), .\Kp[11] (Kp[11]), .\Kp[12] (Kp[12]), .\Ki[12] (Ki[12]), 
            .\Ki[13] (Ki[13]), .\Ki[14] (Ki[14]), .\Ki[15] (Ki[15]), .IntegralLimit({IntegralLimit}), 
            .duty({duty}), .clk32MHz(clk32MHz), .VCC_net(VCC_net), .setpoint({setpoint}), 
            .motor_state({motor_state})) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(289[16] 301[4])
    SB_CARRY add_157_6 (.CI(n38449), .I0(delay_counter[4]), .I1(GND_net), 
            .CO(n38450));
    SB_CARRY add_1006_3 (.CI(n38653), .I0(n4722), .I1(n24), .CO(n38654));
    SB_LUT4 add_1006_2_lut (.I0(GND_net), .I1(n4723), .I2(n4698), .I3(VCC_net), 
            .O(n4508)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1006_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_157_14_lut (.I0(GND_net), .I1(delay_counter[12]), .I2(GND_net), 
            .I3(n38457), .O(n1316)) /* synthesis syn_instantiated=1 */ ;
    defparam add_157_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1006_2 (.CI(VCC_net), .I0(n4723), .I1(n4698), .CO(n38653));
    SB_CARRY add_157_14 (.CI(n38457), .I0(delay_counter[12]), .I1(GND_net), 
            .CO(n38458));
    SB_LUT4 mux_248_i9_3_lut_4_lut (.I0(n27015), .I1(control_mode[1]), .I2(motor_state_23__N_123[8]), 
            .I3(encoder0_position_scaled[8]), .O(motor_state[8]));   // verilog/TinyFPGA_B.v(284[5:22])
    defparam mux_248_i9_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 i15684_3_lut (.I0(\data_out_frame[19] [1]), .I1(displacement[9]), 
            .I2(n24278), .I3(GND_net), .O(n29632));   // verilog/coms.v(128[12] 303[6])
    defparam i15684_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15685_3_lut (.I0(\data_out_frame[19] [0]), .I1(displacement[8]), 
            .I2(n24278), .I3(GND_net), .O(n29633));   // verilog/coms.v(128[12] 303[6])
    defparam i15685_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15203_3_lut (.I0(IntegralLimit[6]), .I1(\data_in_frame[13] [6]), 
            .I2(n28521), .I3(GND_net), .O(n29151));   // verilog/coms.v(128[12] 303[6])
    defparam i15203_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15686_3_lut (.I0(\data_out_frame[18] [7]), .I1(displacement[23]), 
            .I2(n24278), .I3(GND_net), .O(n29634));   // verilog/coms.v(128[12] 303[6])
    defparam i15686_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i1574_3_lut (.I0(n2315), .I1(n2382), 
            .I2(n2346), .I3(GND_net), .O(n2414));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1574_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_248_i10_3_lut_4_lut (.I0(n27015), .I1(control_mode[1]), 
            .I2(motor_state_23__N_123[9]), .I3(encoder0_position_scaled[9]), 
            .O(motor_state[9]));   // verilog/TinyFPGA_B.v(284[5:22])
    defparam mux_248_i10_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 encoder0_position_31__I_0_i1573_3_lut (.I0(n2314), .I1(n2381), 
            .I2(n2346), .I3(GND_net), .O(n2413));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1573_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1577_3_lut (.I0(n2318), .I1(n2385), 
            .I2(n2346), .I3(GND_net), .O(n2417));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1577_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15687_3_lut (.I0(\data_out_frame[18] [6]), .I1(displacement[22]), 
            .I2(n24278), .I3(GND_net), .O(n29635));   // verilog/coms.v(128[12] 303[6])
    defparam i15687_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_17_inv_0_i5_1_lut (.I0(current[4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n21));   // verilog/TinyFPGA_B.v(122[16:24])
    defparam unary_minus_17_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i15688_3_lut (.I0(\data_out_frame[18] [5]), .I1(displacement[21]), 
            .I2(n24278), .I3(GND_net), .O(n29636));   // verilog/coms.v(128[12] 303[6])
    defparam i15688_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i1576_3_lut (.I0(n2317), .I1(n2384), 
            .I2(n2346), .I3(GND_net), .O(n2416));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1576_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_248_i11_3_lut_4_lut (.I0(n27015), .I1(control_mode[1]), 
            .I2(motor_state_23__N_123[10]), .I3(encoder0_position_scaled[10]), 
            .O(motor_state[10]));   // verilog/TinyFPGA_B.v(284[5:22])
    defparam mux_248_i11_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 encoder0_position_31__I_0_i1575_3_lut (.I0(n2316), .I1(n2383), 
            .I2(n2346), .I3(GND_net), .O(n2415));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1575_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1578_3_lut (.I0(n2319), .I1(n2386), 
            .I2(n2346), .I3(GND_net), .O(n2418));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1578_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1590_3_lut (.I0(n2331), .I1(n2398), 
            .I2(n2346), .I3(GND_net), .O(n2430));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1590_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_248_i12_3_lut_4_lut (.I0(n27015), .I1(control_mode[1]), 
            .I2(motor_state_23__N_123[11]), .I3(encoder0_position_scaled[11]), 
            .O(motor_state[11]));   // verilog/TinyFPGA_B.v(284[5:22])
    defparam mux_248_i12_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 encoder0_position_31__I_0_i1589_3_lut (.I0(n2330), .I1(n2397), 
            .I2(n2346), .I3(GND_net), .O(n2429));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1589_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15689_3_lut (.I0(\data_out_frame[18] [4]), .I1(displacement[20]), 
            .I2(n24278), .I3(GND_net), .O(n29637));   // verilog/coms.v(128[12] 303[6])
    defparam i15689_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15690_3_lut (.I0(\data_out_frame[18] [3]), .I1(displacement[19]), 
            .I2(n24278), .I3(GND_net), .O(n29638));   // verilog/coms.v(128[12] 303[6])
    defparam i15690_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_248_i13_3_lut_4_lut (.I0(n27015), .I1(control_mode[1]), 
            .I2(motor_state_23__N_123[12]), .I3(encoder0_position_scaled[12]), 
            .O(motor_state[12]));   // verilog/TinyFPGA_B.v(284[5:22])
    defparam mux_248_i13_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 encoder0_position_31__I_0_i1585_3_lut (.I0(n2326), .I1(n2393), 
            .I2(n2346), .I3(GND_net), .O(n2425));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1585_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 unary_minus_17_inv_0_i6_1_lut (.I0(current[5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n20));   // verilog/TinyFPGA_B.v(122[16:24])
    defparam unary_minus_17_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i15691_3_lut (.I0(\data_out_frame[18] [2]), .I1(displacement[18]), 
            .I2(n24278), .I3(GND_net), .O(n29639));   // verilog/coms.v(128[12] 303[6])
    defparam i15691_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_248_i14_3_lut_4_lut (.I0(n27015), .I1(control_mode[1]), 
            .I2(motor_state_23__N_123[13]), .I3(encoder0_position_scaled[13]), 
            .O(motor_state[13]));   // verilog/TinyFPGA_B.v(284[5:22])
    defparam mux_248_i14_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 i15692_3_lut (.I0(\data_out_frame[18] [1]), .I1(displacement[17]), 
            .I2(n24278), .I3(GND_net), .O(n29640));   // verilog/coms.v(128[12] 303[6])
    defparam i15692_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15693_3_lut (.I0(\data_out_frame[18] [0]), .I1(displacement[16]), 
            .I2(n24278), .I3(GND_net), .O(n29641));   // verilog/coms.v(128[12] 303[6])
    defparam i15693_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15694_3_lut (.I0(\data_out_frame[17] [7]), .I1(pwm_setpoint[7]), 
            .I2(n24278), .I3(GND_net), .O(n29642));   // verilog/coms.v(128[12] 303[6])
    defparam i15694_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_17_inv_0_i7_1_lut (.I0(current[6]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n19));   // verilog/TinyFPGA_B.v(122[16:24])
    defparam unary_minus_17_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_248_i15_3_lut_4_lut (.I0(n27015), .I1(control_mode[1]), 
            .I2(motor_state_23__N_123[14]), .I3(encoder0_position_scaled[14]), 
            .O(motor_state[14]));   // verilog/TinyFPGA_B.v(284[5:22])
    defparam mux_248_i15_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 i15695_3_lut (.I0(\data_out_frame[17] [6]), .I1(pwm_setpoint[6]), 
            .I2(n24278), .I3(GND_net), .O(n29643));   // verilog/coms.v(128[12] 303[6])
    defparam i15695_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_248_i16_3_lut_4_lut (.I0(n27015), .I1(control_mode[1]), 
            .I2(motor_state_23__N_123[15]), .I3(encoder0_position_scaled[15]), 
            .O(motor_state[15]));   // verilog/TinyFPGA_B.v(284[5:22])
    defparam mux_248_i16_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 i15696_3_lut (.I0(\data_out_frame[17] [5]), .I1(pwm_setpoint[5]), 
            .I2(n24278), .I3(GND_net), .O(n29644));   // verilog/coms.v(128[12] 303[6])
    defparam i15696_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15697_3_lut (.I0(\data_out_frame[17] [4]), .I1(pwm_setpoint[4]), 
            .I2(n24278), .I3(GND_net), .O(n29645));   // verilog/coms.v(128[12] 303[6])
    defparam i15697_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15698_3_lut (.I0(\data_out_frame[17] [3]), .I1(pwm_setpoint[3]), 
            .I2(n24278), .I3(GND_net), .O(n29646));   // verilog/coms.v(128[12] 303[6])
    defparam i15698_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i1583_3_lut (.I0(n2324), .I1(n2391), 
            .I2(n2346), .I3(GND_net), .O(n2423));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1583_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1581_3_lut (.I0(n2322), .I1(n2389), 
            .I2(n2346), .I3(GND_net), .O(n2421));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1581_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_248_i17_3_lut_4_lut (.I0(n27015), .I1(control_mode[1]), 
            .I2(motor_state_23__N_123[16]), .I3(encoder0_position_scaled[16]), 
            .O(motor_state[16]));   // verilog/TinyFPGA_B.v(284[5:22])
    defparam mux_248_i17_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 encoder0_position_31__I_0_i1580_3_lut (.I0(n2321), .I1(n2388), 
            .I2(n2346), .I3(GND_net), .O(n2420));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1580_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1579_3_lut (.I0(n2320), .I1(n2387), 
            .I2(n2346), .I3(GND_net), .O(n2419));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1579_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1593_3_lut (.I0(n534), .I1(n2401), 
            .I2(n2346), .I3(GND_net), .O(n2433));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1593_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1592_3_lut (.I0(n2333), .I1(n2400), 
            .I2(n2346), .I3(GND_net), .O(n2432));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1592_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_248_i18_3_lut_4_lut (.I0(n27015), .I1(control_mode[1]), 
            .I2(motor_state_23__N_123[17]), .I3(encoder0_position_scaled[17]), 
            .O(motor_state[17]));   // verilog/TinyFPGA_B.v(284[5:22])
    defparam mux_248_i18_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 i15699_3_lut (.I0(\data_out_frame[17] [2]), .I1(pwm_setpoint[2]), 
            .I2(n24278), .I3(GND_net), .O(n29647));   // verilog/coms.v(128[12] 303[6])
    defparam i15699_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i1591_3_lut (.I0(n2332), .I1(n2399), 
            .I2(n2346), .I3(GND_net), .O(n2431));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1591_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i10_3_lut (.I0(encoder0_position[9]), 
            .I1(n24_adj_5291), .I2(encoder0_position[31]), .I3(GND_net), 
            .O(n535));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_mux_3_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i1588_rep_21_3_lut (.I0(n2329), .I1(n2396), 
            .I2(n2346), .I3(GND_net), .O(n2428));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1588_rep_21_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1582_3_lut (.I0(n2323), .I1(n2390), 
            .I2(n2346), .I3(GND_net), .O(n2422));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1582_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15700_3_lut (.I0(\data_out_frame[17] [1]), .I1(pwm_setpoint[1]), 
            .I2(n24278), .I3(GND_net), .O(n29648));   // verilog/coms.v(128[12] 303[6])
    defparam i15700_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_248_i19_3_lut_4_lut (.I0(n27015), .I1(control_mode[1]), 
            .I2(motor_state_23__N_123[18]), .I3(encoder0_position_scaled[18]), 
            .O(motor_state[18]));   // verilog/TinyFPGA_B.v(284[5:22])
    defparam mux_248_i19_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 mux_248_i20_3_lut_4_lut (.I0(n27015), .I1(control_mode[1]), 
            .I2(motor_state_23__N_123[19]), .I3(encoder0_position_scaled[19]), 
            .O(motor_state[19]));   // verilog/TinyFPGA_B.v(284[5:22])
    defparam mux_248_i20_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 i15701_3_lut (.I0(\data_out_frame[17] [0]), .I1(pwm_setpoint[0]), 
            .I2(n24278), .I3(GND_net), .O(n29649));   // verilog/coms.v(128[12] 303[6])
    defparam i15701_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i35196_1_lut (.I0(n2445), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n50784));
    defparam i35196_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_4_lut_adj_1856 (.I0(n2423), .I1(n2427), .I2(n2425), .I3(n2426), 
            .O(n46993));
    defparam i1_4_lut_adj_1856.LUT_INIT = 16'hfffe;
    SB_LUT4 mux_248_i21_3_lut_4_lut (.I0(n27015), .I1(control_mode[1]), 
            .I2(motor_state_23__N_123[20]), .I3(encoder0_position_scaled[20]), 
            .O(motor_state[20]));   // verilog/TinyFPGA_B.v(284[5:22])
    defparam mux_248_i21_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 mux_248_i22_3_lut_4_lut (.I0(n27015), .I1(control_mode[1]), 
            .I2(motor_state_23__N_123[21]), .I3(encoder0_position_scaled[21]), 
            .O(motor_state[21]));   // verilog/TinyFPGA_B.v(284[5:22])
    defparam mux_248_i22_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 i15702_3_lut (.I0(\data_out_frame[16] [7]), .I1(pwm_setpoint[15]), 
            .I2(n24278), .I3(GND_net), .O(n29650));   // verilog/coms.v(128[12] 303[6])
    defparam i15702_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15703_3_lut (.I0(\data_out_frame[16] [6]), .I1(pwm_setpoint[14]), 
            .I2(n24278), .I3(GND_net), .O(n29651));   // verilog/coms.v(128[12] 303[6])
    defparam i15703_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15580_3_lut (.I0(\data_out_frame[23] [6]), .I1(neopxl_color[22]), 
            .I2(n24278), .I3(GND_net), .O(n29528));   // verilog/coms.v(128[12] 303[6])
    defparam i15580_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15704_3_lut (.I0(\data_out_frame[16] [5]), .I1(pwm_setpoint[13]), 
            .I2(n24278), .I3(GND_net), .O(n29652));   // verilog/coms.v(128[12] 303[6])
    defparam i15704_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_248_i23_3_lut_4_lut (.I0(n27015), .I1(control_mode[1]), 
            .I2(motor_state_23__N_123[22]), .I3(encoder0_position_scaled[22]), 
            .O(motor_state[22]));   // verilog/TinyFPGA_B.v(284[5:22])
    defparam mux_248_i23_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 i15705_3_lut (.I0(\data_out_frame[16] [4]), .I1(pwm_setpoint[12]), 
            .I2(n24278), .I3(GND_net), .O(n29653));   // verilog/coms.v(128[12] 303[6])
    defparam i15705_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1857 (.I0(n2424), .I1(n46993), .I2(n2422), .I3(n2428), 
            .O(n46995));
    defparam i1_4_lut_adj_1857.LUT_INIT = 16'hfffe;
    SB_LUT4 i21517_4_lut (.I0(n535), .I1(n2431), .I2(n2432), .I3(n2433), 
            .O(n35466));
    defparam i21517_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 i1_4_lut_adj_1858 (.I0(n2419), .I1(n2420), .I2(n46995), .I3(n2421), 
            .O(n47001));
    defparam i1_4_lut_adj_1858.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_adj_1859 (.I0(n2429), .I1(n2430), .I2(GND_net), .I3(GND_net), 
            .O(n47195));
    defparam i1_2_lut_adj_1859.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut_adj_1860 (.I0(n2418), .I1(n47195), .I2(n47001), .I3(n35466), 
            .O(n47005));
    defparam i1_4_lut_adj_1860.LUT_INIT = 16'hfefa;
    SB_LUT4 i1_4_lut_adj_1861 (.I0(n2415), .I1(n2416), .I2(n2417), .I3(n47005), 
            .O(n47011));
    defparam i1_4_lut_adj_1861.LUT_INIT = 16'hfffe;
    SB_LUT4 i35199_4_lut (.I0(n2413), .I1(n2412), .I2(n2414), .I3(n47011), 
            .O(n2445));
    defparam i35199_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i15204_4_lut (.I0(CS_MISO_c), .I1(data_adj_5514[5]), .I2(n6_adj_5340), 
            .I3(n27167), .O(n29152));   // verilog/tli4970.v(35[10] 68[6])
    defparam i15204_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 encoder0_position_31__I_0_i1510_3_lut (.I0(n2219), .I1(n2286), 
            .I2(n2247), .I3(GND_net), .O(n2318));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1510_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1509_3_lut (.I0(n2218), .I1(n2285), 
            .I2(n2247), .I3(GND_net), .O(n2317));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1509_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1508_3_lut (.I0(n2217), .I1(n2284), 
            .I2(n2247), .I3(GND_net), .O(n2316));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1508_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_248_i24_3_lut_4_lut (.I0(n27015), .I1(control_mode[1]), 
            .I2(motor_state_23__N_123[23]), .I3(encoder0_position_scaled[23]), 
            .O(motor_state[23]));   // verilog/TinyFPGA_B.v(284[5:22])
    defparam mux_248_i24_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 i12_3_lut_4_lut (.I0(r_SM_Main[1]), .I1(r_SM_Main[2]), .I2(n28562), 
            .I3(rx_data_ready), .O(n43326));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i12_3_lut_4_lut.LUT_INIT = 16'h2f20;
    SB_LUT4 i1_3_lut_3_lut (.I0(\ID_READOUT_FSM.state [0]), .I1(\ID_READOUT_FSM.state [1]), 
            .I2(n27013), .I3(GND_net), .O(n7417));
    defparam i1_3_lut_3_lut.LUT_INIT = 16'h1515;
    SB_LUT4 encoder0_position_31__I_0_i1511_3_lut (.I0(n2220), .I1(n2287), 
            .I2(n2247), .I3(GND_net), .O(n2319));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1511_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i33969_2_lut_3_lut (.I0(n62), .I1(delay_counter[31]), .I2(\ID_READOUT_FSM.state [0]), 
            .I3(GND_net), .O(n49335));
    defparam i33969_2_lut_3_lut.LUT_INIT = 16'hf2f2;
    SB_LUT4 encoder0_position_31__I_0_i1507_3_lut (.I0(n2216), .I1(n2283), 
            .I2(n2247), .I3(GND_net), .O(n2315));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1507_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15581_3_lut (.I0(\data_out_frame[23] [5]), .I1(neopxl_color[21]), 
            .I2(n24278), .I3(GND_net), .O(n29529));   // verilog/coms.v(128[12] 303[6])
    defparam i15581_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29180_4_lut_4_lut_4_lut (.I0(h1), .I1(h3), .I2(h2), .I3(commutation_state[2]), 
            .O(n44694));   // verilog/TinyFPGA_B.v(167[7:23])
    defparam i29180_4_lut_4_lut_4_lut.LUT_INIT = 16'hc544;
    SB_LUT4 i1_2_lut_3_lut (.I0(\ID_READOUT_FSM.state [0]), .I1(\ID_READOUT_FSM.state [1]), 
            .I2(n27013), .I3(GND_net), .O(n27014));   // verilog/TinyFPGA_B.v(393[7:11])
    defparam i1_2_lut_3_lut.LUT_INIT = 16'hfbfb;
    SB_LUT4 encoder0_position_31__I_0_i1505_3_lut (.I0(n2214), .I1(n2281), 
            .I2(n2247), .I3(GND_net), .O(n2313));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1505_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1506_3_lut (.I0(n2215), .I1(n2282), 
            .I2(n2247), .I3(GND_net), .O(n2314));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1506_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1525_3_lut (.I0(n533), .I1(n2301), 
            .I2(n2247), .I3(GND_net), .O(n2333));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1525_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1524_3_lut (.I0(n2233), .I1(n2300), 
            .I2(n2247), .I3(GND_net), .O(n2332));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1524_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1523_3_lut (.I0(n2232), .I1(n2299), 
            .I2(n2247), .I3(GND_net), .O(n2331));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1523_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i11_3_lut (.I0(encoder0_position[10]), 
            .I1(n23_adj_5292), .I2(encoder0_position[31]), .I3(GND_net), 
            .O(n534));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_mux_3_i11_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i1522_3_lut (.I0(n2231), .I1(n2298), 
            .I2(n2247), .I3(GND_net), .O(n2330));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1522_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1521_3_lut (.I0(n2230), .I1(n2297), 
            .I2(n2247), .I3(GND_net), .O(n2329));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1521_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1520_3_lut (.I0(n2229), .I1(n2296), 
            .I2(n2247), .I3(GND_net), .O(n2328));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1520_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1515_rep_39_3_lut (.I0(n2224), .I1(n2291), 
            .I2(n2247), .I3(GND_net), .O(n2323));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1515_rep_39_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1517_3_lut (.I0(n2226), .I1(n2293), 
            .I2(n2247), .I3(GND_net), .O(n2325));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1517_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15582_3_lut (.I0(ID[7]), .I1(data[7]), .I2(n46410), .I3(GND_net), 
            .O(n29530));   // verilog/TinyFPGA_B.v(375[10] 403[6])
    defparam i15582_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1518_3_lut (.I0(n2227), .I1(n2294), 
            .I2(n2247), .I3(GND_net), .O(n2326));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1518_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1513_3_lut (.I0(n2222), .I1(n2289), 
            .I2(n2247), .I3(GND_net), .O(n2321));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1513_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1512_3_lut (.I0(n2221), .I1(n2288), 
            .I2(n2247), .I3(GND_net), .O(n2320));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1512_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1516_3_lut (.I0(n2225), .I1(n2292), 
            .I2(n2247), .I3(GND_net), .O(n2324));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1516_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15212_4_lut (.I0(CS_MISO_c), .I1(data_adj_5514[7]), .I2(n6_adj_5340), 
            .I3(n27180), .O(n29160));   // verilog/tli4970.v(35[10] 68[6])
    defparam i15212_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 encoder0_position_31__I_0_i1519_3_lut (.I0(n2228), .I1(n2295), 
            .I2(n2247), .I3(GND_net), .O(n2327));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1519_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1514_3_lut (.I0(n2223), .I1(n2290), 
            .I2(n2247), .I3(GND_net), .O(n2322));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1514_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i35277_1_lut (.I0(n2346), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n50865));
    defparam i35277_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_4_lut_adj_1862 (.I0(n2326), .I1(n2325), .I2(n2323), .I3(n2328), 
            .O(n46765));
    defparam i1_4_lut_adj_1862.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_3_lut_adj_1863 (.I0(n2322), .I1(n2327), .I2(n2324), .I3(GND_net), 
            .O(n46767));
    defparam i1_3_lut_adj_1863.LUT_INIT = 16'hfefe;
    SB_LUT4 i21519_4_lut (.I0(n534), .I1(n2331), .I2(n2332), .I3(n2333), 
            .O(n35468));
    defparam i21519_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 i1_4_lut_adj_1864 (.I0(n2320), .I1(n2321), .I2(n46767), .I3(n46765), 
            .O(n46773));
    defparam i1_4_lut_adj_1864.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_adj_1865 (.I0(n2329), .I1(n2330), .I2(GND_net), .I3(GND_net), 
            .O(n46969));
    defparam i1_2_lut_adj_1865.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_17_inv_0_i8_1_lut (.I0(current[7]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n18));   // verilog/TinyFPGA_B.v(122[16:24])
    defparam unary_minus_17_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_4_lut_adj_1866 (.I0(n46969), .I1(n2319), .I2(n46773), .I3(n35468), 
            .O(n46777));
    defparam i1_4_lut_adj_1866.LUT_INIT = 16'hfefc;
    SB_LUT4 i1_4_lut_adj_1867 (.I0(n2316), .I1(n2317), .I2(n2318), .I3(n46777), 
            .O(n46783));
    defparam i1_4_lut_adj_1867.LUT_INIT = 16'hfffe;
    SB_LUT4 i35280_4_lut (.I0(n2314), .I1(n2313), .I2(n2315), .I3(n46783), 
            .O(n2346));
    defparam i35280_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i15706_3_lut (.I0(\data_out_frame[16] [3]), .I1(pwm_setpoint[11]), 
            .I2(n24278), .I3(GND_net), .O(n29654));   // verilog/coms.v(128[12] 303[6])
    defparam i15706_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_250_i21_4_lut (.I0(encoder1_position_scaled[20]), .I1(displacement[20]), 
            .I2(n15_adj_5249), .I3(n15_adj_5321), .O(motor_state_23__N_123[20]));   // verilog/TinyFPGA_B.v(285[5] 287[10])
    defparam mux_250_i21_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i15707_3_lut (.I0(\data_out_frame[16] [2]), .I1(pwm_setpoint[10]), 
            .I2(n24278), .I3(GND_net), .O(n29655));   // verilog/coms.v(128[12] 303[6])
    defparam i15707_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15708_3_lut (.I0(\data_out_frame[16] [1]), .I1(pwm_setpoint[9]), 
            .I2(n24278), .I3(GND_net), .O(n29656));   // verilog/coms.v(128[12] 303[6])
    defparam i15708_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15709_3_lut (.I0(\data_out_frame[16] [0]), .I1(pwm_setpoint[8]), 
            .I2(n24278), .I3(GND_net), .O(n29657));   // verilog/coms.v(128[12] 303[6])
    defparam i15709_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15710_3_lut (.I0(\data_out_frame[15] [7]), .I1(pwm_setpoint[23]), 
            .I2(n24278), .I3(GND_net), .O(n29658));   // verilog/coms.v(128[12] 303[6])
    defparam i15710_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i1439_3_lut (.I0(n2116), .I1(n2183), 
            .I2(n2148), .I3(GND_net), .O(n2215));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1439_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1444_3_lut (.I0(n2121), .I1(n2188), 
            .I2(n2148), .I3(GND_net), .O(n2220));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1444_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1443_3_lut (.I0(n2120), .I1(n2187), 
            .I2(n2148), .I3(GND_net), .O(n2219));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1443_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15711_3_lut (.I0(\data_out_frame[15] [6]), .I1(pwm_setpoint[22]), 
            .I2(n24278), .I3(GND_net), .O(n29659));   // verilog/coms.v(128[12] 303[6])
    defparam i15711_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i1457_3_lut (.I0(n532), .I1(n2201), 
            .I2(n2148), .I3(GND_net), .O(n2233));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1457_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1456_3_lut (.I0(n2133), .I1(n2200), 
            .I2(n2148), .I3(GND_net), .O(n2232));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1456_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i12_3_lut (.I0(encoder0_position[11]), 
            .I1(n22_adj_5293), .I2(encoder0_position[31]), .I3(GND_net), 
            .O(n533));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_mux_3_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15712_3_lut (.I0(\data_out_frame[15] [5]), .I1(pwm_setpoint[21]), 
            .I2(n24278), .I3(GND_net), .O(n29660));   // verilog/coms.v(128[12] 303[6])
    defparam i15712_3_lut.LUT_INIT = 16'hcaca;
    pll32MHz pll32MHz_inst (.GND_net(GND_net), .CLK_c(CLK_c), .VCC_net(VCC_net), 
            .clk32MHz(clk32MHz)) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(34[10] 37[2])
    SB_LUT4 i15713_3_lut (.I0(\data_out_frame[15] [4]), .I1(pwm_setpoint[20]), 
            .I2(n24278), .I3(GND_net), .O(n29661));   // verilog/coms.v(128[12] 303[6])
    defparam i15713_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15714_3_lut (.I0(\data_out_frame[15] [3]), .I1(pwm_setpoint[19]), 
            .I2(n24278), .I3(GND_net), .O(n29662));   // verilog/coms.v(128[12] 303[6])
    defparam i15714_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15715_3_lut (.I0(\data_out_frame[15] [2]), .I1(pwm_setpoint[18]), 
            .I2(n24278), .I3(GND_net), .O(n29663));   // verilog/coms.v(128[12] 303[6])
    defparam i15715_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i1449_3_lut (.I0(n2126), .I1(n2193), 
            .I2(n2148), .I3(GND_net), .O(n2225));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1449_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1441_3_lut (.I0(n2118), .I1(n2185), 
            .I2(n2148), .I3(GND_net), .O(n2217));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1441_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1440_3_lut (.I0(n2117), .I1(n2184), 
            .I2(n2148), .I3(GND_net), .O(n2216));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1440_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1451_3_lut (.I0(n2128), .I1(n2195_adj_5401), 
            .I2(n2148), .I3(GND_net), .O(n2227));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1451_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15716_3_lut (.I0(\data_out_frame[15] [1]), .I1(pwm_setpoint[17]), 
            .I2(n24278), .I3(GND_net), .O(n29664));   // verilog/coms.v(128[12] 303[6])
    defparam i15716_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15717_3_lut (.I0(\data_out_frame[15] [0]), .I1(pwm_setpoint[16]), 
            .I2(n24278), .I3(GND_net), .O(n29665));   // verilog/coms.v(128[12] 303[6])
    defparam i15717_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15718_3_lut (.I0(\data_out_frame[14] [7]), .I1(setpoint[7]), 
            .I2(n24278), .I3(GND_net), .O(n29666));   // verilog/coms.v(128[12] 303[6])
    defparam i15718_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i1447_3_lut (.I0(n2124), .I1(n2191), 
            .I2(n2148), .I3(GND_net), .O(n2223));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1447_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1452_3_lut (.I0(n2129), .I1(n2196), 
            .I2(n2148), .I3(GND_net), .O(n2228));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1452_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15719_3_lut (.I0(\data_out_frame[14] [6]), .I1(setpoint[6]), 
            .I2(n24278), .I3(GND_net), .O(n29667));   // verilog/coms.v(128[12] 303[6])
    defparam i15719_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i33862_2_lut_4_lut (.I0(commutation_state[0]), .I1(n4), .I2(commutation_state_prev[0]), 
            .I3(dti_counter[0]), .O(n49334));   // verilog/TinyFPGA_B.v(147[7:48])
    defparam i33862_2_lut_4_lut.LUT_INIT = 16'h2100;
    SB_LUT4 i15720_3_lut (.I0(\data_out_frame[14] [5]), .I1(setpoint[5]), 
            .I2(n24278), .I3(GND_net), .O(n29668));   // verilog/coms.v(128[12] 303[6])
    defparam i15720_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15721_3_lut (.I0(\data_out_frame[14] [4]), .I1(setpoint[4]), 
            .I2(n24278), .I3(GND_net), .O(n29669));   // verilog/coms.v(128[12] 303[6])
    defparam i15721_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i1445_3_lut (.I0(n2122), .I1(n2189), 
            .I2(n2148), .I3(GND_net), .O(n2221));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1445_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15722_3_lut (.I0(\data_out_frame[14] [3]), .I1(setpoint[3]), 
            .I2(n24278), .I3(GND_net), .O(n29670));   // verilog/coms.v(128[12] 303[6])
    defparam i15722_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i1455_3_lut (.I0(n2132), .I1(n2199), 
            .I2(n2148), .I3(GND_net), .O(n2231));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1455_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i33882_2_lut_4_lut (.I0(commutation_state[0]), .I1(n4), .I2(commutation_state_prev[0]), 
            .I3(dti_counter[1]), .O(n49298));   // verilog/TinyFPGA_B.v(147[7:48])
    defparam i33882_2_lut_4_lut.LUT_INIT = 16'h2100;
    SB_LUT4 encoder0_position_31__I_0_i1454_3_lut (.I0(n2131), .I1(n2198), 
            .I2(n2148), .I3(GND_net), .O(n2230));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1454_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15723_3_lut (.I0(\data_out_frame[14] [2]), .I1(setpoint[2]), 
            .I2(n24278), .I3(GND_net), .O(n29671));   // verilog/coms.v(128[12] 303[6])
    defparam i15723_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i1453_3_lut (.I0(n2130), .I1(n2197), 
            .I2(n2148), .I3(GND_net), .O(n2229));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1453_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1448_3_lut (.I0(n2125), .I1(n2192), 
            .I2(n2148), .I3(GND_net), .O(n2224));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1448_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i33881_2_lut_4_lut (.I0(commutation_state[0]), .I1(n4), .I2(commutation_state_prev[0]), 
            .I3(dti_counter[2]), .O(n49297));   // verilog/TinyFPGA_B.v(147[7:48])
    defparam i33881_2_lut_4_lut.LUT_INIT = 16'h2100;
    SB_LUT4 i33880_2_lut_4_lut (.I0(commutation_state[0]), .I1(n4), .I2(commutation_state_prev[0]), 
            .I3(dti_counter[3]), .O(n49296));   // verilog/TinyFPGA_B.v(147[7:48])
    defparam i33880_2_lut_4_lut.LUT_INIT = 16'h2100;
    SB_LUT4 i15724_3_lut (.I0(\data_out_frame[14] [1]), .I1(setpoint[1]), 
            .I2(n24278), .I3(GND_net), .O(n29672));   // verilog/coms.v(128[12] 303[6])
    defparam i15724_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i33879_2_lut_4_lut (.I0(commutation_state[0]), .I1(n4), .I2(commutation_state_prev[0]), 
            .I3(dti_counter[4]), .O(n49295));   // verilog/TinyFPGA_B.v(147[7:48])
    defparam i33879_2_lut_4_lut.LUT_INIT = 16'h2100;
    SB_LUT4 i15725_3_lut (.I0(\data_out_frame[14] [0]), .I1(setpoint[0]), 
            .I2(n24278), .I3(GND_net), .O(n29673));   // verilog/coms.v(128[12] 303[6])
    defparam i15725_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i1450_3_lut (.I0(n2127), .I1(n2194), 
            .I2(n2148), .I3(GND_net), .O(n2226));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1450_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i33878_2_lut_4_lut (.I0(commutation_state[0]), .I1(n4), .I2(commutation_state_prev[0]), 
            .I3(dti_counter[5]), .O(n49294));   // verilog/TinyFPGA_B.v(147[7:48])
    defparam i33878_2_lut_4_lut.LUT_INIT = 16'h2100;
    SB_LUT4 unary_minus_17_inv_0_i9_1_lut (.I0(current[8]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_5253));   // verilog/TinyFPGA_B.v(122[16:24])
    defparam unary_minus_17_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i15726_3_lut (.I0(\data_out_frame[13] [7]), .I1(setpoint[15]), 
            .I2(n24278), .I3(GND_net), .O(n29674));   // verilog/coms.v(128[12] 303[6])
    defparam i15726_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i1442_3_lut (.I0(n2119), .I1(n2186), 
            .I2(n2148), .I3(GND_net), .O(n2218));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1442_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1446_3_lut (.I0(n2123), .I1(n2190), 
            .I2(n2148), .I3(GND_net), .O(n2222));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1446_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i33834_2_lut_4_lut (.I0(commutation_state[0]), .I1(n4), .I2(commutation_state_prev[0]), 
            .I3(dti_counter[6]), .O(n49293));   // verilog/TinyFPGA_B.v(147[7:48])
    defparam i33834_2_lut_4_lut.LUT_INIT = 16'h2100;
    SB_LUT4 i15727_3_lut (.I0(\data_out_frame[13] [6]), .I1(setpoint[14]), 
            .I2(n24278), .I3(GND_net), .O(n29675));   // verilog/coms.v(128[12] 303[6])
    defparam i15727_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i35302_1_lut (.I0(n2247), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n50890));
    defparam i35302_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_4_lut_adj_1868 (.I0(n2222), .I1(n2218), .I2(n2226), .I3(n2224), 
            .O(n46053));
    defparam i1_4_lut_adj_1868.LUT_INIT = 16'hfffe;
    SB_LUT4 i15728_3_lut (.I0(\data_out_frame[13] [5]), .I1(setpoint[13]), 
            .I2(n24278), .I3(GND_net), .O(n29676));   // verilog/coms.v(128[12] 303[6])
    defparam i15728_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15729_3_lut (.I0(\data_out_frame[13] [4]), .I1(setpoint[12]), 
            .I2(n24278), .I3(GND_net), .O(n29677));   // verilog/coms.v(128[12] 303[6])
    defparam i15729_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i21460_3_lut (.I0(n533), .I1(n2232), .I2(n2233), .I3(GND_net), 
            .O(n35408));
    defparam i21460_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i1_4_lut_adj_1869 (.I0(n2221), .I1(n2228), .I2(n2223), .I3(n2227), 
            .O(n46961));
    defparam i1_4_lut_adj_1869.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1870 (.I0(n2229), .I1(n35408), .I2(n2230), .I3(n2231), 
            .O(n44998));
    defparam i1_4_lut_adj_1870.LUT_INIT = 16'ha080;
    SB_LUT4 i15730_3_lut (.I0(\data_out_frame[13] [3]), .I1(setpoint[11]), 
            .I2(n24278), .I3(GND_net), .O(n29678));   // verilog/coms.v(128[12] 303[6])
    defparam i15730_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i33815_2_lut_4_lut (.I0(commutation_state[0]), .I1(n4), .I2(commutation_state_prev[0]), 
            .I3(dti_counter[7]), .O(n49292));   // verilog/TinyFPGA_B.v(147[7:48])
    defparam i33815_2_lut_4_lut.LUT_INIT = 16'h2100;
    SB_LUT4 i1_2_lut_4_lut_adj_1871 (.I0(commutation_state[0]), .I1(n4), 
            .I2(commutation_state_prev[0]), .I3(dti_N_440), .O(n28458));   // verilog/TinyFPGA_B.v(147[7:48])
    defparam i1_2_lut_4_lut_adj_1871.LUT_INIT = 16'hdeff;
    SB_LUT4 i15731_3_lut (.I0(\data_out_frame[13] [2]), .I1(setpoint[10]), 
            .I2(n24278), .I3(GND_net), .O(n29679));   // verilog/coms.v(128[12] 303[6])
    defparam i15731_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29232_4_lut (.I0(n7_adj_5404), .I1(state_adj_5510[0]), .I2(n6_adj_5274), 
            .I3(state_adj_5537[0]), .O(n44748));
    defparam i29232_4_lut.LUT_INIT = 16'hccc8;
    SB_LUT4 i1_4_lut_adj_1872 (.I0(n2216), .I1(n46053), .I2(n2217), .I3(n2225), 
            .O(n46953));
    defparam i1_4_lut_adj_1872.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1873 (.I0(n2219), .I1(n2220), .I2(n44998), .I3(n46961), 
            .O(n46967));
    defparam i1_4_lut_adj_1873.LUT_INIT = 16'hfffe;
    SB_LUT4 i35305_4_lut (.I0(n2214), .I1(n46967), .I2(n46953), .I3(n2215), 
            .O(n2247));
    defparam i35305_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 unary_minus_19_inv_0_i24_1_lut (.I0(duty[23]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(pwm_setpoint_23__N_239));   // verilog/TinyFPGA_B.v(123[25:30])
    defparam unary_minus_19_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_17_inv_0_i10_1_lut (.I0(current[9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n16_adj_5252));   // verilog/TinyFPGA_B.v(122[16:24])
    defparam unary_minus_17_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_4_lut_adj_1874 (.I0(n34717), .I1(n44835), .I2(state_adj_5510[0]), 
            .I3(read), .O(n43386));   // verilog/eeprom.v(26[8] 58[4])
    defparam i1_4_lut_adj_1874.LUT_INIT = 16'h8280;
    SB_LUT4 i509_2_lut (.I0(n1415), .I1(n27013), .I2(GND_net), .I3(GND_net), 
            .O(n2204));   // verilog/TinyFPGA_B.v(394[9] 400[12])
    defparam i509_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 encoder0_position_31__I_0_i1372_3_lut (.I0(n2017), .I1(n2084), 
            .I2(n2049), .I3(GND_net), .O(n2116));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1372_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1378_3_lut (.I0(n2023), .I1(n2090), 
            .I2(n2049), .I3(GND_net), .O(n2122));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1378_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1374_3_lut (.I0(n2019), .I1(n2086), 
            .I2(n2049), .I3(GND_net), .O(n2118));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1374_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1376_3_lut (.I0(n2021), .I1(n2088), 
            .I2(n2049), .I3(GND_net), .O(n2120));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1376_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1375_3_lut (.I0(n2020), .I1(n2087), 
            .I2(n2049), .I3(GND_net), .O(n2119));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1375_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1373_3_lut (.I0(n2018), .I1(n2085), 
            .I2(n2049), .I3(GND_net), .O(n2117));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1373_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1383_3_lut (.I0(n2028), .I1(n2095), 
            .I2(n2049), .I3(GND_net), .O(n2127));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1383_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1384_3_lut (.I0(n2029), .I1(n2096), 
            .I2(n2049), .I3(GND_net), .O(n2128));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1384_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 unary_minus_17_inv_0_i11_1_lut (.I0(current[10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_5251));   // verilog/TinyFPGA_B.v(122[16:24])
    defparam unary_minus_17_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_i1382_3_lut (.I0(n2027), .I1(n2094), 
            .I2(n2049), .I3(GND_net), .O(n2126));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1382_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1381_3_lut (.I0(n2026), .I1(n2093), 
            .I2(n2049), .I3(GND_net), .O(n2125));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1381_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1380_3_lut (.I0(n2025), .I1(n2092), 
            .I2(n2049), .I3(GND_net), .O(n2124));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1380_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1379_3_lut (.I0(n2024), .I1(n2091), 
            .I2(n2049), .I3(GND_net), .O(n2123));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1379_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i33826_4_lut (.I0(n5_adj_5368), .I1(n6_adj_5445), .I2(n7494), 
            .I3(n2204), .O(n49302));   // verilog/TinyFPGA_B.v(375[10] 403[6])
    defparam i33826_4_lut.LUT_INIT = 16'h080c;
    SB_LUT4 i49_4_lut (.I0(n49302), .I1(data_ready), .I2(\ID_READOUT_FSM.state [0]), 
            .I3(n7494), .O(n42724));   // verilog/TinyFPGA_B.v(375[10] 403[6])
    defparam i49_4_lut.LUT_INIT = 16'hfa3a;
    SB_LUT4 encoder0_position_31__I_0_i1377_3_lut (.I0(n2022), .I1(n2089), 
            .I2(n2049), .I3(GND_net), .O(n2121));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1377_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1387_3_lut (.I0(n2032), .I1(n2099), 
            .I2(n2049), .I3(GND_net), .O(n2131));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1387_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1386_3_lut (.I0(n2031), .I1(n2098), 
            .I2(n2049), .I3(GND_net), .O(n2130));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1386_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1385_3_lut (.I0(n2030), .I1(n2097), 
            .I2(n2049), .I3(GND_net), .O(n2129));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1385_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1389_rep_40_3_lut (.I0(n531), .I1(n2101), 
            .I2(n2049), .I3(GND_net), .O(n2133));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1389_rep_40_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1388_3_lut (.I0(n2033), .I1(n2100), 
            .I2(n2049), .I3(GND_net), .O(n2132));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1388_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i13_3_lut (.I0(encoder0_position[12]), 
            .I1(n21_adj_5294), .I2(encoder0_position[31]), .I3(GND_net), 
            .O(n532));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_mux_3_i13_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i35326_1_lut (.I0(n2148), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n50914));
    defparam i35326_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i21462_3_lut (.I0(n532), .I1(n2132), .I2(n2133), .I3(GND_net), 
            .O(n35410));
    defparam i21462_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i1_4_lut_adj_1875 (.I0(n2125), .I1(n2126), .I2(n2128), .I3(n2127), 
            .O(n46849));
    defparam i1_4_lut_adj_1875.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1876 (.I0(n2129), .I1(n35410), .I2(n2130), .I3(n2131), 
            .O(n44972));
    defparam i1_4_lut_adj_1876.LUT_INIT = 16'ha080;
    SB_LUT4 i1_3_lut_adj_1877 (.I0(n2121), .I1(n2123), .I2(n2124), .I3(GND_net), 
            .O(n46815));
    defparam i1_3_lut_adj_1877.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_4_lut_adj_1878 (.I0(n44972), .I1(n2118), .I2(n2122), .I3(n46849), 
            .O(n45989));
    defparam i1_4_lut_adj_1878.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1879 (.I0(n2117), .I1(n2119), .I2(n2120), .I3(n46815), 
            .O(n46821));
    defparam i1_4_lut_adj_1879.LUT_INIT = 16'hfffe;
    SB_LUT4 i35329_4_lut (.I0(n2116), .I1(n2115), .I2(n46821), .I3(n45989), 
            .O(n2148));
    defparam i35329_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 unary_minus_17_inv_0_i12_1_lut (.I0(current[11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n14_adj_5250));   // verilog/TinyFPGA_B.v(122[16:24])
    defparam unary_minus_17_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_250_i22_4_lut (.I0(encoder1_position_scaled[21]), .I1(displacement[21]), 
            .I2(n15_adj_5249), .I3(n15_adj_5321), .O(motor_state_23__N_123[21]));   // verilog/TinyFPGA_B.v(285[5] 287[10])
    defparam mux_250_i22_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i15205_3_lut (.I0(IntegralLimit[5]), .I1(\data_in_frame[13] [5]), 
            .I2(n28521), .I3(GND_net), .O(n29153));   // verilog/coms.v(128[12] 303[6])
    defparam i15205_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5494_3_lut_4_lut_4_lut (.I0(commutation_state[2]), .I1(commutation_state[1]), 
            .I2(dir), .I3(commutation_state[0]), .O(GHA_N_391));   // verilog/TinyFPGA_B.v(180[7] 199[15])
    defparam i5494_3_lut_4_lut_4_lut.LUT_INIT = 16'h12c2;
    SB_LUT4 i15583_3_lut (.I0(ID[6]), .I1(data[6]), .I2(n46410), .I3(GND_net), 
            .O(n29531));   // verilog/TinyFPGA_B.v(375[10] 403[6])
    defparam i15583_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i5496_3_lut_4_lut_4_lut (.I0(commutation_state[2]), .I1(commutation_state[1]), 
            .I2(dir), .I3(commutation_state[0]), .O(GLA_N_408));   // verilog/TinyFPGA_B.v(180[7] 199[15])
    defparam i5496_3_lut_4_lut_4_lut.LUT_INIT = 16'h212c;
    SB_LUT4 i15285_3_lut (.I0(n28972), .I1(r_Bit_Index[0]), .I2(n28666), 
            .I3(GND_net), .O(n29233));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i15285_3_lut.LUT_INIT = 16'h1414;
    SB_LUT4 mux_250_i23_4_lut (.I0(encoder1_position_scaled[22]), .I1(displacement[22]), 
            .I2(n15_adj_5249), .I3(n15_adj_5321), .O(motor_state_23__N_123[22]));   // verilog/TinyFPGA_B.v(285[5] 287[10])
    defparam mux_250_i23_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i1_2_lut_4_lut_adj_1880 (.I0(r_SM_Main[0]), .I1(r_SM_Main[1]), 
            .I2(r_SM_Main[2]), .I3(r_SM_Main_2__N_3706[2]), .O(n43724));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i1_2_lut_4_lut_adj_1880.LUT_INIT = 16'h0800;
    SB_LUT4 i4_4_lut_adj_1881 (.I0(control_mode[3]), .I1(control_mode[5]), 
            .I2(control_mode[4]), .I3(control_mode[7]), .O(n10_adj_5453));   // verilog/TinyFPGA_B.v(285[5:22])
    defparam i4_4_lut_adj_1881.LUT_INIT = 16'hfffe;
    SB_LUT4 i15282_3_lut (.I0(n28970), .I1(r_Bit_Index_adj_5527[0]), .I2(n28662), 
            .I3(GND_net), .O(n29230));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i15282_3_lut.LUT_INIT = 16'h1414;
    SB_LUT4 i5_3_lut_adj_1882 (.I0(control_mode[6]), .I1(n10_adj_5453), 
            .I2(control_mode[2]), .I3(GND_net), .O(n27171));   // verilog/TinyFPGA_B.v(285[5:22])
    defparam i5_3_lut_adj_1882.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_2_lut_adj_1883 (.I0(n27015), .I1(control_mode[1]), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_5321));   // verilog/TinyFPGA_B.v(286[5:22])
    defparam i1_2_lut_adj_1883.LUT_INIT = 16'hbbbb;
    SB_LUT4 i2_3_lut_adj_1884 (.I0(control_mode[0]), .I1(control_mode[1]), 
            .I2(n27171), .I3(GND_net), .O(n15_adj_5249));   // verilog/TinyFPGA_B.v(285[5:22])
    defparam i2_3_lut_adj_1884.LUT_INIT = 16'hfdfd;
    SB_LUT4 mux_250_i24_4_lut (.I0(encoder1_position_scaled[23]), .I1(displacement[23]), 
            .I2(n15_adj_5249), .I3(n15_adj_5321), .O(motor_state_23__N_123[23]));   // verilog/TinyFPGA_B.v(285[5] 287[10])
    defparam mux_250_i24_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i15584_3_lut (.I0(ID[5]), .I1(data[5]), .I2(n46410), .I3(GND_net), 
            .O(n29532));   // verilog/TinyFPGA_B.v(375[10] 403[6])
    defparam i15584_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i35370_1_lut (.I0(n1950), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n50958));
    defparam i35370_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i15585_3_lut (.I0(ID[4]), .I1(data[4]), .I2(n46410), .I3(GND_net), 
            .O(n29533));   // verilog/TinyFPGA_B.v(375[10] 403[6])
    defparam i15585_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15157_3_lut (.I0(\data_out_frame[7] [2]), .I1(encoder0_position_scaled[10]), 
            .I2(n24278), .I3(GND_net), .O(n29105));   // verilog/coms.v(128[12] 303[6])
    defparam i15157_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15158_3_lut (.I0(\data_out_frame[7] [1]), .I1(encoder0_position_scaled[9]), 
            .I2(n24278), .I3(GND_net), .O(n29106));   // verilog/coms.v(128[12] 303[6])
    defparam i15158_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i1305_rep_41_3_lut (.I0(n1918), .I1(n1985), 
            .I2(n1950), .I3(GND_net), .O(n2017));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1305_rep_41_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1318_3_lut (.I0(n1931), .I1(n1998), 
            .I2(n1950), .I3(GND_net), .O(n2030));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1318_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1317_3_lut (.I0(n1930), .I1(n1997), 
            .I2(n1950), .I3(GND_net), .O(n2029));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1317_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1308_3_lut (.I0(n1921), .I1(n1988), 
            .I2(n1950), .I3(GND_net), .O(n2020));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1308_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1306_3_lut (.I0(n1919), .I1(n1986), 
            .I2(n1950), .I3(GND_net), .O(n2018));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1306_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1307_3_lut (.I0(n1920), .I1(n1987), 
            .I2(n1950), .I3(GND_net), .O(n2019));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1307_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i1_1_lut (.I0(encoder1_position_scaled[0]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n25_adj_5314));   // verilog/TinyFPGA_B.v(340[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_i1311_3_lut (.I0(n1924), .I1(n1991), 
            .I2(n1950), .I3(GND_net), .O(n2023));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1311_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1310_3_lut (.I0(n1923), .I1(n1990), 
            .I2(n1950), .I3(GND_net), .O(n2022));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1310_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1309_3_lut (.I0(n1922), .I1(n1989), 
            .I2(n1950), .I3(GND_net), .O(n2021));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1309_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1314_3_lut (.I0(n1927), .I1(n1994), 
            .I2(n1950), .I3(GND_net), .O(n2026));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1314_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1316_3_lut (.I0(n1929), .I1(n1996), 
            .I2(n1950), .I3(GND_net), .O(n2028));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1316_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1313_3_lut (.I0(n1926), .I1(n1993), 
            .I2(n1950), .I3(GND_net), .O(n2025));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1313_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1312_3_lut (.I0(n1925), .I1(n1992), 
            .I2(n1950), .I3(GND_net), .O(n2024));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1312_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1315_3_lut (.I0(n1928), .I1(n1995), 
            .I2(n1950), .I3(GND_net), .O(n2027));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1315_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1321_3_lut (.I0(n530), .I1(n2001), 
            .I2(n1950), .I3(GND_net), .O(n2033));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1321_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i2_1_lut (.I0(encoder1_position_scaled[1]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n24_adj_5315));   // verilog/TinyFPGA_B.v(340[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_i1320_3_lut (.I0(n1933), .I1(n2000), 
            .I2(n1950), .I3(GND_net), .O(n2032));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1320_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1319_3_lut (.I0(n1932), .I1(n1999), 
            .I2(n1950), .I3(GND_net), .O(n2031));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1319_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i14_3_lut (.I0(encoder0_position[13]), 
            .I1(n20_adj_5295), .I2(encoder0_position[31]), .I3(GND_net), 
            .O(n531));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_mux_3_i14_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i35349_1_lut (.I0(n2049), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n50937));
    defparam i35349_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i21525_4_lut (.I0(n531), .I1(n2031), .I2(n2032), .I3(n2033), 
            .O(n35474));
    defparam i21525_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 i1_3_lut_adj_1885 (.I0(n2027), .I1(n2024), .I2(n2025), .I3(GND_net), 
            .O(n46923));
    defparam i1_3_lut_adj_1885.LUT_INIT = 16'hfefe;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i3_1_lut (.I0(encoder1_position_scaled[2]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n23_adj_5316));   // verilog/TinyFPGA_B.v(340[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_2_lut_adj_1886 (.I0(n2028), .I1(n2026), .I2(GND_net), .I3(GND_net), 
            .O(n46935));
    defparam i1_2_lut_adj_1886.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_1887 (.I0(n2021), .I1(n2022), .I2(n2023), .I3(n46935), 
            .O(n46941));
    defparam i1_4_lut_adj_1887.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1888 (.I0(n2029), .I1(n46923), .I2(n35474), .I3(n2030), 
            .O(n46925));
    defparam i1_4_lut_adj_1888.LUT_INIT = 16'heccc;
    SB_LUT4 i1_4_lut_adj_1889 (.I0(n2019), .I1(n2018), .I2(n2020), .I3(n46941), 
            .O(n46250));
    defparam i1_4_lut_adj_1889.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i4_1_lut (.I0(encoder1_position_scaled[3]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n22_adj_5317));   // verilog/TinyFPGA_B.v(340[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i35352_4_lut (.I0(n2017), .I1(n2016), .I2(n46250), .I3(n46925), 
            .O(n2049));
    defparam i35352_4_lut.LUT_INIT = 16'h0001;
    \quadrature_decoder(1,500000)_U0  quad_counter0 (.b_prev(b_prev), .n1891(CLK_c), 
            .encoder0_position({encoder0_position}), .GND_net(GND_net), 
            .a_new({a_new[1], Open_0}), .direction_N_4071(direction_N_4071), 
            .ENCODER0_B_N_keep(ENCODER0_B_N), .ENCODER0_A_N_keep(ENCODER0_A_N), 
            .VCC_net(VCC_net), .n29249(n29249), .n1855(n1855)) /* synthesis lattice_noprune=1 */ ;   // verilog/TinyFPGA_B.v(303[57] 310[6])
    SB_LUT4 encoder0_position_31__I_0_i1239_3_lut (.I0(n1820), .I1(n1887), 
            .I2(n1851), .I3(GND_net), .O(n1919));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1239_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1238_3_lut (.I0(n1819), .I1(n1886), 
            .I2(n1851), .I3(GND_net), .O(n1918));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1238_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1241_3_lut (.I0(n1822), .I1(n1889), 
            .I2(n1851), .I3(GND_net), .O(n1921));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1241_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15586_3_lut (.I0(ID[3]), .I1(data[3]), .I2(n46410), .I3(GND_net), 
            .O(n29534));   // verilog/TinyFPGA_B.v(375[10] 403[6])
    defparam i15586_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1240_3_lut (.I0(n1821), .I1(n1888), 
            .I2(n1851), .I3(GND_net), .O(n1920));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1240_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1253_rep_42_3_lut (.I0(n529), .I1(n1901), 
            .I2(n1851), .I3(GND_net), .O(n1933));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1253_rep_42_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1252_3_lut (.I0(n1833), .I1(n1900), 
            .I2(n1851), .I3(GND_net), .O(n1932));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1252_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i15_3_lut (.I0(encoder0_position[14]), 
            .I1(n19_adj_5296), .I2(encoder0_position[31]), .I3(GND_net), 
            .O(n530));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_mux_3_i15_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i1247_3_lut (.I0(n1828), .I1(n1895), 
            .I2(n1851), .I3(GND_net), .O(n1927));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1247_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15587_3_lut (.I0(ID[2]), .I1(data[2]), .I2(n46410), .I3(GND_net), 
            .O(n29535));   // verilog/TinyFPGA_B.v(375[10] 403[6])
    defparam i15587_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1244_3_lut (.I0(n1825), .I1(n1892), 
            .I2(n1851), .I3(GND_net), .O(n1924));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1244_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1248_3_lut (.I0(n1829), .I1(n1896_adj_5400), 
            .I2(n1851), .I3(GND_net), .O(n1928));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1248_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15588_3_lut (.I0(ID[1]), .I1(data[1]), .I2(n46410), .I3(GND_net), 
            .O(n29536));   // verilog/TinyFPGA_B.v(375[10] 403[6])
    defparam i15588_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1251_3_lut (.I0(n1832), .I1(n1899), 
            .I2(n1851), .I3(GND_net), .O(n1931));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1251_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1250_3_lut (.I0(n1831), .I1(n1898), 
            .I2(n1851), .I3(GND_net), .O(n1930));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1250_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder1_position_scaled_23__I_4_4_lut (.I0(encoder1_position[0]), 
            .I1(encoder1_position[31]), .I2(encoder1_position[1]), .I3(encoder1_position[2]), 
            .O(encoder1_position_scaled_23__N_303));   // verilog/TinyFPGA_B.v(339[33:52])
    defparam encoder1_position_scaled_23__I_4_4_lut.LUT_INIT = 16'hccc8;
    SB_LUT4 encoder0_position_31__I_0_i1249_3_lut (.I0(n1830), .I1(n1897), 
            .I2(n1851), .I3(GND_net), .O(n1929));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1249_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1243_3_lut (.I0(n1824), .I1(n1891_adj_5399), 
            .I2(n1851), .I3(GND_net), .O(n1923));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1243_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1242_3_lut (.I0(n1823), .I1(n1890), 
            .I2(n1851), .I3(GND_net), .O(n1922));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1242_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1246_3_lut (.I0(n1827), .I1(n1894), 
            .I2(n1851), .I3(GND_net), .O(n1926));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1246_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1245_3_lut (.I0(n1826), .I1(n1893), 
            .I2(n1851), .I3(GND_net), .O(n1925));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1245_3_lut.LUT_INIT = 16'hacac;
    \grp_debouncer(3,1000)  debounce (.n29162(n29162), .data_o({h1, h2, 
            h3}), .CLK_c(CLK_c), .n29161(n29161), .reg_B({reg_B}), .n46440(n46440), 
            .data_i({hall1, hall2, hall3}), .n29025(n29025), .GND_net(GND_net), 
            .VCC_net(VCC_net));   // verilog/TinyFPGA_B.v(98[26] 102[3])
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i5_1_lut (.I0(encoder1_position_scaled[4]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n21_adj_5319));   // verilog/TinyFPGA_B.v(340[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_2_lut_adj_1890 (.I0(n1925), .I1(n1926), .I2(GND_net), .I3(GND_net), 
            .O(n46577));
    defparam i1_2_lut_adj_1890.LUT_INIT = 16'heeee;
    SB_LUT4 i1_3_lut_adj_1891 (.I0(n1928), .I1(n1924), .I2(n1927), .I3(GND_net), 
            .O(n46579));
    defparam i1_3_lut_adj_1891.LUT_INIT = 16'hfefe;
    SB_LUT4 i21466_3_lut (.I0(n530), .I1(n1932), .I2(n1933), .I3(GND_net), 
            .O(n35414));
    defparam i21466_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i6_1_lut (.I0(encoder1_position_scaled[5]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n20_adj_5320));   // verilog/TinyFPGA_B.v(340[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_4_lut_adj_1892 (.I0(n1922), .I1(n1923), .I2(n46579), .I3(n46577), 
            .O(n46585));
    defparam i1_4_lut_adj_1892.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1893 (.I0(n1929), .I1(n35414), .I2(n1930), .I3(n1931), 
            .O(n44955));
    defparam i1_4_lut_adj_1893.LUT_INIT = 16'ha080;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i7_1_lut (.I0(encoder1_position_scaled[6]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n19_adj_5322));   // verilog/TinyFPGA_B.v(340[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i8_1_lut (.I0(encoder1_position_scaled[7]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n18_adj_5323));   // verilog/TinyFPGA_B.v(340[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_4_lut_adj_1894 (.I0(n1920), .I1(n44955), .I2(n1921), .I3(n46585), 
            .O(n46591));
    defparam i1_4_lut_adj_1894.LUT_INIT = 16'hfffe;
    SB_LUT4 i35374_4_lut (.I0(n1918), .I1(n1917), .I2(n1919), .I3(n46591), 
            .O(n1950));
    defparam i35374_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_31__I_0_i1172_3_lut (.I0(n1721), .I1(n1788), 
            .I2(n1752), .I3(GND_net), .O(n1820));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1172_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i9_1_lut (.I0(encoder1_position_scaled[8]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n17_adj_5324));   // verilog/TinyFPGA_B.v(340[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_i1171_3_lut (.I0(n1720), .I1(n1787), 
            .I2(n1752), .I3(GND_net), .O(n1819));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1171_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i10_1_lut (.I0(encoder1_position_scaled[9]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n16_adj_5325));   // verilog/TinyFPGA_B.v(340[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_i1174_3_lut (.I0(n1723), .I1(n1790), 
            .I2(n1752), .I3(GND_net), .O(n1822));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1174_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1173_3_lut (.I0(n1722), .I1(n1789), 
            .I2(n1752), .I3(GND_net), .O(n1821));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1173_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1183_3_lut (.I0(n1732), .I1(n1799), 
            .I2(n1752), .I3(GND_net), .O(n1831));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1183_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1182_3_lut (.I0(n1731), .I1(n1798), 
            .I2(n1752), .I3(GND_net), .O(n1830));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1182_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1181_3_lut (.I0(n1730), .I1(n1797), 
            .I2(n1752), .I3(GND_net), .O(n1829));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1181_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1176_3_lut (.I0(n1725), .I1(n1792), 
            .I2(n1752), .I3(GND_net), .O(n1824));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1176_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1175_3_lut (.I0(n1724), .I1(n1791), 
            .I2(n1752), .I3(GND_net), .O(n1823));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1175_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1185_3_lut (.I0(n528), .I1(n1801), 
            .I2(n1752), .I3(GND_net), .O(n1833));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1185_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i11_1_lut (.I0(encoder1_position_scaled[10]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n15_adj_5326));   // verilog/TinyFPGA_B.v(340[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_i1184_3_lut (.I0(n1733), .I1(n1800), 
            .I2(n1752), .I3(GND_net), .O(n1832));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1184_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i16_3_lut (.I0(encoder0_position[15]), 
            .I1(n18_adj_5297), .I2(encoder0_position[31]), .I3(GND_net), 
            .O(n529));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_mux_3_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i1179_3_lut (.I0(n1728), .I1(n1795), 
            .I2(n1752), .I3(GND_net), .O(n1827));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1179_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 unary_minus_19_inv_0_i6_1_lut (.I0(duty[5]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n20_adj_5265));   // verilog/TinyFPGA_B.v(123[25:30])
    defparam unary_minus_19_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_i1178_3_lut (.I0(n1727), .I1(n1794), 
            .I2(n1752), .I3(GND_net), .O(n1826));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1178_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1180_3_lut (.I0(n1729), .I1(n1796), 
            .I2(n1752), .I3(GND_net), .O(n1828));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1180_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i12_1_lut (.I0(encoder1_position_scaled[11]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n14_adj_5327));   // verilog/TinyFPGA_B.v(340[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_i1177_3_lut (.I0(n1726), .I1(n1793), 
            .I2(n1752), .I3(GND_net), .O(n1825));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1177_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15589_3_lut (.I0(\data_out_frame[23] [4]), .I1(neopxl_color[20]), 
            .I2(n24278), .I3(GND_net), .O(n29537));   // verilog/coms.v(128[12] 303[6])
    defparam i15589_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15590_3_lut (.I0(\data_out_frame[23] [3]), .I1(neopxl_color[19]), 
            .I2(n24278), .I3(GND_net), .O(n29538));   // verilog/coms.v(128[12] 303[6])
    defparam i15590_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1895 (.I0(n1825), .I1(n1828), .I2(n1826), .I3(n1827), 
            .O(n46903));
    defparam i1_4_lut_adj_1895.LUT_INIT = 16'hfffe;
    SB_LUT4 i21468_3_lut (.I0(n529), .I1(n1832), .I2(n1833), .I3(GND_net), 
            .O(n35416));
    defparam i21468_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i15591_3_lut (.I0(\data_out_frame[23] [2]), .I1(neopxl_color[18]), 
            .I2(n24278), .I3(GND_net), .O(n29539));   // verilog/coms.v(128[12] 303[6])
    defparam i15591_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i13_1_lut (.I0(encoder1_position_scaled[12]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n13_adj_5328));   // verilog/TinyFPGA_B.v(340[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_3_lut_adj_1896 (.I0(n1823), .I1(n1824), .I2(n46903), .I3(GND_net), 
            .O(n46907));
    defparam i1_3_lut_adj_1896.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_4_lut_adj_1897 (.I0(n1829), .I1(n35416), .I2(n1830), .I3(n1831), 
            .O(n44970));
    defparam i1_4_lut_adj_1897.LUT_INIT = 16'ha080;
    SB_LUT4 i1_4_lut_adj_1898 (.I0(n1821), .I1(n1822), .I2(n44970), .I3(n46907), 
            .O(n46913));
    defparam i1_4_lut_adj_1898.LUT_INIT = 16'hfffe;
    SB_LUT4 i35395_4_lut (.I0(n1819), .I1(n1818), .I2(n1820), .I3(n46913), 
            .O(n1851));
    defparam i35395_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i14_1_lut (.I0(encoder1_position_scaled[13]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n12_adj_5329));   // verilog/TinyFPGA_B.v(340[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_19_inv_0_i7_1_lut (.I0(duty[6]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_5264));   // verilog/TinyFPGA_B.v(123[25:30])
    defparam unary_minus_19_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i15_1_lut (.I0(encoder1_position_scaled[14]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n11_adj_5330));   // verilog/TinyFPGA_B.v(340[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    TLI4970 tli (.n29164(n29164), .\data[8] (data_adj_5514[8]), .n29160(n29160), 
            .\data[7] (data_adj_5514[7]), .n10(n10_adj_5341), .GND_net(GND_net), 
            .n11(n11_adj_5367), .n15(n15_adj_5339), .\state[1] (state_adj_5516[1]), 
            .\state[0] (state_adj_5516[0]), .n29154(n29154), .\data[6] (data_adj_5514[6]), 
            .CLK_c(CLK_c), .n29152(n29152), .\data[5] (data_adj_5514[5]), 
            .n29138(n29138), .\data[4] (data_adj_5514[4]), .n34688(n34688), 
            .VCC_net(VCC_net), .\data[12] (data_adj_5514[12]), .n29103(n29103), 
            .\data[3] (data_adj_5514[3]), .n29073(n29073), .\data[2] (data_adj_5514[2]), 
            .n9(n9_adj_5289), .clk_out(clk_out), .n29057(n29057), .CS_c(CS_c), 
            .n29052(n29052), .\data[1] (data_adj_5514[1]), .n29051(n29051), 
            .\current[0] (current[0]), .n27177(n27177), .n28537(n28537), 
            .\current[15] (current[15]), .\data[15] (data_adj_5514[15]), 
            .n29553(n29553), .\current[1] (current[1]), .n29552(n29552), 
            .\current[2] (current[2]), .n29551(n29551), .\current[3] (current[3]), 
            .n29550(n29550), .\current[4] (current[4]), .n29549(n29549), 
            .\current[5] (current[5]), .n29548(n29548), .\current[6] (current[6]), 
            .n29547(n29547), .\current[7] (current[7]), .n29546(n29546), 
            .\current[8] (current[8]), .n29545(n29545), .\current[9] (current[9]), 
            .n29544(n29544), .\current[10] (current[10]), .state_7__N_4460(state_7__N_4460), 
            .n29543(n29543), .\current[11] (current[11]), .n27143(n27143), 
            .n6(n6), .n29324(n29324), .n29323(n29323), .n29290(n29290), 
            .\data[11] (data_adj_5514[11]), .n29288(n29288), .\data[10] (data_adj_5514[10]), 
            .n29238(n29238), .\data[0] (data_adj_5514[0]), .n29184(n29184), 
            .\data[9] (data_adj_5514[9]), .n34690(n34690), .n27167(n27167), 
            .n27180(n27180), .n6_adj_14(n6_adj_5340), .n27174(n27174), 
            .CS_CLK_c(CS_CLK_c), .n5(n5_adj_5347)) /* synthesis syn_noprune=1, syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(418[11] 424[4])
    SB_LUT4 i15301_3_lut_4_lut (.I0(n1855), .I1(b_prev), .I2(a_new[1]), 
            .I3(direction_N_4071), .O(n29249));   // vhdl/quadrature_decoder.vhd(52[3] 89[10])
    defparam i15301_3_lut_4_lut.LUT_INIT = 16'h3caa;
    SB_LUT4 i15297_3_lut_4_lut (.I0(n1896), .I1(b_prev_adj_5344), .I2(a_new_adj_5490[1]), 
            .I3(direction_N_4071_adj_5345), .O(n29245));   // vhdl/quadrature_decoder.vhd(52[3] 89[10])
    defparam i15297_3_lut_4_lut.LUT_INIT = 16'h3caa;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i16_1_lut (.I0(encoder1_position_scaled[15]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n10_adj_5331));   // verilog/TinyFPGA_B.v(340[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i5498_3_lut_4_lut_4_lut (.I0(commutation_state[2]), .I1(commutation_state[1]), 
            .I2(dir), .I3(commutation_state[0]), .O(GHB_N_413));
    defparam i5498_3_lut_4_lut_4_lut.LUT_INIT = 16'hc121;
    SB_LUT4 mux_1005_i15_3_lut (.I0(duty[14]), .I1(n349), .I2(duty[23]), 
            .I3(GND_net), .O(n4709));   // verilog/TinyFPGA_B.v(118[13] 129[7])
    defparam mux_1005_i15_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n10621_bdd_4_lut (.I0(n10621), .I1(current[15]), .I2(duty[23]), 
            .I3(n4208), .O(n51468));
    defparam n10621_bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i17_1_lut (.I0(encoder1_position_scaled[16]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n9_adj_5332));   // verilog/TinyFPGA_B.v(340[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i18_1_lut (.I0(encoder1_position_scaled[17]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n8_adj_5333));   // verilog/TinyFPGA_B.v(340[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i19_1_lut (.I0(encoder1_position_scaled[18]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n7_adj_5334));   // verilog/TinyFPGA_B.v(340[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i15592_3_lut (.I0(\data_out_frame[23] [1]), .I1(neopxl_color[17]), 
            .I2(n24278), .I3(GND_net), .O(n29540));   // verilog/coms.v(128[12] 303[6])
    defparam i15592_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i20_1_lut (.I0(encoder1_position_scaled[19]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n6_adj_5335));   // verilog/TinyFPGA_B.v(340[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_1005_i16_3_lut (.I0(duty[15]), .I1(n348), .I2(duty[23]), 
            .I3(GND_net), .O(n4708));   // verilog/TinyFPGA_B.v(118[13] 129[7])
    defparam mux_1005_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i21_1_lut (.I0(encoder1_position_scaled[20]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n5_adj_5336));   // verilog/TinyFPGA_B.v(340[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i20621_2_lut (.I0(pwm_out), .I1(GHC), .I2(GND_net), .I3(GND_net), 
            .O(INHC_c_0));   // verilog/TinyFPGA_B.v(84[16:31])
    defparam i20621_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i20620_2_lut (.I0(pwm_out), .I1(GHB), .I2(GND_net), .I3(GND_net), 
            .O(INHB_c_0));   // verilog/TinyFPGA_B.v(82[16:31])
    defparam i20620_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i20712_2_lut (.I0(pwm_out), .I1(GHA), .I2(GND_net), .I3(GND_net), 
            .O(INHA_c_0));   // verilog/TinyFPGA_B.v(80[16:31])
    defparam i20712_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i5500_3_lut_4_lut_4_lut (.I0(commutation_state[2]), .I1(commutation_state[1]), 
            .I2(dir), .I3(commutation_state[0]), .O(GLB_N_422));
    defparam i5500_3_lut_4_lut_4_lut.LUT_INIT = 16'h1c12;
    SB_LUT4 unary_minus_19_inv_0_i8_1_lut (.I0(duty[7]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n18_adj_5263));   // verilog/TinyFPGA_B.v(123[25:30])
    defparam unary_minus_19_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i22_1_lut (.I0(encoder1_position_scaled[21]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n4_adj_5337));   // verilog/TinyFPGA_B.v(340[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i23_1_lut (.I0(encoder1_position_scaled[22]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n3_adj_5338));   // verilog/TinyFPGA_B.v(340[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 LessThan_11_i6_3_lut_3_lut (.I0(duty[2]), .I1(duty[3]), .I2(current[3]), 
            .I3(GND_net), .O(n6_adj_5242));   // verilog/TinyFPGA_B.v(111[10:22])
    defparam LessThan_11_i6_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 LessThan_11_i8_3_lut_3_lut (.I0(duty[4]), .I1(duty[8]), .I2(current[8]), 
            .I3(GND_net), .O(n8_adj_5342));   // verilog/TinyFPGA_B.v(111[10:22])
    defparam LessThan_11_i8_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i24_1_lut (.I0(encoder1_position_scaled[23]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n2_adj_5278));   // verilog/TinyFPGA_B.v(340[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_i1105_3_lut (.I0(n1622), .I1(n1689), 
            .I2(n1653), .I3(GND_net), .O(n1721));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1105_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1104_3_lut (.I0(n1621), .I1(n1688), 
            .I2(n1653), .I3(GND_net), .O(n1720));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1104_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1106_3_lut (.I0(n1623), .I1(n1690), 
            .I2(n1653), .I3(GND_net), .O(n1722));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1106_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1111_3_lut (.I0(n1628), .I1(n1695), 
            .I2(n1653), .I3(GND_net), .O(n1727));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1111_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1109_3_lut (.I0(n1626), .I1(n1693), 
            .I2(n1653), .I3(GND_net), .O(n1725));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1109_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1117_3_lut (.I0(n527), .I1(n1701), 
            .I2(n1653), .I3(GND_net), .O(n1733));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1117_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1116_3_lut (.I0(n1633), .I1(n1700), 
            .I2(n1653), .I3(GND_net), .O(n1732));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1116_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i17_3_lut (.I0(encoder0_position[16]), 
            .I1(n17_adj_5298), .I2(encoder0_position[31]), .I3(GND_net), 
            .O(n528));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_mux_3_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i1115_3_lut (.I0(n1632), .I1(n1699), 
            .I2(n1653), .I3(GND_net), .O(n1731));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1115_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1114_3_lut (.I0(n1631), .I1(n1698), 
            .I2(n1653), .I3(GND_net), .O(n1730));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1114_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1113_3_lut (.I0(n1630), .I1(n1697), 
            .I2(n1653), .I3(GND_net), .O(n1729));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1113_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1110_3_lut (.I0(n1627), .I1(n1694), 
            .I2(n1653), .I3(GND_net), .O(n1726));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1110_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1112_3_lut (.I0(n1629), .I1(n1696), 
            .I2(n1653), .I3(GND_net), .O(n1728));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1112_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1107_3_lut (.I0(n1624), .I1(n1691), 
            .I2(n1653), .I3(GND_net), .O(n1723));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1107_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1108_3_lut (.I0(n1625), .I1(n1692), 
            .I2(n1653), .I3(GND_net), .O(n1724));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1108_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i21470_3_lut (.I0(n528), .I1(n1732), .I2(n1733), .I3(GND_net), 
            .O(n35418));
    defparam i21470_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i1_2_lut_adj_1899 (.I0(n1725), .I1(n1727), .I2(GND_net), .I3(GND_net), 
            .O(n46801));
    defparam i1_2_lut_adj_1899.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_1900 (.I0(n1724), .I1(n1723), .I2(n1728), .I3(n1726), 
            .O(n45982));
    defparam i1_4_lut_adj_1900.LUT_INIT = 16'hfffe;
    SB_LUT4 LessThan_11_i10_3_lut_3_lut (.I0(duty[5]), .I1(duty[6]), .I2(current[6]), 
            .I3(GND_net), .O(n10_adj_5275));   // verilog/TinyFPGA_B.v(111[10:22])
    defparam LessThan_11_i10_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i1_4_lut_adj_1901 (.I0(n1729), .I1(n35418), .I2(n1730), .I3(n1731), 
            .O(n44929));
    defparam i1_4_lut_adj_1901.LUT_INIT = 16'ha080;
    SB_LUT4 i1_4_lut_adj_1902 (.I0(n1722), .I1(n44929), .I2(n45982), .I3(n46801), 
            .O(n46807));
    defparam i1_4_lut_adj_1902.LUT_INIT = 16'hfffe;
    SB_LUT4 i35415_4_lut (.I0(n1720), .I1(n1719), .I2(n1721), .I3(n46807), 
            .O(n1752));
    defparam i35415_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_31__I_0_i1038_3_lut (.I0(n1523), .I1(n1590), 
            .I2(n1554), .I3(GND_net), .O(n1622));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1038_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_1005_i17_3_lut (.I0(duty[16]), .I1(n347), .I2(duty[23]), 
            .I3(GND_net), .O(n4707));   // verilog/TinyFPGA_B.v(118[13] 129[7])
    defparam mux_1005_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i1037_3_lut (.I0(n1522), .I1(n1589), 
            .I2(n1554), .I3(GND_net), .O(n1621));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1037_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1040_3_lut (.I0(n1525), .I1(n1592), 
            .I2(n1554), .I3(GND_net), .O(n1624));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1040_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 unary_minus_19_inv_0_i9_1_lut (.I0(duty[8]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_5262));   // verilog/TinyFPGA_B.v(123[25:30])
    defparam unary_minus_19_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_i1039_3_lut (.I0(n1524), .I1(n1591), 
            .I2(n1554), .I3(GND_net), .O(n1623));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1039_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_1005_i18_3_lut (.I0(duty[17]), .I1(n346), .I2(duty[23]), 
            .I3(GND_net), .O(n4706));   // verilog/TinyFPGA_B.v(118[13] 129[7])
    defparam mux_1005_i18_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i1047_3_lut (.I0(n1532), .I1(n1599), 
            .I2(n1554), .I3(GND_net), .O(n1631));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1047_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1046_3_lut (.I0(n1531), .I1(n1598), 
            .I2(n1554), .I3(GND_net), .O(n1630));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1046_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1045_3_lut (.I0(n1530), .I1(n1597), 
            .I2(n1554), .I3(GND_net), .O(n1629));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1045_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1043_3_lut (.I0(n1528), .I1(n1595), 
            .I2(n1554), .I3(GND_net), .O(n1627));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1043_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1042_3_lut (.I0(n1527), .I1(n1594), 
            .I2(n1554), .I3(GND_net), .O(n1626));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1042_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1044_3_lut (.I0(n1529), .I1(n1596), 
            .I2(n1554), .I3(GND_net), .O(n1628));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1044_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1041_3_lut (.I0(n1526), .I1(n1593), 
            .I2(n1554), .I3(GND_net), .O(n1625));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1041_3_lut.LUT_INIT = 16'hacac;
    coms neopxl_color_23__I_0 (.\data_out_frame[13] ({\data_out_frame[13] }), 
         .GND_net(GND_net), .\data_out_frame[20] ({\data_out_frame[20] }), 
         .\data_out_frame[23] ({\data_out_frame[23] }), .CLK_c(CLK_c), .\data_in_frame[3] ({\data_in_frame[3] }), 
         .\data_out_frame[25] ({\data_out_frame[25] }), .\data_in_frame[5] ({\data_in_frame[5] }), 
         .rx_data({rx_data}), .\data_out_frame[10] ({\data_out_frame[10] }), 
         .\data_out_frame[6] ({\data_out_frame[6] }), .\data_out_frame[8] ({\data_out_frame[8] }), 
         .\data_out_frame[17] ({\data_out_frame[17] }), .\data_out_frame[15] ({\data_out_frame[15] }), 
         .\data_out_frame[16] ({\data_out_frame[16] }), .\data_out_frame[19] ({\data_out_frame[19] }), 
         .\data_out_frame[21] ({\data_out_frame[21] }), .\data_out_frame[12] ({\data_out_frame[12] }), 
         .\data_out_frame[14] ({\data_out_frame[14] }), .\data_out_frame[5] ({\data_out_frame[5] }), 
         .\data_out_frame[4] ({\data_out_frame[4] }), .\data_in_frame[11] ({\data_in_frame[11] }), 
         .\data_in_frame[14] ({\data_in_frame[14] }), .\data_in_frame[13] ({\data_in_frame[13] }), 
         .\data_out_frame[11] ({\data_out_frame[11] }), .\data_out_frame[9] ({\data_out_frame[9] }), 
         .\data_out_frame[7] ({\data_out_frame[7] }), .\data_in_frame[10] ({\data_in_frame[10] }), 
         .\data_in_frame[12] ({\data_in_frame[12] }), .\data_out_frame[18] ({\data_out_frame[18] }), 
         .\data_out_frame[22] ({\data_out_frame[22] }), .\data_in_frame[1] ({\data_in_frame[1] }), 
         .n29158(n29158), .IntegralLimit({IntegralLimit}), .\data_in[1] ({\data_in[1] }), 
         .\data_in[3] ({\data_in[3] }), .\data_in[0] ({\data_in[0] }), .\data_in_frame[21] ({\data_in_frame[21] }), 
         .n29157(n29157), .n29156(n29156), .n29155(n29155), .\data_in_frame[2] ({\data_in_frame[2] }), 
         .\data_in_frame[20] ({\data_in_frame[20] }), .\data_in_frame[9] ({\data_in_frame[9] }), 
         .\data_in_frame[4] ({\data_in_frame[4] }), .rx_data_ready(rx_data_ready), 
         .setpoint({setpoint}), .\data_in_frame[6] ({\data_in_frame[6] }), 
         .n29153(n29153), .n29151(n29151), .n29018(n29018), .n29150(n29150), 
         .n29149(n29149), .n29148(n29148), .n29147(n29147), .n29145(n29145), 
         .n29144(n29144), .n29143(n29143), .n29142(n29142), .n29141(n29141), 
         .n29140(n29140), .n29139(n29139), .n29137(n29137), .n29136(n29136), 
         .n29135(n29135), .n29134(n29134), .n29133(n29133), .n29132(n29132), 
         .n29131(n29131), .n29130(n29130), .n29129(n29129), .ID({ID}), 
         .n29128(n29128), .n29127(n29127), .\data_in_frame[8] ({\data_in_frame[8] }), 
         .\data_out_frame[24] ({\data_out_frame[24] }), .n29126(n29126), 
         .n29125(n29125), .\data_in_frame[22] ({\data_in_frame[22] }), .n29124(n29124), 
         .n29123(n29123), .n29122(n29122), .n29121(n29121), .n29120(n29120), 
         .n29119(n29119), .n29118(n29118), .n29117(n29117), .n29116(n29116), 
         .n29115(n29115), .n29114(n29114), .n29113(n29113), .n29112(n29112), 
         .n29111(n29111), .n29110(n29110), .n29109(n29109), .n29108(n29108), 
         .n29107(n29107), .n28521(n28521), .n29106(n29106), .n29105(n29105), 
         .\data_in[2] ({\data_in[2] }), .n29679(n29679), .n29678(n29678), 
         .n29677(n29677), .n29676(n29676), .n29675(n29675), .n29674(n29674), 
         .n29673(n29673), .n29672(n29672), .n29671(n29671), .n29670(n29670), 
         .n29669(n29669), .n29668(n29668), .n29667(n29667), .n29666(n29666), 
         .n29665(n29665), .n29664(n29664), .n29663(n29663), .n29662(n29662), 
         .n29661(n29661), .n29660(n29660), .n29659(n29659), .n29658(n29658), 
         .n29657(n29657), .n29656(n29656), .n29655(n29655), .n29654(n29654), 
         .n29653(n29653), .n29652(n29652), .n29651(n29651), .n29650(n29650), 
         .n29649(n29649), .n29648(n29648), .n29647(n29647), .n29646(n29646), 
         .n29645(n29645), .n29644(n29644), .n29643(n29643), .n29642(n29642), 
         .n29641(n29641), .n29640(n29640), .n29639(n29639), .n29638(n29638), 
         .n29637(n29637), .n29636(n29636), .n29635(n29635), .n29634(n29634), 
         .n29633(n29633), .n29632(n29632), .n29631(n29631), .n29630(n29630), 
         .n29629(n29629), .n29628(n29628), .n29104(n29104), .n29102(n29102), 
         .n29101(n29101), .n29100(n29100), .n29099(n29099), .n29098(n29098), 
         .n29097(n29097), .n29096(n29096), .n29095(n29095), .n29094(n29094), 
         .n29093(n29093), .n29092(n29092), .n29091(n29091), .n29090(n29090), 
         .n29089(n29089), .n29088(n29088), .n29087(n29087), .n29086(n29086), 
         .n29085(n29085), .n29084(n29084), .n29083(n29083), .n29082(n29082), 
         .n29081(n29081), .n29080(n29080), .n29079(n29079), .n29078(n29078), 
         .n29077(n29077), .n29076(n29076), .n29075(n29075), .n29074(n29074), 
         .DE_c(DE_c), .n29067(n29067), .n29065(n29065), .n29064(n29064), 
         .n29063(n29063), .n29062(n29062), .n29061(n29061), .n29060(n29060), 
         .n29056(n29056), .n29627(n29627), .LED_c(LED_c), .n29626(n29626), 
         .n29625(n29625), .n29624(n29624), .n29623(n29623), .n29622(n29622), 
         .n29621(n29621), .n29620(n29620), .n29619(n29619), .n29618(n29618), 
         .n29617(n29617), .n29616(n29616), .n29615(n29615), .n29614(n29614), 
         .n29613(n29613), .n29612(n29612), .n29611(n29611), .n29610(n29610), 
         .n29609(n29609), .n29608(n29608), .n29607(n29607), .n29606(n29606), 
         .n29605(n29605), .n29604(n29604), .n29602(n29602), .n29599(n29599), 
         .control_mode({control_mode}), .n29598(n29598), .n29597(n29597), 
         .n29596(n29596), .n29595(n29595), .n29055(n29055), .n29050(n29050), 
         .n29049(n29049), .n29047(n29047), .PWMLimit({PWMLimit}), .n29046(n29046), 
         .current_limit({current_limit}), .n29045(n29045), .n29043(n29043), 
         .neopxl_color({neopxl_color}), .n29042(n29042), .\Ki[0] (Ki[0]), 
         .n29041(n29041), .\Kp[0] (Kp[0]), .n29040(n29040), .n29026(n29026), 
         .n29594(n29594), .n29593(n29593), .n29592(n29592), .n29591(n29591), 
         .n29590(n29590), .n29024(n29024), .n29589(n29589), .n29023(n29023), 
         .n29588(n29588), .n29587(n29587), .n29586(n29586), .n29585(n29585), 
         .n29584(n29584), .n29583(n29583), .n29582(n29582), .n29581(n29581), 
         .n29580(n29580), .n29579(n29579), .n29578(n29578), .n29577(n29577), 
         .n29576(n29576), .n29575(n29575), .n29574(n29574), .n29573(n29573), 
         .n43838(n43838), .n29572(n29572), .n29571(n29571), .n29570(n29570), 
         .n29569(n29569), .n29568(n29568), .n43847(n43847), .n43822(n43822), 
         .n29567(n29567), .n29566(n29566), .n29021(n29021), .n29565(n29565), 
         .n29564(n29564), .n29563(n29563), .n29562(n29562), .n29561(n29561), 
         .n29560(n29560), .n29559(n29559), .n29558(n29558), .n29557(n29557), 
         .n29556(n29556), .n29555(n29555), .n24278(n24278), .n29020(n29020), 
         .n29542(n29542), .n29541(n29541), .n29540(n29540), .n29539(n29539), 
         .n29538(n29538), .n29537(n29537), .n29529(n29529), .n29528(n29528), 
         .n29527(n29527), .n29526(n29526), .n29525(n29525), .n29523(n29523), 
         .n29522(n29522), .n29521(n29521), .n29520(n29520), .n29519(n29519), 
         .n29518(n29518), .n29517(n29517), .n29506(n29506), .n29505(n29505), 
         .n29504(n29504), .n29503(n29503), .n29501(n29501), .n29500(n29500), 
         .n29499(n29499), .n29466(n29466), .n29465(n29465), .n29464(n29464), 
         .n29463(n29463), .n29462(n29462), .n29461(n29461), .n29460(n29460), 
         .n29459(n29459), .n29458(n29458), .n29457(n29457), .n29456(n29456), 
         .n29455(n29455), .n29454(n29454), .n29453(n29453), .n29452(n29452), 
         .n29451(n29451), .n29450(n29450), .n29449(n29449), .n29448(n29448), 
         .n29447(n29447), .n29446(n29446), .n29445(n29445), .n29444(n29444), 
         .n28522(n28522), .n29403(n29403), .n29402(n29402), .n29401(n29401), 
         .n29400(n29400), .n29399(n29399), .n29398(n29398), .n29397(n29397), 
         .n29396(n29396), .n29395(n29395), .n29394(n29394), .n29393(n29393), 
         .n29392(n29392), .n29391(n29391), .n29390(n29390), .n29389(n29389), 
         .n29388(n29388), .n29339(n29339), .n29338(n29338), .n29336(n29336), 
         .n29335(n29335), .n29334(n29334), .n29333(n29333), .n29332(n29332), 
         .n29331(n29331), .n29330(n29330), .n29329(n29329), .n29328(n29328), 
         .n29327(n29327), .n29326(n29326), .n29325(n29325), .n29322(n29322), 
         .n29321(n29321), .n29270(n29270), .n29269(n29269), .n29268(n29268), 
         .n29267(n29267), .n29266(n29266), .n29265(n29265), .n29264(n29264), 
         .n29263(n29263), .n29262(n29262), .n29261(n29261), .n29260(n29260), 
         .n29259(n29259), .n29258(n29258), .n29257(n29257), .n29256(n29256), 
         .n29255(n29255), .n29244(n29244), .n29243(n29243), .n29242(n29242), 
         .n29241(n29241), .n29240(n29240), .n29239(n29239), .n29225(n29225), 
         .n29224(n29224), .n29223(n29223), .n29221(n29221), .n29220(n29220), 
         .n29219(n29219), .n29218(n29218), .n29217(n29217), .n29216(n29216), 
         .n29215(n29215), .n29214(n29214), .n29213(n29213), .n29212(n29212), 
         .n29211(n29211), .n29210(n29210), .n29209(n29209), .n29208(n29208), 
         .n29207(n29207), .n29206(n29206), .n29205(n29205), .n29204(n29204), 
         .n29203(n29203), .n29202(n29202), .n29201(n29201), .n29200(n29200), 
         .n29199(n29199), .\Kp[1] (Kp[1]), .n29198(n29198), .\Kp[2] (Kp[2]), 
         .n29197(n29197), .\Kp[3] (Kp[3]), .n29196(n29196), .\Kp[4] (Kp[4]), 
         .n29195(n29195), .\Kp[5] (Kp[5]), .n29194(n29194), .\Kp[6] (Kp[6]), 
         .n29193(n29193), .\Kp[7] (Kp[7]), .n29192(n29192), .\Kp[8] (Kp[8]), 
         .n29191(n29191), .\Kp[9] (Kp[9]), .n29190(n29190), .\Kp[10] (Kp[10]), 
         .n29189(n29189), .\Kp[11] (Kp[11]), .n29188(n29188), .\Kp[12] (Kp[12]), 
         .n29187(n29187), .\Kp[13] (Kp[13]), .n29183(n29183), .\Kp[14] (Kp[14]), 
         .n29182(n29182), .\Kp[15] (Kp[15]), .n29181(n29181), .\Ki[1] (Ki[1]), 
         .n29180(n29180), .\Ki[2] (Ki[2]), .n29179(n29179), .\Ki[3] (Ki[3]), 
         .n29178(n29178), .\Ki[4] (Ki[4]), .n29177(n29177), .\Ki[5] (Ki[5]), 
         .n29176(n29176), .\Ki[6] (Ki[6]), .n29175(n29175), .\Ki[7] (Ki[7]), 
         .n29174(n29174), .\Ki[8] (Ki[8]), .n29173(n29173), .\Ki[9] (Ki[9]), 
         .n29172(n29172), .\Ki[10] (Ki[10]), .n29171(n29171), .\Ki[11] (Ki[11]), 
         .n29019(n29019), .n29170(n29170), .\Ki[12] (Ki[12]), .n29169(n29169), 
         .\Ki[13] (Ki[13]), .n29168(n29168), .\Ki[14] (Ki[14]), .n29167(n29167), 
         .\Ki[15] (Ki[15]), .\state[0] (state_adj_5537[0]), .\state[2] (state_adj_5537[2]), 
         .\state[3] (state_adj_5537[3]), .n7754(n7754), .n43824(n43824), 
         .n43848(n43848), .n43839(n43839), .tx_active(tx_active), .\r_Bit_Index[0] (r_Bit_Index_adj_5527[0]), 
         .tx_o(tx_o), .r_SM_Main({r_SM_Main_adj_5525}), .VCC_net(VCC_net), 
         .\r_SM_Main_2__N_3777[1] (r_SM_Main_2__N_3777[1]), .n29230(n29230), 
         .n51602(n51602), .n29066(n29066), .n28662(n28662), .n28970(n28970), 
         .n19541(n19541), .n4(n4_adj_5272), .tx_enable(tx_enable), .\r_SM_Main_2__N_3706[2] (r_SM_Main_2__N_3706[2]), 
         .n4_adj_6(n4_adj_5287), .r_SM_Main_adj_13({r_SM_Main}), .r_Rx_Data(r_Rx_Data), 
         .RX_N_10(RX_N_10), .\r_Bit_Index[0]_adj_10 (r_Bit_Index[0]), .n4_adj_11(n4_adj_5245), 
         .n4_adj_12(n4_adj_5362), .n34695(n34695), .n29233(n29233), .n43326(n43326), 
         .n28666(n28666), .n28972(n28972), .n28562(n28562), .n29524(n29524), 
         .n29516(n29516), .n29510(n29510), .n29508(n29508), .n29502(n29502), 
         .n29467(n29467), .n29404(n29404), .n43724(n43724), .n29237(n29237), 
         .n27131(n27131), .n27126(n27126)) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(255[8] 279[4])
    SB_LUT4 encoder0_position_31__I_0_i1049_3_lut (.I0(n526), .I1(n1601), 
            .I2(n1554), .I3(GND_net), .O(n1633));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1049_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1048_3_lut (.I0(n1533), .I1(n1600), 
            .I2(n1554), .I3(GND_net), .O(n1632));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i1048_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i18_3_lut (.I0(encoder0_position[17]), 
            .I1(n16_adj_5299), .I2(encoder0_position[31]), .I3(GND_net), 
            .O(n527));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_mux_3_i18_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i21472_3_lut (.I0(n527), .I1(n1632), .I2(n1633), .I3(GND_net), 
            .O(n35420));
    defparam i21472_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i1_4_lut_adj_1903 (.I0(n1625), .I1(n1628), .I2(n1626), .I3(n1627), 
            .O(n46881));
    defparam i1_4_lut_adj_1903.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1904 (.I0(n1629), .I1(n35420), .I2(n1630), .I3(n1631), 
            .O(n44933));
    defparam i1_4_lut_adj_1904.LUT_INIT = 16'ha080;
    SB_LUT4 i1_4_lut_adj_1905 (.I0(n1623), .I1(n44933), .I2(n1624), .I3(n46881), 
            .O(n46887));
    defparam i1_4_lut_adj_1905.LUT_INIT = 16'hfffe;
    SB_LUT4 i35434_4_lut (.I0(n1621), .I1(n1620), .I2(n1622), .I3(n46887), 
            .O(n1653));
    defparam i35434_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_31__I_0_i971_3_lut (.I0(n1424), .I1(n1491), 
            .I2(n1455), .I3(GND_net), .O(n1523));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i971_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i970_3_lut (.I0(n1423), .I1(n1490), 
            .I2(n1455), .I3(GND_net), .O(n1522));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i970_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_1005_i19_3_lut (.I0(duty[18]), .I1(n345), .I2(duty[23]), 
            .I3(GND_net), .O(n4705));   // verilog/TinyFPGA_B.v(118[13] 129[7])
    defparam mux_1005_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i978_3_lut (.I0(n1431), .I1(n1498), 
            .I2(n1455), .I3(GND_net), .O(n1530));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i978_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i977_3_lut (.I0(n1430), .I1(n1497), 
            .I2(n1455), .I3(GND_net), .O(n1529));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i977_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_1005_i20_3_lut (.I0(duty[19]), .I1(n344), .I2(duty[23]), 
            .I3(GND_net), .O(n4704));   // verilog/TinyFPGA_B.v(118[13] 129[7])
    defparam mux_1005_i20_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i974_3_lut (.I0(n1427), .I1(n1494), 
            .I2(n1455), .I3(GND_net), .O(n1526));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i974_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i973_3_lut (.I0(n1426), .I1(n1493), 
            .I2(n1455), .I3(GND_net), .O(n1525));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i973_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i972_3_lut (.I0(n1425), .I1(n1492), 
            .I2(n1455), .I3(GND_net), .O(n1524));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i972_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i981_3_lut (.I0(n525), .I1(n1501), 
            .I2(n1455), .I3(GND_net), .O(n1533));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i981_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i980_3_lut (.I0(n1433), .I1(n1500), 
            .I2(n1455), .I3(GND_net), .O(n1532));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i980_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i979_3_lut (.I0(n1432), .I1(n1499), 
            .I2(n1455), .I3(GND_net), .O(n1531));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i979_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i19_3_lut (.I0(encoder0_position[18]), 
            .I1(n15_adj_5300), .I2(encoder0_position[31]), .I3(GND_net), 
            .O(n526));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_mux_3_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i975_3_lut (.I0(n1428), .I1(n1495), 
            .I2(n1455), .I3(GND_net), .O(n1527));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i975_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i976_3_lut (.I0(n1429), .I1(n1496), 
            .I2(n1455), .I3(GND_net), .O(n1528));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i976_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 unary_minus_19_inv_0_i10_1_lut (.I0(duty[9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n16_adj_5261));   // verilog/TinyFPGA_B.v(123[25:30])
    defparam unary_minus_19_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_2_lut_adj_1906 (.I0(n1528), .I1(n1527), .I2(GND_net), .I3(GND_net), 
            .O(n46603));
    defparam i1_2_lut_adj_1906.LUT_INIT = 16'heeee;
    SB_LUT4 i21535_4_lut (.I0(n526), .I1(n1531), .I2(n1532), .I3(n1533), 
            .O(n35484));
    defparam i21535_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 i1_4_lut_adj_1907 (.I0(n1524), .I1(n1525), .I2(n1526), .I3(n46603), 
            .O(n46609));
    defparam i1_4_lut_adj_1907.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1908 (.I0(n1529), .I1(n46609), .I2(n35484), .I3(n1530), 
            .O(n46611));
    defparam i1_4_lut_adj_1908.LUT_INIT = 16'heccc;
    SB_LUT4 i35452_4_lut (.I0(n1522), .I1(n1521), .I2(n46611), .I3(n1523), 
            .O(n1554));
    defparam i35452_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 LessThan_15_i6_3_lut_3_lut (.I0(current_limit[2]), .I1(current_limit[3]), 
            .I2(current[3]), .I3(GND_net), .O(n6_adj_5364));   // verilog/TinyFPGA_B.v(119[9:30])
    defparam LessThan_15_i6_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i33828_2_lut_4_lut (.I0(current[8]), .I1(current_limit[8]), 
            .I2(current[4]), .I3(current_limit[4]), .O(n49415));
    defparam i33828_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 LessThan_15_i8_3_lut_3_lut (.I0(current_limit[4]), .I1(current_limit[8]), 
            .I2(current[8]), .I3(GND_net), .O(n8_adj_5350));   // verilog/TinyFPGA_B.v(119[9:30])
    defparam LessThan_15_i8_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i20719_1_lut_2_lut (.I0(n24462), .I1(dti), .I2(GND_net), .I3(GND_net), 
            .O(n2195));
    defparam i20719_1_lut_2_lut.LUT_INIT = 16'h7777;
    \quadrature_decoder(1,500000)  quad_counter1 (.n1891(CLK_c), .b_prev(b_prev_adj_5344), 
            .GND_net(GND_net), .a_new({a_new_adj_5490[1], Open_1}), .direction_N_4071(direction_N_4071_adj_5345), 
            .ENCODER1_B_N_keep(ENCODER1_B_N), .ENCODER1_A_N_keep(ENCODER1_A_N), 
            .encoder1_position({encoder1_position}), .VCC_net(VCC_net), 
            .n29245(n29245), .n1896(n1896)) /* synthesis lattice_noprune=1 */ ;   // verilog/TinyFPGA_B.v(312[57] 319[6])
    SB_LUT4 i15206_4_lut (.I0(CS_MISO_c), .I1(data_adj_5514[6]), .I2(n6_adj_5340), 
            .I3(n27177), .O(n29154));   // verilog/tli4970.v(35[10] 68[6])
    defparam i15206_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 encoder0_position_31__I_0_i903_3_lut (.I0(n1324_adj_5394), .I1(n1391), 
            .I2(n1356), .I3(GND_net), .O(n1423));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i903_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i906_3_lut (.I0(n1327_adj_5397), .I1(n1394), 
            .I2(n1356), .I3(GND_net), .O(n1426));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i906_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i905_3_lut (.I0(n1326_adj_5396), .I1(n1393), 
            .I2(n1356), .I3(GND_net), .O(n1425));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i905_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i904_3_lut (.I0(n1325_adj_5395), .I1(n1392), 
            .I2(n1356), .I3(GND_net), .O(n1424));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i904_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i908_3_lut (.I0(n1329), .I1(n1396), 
            .I2(n1356), .I3(GND_net), .O(n1428));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i908_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i907_3_lut (.I0(n1328_adj_5398), .I1(n1395), 
            .I2(n1356), .I3(GND_net), .O(n1427));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i907_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i911_3_lut (.I0(n1332), .I1(n1399), 
            .I2(n1356), .I3(GND_net), .O(n1431));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i911_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i910_3_lut (.I0(n1331), .I1(n1398), 
            .I2(n1356), .I3(GND_net), .O(n1430));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i910_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i909_3_lut (.I0(n1330), .I1(n1397), 
            .I2(n1356), .I3(GND_net), .O(n1429));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i909_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i913_3_lut (.I0(n938), .I1(n1401), 
            .I2(n1356), .I3(GND_net), .O(n1433));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i913_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i912_3_lut (.I0(n1333), .I1(n1400), 
            .I2(n1356), .I3(GND_net), .O(n1432));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i912_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i20_3_lut (.I0(encoder0_position[19]), 
            .I1(n14_adj_5301), .I2(encoder0_position[31]), .I3(GND_net), 
            .O(n525));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_mux_3_i20_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i21476_3_lut (.I0(n525), .I1(n1432), .I2(n1433), .I3(GND_net), 
            .O(n35424));
    defparam i21476_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i1_2_lut_adj_1909 (.I0(n1427), .I1(n1428), .I2(GND_net), .I3(GND_net), 
            .O(n46857));
    defparam i1_2_lut_adj_1909.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_1910 (.I0(n1429), .I1(n35424), .I2(n1430), .I3(n1431), 
            .O(n44924));
    defparam i1_4_lut_adj_1910.LUT_INIT = 16'ha080;
    SB_LUT4 i1_4_lut_adj_1911 (.I0(n1424), .I1(n1425), .I2(n1426), .I3(n46857), 
            .O(n46863));
    defparam i1_4_lut_adj_1911.LUT_INIT = 16'hfffe;
    SB_LUT4 i35469_4_lut (.I0(n1423), .I1(n1422), .I2(n46863), .I3(n44924), 
            .O(n1455));
    defparam i35469_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_31__I_0_i836_3_lut (.I0(n1225), .I1(n1292), 
            .I2(n1257), .I3(GND_net), .O(n1324_adj_5394));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i836_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i843_3_lut (.I0(n1232), .I1(n1299_adj_5390), 
            .I2(n1257), .I3(GND_net), .O(n1331));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i843_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i842_3_lut (.I0(n1231), .I1(n1298_adj_5389), 
            .I2(n1257), .I3(GND_net), .O(n1330));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i842_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i841_3_lut (.I0(n1230), .I1(n1297_adj_5388), 
            .I2(n1257), .I3(GND_net), .O(n1329));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i841_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i840_3_lut (.I0(n1229), .I1(n1296), 
            .I2(n1257), .I3(GND_net), .O(n1328_adj_5398));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i840_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i839_3_lut (.I0(n1228), .I1(n1295), 
            .I2(n1257), .I3(GND_net), .O(n1327_adj_5397));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i839_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i838_3_lut (.I0(n1227), .I1(n1294), 
            .I2(n1257), .I3(GND_net), .O(n1326_adj_5396));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i838_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i837_3_lut (.I0(n1226), .I1(n1293), 
            .I2(n1257), .I3(GND_net), .O(n1325_adj_5395));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i837_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i845_3_lut (.I0(n937), .I1(n1301_adj_5392), 
            .I2(n1257), .I3(GND_net), .O(n1333));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i845_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i844_3_lut (.I0(n1233), .I1(n1300_adj_5391), 
            .I2(n1257), .I3(GND_net), .O(n1332));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i844_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i21_3_lut (.I0(encoder0_position[20]), 
            .I1(n13_adj_5302), .I2(encoder0_position[31]), .I3(GND_net), 
            .O(n938));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_mux_3_i21_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i21478_3_lut (.I0(n938), .I1(n1332), .I2(n1333), .I3(GND_net), 
            .O(n35426));
    defparam i21478_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i1_4_lut_adj_1912 (.I0(n1325_adj_5395), .I1(n1326_adj_5396), 
            .I2(n1327_adj_5397), .I3(n1328_adj_5398), .O(n46793));
    defparam i1_4_lut_adj_1912.LUT_INIT = 16'hfffe;
    SB_LUT4 unary_minus_19_inv_0_i11_1_lut (.I0(duty[10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_5260));   // verilog/TinyFPGA_B.v(123[25:30])
    defparam unary_minus_19_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_4_lut_adj_1913 (.I0(n1329), .I1(n35426), .I2(n1330), .I3(n1331), 
            .O(n44905));
    defparam i1_4_lut_adj_1913.LUT_INIT = 16'ha080;
    SB_LUT4 i35485_4_lut (.I0(n44905), .I1(n1323_adj_5393), .I2(n1324_adj_5394), 
            .I3(n46793), .O(n1356));
    defparam i35485_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_31__I_0_i775_3_lut (.I0(n1132), .I1(n1199), 
            .I2(n1158), .I3(GND_net), .O(n1231));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i775_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i774_3_lut (.I0(n1131), .I1(n1198), 
            .I2(n1158), .I3(GND_net), .O(n1230));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i774_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i773_3_lut (.I0(n1130), .I1(n1197), 
            .I2(n1158), .I3(GND_net), .O(n1229));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i773_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i772_3_lut (.I0(n1129), .I1(n1196), 
            .I2(n1158), .I3(GND_net), .O(n1228));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i772_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i771_3_lut (.I0(n1128), .I1(n1195), 
            .I2(n1158), .I3(GND_net), .O(n1227));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i771_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i770_3_lut (.I0(n1127), .I1(n1194), 
            .I2(n1158), .I3(GND_net), .O(n1226));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i770_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i769_3_lut (.I0(n1126), .I1(n1193), 
            .I2(n1158), .I3(GND_net), .O(n1225));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i769_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i777_3_lut (.I0(n522), .I1(n1201), 
            .I2(n1158), .I3(GND_net), .O(n1233));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i777_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_1005_i21_3_lut (.I0(duty[20]), .I1(n343), .I2(duty[23]), 
            .I3(GND_net), .O(n4703));   // verilog/TinyFPGA_B.v(118[13] 129[7])
    defparam mux_1005_i21_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1005_i22_3_lut (.I0(duty[21]), .I1(n342), .I2(duty[23]), 
            .I3(GND_net), .O(n4702));   // verilog/TinyFPGA_B.v(118[13] 129[7])
    defparam mux_1005_i22_3_lut.LUT_INIT = 16'hcaca;
    EEPROM eeprom (.GND_net(GND_net), .CLK_c(CLK_c), .n6129({n6130}), 
           .\state[1] (state_adj_5510[1]), .\state[0] (state_adj_5510[0]), 
           .n43386(n43386), .read(read), .\state[2] (state_adj_5537[2]), 
           .n7(n7_adj_5404), .n29054(n29054), .rw(rw), .n43506(n43506), 
           .data_ready(data_ready), .enable_slow_N_4354(enable_slow_N_4354), 
           .n43380(n43380), .n34717(n34717), .n44748(n44748), .n44835(n44835), 
           .\state[3] (state_adj_5537[3]), .n6(n6_adj_5274), .n29159(n29159), 
           .data({data}), .\state_7__N_4251[0] (state_7__N_4251[0]), .n7210(n7210), 
           .sda_enable(sda_enable), .n29146(n29146), .\saved_addr[0] (saved_addr[0]), 
           .scl_enable(scl_enable), .\state_7__N_4267[3] (state_7__N_4267[3]), 
           .\state[0]_adj_2 (state_adj_5537[0]), .n4(n4_adj_5346), .n4_adj_3(n4_adj_5248), 
           .n27152(n27152), .n34660(n34660), .scl(scl), .n10(n10_adj_5410), 
           .n29033(n29033), .n29032(n29032), .n29031(n29031), .n29030(n29030), 
           .n29029(n29029), .n29028(n29028), .n29027(n29027), .n7754(n7754), 
           .sda_out(sda_out), .VCC_net(VCC_net), .n27147(n27147), .n8(n8), 
           .n49357(n49357), .n34664(n34664)) /* synthesis syn_noprune=1, syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(405[10] 416[6])
    SB_LUT4 encoder0_position_31__I_0_i776_3_lut (.I0(n1133), .I1(n1200), 
            .I2(n1158), .I3(GND_net), .O(n1232));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_i776_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i22_3_lut (.I0(encoder0_position[21]), 
            .I1(n12_adj_5303), .I2(encoder0_position[31]), .I3(GND_net), 
            .O(n937));   // verilog/TinyFPGA_B.v(338[33:53])
    defparam encoder0_position_31__I_0_mux_3_i22_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15391_3_lut (.I0(\data_in_frame[13] [0]), .I1(rx_data[0]), 
            .I2(n43847), .I3(GND_net), .O(n29339));   // verilog/coms.v(128[12] 303[6])
    defparam i15391_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i21480_3_lut (.I0(n937), .I1(n1232), .I2(n1233), .I3(GND_net), 
            .O(n35428));
    defparam i21480_3_lut.LUT_INIT = 16'hc8c8;
    pwm PWM (.pwm_out(pwm_out), .clk32MHz(clk32MHz), .GND_net(GND_net), 
        .pwm_setpoint({pwm_setpoint}), .VCC_net(VCC_net)) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(89[6] 94[3])
    
endmodule
//
// Verilog Description of module \neopixel(CLOCK_SPEED_HZ=16000000) 
//

module \neopixel(CLOCK_SPEED_HZ=16000000)  (GND_net, timer, CLK_c, \neo_pixel_transmitter.t0 , 
            neopxl_color, VCC_net, \state[1] , n42404, \state_3__N_552[1] , 
            LED_c, n29069, n28592, n44637, n29022, n29498, n29497, 
            n29496, n29495, n29494, n29493, n29492, n29491, n29490, 
            n29489, n29488, n29487, n29486, n29485, n29484, n29483, 
            n29482, n29481, n29480, n29479, n29478, n29477, n29476, 
            n29475, n29474, n29473, n29472, n29471, n29470, n29469, 
            n29468, NEOPXL_c) /* synthesis syn_module_defined=1 */ ;
    input GND_net;
    output [31:0]timer;
    input CLK_c;
    output [31:0]\neo_pixel_transmitter.t0 ;
    input [23:0]neopxl_color;
    input VCC_net;
    output \state[1] ;
    output n42404;
    output \state_3__N_552[1] ;
    input LED_c;
    input n29069;
    output n28592;
    output n44637;
    input n29022;
    input n29498;
    input n29497;
    input n29496;
    input n29495;
    input n29494;
    input n29493;
    input n29492;
    input n29491;
    input n29490;
    input n29489;
    input n29488;
    input n29487;
    input n29486;
    input n29485;
    input n29484;
    input n29483;
    input n29482;
    input n29481;
    input n29480;
    input n29479;
    input n29478;
    input n29477;
    input n29476;
    input n29475;
    input n29474;
    input n29473;
    input n29472;
    input n29471;
    input n29470;
    input n29469;
    input n29468;
    output NEOPXL_c;
    
    wire CLK_c /* synthesis SET_AS_NETWORK=CLK_c, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(3[9:12])
    
    wire n39323, n39324;
    wire [31:0]n133;
    
    wire n39322, n39321, \neo_pixel_transmitter.done_N_760 , n51587, 
        \neo_pixel_transmitter.done , n39320, start_N_751, n7, start;
    wire [31:0]n1;
    
    wire n39319;
    wire [31:0]n282;
    wire [31:0]bit_ctr;   // verilog/neopixel.v(18[12:19])
    
    wire n38523, n38524, n38522, n39318, n39317, n39316, n39315, 
        n48167, n48168, n48057, n39314, n48056, n28484, n28887, 
        n40044, n44736;
    wire [3:0]state;   // verilog/neopixel.v(16[20:25])
    
    wire n49717, n49277, n35348, n27032, n44845, n49718, n44865, 
        \neo_pixel_transmitter.done_N_766 , n38521, n38520, n38519, 
        n39326, n39327, n38518, n38517, n38516, n38515, n27184, 
        n38706, n47713, n38705, n47711, n38704, n47709, n38514, 
        n44791, n7_adj_5236, n27160, n35336, n30_adj_5237, n48, 
        n46, n47, n45, n44, n43, n54, n38513, n38703, n47707, 
        n38512, n38702, n47705, n51327, n51561;
    wire [31:0]color_bit_N_746;
    
    wire n50148, n35253, n40743, n38511, n38701, n47703, n38700, 
        n47701, n51285, n50230, n51219, n49348, n38699, n47699;
    wire [3:0]state_3__N_552;
    
    wire n39325, n38510, n38698, n47697, n38697, n47695, n38509, 
        n38696, n47693, n49, n38695, n47691, n38508, n38694, n47689, 
        n38507, n38506, n2208, n35127, n7565, n49346;
    wire [31:0]one_wire_N_703;
    
    wire n38693, n47687, n38505, n38692, n47685, n38691, n47683, 
        n4_adj_5239, n47663, n47669, n49283, n44801, n43815, n44732, 
        n103, n16_adj_5240, n6_adj_5241, n48173, n48174, n51282, 
        n48099, n48098, n51558, n38690, n47681, n38689, n47679, 
        n38504, n38688, n47677, n38503, n2222, n44630, n49279, 
        n38687, n38686, n38502, n38685, n38501, n38684, n38683, 
        n38500, n38682, n38681, n51324, n38680, n38679, n38678, 
        n38677, n38676, n39344, n39343, n39342, n39341, n39340, 
        n39339, n39338, n39337, n39336, n39335, n39334, n39333, 
        n39332, n39331, n39330, n39329, n38530, n38529, n39328, 
        n38528, n38527, n38526, n46519, n38525, n51216;
    
    SB_CARRY timer_2245_add_4_12 (.CI(n39323), .I0(GND_net), .I1(timer[10]), 
            .CO(n39324));
    SB_LUT4 timer_2245_add_4_11_lut (.I0(GND_net), .I1(GND_net), .I2(timer[9]), 
            .I3(n39322), .O(n133[9])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2245_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2245_add_4_11 (.CI(n39322), .I0(GND_net), .I1(timer[9]), 
            .CO(n39323));
    SB_LUT4 timer_2245_add_4_10_lut (.I0(GND_net), .I1(GND_net), .I2(timer[8]), 
            .I3(n39321), .O(n133[8])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2245_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2245_add_4_10 (.CI(n39321), .I0(GND_net), .I1(timer[8]), 
            .CO(n39322));
    SB_DFFE \neo_pixel_transmitter.done_104  (.Q(\neo_pixel_transmitter.done ), 
            .C(CLK_c), .E(n51587), .D(\neo_pixel_transmitter.done_N_760 ));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 timer_2245_add_4_9_lut (.I0(GND_net), .I1(GND_net), .I2(timer[7]), 
            .I3(n39320), .O(n133[7])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2245_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_DFFE start_103 (.Q(start), .C(CLK_c), .E(n7), .D(start_N_751));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 sub_14_inv_0_i1_1_lut (.I0(\neo_pixel_transmitter.t0 [0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[0]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i2_1_lut (.I0(\neo_pixel_transmitter.t0 [1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[1]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY timer_2245_add_4_9 (.CI(n39320), .I0(GND_net), .I1(timer[7]), 
            .CO(n39321));
    SB_LUT4 timer_2245_add_4_8_lut (.I0(GND_net), .I1(GND_net), .I2(timer[6]), 
            .I3(n39319), .O(n133[6])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2245_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_21_26_lut (.I0(GND_net), .I1(bit_ctr[24]), .I2(GND_net), 
            .I3(n38523), .O(n282[24])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2245_add_4_8 (.CI(n39319), .I0(GND_net), .I1(timer[6]), 
            .CO(n39320));
    SB_LUT4 sub_14_inv_0_i3_1_lut (.I0(\neo_pixel_transmitter.t0 [2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[2]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i4_1_lut (.I0(\neo_pixel_transmitter.t0 [3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[3]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_21_26 (.CI(n38523), .I0(bit_ctr[24]), .I1(GND_net), .CO(n38524));
    SB_LUT4 add_21_25_lut (.I0(GND_net), .I1(bit_ctr[23]), .I2(GND_net), 
            .I3(n38522), .O(n282[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 timer_2245_add_4_7_lut (.I0(GND_net), .I1(GND_net), .I2(timer[5]), 
            .I3(n39318), .O(n133[5])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2245_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2245_add_4_7 (.CI(n39318), .I0(GND_net), .I1(timer[5]), 
            .CO(n39319));
    SB_LUT4 sub_14_inv_0_i5_1_lut (.I0(\neo_pixel_transmitter.t0 [4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[4]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i6_1_lut (.I0(\neo_pixel_transmitter.t0 [5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[5]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i7_1_lut (.I0(\neo_pixel_transmitter.t0 [6]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[6]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 timer_2245_add_4_6_lut (.I0(GND_net), .I1(GND_net), .I2(timer[4]), 
            .I3(n39317), .O(n133[4])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2245_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2245_add_4_6 (.CI(n39317), .I0(GND_net), .I1(timer[4]), 
            .CO(n39318));
    SB_LUT4 timer_2245_add_4_5_lut (.I0(GND_net), .I1(GND_net), .I2(timer[3]), 
            .I3(n39316), .O(n133[3])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2245_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2245_add_4_5 (.CI(n39316), .I0(GND_net), .I1(timer[3]), 
            .CO(n39317));
    SB_LUT4 timer_2245_add_4_4_lut (.I0(GND_net), .I1(GND_net), .I2(timer[2]), 
            .I3(n39315), .O(n133[2])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2245_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i32580_3_lut (.I0(neopxl_color[16]), .I1(neopxl_color[17]), 
            .I2(bit_ctr[0]), .I3(GND_net), .O(n48167));
    defparam i32580_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY timer_2245_add_4_4 (.CI(n39315), .I0(GND_net), .I1(timer[2]), 
            .CO(n39316));
    SB_LUT4 i32581_3_lut (.I0(neopxl_color[18]), .I1(neopxl_color[19]), 
            .I2(bit_ctr[0]), .I3(GND_net), .O(n48168));
    defparam i32581_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i32470_3_lut (.I0(neopxl_color[22]), .I1(neopxl_color[23]), 
            .I2(bit_ctr[0]), .I3(GND_net), .O(n48057));
    defparam i32470_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 timer_2245_add_4_3_lut (.I0(GND_net), .I1(GND_net), .I2(timer[1]), 
            .I3(n39314), .O(n133[1])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2245_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2245_add_4_3 (.CI(n39314), .I0(GND_net), .I1(timer[1]), 
            .CO(n39315));
    SB_LUT4 i32469_3_lut (.I0(neopxl_color[20]), .I1(neopxl_color[21]), 
            .I2(bit_ctr[0]), .I3(GND_net), .O(n48056));
    defparam i32469_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 sub_14_inv_0_i8_1_lut (.I0(\neo_pixel_transmitter.t0 [7]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[7]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i9_1_lut (.I0(\neo_pixel_transmitter.t0 [8]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[8]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_DFFESR bit_ctr_i0_i1 (.Q(bit_ctr[1]), .C(CLK_c), .E(n28484), .D(n282[1]), 
            .R(n28887));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i2 (.Q(bit_ctr[2]), .C(CLK_c), .E(n28484), .D(n282[2]), 
            .R(n28887));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i3 (.Q(bit_ctr[3]), .C(CLK_c), .E(n28484), .D(n282[3]), 
            .R(n28887));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i4 (.Q(bit_ctr[4]), .C(CLK_c), .E(n28484), .D(n282[4]), 
            .R(n28887));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i5 (.Q(bit_ctr[5]), .C(CLK_c), .E(n28484), .D(n282[5]), 
            .R(n28887));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i6 (.Q(bit_ctr[6]), .C(CLK_c), .E(n28484), .D(n282[6]), 
            .R(n28887));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i7 (.Q(bit_ctr[7]), .C(CLK_c), .E(n28484), .D(n282[7]), 
            .R(n28887));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i8 (.Q(bit_ctr[8]), .C(CLK_c), .E(n28484), .D(n282[8]), 
            .R(n28887));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i9 (.Q(bit_ctr[9]), .C(CLK_c), .E(n28484), .D(n282[9]), 
            .R(n28887));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i10 (.Q(bit_ctr[10]), .C(CLK_c), .E(n28484), 
            .D(n282[10]), .R(n28887));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i11 (.Q(bit_ctr[11]), .C(CLK_c), .E(n28484), 
            .D(n282[11]), .R(n28887));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i12 (.Q(bit_ctr[12]), .C(CLK_c), .E(n28484), 
            .D(n282[12]), .R(n28887));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i13 (.Q(bit_ctr[13]), .C(CLK_c), .E(n28484), 
            .D(n282[13]), .R(n28887));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i14 (.Q(bit_ctr[14]), .C(CLK_c), .E(n28484), 
            .D(n282[14]), .R(n28887));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i15 (.Q(bit_ctr[15]), .C(CLK_c), .E(n28484), 
            .D(n282[15]), .R(n28887));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i16 (.Q(bit_ctr[16]), .C(CLK_c), .E(n28484), 
            .D(n282[16]), .R(n28887));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i17 (.Q(bit_ctr[17]), .C(CLK_c), .E(n28484), 
            .D(n282[17]), .R(n28887));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i18 (.Q(bit_ctr[18]), .C(CLK_c), .E(n28484), 
            .D(n282[18]), .R(n28887));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i19 (.Q(bit_ctr[19]), .C(CLK_c), .E(n28484), 
            .D(n282[19]), .R(n28887));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 sub_14_inv_0_i10_1_lut (.I0(\neo_pixel_transmitter.t0 [9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[9]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_DFFESR bit_ctr_i0_i20 (.Q(bit_ctr[20]), .C(CLK_c), .E(n28484), 
            .D(n282[20]), .R(n28887));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i21 (.Q(bit_ctr[21]), .C(CLK_c), .E(n28484), 
            .D(n282[21]), .R(n28887));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 sub_14_inv_0_i11_1_lut (.I0(\neo_pixel_transmitter.t0 [10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[10]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_DFFESR bit_ctr_i0_i22 (.Q(bit_ctr[22]), .C(CLK_c), .E(n28484), 
            .D(n282[22]), .R(n28887));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i23 (.Q(bit_ctr[23]), .C(CLK_c), .E(n28484), 
            .D(n282[23]), .R(n28887));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i24 (.Q(bit_ctr[24]), .C(CLK_c), .E(n28484), 
            .D(n282[24]), .R(n28887));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i25 (.Q(bit_ctr[25]), .C(CLK_c), .E(n28484), 
            .D(n282[25]), .R(n28887));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i26 (.Q(bit_ctr[26]), .C(CLK_c), .E(n28484), 
            .D(n282[26]), .R(n28887));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i27 (.Q(bit_ctr[27]), .C(CLK_c), .E(n28484), 
            .D(n282[27]), .R(n28887));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i28 (.Q(bit_ctr[28]), .C(CLK_c), .E(n28484), 
            .D(n282[28]), .R(n28887));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i29 (.Q(bit_ctr[29]), .C(CLK_c), .E(n28484), 
            .D(n282[29]), .R(n28887));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i30 (.Q(bit_ctr[30]), .C(CLK_c), .E(n28484), 
            .D(n282[30]), .R(n28887));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i31 (.Q(bit_ctr[31]), .C(CLK_c), .E(n28484), 
            .D(n282[31]), .R(n28887));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 timer_2245_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(timer[0]), 
            .I3(VCC_net), .O(n133[0])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2245_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2245_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(timer[0]), 
            .CO(n39314));
    SB_LUT4 sub_14_inv_0_i12_1_lut (.I0(\neo_pixel_transmitter.t0 [11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[11]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i13_1_lut (.I0(\neo_pixel_transmitter.t0 [12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[12]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i30_1_lut (.I0(\neo_pixel_transmitter.t0 [29]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[29]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i30_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i31_1_lut (.I0(\neo_pixel_transmitter.t0 [30]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[30]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i31_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i32_1_lut (.I0(\neo_pixel_transmitter.t0 [31]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[31]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i32_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i34429_4_lut (.I0(n40044), .I1(n44736), .I2(\neo_pixel_transmitter.done ), 
            .I3(state[0]), .O(n49717));
    defparam i34429_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i53_4_lut (.I0(n49277), .I1(n35348), .I2(\state[1] ), .I3(n27032), 
            .O(n44845));
    defparam i53_4_lut.LUT_INIT = 16'hcfca;
    SB_LUT4 i52_4_lut (.I0(n44845), .I1(n49718), .I2(state[0]), .I3(\neo_pixel_transmitter.done ), 
            .O(n44865));
    defparam i52_4_lut.LUT_INIT = 16'h3335;
    SB_LUT4 i3_1_lut (.I0(\neo_pixel_transmitter.done ), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(\neo_pixel_transmitter.done_N_766 ));   // verilog/neopixel.v(35[12] 117[6])
    defparam i3_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_21_25 (.CI(n38522), .I0(bit_ctr[23]), .I1(GND_net), .CO(n38523));
    SB_LUT4 sub_14_inv_0_i14_1_lut (.I0(\neo_pixel_transmitter.t0 [13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[13]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_21_24_lut (.I0(GND_net), .I1(bit_ctr[22]), .I2(GND_net), 
            .I3(n38521), .O(n282[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_21_24 (.CI(n38521), .I0(bit_ctr[22]), .I1(GND_net), .CO(n38522));
    SB_LUT4 add_21_23_lut (.I0(GND_net), .I1(bit_ctr[21]), .I2(GND_net), 
            .I3(n38520), .O(n282[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_21_23 (.CI(n38520), .I0(bit_ctr[21]), .I1(GND_net), .CO(n38521));
    SB_LUT4 add_21_22_lut (.I0(GND_net), .I1(bit_ctr[20]), .I2(GND_net), 
            .I3(n38519), .O(n282[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_14_inv_0_i15_1_lut (.I0(\neo_pixel_transmitter.t0 [14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[14]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_21_22 (.CI(n38519), .I0(bit_ctr[20]), .I1(GND_net), .CO(n38520));
    SB_CARRY timer_2245_add_4_15 (.CI(n39326), .I0(GND_net), .I1(timer[13]), 
            .CO(n39327));
    SB_LUT4 add_21_21_lut (.I0(GND_net), .I1(bit_ctr[19]), .I2(GND_net), 
            .I3(n38518), .O(n282[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_21_21 (.CI(n38518), .I0(bit_ctr[19]), .I1(GND_net), .CO(n38519));
    SB_LUT4 add_21_20_lut (.I0(GND_net), .I1(bit_ctr[18]), .I2(GND_net), 
            .I3(n38517), .O(n282[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_21_20 (.CI(n38517), .I0(bit_ctr[18]), .I1(GND_net), .CO(n38518));
    SB_LUT4 add_21_19_lut (.I0(GND_net), .I1(bit_ctr[17]), .I2(GND_net), 
            .I3(n38516), .O(n282[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_21_19 (.CI(n38516), .I0(bit_ctr[17]), .I1(GND_net), .CO(n38517));
    SB_LUT4 add_21_18_lut (.I0(GND_net), .I1(bit_ctr[16]), .I2(GND_net), 
            .I3(n38515), .O(n282[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_14_add_2_33_lut (.I0(n47713), .I1(timer[31]), .I2(n1[31]), 
            .I3(n38706), .O(n27184)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_33_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 sub_14_add_2_32_lut (.I0(n47711), .I1(timer[30]), .I2(n1[30]), 
            .I3(n38705), .O(n47713)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_32_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_14_add_2_32 (.CI(n38705), .I0(timer[30]), .I1(n1[30]), 
            .CO(n38706));
    SB_LUT4 sub_14_add_2_31_lut (.I0(n47709), .I1(timer[29]), .I2(n1[29]), 
            .I3(n38704), .O(n47711)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_31_lut.LUT_INIT = 16'hebbe;
    SB_CARRY add_21_18 (.CI(n38515), .I0(bit_ctr[16]), .I1(GND_net), .CO(n38516));
    SB_DFF timer_2245__i31 (.Q(timer[31]), .C(CLK_c), .D(n133[31]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2245__i30 (.Q(timer[30]), .C(CLK_c), .D(n133[30]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2245__i29 (.Q(timer[29]), .C(CLK_c), .D(n133[29]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2245__i28 (.Q(timer[28]), .C(CLK_c), .D(n133[28]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2245__i27 (.Q(timer[27]), .C(CLK_c), .D(n133[27]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2245__i26 (.Q(timer[26]), .C(CLK_c), .D(n133[26]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2245__i25 (.Q(timer[25]), .C(CLK_c), .D(n133[25]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2245__i24 (.Q(timer[24]), .C(CLK_c), .D(n133[24]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2245__i23 (.Q(timer[23]), .C(CLK_c), .D(n133[23]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2245__i22 (.Q(timer[22]), .C(CLK_c), .D(n133[22]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2245__i21 (.Q(timer[21]), .C(CLK_c), .D(n133[21]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2245__i20 (.Q(timer[20]), .C(CLK_c), .D(n133[20]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2245__i19 (.Q(timer[19]), .C(CLK_c), .D(n133[19]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2245__i18 (.Q(timer[18]), .C(CLK_c), .D(n133[18]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2245__i17 (.Q(timer[17]), .C(CLK_c), .D(n133[17]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2245__i16 (.Q(timer[16]), .C(CLK_c), .D(n133[16]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2245__i15 (.Q(timer[15]), .C(CLK_c), .D(n133[15]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2245__i14 (.Q(timer[14]), .C(CLK_c), .D(n133[14]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2245__i13 (.Q(timer[13]), .C(CLK_c), .D(n133[13]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2245__i12 (.Q(timer[12]), .C(CLK_c), .D(n133[12]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2245__i11 (.Q(timer[11]), .C(CLK_c), .D(n133[11]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2245__i10 (.Q(timer[10]), .C(CLK_c), .D(n133[10]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2245__i9 (.Q(timer[9]), .C(CLK_c), .D(n133[9]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2245__i8 (.Q(timer[8]), .C(CLK_c), .D(n133[8]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2245__i7 (.Q(timer[7]), .C(CLK_c), .D(n133[7]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2245__i6 (.Q(timer[6]), .C(CLK_c), .D(n133[6]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2245__i5 (.Q(timer[5]), .C(CLK_c), .D(n133[5]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2245__i4 (.Q(timer[4]), .C(CLK_c), .D(n133[4]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2245__i3 (.Q(timer[3]), .C(CLK_c), .D(n133[3]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2245__i2 (.Q(timer[2]), .C(CLK_c), .D(n133[2]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2245__i1 (.Q(timer[1]), .C(CLK_c), .D(n133[1]));   // verilog/neopixel.v(12[12:21])
    SB_LUT4 add_21_17_lut (.I0(GND_net), .I1(bit_ctr[15]), .I2(GND_net), 
            .I3(n38514), .O(n282[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i29273_4_lut (.I0(n27032), .I1(n44736), .I2(n40044), .I3(state[0]), 
            .O(n44791));
    defparam i29273_4_lut.LUT_INIT = 16'hfaee;
    SB_LUT4 i20_4_lut (.I0(\neo_pixel_transmitter.done ), .I1(\state[1] ), 
            .I2(start), .I3(n44791), .O(n7_adj_5236));
    defparam i20_4_lut.LUT_INIT = 16'hcecf;
    SB_LUT4 i1_4_lut (.I0(n27160), .I1(n7_adj_5236), .I2(n35336), .I3(\state[1] ), 
            .O(n42404));
    defparam i1_4_lut.LUT_INIT = 16'hcc8c;
    SB_LUT4 sub_14_inv_0_i16_1_lut (.I0(\neo_pixel_transmitter.t0 [15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[15]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i2_2_lut (.I0(bit_ctr[22]), .I1(bit_ctr[17]), .I2(GND_net), 
            .I3(GND_net), .O(n30_adj_5237));
    defparam i2_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i20_4_lut_adj_1730 (.I0(bit_ctr[20]), .I1(bit_ctr[7]), .I2(bit_ctr[16]), 
            .I3(bit_ctr[30]), .O(n48));
    defparam i20_4_lut_adj_1730.LUT_INIT = 16'hfffe;
    SB_LUT4 i18_4_lut (.I0(bit_ctr[25]), .I1(bit_ctr[10]), .I2(bit_ctr[9]), 
            .I3(bit_ctr[27]), .O(n46));
    defparam i18_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i19_4_lut (.I0(bit_ctr[15]), .I1(bit_ctr[29]), .I2(bit_ctr[12]), 
            .I3(bit_ctr[23]), .O(n47));
    defparam i19_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_4_lut (.I0(bit_ctr[19]), .I1(bit_ctr[21]), .I2(bit_ctr[31]), 
            .I3(bit_ctr[14]), .O(n45));
    defparam i17_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut (.I0(bit_ctr[11]), .I1(bit_ctr[5]), .I2(bit_ctr[28]), 
            .I3(bit_ctr[6]), .O(n44));
    defparam i16_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut (.I0(bit_ctr[3]), .I1(n30_adj_5237), .I2(bit_ctr[13]), 
            .I3(bit_ctr[4]), .O(n43));
    defparam i15_4_lut.LUT_INIT = 16'hfefc;
    SB_LUT4 i26_4_lut (.I0(n45), .I1(n47), .I2(n46), .I3(n48), .O(n54));
    defparam i26_4_lut.LUT_INIT = 16'hfffe;
    SB_CARRY add_21_17 (.CI(n38514), .I0(bit_ctr[15]), .I1(GND_net), .CO(n38515));
    SB_LUT4 add_21_16_lut (.I0(GND_net), .I1(bit_ctr[14]), .I2(GND_net), 
            .I3(n38513), .O(n282[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_31 (.CI(n38704), .I0(timer[29]), .I1(n1[29]), 
            .CO(n38705));
    SB_LUT4 sub_14_add_2_30_lut (.I0(n47707), .I1(timer[28]), .I2(n1[28]), 
            .I3(n38703), .O(n47709)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_30_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_14_add_2_30 (.CI(n38703), .I0(timer[28]), .I1(n1[28]), 
            .CO(n38704));
    SB_CARRY add_21_16 (.CI(n38513), .I0(bit_ctr[14]), .I1(GND_net), .CO(n38514));
    SB_LUT4 add_21_15_lut (.I0(GND_net), .I1(bit_ctr[13]), .I2(GND_net), 
            .I3(n38512), .O(n282[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_21_15 (.CI(n38512), .I0(bit_ctr[13]), .I1(GND_net), .CO(n38513));
    SB_LUT4 sub_14_add_2_29_lut (.I0(n47705), .I1(timer[27]), .I2(n1[27]), 
            .I3(n38702), .O(n47707)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_29_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 i34560_3_lut (.I0(n51327), .I1(n51561), .I2(color_bit_N_746[2]), 
            .I3(GND_net), .O(n50148));
    defparam i34560_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_3_lut (.I0(bit_ctr[4]), .I1(bit_ctr[3]), .I2(n35253), .I3(GND_net), 
            .O(n40743));
    defparam i1_3_lut.LUT_INIT = 16'h6a6a;
    SB_CARRY sub_14_add_2_29 (.CI(n38702), .I0(timer[27]), .I1(n1[27]), 
            .CO(n38703));
    SB_LUT4 add_21_14_lut (.I0(GND_net), .I1(bit_ctr[12]), .I2(GND_net), 
            .I3(n38511), .O(n282[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_21_14 (.CI(n38511), .I0(bit_ctr[12]), .I1(GND_net), .CO(n38512));
    SB_LUT4 sub_14_add_2_28_lut (.I0(n47703), .I1(timer[26]), .I2(n1[26]), 
            .I3(n38701), .O(n47705)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_28_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_14_add_2_28 (.CI(n38701), .I0(timer[26]), .I1(n1[26]), 
            .CO(n38702));
    SB_LUT4 sub_14_add_2_27_lut (.I0(n47701), .I1(timer[25]), .I2(n1[25]), 
            .I3(n38700), .O(n47703)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_27_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_14_add_2_27 (.CI(n38700), .I0(timer[25]), .I1(n1[25]), 
            .CO(n38701));
    SB_LUT4 i34642_4_lut (.I0(n50148), .I1(n51285), .I2(bit_ctr[3]), .I3(n35253), 
            .O(n50230));   // verilog/neopixel.v(22[26:38])
    defparam i34642_4_lut.LUT_INIT = 16'hacca;
    SB_LUT4 i33823_3_lut (.I0(n51219), .I1(bit_ctr[3]), .I2(n35253), .I3(GND_net), 
            .O(n49348));
    defparam i33823_3_lut.LUT_INIT = 16'h2828;
    SB_LUT4 sub_14_add_2_26_lut (.I0(n47699), .I1(timer[24]), .I2(n1[24]), 
            .I3(n38699), .O(n47701)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_26_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 i20622_4_lut (.I0(n49348), .I1(\state_3__N_552[1] ), .I2(n50230), 
            .I3(n40743), .O(state_3__N_552[0]));   // verilog/neopixel.v(40[18] 45[12])
    defparam i20622_4_lut.LUT_INIT = 16'h3022;
    SB_CARRY timer_2245_add_4_14 (.CI(n39325), .I0(GND_net), .I1(timer[12]), 
            .CO(n39326));
    SB_CARRY sub_14_add_2_26 (.CI(n38699), .I0(timer[24]), .I1(n1[24]), 
            .CO(n38700));
    SB_LUT4 add_21_13_lut (.I0(GND_net), .I1(bit_ctr[11]), .I2(GND_net), 
            .I3(n38510), .O(n282[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 timer_2245_add_4_13_lut (.I0(GND_net), .I1(GND_net), .I2(timer[11]), 
            .I3(n39324), .O(n133[11])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2245_add_4_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_21_13 (.CI(n38510), .I0(bit_ctr[11]), .I1(GND_net), .CO(n38511));
    SB_LUT4 sub_14_add_2_25_lut (.I0(n47697), .I1(timer[23]), .I2(n1[23]), 
            .I3(n38698), .O(n47699)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_25_lut.LUT_INIT = 16'hebbe;
    SB_CARRY timer_2245_add_4_13 (.CI(n39324), .I0(GND_net), .I1(timer[11]), 
            .CO(n39325));
    SB_CARRY sub_14_add_2_25 (.CI(n38698), .I0(timer[23]), .I1(n1[23]), 
            .CO(n38699));
    SB_LUT4 sub_14_add_2_24_lut (.I0(n47695), .I1(timer[22]), .I2(n1[22]), 
            .I3(n38697), .O(n47697)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_24_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_14_add_2_24 (.CI(n38697), .I0(timer[22]), .I1(n1[22]), 
            .CO(n38698));
    SB_LUT4 add_21_12_lut (.I0(GND_net), .I1(bit_ctr[10]), .I2(GND_net), 
            .I3(n38509), .O(n282[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_14_add_2_23_lut (.I0(n47693), .I1(timer[21]), .I2(n1[21]), 
            .I3(n38696), .O(n47695)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_23_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 i21_4_lut (.I0(bit_ctr[24]), .I1(bit_ctr[8]), .I2(bit_ctr[18]), 
            .I3(bit_ctr[26]), .O(n49));
    defparam i21_4_lut.LUT_INIT = 16'hfffe;
    SB_CARRY add_21_12 (.CI(n38509), .I0(bit_ctr[10]), .I1(GND_net), .CO(n38510));
    SB_CARRY sub_14_add_2_23 (.CI(n38696), .I0(timer[21]), .I1(n1[21]), 
            .CO(n38697));
    SB_LUT4 sub_14_add_2_22_lut (.I0(n47691), .I1(timer[20]), .I2(n1[20]), 
            .I3(n38695), .O(n47693)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_22_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_14_add_2_22 (.CI(n38695), .I0(timer[20]), .I1(n1[20]), 
            .CO(n38696));
    SB_LUT4 add_21_11_lut (.I0(GND_net), .I1(bit_ctr[9]), .I2(GND_net), 
            .I3(n38508), .O(n282[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_14_add_2_21_lut (.I0(n47689), .I1(timer[19]), .I2(n1[19]), 
            .I3(n38694), .O(n47691)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_21_lut.LUT_INIT = 16'hebbe;
    SB_CARRY add_21_11 (.CI(n38508), .I0(bit_ctr[9]), .I1(GND_net), .CO(n38509));
    SB_LUT4 i27_4_lut (.I0(n49), .I1(n54), .I2(n43), .I3(n44), .O(\state_3__N_552[1] ));
    defparam i27_4_lut.LUT_INIT = 16'hfffe;
    SB_CARRY sub_14_add_2_21 (.CI(n38694), .I0(timer[19]), .I1(n1[19]), 
            .CO(n38695));
    SB_LUT4 i1_2_lut (.I0(start), .I1(\neo_pixel_transmitter.done ), .I2(GND_net), 
            .I3(GND_net), .O(n27160));   // verilog/neopixel.v(52[18] 72[12])
    defparam i1_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 add_21_10_lut (.I0(GND_net), .I1(bit_ctr[8]), .I2(GND_net), 
            .I3(n38507), .O(n282[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_21_10 (.CI(n38507), .I0(bit_ctr[8]), .I1(GND_net), .CO(n38508));
    SB_LUT4 add_21_9_lut (.I0(GND_net), .I1(bit_ctr[7]), .I2(GND_net), 
            .I3(n38506), .O(n282[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i513_2_lut (.I0(LED_c), .I1(\state_3__N_552[1] ), .I2(GND_net), 
            .I3(GND_net), .O(n2208));   // verilog/neopixel.v(40[18] 45[12])
    defparam i513_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i4631_4_lut (.I0(n35127), .I1(n2208), .I2(\state[1] ), .I3(n27160), 
            .O(n7565));
    defparam i4631_4_lut.LUT_INIT = 16'h3f35;
    SB_LUT4 i33816_3_lut (.I0(n40044), .I1(n27160), .I2(n27032), .I3(GND_net), 
            .O(n49346));
    defparam i33816_3_lut.LUT_INIT = 16'hcdcd;
    SB_LUT4 i34918_4_lut (.I0(\state[1] ), .I1(n49346), .I2(n7565), .I3(state[0]), 
            .O(n28484));
    defparam i34918_4_lut.LUT_INIT = 16'h0f11;
    SB_LUT4 i21402_4_lut (.I0(one_wire_N_703[8]), .I1(n27184), .I2(one_wire_N_703[10]), 
            .I3(one_wire_N_703[9]), .O(n35348));
    defparam i21402_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 sub_14_add_2_20_lut (.I0(n47687), .I1(timer[18]), .I2(n1[18]), 
            .I3(n38693), .O(n47689)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_20_lut.LUT_INIT = 16'hebbe;
    SB_CARRY add_21_9 (.CI(n38506), .I0(bit_ctr[7]), .I1(GND_net), .CO(n38507));
    SB_LUT4 add_21_8_lut (.I0(GND_net), .I1(bit_ctr[6]), .I2(GND_net), 
            .I3(n38505), .O(n282[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_20 (.CI(n38693), .I0(timer[18]), .I1(n1[18]), 
            .CO(n38694));
    SB_LUT4 sub_14_add_2_19_lut (.I0(n47685), .I1(timer[17]), .I2(n1[17]), 
            .I3(n38692), .O(n47687)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_19_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_14_add_2_19 (.CI(n38692), .I0(timer[17]), .I1(n1[17]), 
            .CO(n38693));
    SB_LUT4 sub_14_add_2_18_lut (.I0(n47683), .I1(timer[16]), .I2(n1[16]), 
            .I3(n38691), .O(n47685)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_18_lut.LUT_INIT = 16'hebbe;
    SB_DFF timer_2245__i0 (.Q(timer[0]), .C(CLK_c), .D(n133[0]));   // verilog/neopixel.v(12[12:21])
    SB_DFFE state_i1 (.Q(\state[1] ), .C(CLK_c), .E(VCC_net), .D(n29069));   // verilog/neopixel.v(35[12] 117[6])
    SB_CARRY sub_14_add_2_18 (.CI(n38691), .I0(timer[16]), .I1(n1[16]), 
            .CO(n38692));
    SB_LUT4 i29220_2_lut (.I0(one_wire_N_703[3]), .I1(one_wire_N_703[2]), 
            .I2(GND_net), .I3(GND_net), .O(n44736));
    defparam i29220_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i2_2_lut_adj_1731 (.I0(one_wire_N_703[2]), .I1(n4_adj_5239), 
            .I2(GND_net), .I3(GND_net), .O(n40044));
    defparam i2_2_lut_adj_1731.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1732 (.I0(one_wire_N_703[5]), .I1(one_wire_N_703[4]), 
            .I2(GND_net), .I3(GND_net), .O(n47663));   // verilog/neopixel.v(104[14:39])
    defparam i1_2_lut_adj_1732.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_1733 (.I0(one_wire_N_703[8]), .I1(one_wire_N_703[7]), 
            .I2(one_wire_N_703[6]), .I3(n47663), .O(n47669));   // verilog/neopixel.v(104[14:39])
    defparam i1_4_lut_adj_1733.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1734 (.I0(one_wire_N_703[10]), .I1(n27184), .I2(one_wire_N_703[9]), 
            .I3(n47669), .O(n27032));   // verilog/neopixel.v(104[14:39])
    defparam i1_4_lut_adj_1734.LUT_INIT = 16'hfffe;
    SB_LUT4 i29277_4_lut (.I0(n27032), .I1(n40044), .I2(n44736), .I3(state[0]), 
            .O(n35336));
    defparam i29277_4_lut.LUT_INIT = 16'hfaee;
    SB_LUT4 i33918_2_lut (.I0(\neo_pixel_transmitter.done ), .I1(state[0]), 
            .I2(GND_net), .I3(GND_net), .O(n49283));
    defparam i33918_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i29281_3_lut (.I0(\neo_pixel_transmitter.done ), .I1(start), 
            .I2(n35336), .I3(GND_net), .O(n44801));
    defparam i29281_3_lut.LUT_INIT = 16'hecec;
    SB_LUT4 i15_4_lut_adj_1735 (.I0(n44801), .I1(n49283), .I2(\state[1] ), 
            .I3(n35348), .O(n7));
    defparam i15_4_lut_adj_1735.LUT_INIT = 16'h3a0a;
    SB_LUT4 i35545_2_lut (.I0(start), .I1(\state[1] ), .I2(GND_net), .I3(GND_net), 
            .O(start_N_751));   // verilog/neopixel.v(36[4] 116[11])
    defparam i35545_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 i34887_2_lut (.I0(\neo_pixel_transmitter.done ), .I1(state[0]), 
            .I2(GND_net), .I3(GND_net), .O(n43815));
    defparam i34887_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i29216_2_lut (.I0(start), .I1(\state[1] ), .I2(GND_net), .I3(GND_net), 
            .O(n44732));
    defparam i29216_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_1736 (.I0(one_wire_N_703[2]), .I1(n43815), .I2(one_wire_N_703[3]), 
            .I3(n4_adj_5239), .O(n103));
    defparam i1_4_lut_adj_1736.LUT_INIT = 16'h45cd;
    SB_LUT4 i6_4_lut (.I0(one_wire_N_703[7]), .I1(one_wire_N_703[9]), .I2(n44732), 
            .I3(n103), .O(n16_adj_5240));
    defparam i6_4_lut.LUT_INIT = 16'h0100;
    SB_LUT4 i1_4_lut_adj_1737 (.I0(one_wire_N_703[8]), .I1(one_wire_N_703[4]), 
            .I2(n16_adj_5240), .I3(n27184), .O(n6_adj_5241));
    defparam i1_4_lut_adj_1737.LUT_INIT = 16'hffef;
    SB_LUT4 i4_4_lut (.I0(one_wire_N_703[6]), .I1(one_wire_N_703[10]), .I2(one_wire_N_703[5]), 
            .I3(n6_adj_5241), .O(n51587));
    defparam i4_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 mux_1305_Mux_0_i3_3_lut (.I0(start), .I1(\neo_pixel_transmitter.done ), 
            .I2(\state[1] ), .I3(GND_net), .O(\neo_pixel_transmitter.done_N_760 ));   // verilog/neopixel.v(36[4] 116[11])
    defparam mux_1305_Mux_0_i3_3_lut.LUT_INIT = 16'hc1c1;
    SB_LUT4 color_bit_N_746_1__bdd_4_lut (.I0(color_bit_N_746[1]), .I1(n48173), 
            .I2(n48174), .I3(color_bit_N_746[2]), .O(n51282));
    defparam color_bit_N_746_1__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n51282_bdd_4_lut (.I0(n51282), .I1(n48099), .I2(n48098), .I3(color_bit_N_746[2]), 
            .O(n51285));
    defparam n51282_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n51558_bdd_4_lut (.I0(n51558), .I1(neopxl_color[9]), .I2(neopxl_color[8]), 
            .I3(color_bit_N_746[1]), .O(n51561));
    defparam n51558_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFFESS state_i0 (.Q(state[0]), .C(CLK_c), .E(n28592), .D(state_3__N_552[0]), 
            .S(n44637));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 sub_14_add_2_17_lut (.I0(n47681), .I1(timer[15]), .I2(n1[15]), 
            .I3(n38690), .O(n47683)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_17_lut.LUT_INIT = 16'hebbe;
    SB_DFF \neo_pixel_transmitter.t0_i0_i0  (.Q(\neo_pixel_transmitter.t0 [0]), 
           .C(CLK_c), .D(n29022));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i0 (.Q(bit_ctr[0]), .C(CLK_c), .E(n28484), .D(n282[0]), 
            .R(n28887));   // verilog/neopixel.v(35[12] 117[6])
    SB_CARRY add_21_8 (.CI(n38505), .I0(bit_ctr[6]), .I1(GND_net), .CO(n38506));
    SB_CARRY sub_14_add_2_17 (.CI(n38690), .I0(timer[15]), .I1(n1[15]), 
            .CO(n38691));
    SB_LUT4 i32511_3_lut (.I0(neopxl_color[0]), .I1(neopxl_color[1]), .I2(bit_ctr[0]), 
            .I3(GND_net), .O(n48098));
    defparam i32511_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i32512_3_lut (.I0(neopxl_color[2]), .I1(neopxl_color[3]), .I2(bit_ctr[0]), 
            .I3(GND_net), .O(n48099));
    defparam i32512_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i32587_3_lut (.I0(neopxl_color[6]), .I1(neopxl_color[7]), .I2(bit_ctr[0]), 
            .I3(GND_net), .O(n48174));
    defparam i32587_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i32586_3_lut (.I0(neopxl_color[4]), .I1(neopxl_color[5]), .I2(bit_ctr[0]), 
            .I3(GND_net), .O(n48173));
    defparam i32586_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 sub_14_add_2_16_lut (.I0(n47679), .I1(timer[14]), .I2(n1[14]), 
            .I3(n38689), .O(n47681)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_16_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_14_add_2_16 (.CI(n38689), .I0(timer[14]), .I1(n1[14]), 
            .CO(n38690));
    SB_LUT4 add_21_7_lut (.I0(GND_net), .I1(bit_ctr[5]), .I2(GND_net), 
            .I3(n38504), .O(n282[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_14_add_2_15_lut (.I0(n47677), .I1(timer[13]), .I2(n1[13]), 
            .I3(n38688), .O(n47679)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_15_lut.LUT_INIT = 16'hebbe;
    SB_CARRY add_21_7 (.CI(n38504), .I0(bit_ctr[5]), .I1(GND_net), .CO(n38505));
    SB_LUT4 add_21_6_lut (.I0(GND_net), .I1(bit_ctr[4]), .I2(GND_net), 
            .I3(n38503), .O(n282[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_21_6 (.CI(n38503), .I0(bit_ctr[4]), .I1(GND_net), .CO(n38504));
    SB_CARRY sub_14_add_2_15 (.CI(n38688), .I0(timer[13]), .I1(n1[13]), 
            .CO(n38689));
    SB_LUT4 i527_2_lut (.I0(n35348), .I1(\neo_pixel_transmitter.done ), 
            .I2(GND_net), .I3(GND_net), .O(n2222));   // verilog/neopixel.v(103[9] 111[12])
    defparam i527_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 i1_4_lut_adj_1738 (.I0(\state[1] ), .I1(n44630), .I2(n2222), 
            .I3(state[0]), .O(n28592));
    defparam i1_4_lut_adj_1738.LUT_INIT = 16'hee4e;
    SB_LUT4 i15_4_lut_adj_1739 (.I0(n35336), .I1(n49279), .I2(\state[1] ), 
            .I3(n27160), .O(n44637));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15_4_lut_adj_1739.LUT_INIT = 16'h303a;
    SB_LUT4 i1_2_lut_adj_1740 (.I0(bit_ctr[1]), .I1(bit_ctr[0]), .I2(GND_net), 
            .I3(GND_net), .O(color_bit_N_746[1]));
    defparam i1_2_lut_adj_1740.LUT_INIT = 16'h6666;
    SB_LUT4 sub_14_add_2_14_lut (.I0(one_wire_N_703[11]), .I1(timer[12]), 
            .I2(n1[12]), .I3(n38687), .O(n47677)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_14_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_14_add_2_14 (.CI(n38687), .I0(timer[12]), .I1(n1[12]), 
            .CO(n38688));
    SB_LUT4 sub_14_add_2_13_lut (.I0(GND_net), .I1(timer[11]), .I2(n1[11]), 
            .I3(n38686), .O(one_wire_N_703[11])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_21_5_lut (.I0(GND_net), .I1(bit_ctr[3]), .I2(GND_net), 
            .I3(n38502), .O(n282[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_13 (.CI(n38686), .I0(timer[11]), .I1(n1[11]), 
            .CO(n38687));
    SB_CARRY add_21_5 (.CI(n38502), .I0(bit_ctr[3]), .I1(GND_net), .CO(n38503));
    SB_LUT4 sub_14_add_2_12_lut (.I0(GND_net), .I1(timer[10]), .I2(n1[10]), 
            .I3(n38685), .O(one_wire_N_703[10])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_12 (.CI(n38685), .I0(timer[10]), .I1(n1[10]), 
            .CO(n38686));
    SB_LUT4 add_21_4_lut (.I0(GND_net), .I1(bit_ctr[2]), .I2(GND_net), 
            .I3(n38501), .O(n282[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_14_add_2_11_lut (.I0(GND_net), .I1(timer[9]), .I2(n1[9]), 
            .I3(n38684), .O(one_wire_N_703[9])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_11 (.CI(n38684), .I0(timer[9]), .I1(n1[9]), 
            .CO(n38685));
    SB_CARRY add_21_4 (.CI(n38501), .I0(bit_ctr[2]), .I1(GND_net), .CO(n38502));
    SB_LUT4 sub_14_add_2_10_lut (.I0(GND_net), .I1(timer[8]), .I2(n1[8]), 
            .I3(n38683), .O(one_wire_N_703[8])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_21_3_lut (.I0(GND_net), .I1(bit_ctr[1]), .I2(GND_net), 
            .I3(n38500), .O(n282[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_10 (.CI(n38683), .I0(timer[8]), .I1(n1[8]), 
            .CO(n38684));
    SB_CARRY add_21_3 (.CI(n38500), .I0(bit_ctr[1]), .I1(GND_net), .CO(n38501));
    SB_LUT4 sub_14_add_2_9_lut (.I0(GND_net), .I1(timer[7]), .I2(n1[7]), 
            .I3(n38682), .O(one_wire_N_703[7])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_9 (.CI(n38682), .I0(timer[7]), .I1(n1[7]), .CO(n38683));
    SB_LUT4 add_21_2_lut (.I0(GND_net), .I1(bit_ctr[0]), .I2(GND_net), 
            .I3(VCC_net), .O(n282[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_21_2 (.CI(VCC_net), .I0(bit_ctr[0]), .I1(GND_net), .CO(n38500));
    SB_LUT4 sub_14_add_2_8_lut (.I0(GND_net), .I1(timer[6]), .I2(n1[6]), 
            .I3(n38681), .O(one_wire_N_703[6])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_8 (.CI(n38681), .I0(timer[6]), .I1(n1[6]), .CO(n38682));
    SB_LUT4 bit_ctr_0__bdd_4_lut_35908_4_lut_4_lut (.I0(bit_ctr[1]), .I1(bit_ctr[0]), 
            .I2(neopxl_color[13]), .I3(neopxl_color[12]), .O(n51324));   // verilog/neopixel.v(19[6:15])
    defparam bit_ctr_0__bdd_4_lut_35908_4_lut_4_lut.LUT_INIT = 16'hd5c4;
    SB_LUT4 sub_14_add_2_7_lut (.I0(GND_net), .I1(timer[5]), .I2(n1[5]), 
            .I3(n38680), .O(one_wire_N_703[5])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_7 (.CI(n38680), .I0(timer[5]), .I1(n1[5]), .CO(n38681));
    SB_LUT4 sub_14_add_2_6_lut (.I0(GND_net), .I1(timer[4]), .I2(n1[4]), 
            .I3(n38679), .O(one_wire_N_703[4])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_6 (.CI(n38679), .I0(timer[4]), .I1(n1[4]), .CO(n38680));
    SB_LUT4 sub_14_add_2_5_lut (.I0(GND_net), .I1(timer[3]), .I2(n1[3]), 
            .I3(n38678), .O(one_wire_N_703[3])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_5 (.CI(n38678), .I0(timer[3]), .I1(n1[3]), .CO(n38679));
    SB_LUT4 sub_14_add_2_4_lut (.I0(GND_net), .I1(timer[2]), .I2(n1[2]), 
            .I3(n38677), .O(one_wire_N_703[2])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_4 (.CI(n38677), .I0(timer[2]), .I1(n1[2]), .CO(n38678));
    SB_LUT4 sub_14_add_2_3_lut (.I0(one_wire_N_703[3]), .I1(timer[1]), .I2(n1[1]), 
            .I3(n38676), .O(n4_adj_5239)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_3_lut.LUT_INIT = 16'h8228;
    SB_CARRY sub_14_add_2_3 (.CI(n38676), .I0(timer[1]), .I1(n1[1]), .CO(n38677));
    SB_CARRY sub_14_add_2_2 (.CI(VCC_net), .I0(timer[0]), .I1(n1[0]), 
            .CO(n38676));
    SB_LUT4 timer_2245_add_4_33_lut (.I0(GND_net), .I1(GND_net), .I2(timer[31]), 
            .I3(n39344), .O(n133[31])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2245_add_4_33_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 timer_2245_add_4_32_lut (.I0(GND_net), .I1(GND_net), .I2(timer[30]), 
            .I3(n39343), .O(n133[30])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2245_add_4_32_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2245_add_4_32 (.CI(n39343), .I0(GND_net), .I1(timer[30]), 
            .CO(n39344));
    SB_LUT4 timer_2245_add_4_31_lut (.I0(GND_net), .I1(GND_net), .I2(timer[29]), 
            .I3(n39342), .O(n133[29])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2245_add_4_31_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2245_add_4_31 (.CI(n39342), .I0(GND_net), .I1(timer[29]), 
            .CO(n39343));
    SB_LUT4 timer_2245_add_4_30_lut (.I0(GND_net), .I1(GND_net), .I2(timer[28]), 
            .I3(n39341), .O(n133[28])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2245_add_4_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2245_add_4_30 (.CI(n39341), .I0(GND_net), .I1(timer[28]), 
            .CO(n39342));
    SB_LUT4 timer_2245_add_4_29_lut (.I0(GND_net), .I1(GND_net), .I2(timer[27]), 
            .I3(n39340), .O(n133[27])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2245_add_4_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2245_add_4_29 (.CI(n39340), .I0(GND_net), .I1(timer[27]), 
            .CO(n39341));
    SB_LUT4 timer_2245_add_4_28_lut (.I0(GND_net), .I1(GND_net), .I2(timer[26]), 
            .I3(n39339), .O(n133[26])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2245_add_4_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2245_add_4_28 (.CI(n39339), .I0(GND_net), .I1(timer[26]), 
            .CO(n39340));
    SB_LUT4 timer_2245_add_4_27_lut (.I0(GND_net), .I1(GND_net), .I2(timer[25]), 
            .I3(n39338), .O(n133[25])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2245_add_4_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2245_add_4_27 (.CI(n39338), .I0(GND_net), .I1(timer[25]), 
            .CO(n39339));
    SB_LUT4 timer_2245_add_4_26_lut (.I0(GND_net), .I1(GND_net), .I2(timer[24]), 
            .I3(n39337), .O(n133[24])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2245_add_4_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2245_add_4_26 (.CI(n39337), .I0(GND_net), .I1(timer[24]), 
            .CO(n39338));
    SB_LUT4 timer_2245_add_4_25_lut (.I0(GND_net), .I1(GND_net), .I2(timer[23]), 
            .I3(n39336), .O(n133[23])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2245_add_4_25_lut.LUT_INIT = 16'hC33C;
    SB_DFF \neo_pixel_transmitter.t0_i0_i1  (.Q(\neo_pixel_transmitter.t0 [1]), 
           .C(CLK_c), .D(n29498));   // verilog/neopixel.v(35[12] 117[6])
    SB_CARRY timer_2245_add_4_25 (.CI(n39336), .I0(GND_net), .I1(timer[23]), 
            .CO(n39337));
    SB_DFF \neo_pixel_transmitter.t0_i0_i2  (.Q(\neo_pixel_transmitter.t0 [2]), 
           .C(CLK_c), .D(n29497));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i3  (.Q(\neo_pixel_transmitter.t0 [3]), 
           .C(CLK_c), .D(n29496));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i4  (.Q(\neo_pixel_transmitter.t0 [4]), 
           .C(CLK_c), .D(n29495));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i5  (.Q(\neo_pixel_transmitter.t0 [5]), 
           .C(CLK_c), .D(n29494));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i6  (.Q(\neo_pixel_transmitter.t0 [6]), 
           .C(CLK_c), .D(n29493));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i7  (.Q(\neo_pixel_transmitter.t0 [7]), 
           .C(CLK_c), .D(n29492));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i8  (.Q(\neo_pixel_transmitter.t0 [8]), 
           .C(CLK_c), .D(n29491));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i9  (.Q(\neo_pixel_transmitter.t0 [9]), 
           .C(CLK_c), .D(n29490));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i10  (.Q(\neo_pixel_transmitter.t0 [10]), 
           .C(CLK_c), .D(n29489));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i11  (.Q(\neo_pixel_transmitter.t0 [11]), 
           .C(CLK_c), .D(n29488));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i12  (.Q(\neo_pixel_transmitter.t0 [12]), 
           .C(CLK_c), .D(n29487));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 timer_2245_add_4_24_lut (.I0(GND_net), .I1(GND_net), .I2(timer[22]), 
            .I3(n39335), .O(n133[22])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2245_add_4_24_lut.LUT_INIT = 16'hC33C;
    SB_DFF \neo_pixel_transmitter.t0_i0_i13  (.Q(\neo_pixel_transmitter.t0 [13]), 
           .C(CLK_c), .D(n29486));   // verilog/neopixel.v(35[12] 117[6])
    SB_CARRY timer_2245_add_4_24 (.CI(n39335), .I0(GND_net), .I1(timer[22]), 
            .CO(n39336));
    SB_DFF \neo_pixel_transmitter.t0_i0_i14  (.Q(\neo_pixel_transmitter.t0 [14]), 
           .C(CLK_c), .D(n29485));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 timer_2245_add_4_23_lut (.I0(GND_net), .I1(GND_net), .I2(timer[21]), 
            .I3(n39334), .O(n133[21])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2245_add_4_23_lut.LUT_INIT = 16'hC33C;
    SB_DFF \neo_pixel_transmitter.t0_i0_i15  (.Q(\neo_pixel_transmitter.t0 [15]), 
           .C(CLK_c), .D(n29484));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i16  (.Q(\neo_pixel_transmitter.t0 [16]), 
           .C(CLK_c), .D(n29483));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i17  (.Q(\neo_pixel_transmitter.t0 [17]), 
           .C(CLK_c), .D(n29482));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i18  (.Q(\neo_pixel_transmitter.t0 [18]), 
           .C(CLK_c), .D(n29481));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i19  (.Q(\neo_pixel_transmitter.t0 [19]), 
           .C(CLK_c), .D(n29480));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i20  (.Q(\neo_pixel_transmitter.t0 [20]), 
           .C(CLK_c), .D(n29479));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i21  (.Q(\neo_pixel_transmitter.t0 [21]), 
           .C(CLK_c), .D(n29478));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i22  (.Q(\neo_pixel_transmitter.t0 [22]), 
           .C(CLK_c), .D(n29477));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i23  (.Q(\neo_pixel_transmitter.t0 [23]), 
           .C(CLK_c), .D(n29476));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i24  (.Q(\neo_pixel_transmitter.t0 [24]), 
           .C(CLK_c), .D(n29475));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i25  (.Q(\neo_pixel_transmitter.t0 [25]), 
           .C(CLK_c), .D(n29474));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i26  (.Q(\neo_pixel_transmitter.t0 [26]), 
           .C(CLK_c), .D(n29473));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i27  (.Q(\neo_pixel_transmitter.t0 [27]), 
           .C(CLK_c), .D(n29472));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i28  (.Q(\neo_pixel_transmitter.t0 [28]), 
           .C(CLK_c), .D(n29471));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i29  (.Q(\neo_pixel_transmitter.t0 [29]), 
           .C(CLK_c), .D(n29470));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i30  (.Q(\neo_pixel_transmitter.t0 [30]), 
           .C(CLK_c), .D(n29469));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i31  (.Q(\neo_pixel_transmitter.t0 [31]), 
           .C(CLK_c), .D(n29468));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 sub_14_inv_0_i17_1_lut (.I0(\neo_pixel_transmitter.t0 [16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[16]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY timer_2245_add_4_23 (.CI(n39334), .I0(GND_net), .I1(timer[21]), 
            .CO(n39335));
    SB_LUT4 timer_2245_add_4_22_lut (.I0(GND_net), .I1(GND_net), .I2(timer[20]), 
            .I3(n39333), .O(n133[20])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2245_add_4_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2245_add_4_22 (.CI(n39333), .I0(GND_net), .I1(timer[20]), 
            .CO(n39334));
    SB_LUT4 timer_2245_add_4_21_lut (.I0(GND_net), .I1(GND_net), .I2(timer[19]), 
            .I3(n39332), .O(n133[19])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2245_add_4_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2245_add_4_21 (.CI(n39332), .I0(GND_net), .I1(timer[19]), 
            .CO(n39333));
    SB_LUT4 timer_2245_add_4_20_lut (.I0(GND_net), .I1(GND_net), .I2(timer[18]), 
            .I3(n39331), .O(n133[18])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2245_add_4_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2245_add_4_20 (.CI(n39331), .I0(GND_net), .I1(timer[18]), 
            .CO(n39332));
    SB_LUT4 timer_2245_add_4_19_lut (.I0(GND_net), .I1(GND_net), .I2(timer[17]), 
            .I3(n39330), .O(n133[17])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2245_add_4_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2245_add_4_19 (.CI(n39330), .I0(GND_net), .I1(timer[17]), 
            .CO(n39331));
    SB_LUT4 timer_2245_add_4_18_lut (.I0(GND_net), .I1(GND_net), .I2(timer[16]), 
            .I3(n39329), .O(n133[16])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2245_add_4_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2245_add_4_18 (.CI(n39329), .I0(GND_net), .I1(timer[16]), 
            .CO(n39330));
    SB_LUT4 add_21_33_lut (.I0(GND_net), .I1(bit_ctr[31]), .I2(GND_net), 
            .I3(n38530), .O(n282[31])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_33_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_21_32_lut (.I0(GND_net), .I1(bit_ctr[30]), .I2(GND_net), 
            .I3(n38529), .O(n282[30])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_32_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 timer_2245_add_4_17_lut (.I0(GND_net), .I1(GND_net), .I2(timer[15]), 
            .I3(n39328), .O(n133[15])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2245_add_4_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2245_add_4_17 (.CI(n39328), .I0(GND_net), .I1(timer[15]), 
            .CO(n39329));
    SB_CARRY add_21_32 (.CI(n38529), .I0(bit_ctr[30]), .I1(GND_net), .CO(n38530));
    SB_LUT4 add_21_31_lut (.I0(GND_net), .I1(bit_ctr[29]), .I2(GND_net), 
            .I3(n38528), .O(n282[29])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_31_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 timer_2245_add_4_14_lut (.I0(GND_net), .I1(GND_net), .I2(timer[12]), 
            .I3(n39325), .O(n133[12])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2245_add_4_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 timer_2245_add_4_16_lut (.I0(GND_net), .I1(GND_net), .I2(timer[14]), 
            .I3(n39327), .O(n133[14])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2245_add_4_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2245_add_4_16 (.CI(n39327), .I0(GND_net), .I1(timer[14]), 
            .CO(n39328));
    SB_LUT4 timer_2245_add_4_15_lut (.I0(GND_net), .I1(GND_net), .I2(timer[13]), 
            .I3(n39326), .O(n133[13])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2245_add_4_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 timer_2245_add_4_12_lut (.I0(GND_net), .I1(GND_net), .I2(timer[10]), 
            .I3(n39323), .O(n133[10])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2245_add_4_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_21_31 (.CI(n38528), .I0(bit_ctr[29]), .I1(GND_net), .CO(n38529));
    SB_LUT4 add_21_30_lut (.I0(GND_net), .I1(bit_ctr[28]), .I2(GND_net), 
            .I3(n38527), .O(n282[28])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_21_30 (.CI(n38527), .I0(bit_ctr[28]), .I1(GND_net), .CO(n38528));
    SB_LUT4 add_21_29_lut (.I0(GND_net), .I1(bit_ctr[27]), .I2(GND_net), 
            .I3(n38526), .O(n282[27])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_21_29 (.CI(n38526), .I0(bit_ctr[27]), .I1(GND_net), .CO(n38527));
    SB_DFFESR one_wire_108 (.Q(NEOPXL_c), .C(CLK_c), .E(n44865), .D(\neo_pixel_transmitter.done_N_766 ), 
            .R(n46519));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 add_21_28_lut (.I0(GND_net), .I1(bit_ctr[26]), .I2(GND_net), 
            .I3(n38525), .O(n282[26])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_21_28 (.CI(n38525), .I0(bit_ctr[26]), .I1(GND_net), .CO(n38526));
    SB_LUT4 add_21_27_lut (.I0(GND_net), .I1(bit_ctr[25]), .I2(GND_net), 
            .I3(n38524), .O(n282[25])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_21_27 (.CI(n38524), .I0(bit_ctr[25]), .I1(GND_net), .CO(n38525));
    SB_LUT4 sub_14_inv_0_i18_1_lut (.I0(\neo_pixel_transmitter.t0 [17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[17]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i33805_2_lut_3_lut (.I0(n35348), .I1(\neo_pixel_transmitter.done ), 
            .I2(state[0]), .I3(GND_net), .O(n49279));   // verilog/neopixel.v(35[12] 117[6])
    defparam i33805_2_lut_3_lut.LUT_INIT = 16'hfdfd;
    SB_LUT4 i1_2_lut_3_lut (.I0(n35336), .I1(start), .I2(\neo_pixel_transmitter.done ), 
            .I3(GND_net), .O(n44630));
    defparam i1_2_lut_3_lut.LUT_INIT = 16'h2020;
    SB_LUT4 bit_ctr_0__bdd_4_lut_4_lut (.I0(bit_ctr[0]), .I1(neopxl_color[10]), 
            .I2(neopxl_color[11]), .I3(bit_ctr[1]), .O(n51558));
    defparam bit_ctr_0__bdd_4_lut_4_lut.LUT_INIT = 16'heea0;
    SB_LUT4 i2_2_lut_3_lut (.I0(n27032), .I1(one_wire_N_703[3]), .I2(one_wire_N_703[2]), 
            .I3(GND_net), .O(n35127));
    defparam i2_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i2_3_lut_4_lut (.I0(state[0]), .I1(\state[1] ), .I2(LED_c), 
            .I3(\state_3__N_552[1] ), .O(n28887));   // verilog/neopixel.v(35[12] 117[6])
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 n51324_bdd_4_lut_4_lut (.I0(color_bit_N_746[1]), .I1(neopxl_color[14]), 
            .I2(neopxl_color[15]), .I3(n51324), .O(n51327));   // verilog/neopixel.v(19[6:15])
    defparam n51324_bdd_4_lut_4_lut.LUT_INIT = 16'hf588;
    SB_LUT4 sub_14_inv_0_i19_1_lut (.I0(\neo_pixel_transmitter.t0 [18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[18]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i21312_2_lut_3_lut (.I0(bit_ctr[1]), .I1(bit_ctr[0]), .I2(bit_ctr[2]), 
            .I3(GND_net), .O(n35253));
    defparam i21312_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_2_lut_3_lut_adj_1741 (.I0(bit_ctr[1]), .I1(bit_ctr[0]), .I2(bit_ctr[2]), 
            .I3(GND_net), .O(color_bit_N_746[2]));
    defparam i1_2_lut_3_lut_adj_1741.LUT_INIT = 16'h1e1e;
    SB_LUT4 sub_14_inv_0_i20_1_lut (.I0(\neo_pixel_transmitter.t0 [19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[19]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i21_1_lut (.I0(\neo_pixel_transmitter.t0 [20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[20]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i22_1_lut (.I0(\neo_pixel_transmitter.t0 [21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[21]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i23_1_lut (.I0(\neo_pixel_transmitter.t0 [22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[22]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i24_1_lut (.I0(\neo_pixel_transmitter.t0 [23]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[23]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i25_1_lut (.I0(\neo_pixel_transmitter.t0 [24]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[24]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i25_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i26_1_lut (.I0(\neo_pixel_transmitter.t0 [25]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[25]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i26_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i27_1_lut (.I0(\neo_pixel_transmitter.t0 [26]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[26]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i27_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i28_1_lut (.I0(\neo_pixel_transmitter.t0 [27]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[27]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i28_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i34130_3_lut_4_lut (.I0(n27032), .I1(n49717), .I2(start), 
            .I3(\state[1] ), .O(n49718));
    defparam i34130_3_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i33935_2_lut_3_lut (.I0(one_wire_N_703[3]), .I1(one_wire_N_703[2]), 
            .I2(start), .I3(GND_net), .O(n49277));
    defparam i33935_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i3_4_lut_4_lut (.I0(n35348), .I1(\state[1] ), .I2(state[0]), 
            .I3(\neo_pixel_transmitter.done ), .O(n46519));
    defparam i3_4_lut_4_lut.LUT_INIT = 16'h0004;
    SB_LUT4 sub_14_inv_0_i29_1_lut (.I0(\neo_pixel_transmitter.t0 [28]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[28]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i29_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 color_bit_N_746_1__bdd_4_lut_35681 (.I0(color_bit_N_746[1]), .I1(n48056), 
            .I2(n48057), .I3(color_bit_N_746[2]), .O(n51216));
    defparam color_bit_N_746_1__bdd_4_lut_35681.LUT_INIT = 16'he4aa;
    SB_LUT4 n51216_bdd_4_lut (.I0(n51216), .I1(n48168), .I2(n48167), .I3(color_bit_N_746[2]), 
            .O(n51219));
    defparam n51216_bdd_4_lut.LUT_INIT = 16'haad8;
    
endmodule
//
// Verilog Description of module motorControl
//

module motorControl (\Kp[13] , GND_net, \Kp[14] , \Kp[1] , \Kp[0] , 
            \Kp[15] , \Ki[6] , \Ki[3] , \Ki[4] , \Kp[2] , \Kp[3] , 
            \Ki[5] , \Kp[4] , PWMLimit, \Kp[5] , \Ki[7] , \Kp[9] , 
            \Ki[8] , \Kp[6] , \Ki[2] , \Ki[9] , \Ki[10] , \Ki[1] , 
            \Ki[0] , \Ki[11] , \Kp[10] , \Kp[7] , \Kp[8] , \Kp[11] , 
            \Kp[12] , \Ki[12] , \Ki[13] , \Ki[14] , \Ki[15] , IntegralLimit, 
            duty, clk32MHz, VCC_net, setpoint, motor_state) /* synthesis syn_module_defined=1 */ ;
    input \Kp[13] ;
    input GND_net;
    input \Kp[14] ;
    input \Kp[1] ;
    input \Kp[0] ;
    input \Kp[15] ;
    input \Ki[6] ;
    input \Ki[3] ;
    input \Ki[4] ;
    input \Kp[2] ;
    input \Kp[3] ;
    input \Ki[5] ;
    input \Kp[4] ;
    input [23:0]PWMLimit;
    input \Kp[5] ;
    input \Ki[7] ;
    input \Kp[9] ;
    input \Ki[8] ;
    input \Kp[6] ;
    input \Ki[2] ;
    input \Ki[9] ;
    input \Ki[10] ;
    input \Ki[1] ;
    input \Ki[0] ;
    input \Ki[11] ;
    input \Kp[10] ;
    input \Kp[7] ;
    input \Kp[8] ;
    input \Kp[11] ;
    input \Kp[12] ;
    input \Ki[12] ;
    input \Ki[13] ;
    input \Ki[14] ;
    input \Ki[15] ;
    input [23:0]IntegralLimit;
    output [23:0]duty;
    input clk32MHz;
    input VCC_net;
    input [23:0]setpoint;
    input [23:0]motor_state;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    wire [23:0]n1;
    
    wire n968, n1041, n116, n38733;
    wire [23:0]n1_adj_5234;
    
    wire n38734, n47, n1114;
    wire [23:0]\PID_CONTROLLER.integral_23__N_3836 ;
    
    wire n463, n256, n329, n189, n262, n89, n20_adj_4815, n402, 
        n335, n475, n39716;
    wire [20:0]n12180;
    
    wire n296, n39717;
    wire [23:0]n1_adj_5235;
    
    wire n408, n7, n38732;
    wire [23:0]\PID_CONTROLLER.integral ;   // verilog/motorControl.v(23[23:31])
    
    wire n548, n697;
    wire [14:0]n16544;
    wire [13:0]n17024;
    
    wire n974, n39582, n621, n481, n177, n694, n767, n95, n26, 
        n840, n770, n554, n627, n162, n235, n308, n700, n381, 
        n454, n89_adj_4816, n20_adj_4817, n74, n5, n162_adj_4818, 
        n527, n600, n673, n746, n5_adj_4819, n38731, n39583;
    wire [21:0]n11163;
    
    wire n223, n39715, n901, n39581, n819, n892, n147, n828, 
        n39580, n965, n1038, n1111, n116_adj_4820, n47_adj_4821, 
        n189_adj_4822, n220, n262_adj_4823, n335_adj_4824, n235_adj_4825, 
        n408_adj_4826, n481_adj_4827, n308_adj_4828, n554_adj_4829, 
        n293, n366, n627_adj_4830, n700_adj_4831, n381_adj_4832, n86, 
        n17, n159, n439, n536, n609, n512, n454_adj_4834, n232, 
        n305, n527_adj_4835, n600_adj_4836, n585, n673_adj_4837, n378, 
        n451, n524, n597, n670, n743, n816, n658, n746_adj_4838, 
        n889, n819_adj_4839, n892_adj_4840, n962, n1035, n965_adj_4841, 
        n1108, n731, n1038_adj_4842, n804, n3, n38730, n83, n14_adj_4844, 
        n156, n1111_adj_4845, n877, n229, n302, n375, n448, n86_adj_4846, 
        n17_adj_4847, n521, n755, n39579, n159_adj_4848, n369, n1047, 
        n232_adj_4849, n950, n305_adj_4851, n378_adj_4852, n1120, 
        n442, n594, n667, n740, n813, n886, n959, n1023, n515, 
        n1032, n250, n1105, n451_adj_4854, n323, n83_adj_4855, n14_adj_4856, 
        n156_adj_4857, n396, n588, n229_adj_4858, n661, n302_adj_4859, 
        \PID_CONTROLLER.integral_23__N_3884 ;
    wire [23:0]n4751;
    
    wire n1096, n469, n150, n39714, n542, n682, n39578, n375_adj_4861, 
        n448_adj_4862, n734, n119, n615, n50, n807, n521_adj_4865, 
        n880, n953, n1026, n8, n77;
    wire [19:0]n13104;
    
    wire n39713, n688, n192, n39577, n39712, n761, n1099, n110, 
        n41, n39576, n183, n39711, n834, n39710, n256_adj_4873, 
        n594_adj_4874, n39575, n907, n265, n329_adj_4877, n980, 
        n667_adj_4879, n122, n53, n402_adj_4881, n740_adj_4882, n195, 
        n813_adj_4885, n268, n341, n414, n886_adj_4887, n487, n959_adj_4888, 
        n338, n1032_adj_4890, n560, n1105_adj_4891, n101, n32, n174, 
        n247, n320, n393, n80, n11_adj_4897, n80_adj_4898, n11_adj_4899, 
        n153, n466, n226, n539;
    wire [23:0]duty_23__N_3812;
    
    wire n612, n299;
    wire [23:0]\PID_CONTROLLER.integral_23__N_3887 ;
    
    wire n38729, n38728, n153_adj_4904, n17_adj_4905, n9_adj_4906, 
        n11_adj_4907, n38727, n49653, n49651, n226_adj_4908, n51808, 
        n50178, n49959, n51790, n49957, n39709, n49955, n38726, 
        n51784, n27, n15_adj_4909, n13_adj_4910, n11_adj_4911, n49600, 
        n21_adj_4912, n19_adj_4913, n17_adj_4914, n9_adj_4915, n49606, 
        n43, n16_adj_4916, n49583, n411, n8_adj_4917, n45, n24_adj_4918, 
        n299_adj_4919, n49619, n49931, n49927, n25_adj_4920, n23_adj_4921, 
        n50354, n372, n31, n29, n50152, n37, n35, n33, n50416, 
        n49961, n524_adj_4923, n51777, n49949, n51772, n12_adj_4924, 
        n49631, n51795, n10_adj_4925, n30, n50300, n49639, n51775, 
        n445, n518, n591, n664, n50172, n51801, n390, n39574, 
        n50360, n51766, n317, n39573, n244, n39572, n171, n39571, 
        n29_adj_4927, n98, n50446, n51763, n16_adj_4928;
    wire [12:0]n17444;
    
    wire n1050, n39570, n39708, n49621, n737, n38725, n810, n883, 
        n956, n1029, n24_adj_4929, n6_adj_4930, n1102, n50246, n77_adj_4932, 
        n8_adj_4933, n50247, n150_adj_4934, n1102_adj_4935, n39707, 
        n1029_adj_4936, n39706, n956_adj_4937, n39705, n49623, n223_adj_4938, 
        n296_adj_4939, n977, n39569, n883_adj_4940, n39704, n8_adj_4941, 
        n51761, n50248, n369_adj_4942, n442_adj_4943, n49764, n515_adj_4944, 
        n4_adj_4945, n588_adj_4946, n50274, n50275, n661_adj_4947, 
        n12_adj_4949, n49594, n10_adj_4950, n734_adj_4951, n807_adj_4952, 
        n30_adj_4953, n49596, n50382, n49776, n50460, n50461, n904, 
        n39568, n38724, n39, n50439, n6_adj_4954, n880_adj_4955, 
        n953_adj_4957, n1026_adj_4958, n810_adj_4959, n39703, n737_adj_4960, 
        n39702, n831, n39567, n1099_adj_4961, n50278, n50279, n49585, 
        n50250, n49774, n41_adj_4962, n49587, n74_adj_4964, n38723, 
        n5_adj_4965, n147_adj_4966, n484, n50396, n220_adj_4967, n293_adj_4968, 
        n664_adj_4969, n39701, n758, n39566, n49782, n50398, n4_adj_4970, 
        n50284, n50285, n49633, n50380, n49766, n50458, n475_adj_4971, 
        n50459, n50443, n366_adj_4972, n49625, n439_adj_4973, n50392, 
        n49772, n548_adj_4975, n512_adj_4976, n585_adj_4977, n591_adj_4978, 
        n39700, n685, n39565, n658_adj_4979, \PID_CONTROLLER.integral_23__N_3886 , 
        n50394, n621_adj_4980, n518_adj_4981, n39699, n731_adj_4982, 
        n445_adj_4983, n39698, n372_adj_4984, n39697, n694_adj_4985, 
        n804_adj_4986, n877_adj_4987, n950_adj_4988, n38637, n38722, 
        n39696, n1023_adj_4989, n1096_adj_4990, n557, n39564, n39563, 
        n39695, n39562, n767_adj_4991, n597_adj_4992, n39694, n38636, 
        n38721;
    wire [18:0]n13944;
    
    wire n39693, n39561, n39692, n630, n840_adj_4994, n39691, n107, 
        n38, n39560, n39690, n38635, n39559, n180, n38720, n39689, 
        n38634, n38719, n39558;
    wire [23:0]duty_23__N_3936;
    wire [23:0]n257;
    
    wire n256_adj_4995;
    wire [23:0]duty_23__N_3911;
    
    wire duty_23__N_3935, n38718, n39688, n253;
    wire [6:0]n18991;
    wire [5:0]n19088;
    
    wire n39557, n326, n39687, n39686, n39556, n39685, n39555, 
        n39554, n38633, n38717, n39553, n38716, n39684, n399, 
        n38632, n38715, n38631, n38714, n39552, n39683, n38713, 
        n39682;
    wire [11:0]n17808;
    
    wire n39551, n38630, n39550, n38629, n38712, n38628, n38711, 
        n39681, n39549, n38710, n39548, n38709, n39547, n38627, 
        n38708, n38707, n39680, n39546, n38626, n39679, n39678, 
        n39545, n39544, n38625, n39677, n472, n39676, n39543, 
        n39675, n39542, n39541, n545, n618;
    wire [9:0]n18504;
    wire [8:0]n18703;
    
    wire n39674, n39540, n691, n39673, n168, n624, n39672, n38624, 
        n35_adj_5004, n104, n551, n39671, n38623, n478, n39670;
    wire [10:0]n18120;
    
    wire n910, n39539, n241, n837, n39538, n38622, n405, n39669, 
        n38621, n38620, n38619, n38618, n764, n39537, n332, n39668, 
        n38617, n691_adj_5005, n39536, n259_adj_5006, n39667, n38616, 
        n186, n39666, n618_adj_5007, n39535, n38615, n44, n113, 
        n545_adj_5008, n39534;
    wire [17:0]n14704;
    
    wire n39665, n39664, n472_adj_5009, n39533, n39663, n399_adj_5010, 
        n39532, n39662, n326_adj_5011, n39531, n253_adj_5012, n39530, 
        n314, n670_adj_5013, n180_adj_5014, n39529, n38_adj_5015, 
        n107_adj_5016, n764_adj_5017, n837_adj_5018, n910_adj_5019, 
        n387, n460, n125, n56, n45851, n490, n39528, n1108_adj_5020, 
        n39661, n198, n271_adj_5022, n344, n417, n6_adj_5023;
    wire [3:0]n19184;
    wire [4:0]n19124;
    wire [4:0]n19159;
    
    wire n417_adj_5024, n39527, n1035_adj_5025, n39660, n962_adj_5026, 
        n39659, n889_adj_5027, n39658, n344_adj_5028, n39526, n271_adj_5029, 
        n39525, n198_adj_5030, n39524, n816_adj_5031, n39657, n56_adj_5032, 
        n125_adj_5033, n743_adj_5034, n39656;
    wire [0:0]n11187;
    wire [0:0]n10656;
    
    wire n38614, n39655;
    wire [47:0]n106;
    wire [47:0]n155;
    
    wire n38613, n4_adj_5035;
    wire [2:0]n19224;
    wire [1:0]n19248;
    
    wire n490_adj_5036, n12_adj_5037, n8_adj_5038, n11_adj_5039, n6_adj_5040, 
        n38389, n39654, n18_adj_5041, n13_adj_5042, n4_adj_5043, n46355, 
        n49485, n49506;
    wire [21:0]n11694;
    
    wire n39990, n39989, n39988, n39987, n39986, n104_adj_5044, 
        n39985, n39984, n39983, n39982, n39981, n35_adj_5045, n39980, 
        n39979, n177_adj_5046, n39978, n39977, n39976, n39975, n39974, 
        n39973, n250_adj_5048, n323_adj_5049, n39972, n49544, n396_adj_5050, 
        n469_adj_5051, n533, n39971, n39970, n39969, n542_adj_5055;
    wire [20:0]n12663;
    
    wire n39968, n39967, n39966, n39965, n615_adj_5056, n39964, 
        n39963, n688_adj_5057, n39962, n606, n761_adj_5058, n39961, 
        n39960, n39959, n39958, n834_adj_5059, n39957, n39956, n39955, 
        n39954, n39953, n39952, n39951, n39950, n49557, n907_adj_5061, 
        n39949, n39948;
    wire [19:0]n13544;
    
    wire n39947, n39946, n39945, n980_adj_5063, n39944, n39943, 
        n101_adj_5064, n32_adj_5065, n174_adj_5066, n39942, n39941, 
        n39940, n39939, n39938, n39937, n247_adj_5067, n39936, n39935, 
        n39934, n39933, n39932, n320_adj_5069, n38612, n393_adj_5071, 
        n38611, n466_adj_5073, n539_adj_5074, n679, n612_adj_5075, 
        n39653, n39931, n39930, n39929, n39928;
    wire [18:0]n14343;
    
    wire n39927, n685_adj_5078, n39926, n39652, n38610, n758_adj_5079, 
        n39925, n39924, n39923, n39922, n39921, n38609, n39920, 
        n39919, n39918, n39917, n39916, n39915, n39651, n39650, 
        n39649, n39648, n39914, n39913, n39912, n39911, n39910;
    wire [16:0]n15388;
    
    wire n39647, n39646, n38608, n752, n39645, n38607, n39644, 
        n39909;
    wire [17:0]n15064;
    
    wire n39908, n39907, n39906, n38606, n39643, n38605, n38604, 
        n39905, n39904, n39642, n39903, n39902, n39641, n39640, 
        n39901, n39639, n39900, n39899, n38603, n39898, n39897, 
        n39896, n39895, n39894, n39638, n39637, n38602, n39636, 
        n39893, n39892, n39635, n831_adj_5083, n904_adj_5084, n39891, 
        n39634;
    wire [8:0]n18604;
    wire [7:0]n18784;
    
    wire n39890, n39889, n38601, n38600, n39888, n39633, n39887, 
        n39886, n38599, n39632, n39885, n39884, n39883;
    wire [16:0]n15711;
    
    wire n39882, n39881, n39880, n39879, n39878, n39877, n38598, 
        n39876, n39875, n39874, n39873, n39872, n39871, n39631, 
        n39870, n39869;
    wire [7:0]n18864;
    
    wire n39630, n38597, n39868, n39867, n825, n39866, n39629, 
        n39628;
    wire [9:0]n18384;
    
    wire n39492, n39491, n39490, n39627, n38596, n39489, n39488, 
        n39626, n39487, n39625, n39486;
    wire [15:0]n16288;
    
    wire n39865, n39864, n39624, n39623, n39485, n39484, n39863, 
        n39862, n39861, n895, n39860, n822, n39859, n38595, n749, 
        n39858, n676, n39857, n603, n39856, n530, n39855, n457, 
        n39854, n384, n39853, n183_adj_5087, n39483, n311, n39852, 
        n238, n39851, n165, n39850, n23_adj_5088, n92;
    wire [6:0]n18928;
    
    wire n630_adj_5089, n39849, n38594;
    wire [15:0]n16000;
    
    wire n39622, n557_adj_5090, n39848, n484_adj_5091, n39847, n411_adj_5092, 
        n39846, n338_adj_5093, n39845, n265_adj_5094, n39844, n770_adj_5095, 
        n38820, n192_adj_5096, n39843, n38593, n39621, n41_adj_5097, 
        n110_adj_5098, n697_adj_5099, n38819, n50_adj_5100, n119_adj_5101, 
        n38592, n1114_adj_5102, n39620, n624_adj_5103, n38818, n1041_adj_5104, 
        n39619;
    wire [14:0]n16799;
    
    wire n39842, n1117, n39841, n1044, n39840, n551_adj_5105, n38817, 
        n478_adj_5106, n38816, n405_adj_5107, n38815, n968_adj_5108, 
        n39618, n971, n39839, n332_adj_5109, n38814, n898, n39838, 
        n259_adj_5110, n38813, n825_adj_5111, n39837, n752_adj_5112, 
        n39836, n186_adj_5113, n38812, n44_adj_5114, n113_adj_5115, 
        n895_adj_5116, n39617, n822_adj_5117, n39616, n679_adj_5118, 
        n39835, n749_adj_5119, n39615, n676_adj_5120, n39614, n603_adj_5121, 
        n39613, n530_adj_5122, n39612, n606_adj_5123, n39834, n533_adj_5124, 
        n39833, n460_adj_5125, n39832, n387_adj_5126, n39831, n314_adj_5127, 
        n39830, n241_adj_5128, n39829, n457_adj_5129, n39611, n168_adj_5130, 
        n39828, n384_adj_5131, n39610, n26_adj_5132, n95_adj_5133;
    wire [13:0]n17248;
    
    wire n1120_adj_5134, n39827, n1047_adj_5135, n39826, n974_adj_5136, 
        n39825, n901_adj_5137, n39824, n828_adj_5138, n39823, n755_adj_5139, 
        n39822, n682_adj_5140, n39821, n311_adj_5141, n39609, n609_adj_5142, 
        n39820, n49542, n238_adj_5143, n39608, n536_adj_5144, n39819, 
        n463_adj_5145, n39818, n390_adj_5146, n39817, n317_adj_5147, 
        n39816, n244_adj_5148, n39815, n171_adj_5149, n39814, n29_adj_5150, 
        n98_adj_5151;
    wire [5:0]n19040;
    
    wire n560_adj_5152, n39813, n487_adj_5153, n39812, n6_adj_5154, 
        n898_adj_5155, n414_adj_5156, n39811, n341_adj_5157, n39810, 
        n268_adj_5158, n39809, n165_adj_5159, n39607, n195_adj_5160, 
        n39808, n53_adj_5161, n122_adj_5162;
    wire [12:0]n17639;
    
    wire n1050_adj_5163, n39807, n977_adj_5164, n39806, n49581, n23_adj_5165, 
        n92_adj_5166, n39606, n1117_adj_5167, n39605, n1044_adj_5168, 
        n39604, n971_adj_5169, n39603, n39602, n39601, n39805, n39804, 
        n39600, n39803, n39802, n6_adj_5170, n38775, n38774, n39801, 
        n39599, n39800, n39799, n39798, n38773, n39797, n38772, 
        n39796, n39795;
    wire [11:0]n17976;
    
    wire n39794, n38771, n39793, n38770, n39792, n39791, n39598, 
        n39790, n39789, n39788, n39597, n38769, n39787, n39786, 
        n39785, n39784, n39783, n39782, n39781, n39780, n39779, 
        n38768, n39778, n39596, n39595;
    wire [10:0]n18263;
    
    wire n39777, n39776, n39775, n39594, n39593, n38767, n39592, 
        n39774, n39773, n39772, n39771, n39770, n39769, n39768, 
        n39767, n39766, n39765, n39764, n39763, n39762, n39761, 
        n38766, n38765, n38764, n39760, n39759, n39758, n39757, 
        n39756, n39755, n39754, n39753, n39752, n39751, n39750, 
        n39749, n39748, n39747, n39746, n39745, n39744, n39743, 
        n39742, n39741, n39740, n39739, n39738, n39737, n39736, 
        n39735, n39734, n38763, n39733, n39732, n38762, n6_adj_5171;
    wire [3:0]n19208;
    
    wire n38761, n39731, n39591, n38760, n39590, n38759, n39730, 
        n39589, n38758, n39729, n38757, n39588, n38756, n38755, 
        n38754, n39728, n39587, n38753, n38752, n38751, n38750, 
        n39586, n38749, n38748, n38747, n38746, n38745, n39727, 
        n39585, n38744, n38743, n38742, n38741, n39726, n38740, 
        n39725, n38739, n39724, n39723, n38738, n39722, n39721, 
        n39720, n38737, n39719, n38736, n39718, n38735, n39584;
    wire [1:0]n19256;
    
    wire n4_adj_5172;
    wire [2:0]n19239;
    
    wire n12_adj_5173, n8_adj_5174, n11_adj_5175, n6_adj_5176, n38216, 
        n4_adj_5177, n18_adj_5178, n13_adj_5179, n4_adj_5180, n38355, 
        n38323, n38405, n38232, n38191, n4_adj_5181, n38273, n41_adj_5182, 
        n39_adj_5183, n45_adj_5184, n37_adj_5185, n23_adj_5186, n25_adj_5187, 
        n43_adj_5188, n29_adj_5189, n31_adj_5190, n35_adj_5191, n11_adj_5192, 
        n13_adj_5193, n15_adj_5194, n27_adj_5195, n33_adj_5196, n9_adj_5197, 
        n17_adj_5198, n19_adj_5199, n21_adj_5200, n49571, n49563, 
        n12_adj_5201, n10_adj_5202, n30_adj_5203, n49897, n49893, 
        n50342, n50104, n50410, n16_adj_5204, n50136, n50137, n8_adj_5205, 
        n24_adj_5206, n49546, n50252, n49784, n4_adj_5207, n50122, 
        n50123, n49559, n50330, n49786, n50436, n50437, n50415, 
        n49548, n50400, n49792, n50402, n39_adj_5208, n41_adj_5209, 
        n45_adj_5210, n37_adj_5211, n29_adj_5212, n31_adj_5213, n23_adj_5214, 
        n25_adj_5215, n43_adj_5216, n35_adj_5217, n33_adj_5218, n11_adj_5219, 
        n13_adj_5220, n15_adj_5221, n27_adj_5222, n9_adj_5223, n17_adj_5224, 
        n19_adj_5225, n21_adj_5226, n49531, n49520, n12_adj_5227, 
        n10_adj_5228, n30_adj_5229, n49865, n49861, n50334, n50088, 
        n50408, n16_adj_5230, n50112, n50113, n8_adj_5231, n24_adj_5232, 
        n49489, n50254, n49794, n4_adj_5233, n50108, n50109, n49511, 
        n50336, n49796, n50432, n50433, n50413, n49491, n50404, 
        n49802, n50406;
    
    SB_LUT4 mult_10_i651_2_lut (.I0(\Kp[13] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n968));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i651_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i700_2_lut (.I0(\Kp[14] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n1041));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i700_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i79_2_lut (.I0(\Kp[1] ), .I1(n1[14]), .I2(GND_net), 
            .I3(GND_net), .O(n116));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i79_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY unary_minus_5_add_3_6 (.CI(n38733), .I0(GND_net), .I1(n1_adj_5234[4]), 
            .CO(n38734));
    SB_LUT4 mult_10_i32_2_lut (.I0(\Kp[0] ), .I1(n1[15]), .I2(GND_net), 
            .I3(GND_net), .O(n47));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i32_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i749_2_lut (.I0(\Kp[15] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n1114));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i749_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i312_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n463));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i312_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i173_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n256));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i173_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i222_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n329));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i222_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i128_2_lut (.I0(\Kp[2] ), .I1(n1[14]), .I2(GND_net), 
            .I3(GND_net), .O(n189));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i128_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i177_2_lut (.I0(\Kp[3] ), .I1(n1[14]), .I2(GND_net), 
            .I3(GND_net), .O(n262));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i177_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i61_2_lut (.I0(\Kp[1] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n89));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i61_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i14_2_lut (.I0(\Kp[0] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n20_adj_4815));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i14_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i271_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n402));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i271_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i226_2_lut (.I0(\Kp[4] ), .I1(n1[14]), .I2(GND_net), 
            .I3(GND_net), .O(n335));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i226_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i320_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n475));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i320_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4955_5 (.CI(n39716), .I0(n12180[2]), .I1(n296), .CO(n39717));
    SB_LUT4 unary_minus_16_inv_0_i10_1_lut (.I0(PWMLimit[9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5235[9]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i275_2_lut (.I0(\Kp[5] ), .I1(n1[14]), .I2(GND_net), 
            .I3(GND_net), .O(n408));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i275_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_add_3_5_lut (.I0(\PID_CONTROLLER.integral [3]), 
            .I1(GND_net), .I2(n1_adj_5234[3]), .I3(n38732), .O(n7)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_5_lut.LUT_INIT = 16'h6996;
    SB_CARRY unary_minus_5_add_3_5 (.CI(n38732), .I0(GND_net), .I1(n1_adj_5234[3]), 
            .CO(n38733));
    SB_LUT4 mult_11_i369_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n548));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i369_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i469_2_lut (.I0(\Kp[9] ), .I1(n1[13]), .I2(GND_net), 
            .I3(GND_net), .O(n697));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i469_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5216_14_lut (.I0(GND_net), .I1(n17024[11]), .I2(n974), 
            .I3(n39582), .O(n16544[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5216_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i418_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n621));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i418_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i324_2_lut (.I0(\Kp[6] ), .I1(n1[14]), .I2(GND_net), 
            .I3(GND_net), .O(n481));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i324_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i120_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n177));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i120_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i467_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n694));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i467_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i11_1_lut (.I0(PWMLimit[10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5235[10]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i516_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n767));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i516_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i65_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n95));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i65_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i18_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n26));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i18_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i565_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n840));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i565_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i518_2_lut (.I0(\Kp[10] ), .I1(n1[13]), .I2(GND_net), 
            .I3(GND_net), .O(n770));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i518_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i373_2_lut (.I0(\Kp[7] ), .I1(n1[14]), .I2(GND_net), 
            .I3(GND_net), .O(n554));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i373_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i422_2_lut (.I0(\Kp[8] ), .I1(n1[14]), .I2(GND_net), 
            .I3(GND_net), .O(n627));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i422_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i110_2_lut (.I0(\Kp[2] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n162));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i110_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i159_2_lut (.I0(\Kp[3] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n235));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i159_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i12_1_lut (.I0(PWMLimit[11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5235[11]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i208_2_lut (.I0(\Kp[4] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n308));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i208_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i471_2_lut (.I0(\Kp[9] ), .I1(n1[14]), .I2(GND_net), 
            .I3(GND_net), .O(n700));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i471_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i257_2_lut (.I0(\Kp[5] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n381));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i257_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i306_2_lut (.I0(\Kp[6] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n454));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i306_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i61_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n89_adj_4816));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i61_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i14_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n20_adj_4817));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i14_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i51_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n74));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i51_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i4_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n5));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i4_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i110_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n162_adj_4818));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i110_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i355_2_lut (.I0(\Kp[7] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n527));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i355_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i404_2_lut (.I0(\Kp[8] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n600));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i404_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i453_2_lut (.I0(\Kp[9] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n673));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i453_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i502_2_lut (.I0(\Kp[10] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n746));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i502_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_add_3_4_lut (.I0(\PID_CONTROLLER.integral [2]), 
            .I1(GND_net), .I2(n1_adj_5234[2]), .I3(n38731), .O(n5_adj_4819)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_4_lut.LUT_INIT = 16'h6996;
    SB_CARRY add_5216_14 (.CI(n39582), .I0(n17024[11]), .I1(n974), .CO(n39583));
    SB_LUT4 add_4955_4_lut (.I0(GND_net), .I1(n12180[1]), .I2(n223), .I3(n39715), 
            .O(n11163[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4955_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5216_13_lut (.I0(GND_net), .I1(n17024[10]), .I2(n901), 
            .I3(n39581), .O(n16544[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5216_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i551_2_lut (.I0(\Kp[11] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n819));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i551_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i600_2_lut (.I0(\Kp[12] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n892));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i600_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i100_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n147));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i100_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4955_4 (.CI(n39715), .I0(n12180[1]), .I1(n223), .CO(n39716));
    SB_CARRY add_5216_13 (.CI(n39581), .I0(n17024[10]), .I1(n901), .CO(n39582));
    SB_LUT4 add_5216_12_lut (.I0(GND_net), .I1(n17024[9]), .I2(n828), 
            .I3(n39580), .O(n16544[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5216_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i649_2_lut (.I0(\Kp[13] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n965));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i649_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i698_2_lut (.I0(\Kp[14] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n1038));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i698_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i747_2_lut (.I0(\Kp[15] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n1111));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i747_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i79_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [14]), 
            .I2(GND_net), .I3(GND_net), .O(n116_adj_4820));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i79_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i32_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [15]), 
            .I2(GND_net), .I3(GND_net), .O(n47_adj_4821));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i32_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i128_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [14]), 
            .I2(GND_net), .I3(GND_net), .O(n189_adj_4822));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i128_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i149_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n220));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i149_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i177_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [14]), 
            .I2(GND_net), .I3(GND_net), .O(n262_adj_4823));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i177_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i226_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [14]), 
            .I2(GND_net), .I3(GND_net), .O(n335_adj_4824));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i226_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i159_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n235_adj_4825));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i159_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i275_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [14]), 
            .I2(GND_net), .I3(GND_net), .O(n408_adj_4826));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i275_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i324_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [14]), 
            .I2(GND_net), .I3(GND_net), .O(n481_adj_4827));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i324_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i208_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n308_adj_4828));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i208_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i373_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [14]), 
            .I2(GND_net), .I3(GND_net), .O(n554_adj_4829));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i373_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i198_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n293));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i198_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i247_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n366));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i247_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i422_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [14]), 
            .I2(GND_net), .I3(GND_net), .O(n627_adj_4830));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i422_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i471_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [14]), 
            .I2(GND_net), .I3(GND_net), .O(n700_adj_4831));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i471_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i257_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n381_adj_4832));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i257_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i59_2_lut (.I0(\Kp[1] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n86));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i59_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i12_2_lut (.I0(\Kp[0] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n17));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i12_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i108_2_lut (.I0(\Kp[2] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n159));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i108_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i296_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n439));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i296_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i361_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n536));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i361_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i410_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n609));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i410_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i345_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n512));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i345_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i306_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n454_adj_4834));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i306_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i157_2_lut (.I0(\Kp[3] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n232));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i157_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i206_2_lut (.I0(\Kp[4] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n305));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i206_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i355_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n527_adj_4835));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i355_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i404_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n600_adj_4836));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i404_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i394_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n585));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i394_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i453_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n673_adj_4837));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i453_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i255_2_lut (.I0(\Kp[5] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n378));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i255_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i304_2_lut (.I0(\Kp[6] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n451));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i304_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i353_2_lut (.I0(\Kp[7] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n524));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i353_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i402_2_lut (.I0(\Kp[8] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n597));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i402_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i451_2_lut (.I0(\Kp[9] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n670));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i451_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i500_2_lut (.I0(\Kp[10] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n743));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i500_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i549_2_lut (.I0(\Kp[11] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n816));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i549_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i443_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n658));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i443_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i502_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n746_adj_4838));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i502_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i598_2_lut (.I0(\Kp[12] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n889));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i598_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i551_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n819_adj_4839));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i551_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i600_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n892_adj_4840));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i600_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i647_2_lut (.I0(\Kp[13] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n962));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i647_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i696_2_lut (.I0(\Kp[14] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n1035));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i696_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i649_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n965_adj_4841));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i649_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i745_2_lut (.I0(\Kp[15] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n1108));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i745_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i492_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n731));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i492_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i698_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n1038_adj_4842));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i698_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i541_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n804));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i541_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5216_12 (.CI(n39580), .I0(n17024[9]), .I1(n828), .CO(n39581));
    SB_CARRY unary_minus_5_add_3_4 (.CI(n38731), .I0(GND_net), .I1(n1_adj_5234[2]), 
            .CO(n38732));
    SB_LUT4 unary_minus_5_add_3_3_lut (.I0(\PID_CONTROLLER.integral [1]), 
            .I1(GND_net), .I2(n1_adj_5234[1]), .I3(n38730), .O(n3)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_3_lut.LUT_INIT = 16'h6996;
    SB_LUT4 mult_10_i57_2_lut (.I0(\Kp[1] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n83));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i57_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i10_2_lut (.I0(\Kp[0] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n14_adj_4844));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i10_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i106_2_lut (.I0(\Kp[2] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n156));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i106_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i747_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n1111_adj_4845));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i747_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i590_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n877));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i590_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i155_2_lut (.I0(\Kp[3] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n229));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i155_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i204_2_lut (.I0(\Kp[4] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n302));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i204_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i253_2_lut (.I0(\Kp[5] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n375));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i253_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i302_2_lut (.I0(\Kp[6] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n448));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i302_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i59_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n86_adj_4846));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i59_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i12_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_4847));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i12_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i351_2_lut (.I0(\Kp[7] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n521));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i351_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5216_11_lut (.I0(GND_net), .I1(n17024[8]), .I2(n755), 
            .I3(n39579), .O(n16544[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5216_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i108_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n159_adj_4848));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i108_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i249_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n369));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i249_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i704_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n1047));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i704_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i157_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n232_adj_4849));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i157_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i639_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n950));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i639_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i6_1_lut (.I0(IntegralLimit[5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5234[5]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i206_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n305_adj_4851));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i206_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i255_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n378_adj_4852));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i255_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i753_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n1120));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i753_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i7_1_lut (.I0(IntegralLimit[6]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5234[6]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i298_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n442));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i298_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i400_2_lut (.I0(\Kp[8] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n594));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i400_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i449_2_lut (.I0(\Kp[9] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n667));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i449_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i8_1_lut (.I0(IntegralLimit[7]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5234[7]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i498_2_lut (.I0(\Kp[10] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n740));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i498_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i547_2_lut (.I0(\Kp[11] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n813));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i547_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i596_2_lut (.I0(\Kp[12] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n886));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i596_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i645_2_lut (.I0(\Kp[13] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n959));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i645_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i688_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n1023));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i688_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i347_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n515));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i347_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i9_1_lut (.I0(IntegralLimit[8]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5234[8]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i694_2_lut (.I0(\Kp[14] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n1032));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i694_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i169_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n250));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i169_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i743_2_lut (.I0(\Kp[15] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n1105));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i743_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i304_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n451_adj_4854));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i304_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i218_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n323));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i218_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i57_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n83_adj_4855));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i57_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i10_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n14_adj_4856));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i10_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i106_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n156_adj_4857));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i106_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i267_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n396));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i267_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i396_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n588));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i396_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i155_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n229_adj_4858));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i155_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i445_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n661));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i445_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i204_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n302_adj_4859));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i204_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i20918_2_lut (.I0(n1[11]), .I1(\PID_CONTROLLER.integral_23__N_3884 ), 
            .I2(GND_net), .I3(GND_net), .O(n4751[11]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i20918_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i737_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n1096));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i737_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i316_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n469));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i316_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4955_3_lut (.I0(GND_net), .I1(n12180[0]), .I2(n150), .I3(n39714), 
            .O(n11163[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4955_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5216_11 (.CI(n39579), .I0(n17024[8]), .I1(n755), .CO(n39580));
    SB_LUT4 mult_11_i365_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n542));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i365_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5216_10_lut (.I0(GND_net), .I1(n17024[7]), .I2(n682), 
            .I3(n39578), .O(n16544[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5216_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i253_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n375_adj_4861));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i253_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i302_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n448_adj_4862));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i302_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i494_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n734));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i494_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i10_1_lut (.I0(IntegralLimit[9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5234[9]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i20917_2_lut (.I0(n1[12]), .I1(\PID_CONTROLLER.integral_23__N_3884 ), 
            .I2(GND_net), .I3(GND_net), .O(n4751[12]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i20917_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i81_2_lut (.I0(\Kp[1] ), .I1(n1[15]), .I2(GND_net), 
            .I3(GND_net), .O(n119));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i81_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i414_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n615));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i414_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i34_2_lut (.I0(\Kp[0] ), .I1(n1[16]), .I2(GND_net), 
            .I3(GND_net), .O(n50));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i34_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i543_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n807));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i543_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i351_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n521_adj_4865));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i351_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i592_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n880));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i592_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i11_1_lut (.I0(IntegralLimit[10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5234[10]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i641_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n953));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i641_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i12_1_lut (.I0(IntegralLimit[11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5234[11]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i690_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n1026));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i690_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i13_1_lut (.I0(IntegralLimit[12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5234[12]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_5_inv_0_i14_1_lut (.I0(IntegralLimit[13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5234[13]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_4955_3 (.CI(n39714), .I0(n12180[0]), .I1(n150), .CO(n39715));
    SB_LUT4 add_4955_2_lut (.I0(GND_net), .I1(n8), .I2(n77), .I3(GND_net), 
            .O(n11163[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4955_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4955_2 (.CI(GND_net), .I0(n8), .I1(n77), .CO(n39714));
    SB_LUT4 add_5000_22_lut (.I0(GND_net), .I1(n13104[19]), .I2(GND_net), 
            .I3(n39713), .O(n12180[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5000_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_inv_0_i15_1_lut (.I0(IntegralLimit[14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5234[14]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_5216_10 (.CI(n39578), .I0(n17024[7]), .I1(n682), .CO(n39579));
    SB_LUT4 i20916_2_lut (.I0(n1[13]), .I1(\PID_CONTROLLER.integral_23__N_3884 ), 
            .I2(GND_net), .I3(GND_net), .O(n4751[13]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i20916_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i16_1_lut (.I0(IntegralLimit[15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5234[15]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i463_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n688));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i463_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i130_2_lut (.I0(\Kp[2] ), .I1(n1[15]), .I2(GND_net), 
            .I3(GND_net), .O(n192));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i130_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5216_9_lut (.I0(GND_net), .I1(n17024[6]), .I2(n609), .I3(n39577), 
            .O(n16544[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5216_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5000_21_lut (.I0(GND_net), .I1(n13104[18]), .I2(GND_net), 
            .I3(n39712), .O(n12180[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5000_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5000_21 (.CI(n39712), .I0(n13104[18]), .I1(GND_net), 
            .CO(n39713));
    SB_LUT4 mult_11_i512_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n761));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i512_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i739_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n1099));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i739_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i75_2_lut (.I0(\Kp[1] ), .I1(n1[12]), .I2(GND_net), 
            .I3(GND_net), .O(n110));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i75_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i17_1_lut (.I0(IntegralLimit[16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5234[16]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i28_2_lut (.I0(\Kp[0] ), .I1(n1[13]), .I2(GND_net), 
            .I3(GND_net), .O(n41));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i28_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5216_9 (.CI(n39577), .I0(n17024[6]), .I1(n609), .CO(n39578));
    SB_LUT4 add_5216_8_lut (.I0(GND_net), .I1(n17024[5]), .I2(n536), .I3(n39576), 
            .O(n16544[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5216_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5216_8 (.CI(n39576), .I0(n17024[5]), .I1(n536), .CO(n39577));
    SB_LUT4 mult_10_i124_2_lut (.I0(\Kp[2] ), .I1(n1[12]), .I2(GND_net), 
            .I3(GND_net), .O(n183));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i124_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5000_20_lut (.I0(GND_net), .I1(n13104[17]), .I2(GND_net), 
            .I3(n39711), .O(n12180[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5000_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_inv_0_i18_1_lut (.I0(IntegralLimit[17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5234[17]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i561_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n834));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i561_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5000_20 (.CI(n39711), .I0(n13104[17]), .I1(GND_net), 
            .CO(n39712));
    SB_LUT4 add_5000_19_lut (.I0(GND_net), .I1(n13104[16]), .I2(GND_net), 
            .I3(n39710), .O(n12180[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5000_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i173_2_lut (.I0(\Kp[3] ), .I1(n1[12]), .I2(GND_net), 
            .I3(GND_net), .O(n256_adj_4873));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i173_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i400_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n594_adj_4874));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i400_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i19_1_lut (.I0(IntegralLimit[18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5234[18]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i20915_2_lut (.I0(n1[14]), .I1(\PID_CONTROLLER.integral_23__N_3884 ), 
            .I2(GND_net), .I3(GND_net), .O(n4751[14]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i20915_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5216_7_lut (.I0(GND_net), .I1(n17024[4]), .I2(n463), .I3(n39575), 
            .O(n16544[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5216_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i20914_2_lut (.I0(n1[15]), .I1(\PID_CONTROLLER.integral_23__N_3884 ), 
            .I2(GND_net), .I3(GND_net), .O(n4751[15]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i20914_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i610_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n907));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i610_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i20_1_lut (.I0(IntegralLimit[19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5234[19]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i20913_2_lut (.I0(n1[16]), .I1(\PID_CONTROLLER.integral_23__N_3884 ), 
            .I2(GND_net), .I3(GND_net), .O(n4751[16]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i20913_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i21_1_lut (.I0(IntegralLimit[20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5234[20]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i179_2_lut (.I0(\Kp[3] ), .I1(n1[15]), .I2(GND_net), 
            .I3(GND_net), .O(n265));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i179_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i22_1_lut (.I0(IntegralLimit[21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5234[21]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i222_2_lut (.I0(\Kp[4] ), .I1(n1[12]), .I2(GND_net), 
            .I3(GND_net), .O(n329_adj_4877));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i222_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i23_1_lut (.I0(IntegralLimit[22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5234[22]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i659_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n980));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i659_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i449_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n667_adj_4879));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i449_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i83_2_lut (.I0(\Kp[1] ), .I1(n1[16]), .I2(GND_net), 
            .I3(GND_net), .O(n122));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i83_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i36_2_lut (.I0(\Kp[0] ), .I1(n1[17]), .I2(GND_net), 
            .I3(GND_net), .O(n53));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i36_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i271_2_lut (.I0(\Kp[5] ), .I1(n1[12]), .I2(GND_net), 
            .I3(GND_net), .O(n402_adj_4881));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i271_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i498_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n740_adj_4882));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i498_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i24_1_lut (.I0(IntegralLimit[23]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5234[23]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i132_2_lut (.I0(\Kp[2] ), .I1(n1[16]), .I2(GND_net), 
            .I3(GND_net), .O(n195));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i132_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i20912_2_lut (.I0(n1[17]), .I1(\PID_CONTROLLER.integral_23__N_3884 ), 
            .I2(GND_net), .I3(GND_net), .O(n4751[17]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i20912_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i1_1_lut (.I0(PWMLimit[0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5235[0]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i20911_2_lut (.I0(n1[18]), .I1(\PID_CONTROLLER.integral_23__N_3884 ), 
            .I2(GND_net), .I3(GND_net), .O(n4751[18]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i20911_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i2_1_lut (.I0(PWMLimit[1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5235[1]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i547_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n813_adj_4885));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i547_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i181_2_lut (.I0(\Kp[3] ), .I1(n1[16]), .I2(GND_net), 
            .I3(GND_net), .O(n268));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i181_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i53_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n77));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i53_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i6_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n8));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i6_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i20910_2_lut (.I0(n1[19]), .I1(\PID_CONTROLLER.integral_23__N_3884 ), 
            .I2(GND_net), .I3(GND_net), .O(n4751[19]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i20910_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i459_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n682));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i459_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i230_2_lut (.I0(\Kp[4] ), .I1(n1[16]), .I2(GND_net), 
            .I3(GND_net), .O(n341));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i230_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i102_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n150));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i102_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i279_2_lut (.I0(\Kp[5] ), .I1(n1[16]), .I2(GND_net), 
            .I3(GND_net), .O(n414));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i279_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i596_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n886_adj_4887));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i596_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i328_2_lut (.I0(\Kp[6] ), .I1(n1[16]), .I2(GND_net), 
            .I3(GND_net), .O(n487));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i328_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i645_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n959_adj_4888));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i645_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i228_2_lut (.I0(\Kp[4] ), .I1(n1[15]), .I2(GND_net), 
            .I3(GND_net), .O(n338));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i228_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i13_1_lut (.I0(PWMLimit[12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5235[12]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i694_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n1032_adj_4890));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i694_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i377_2_lut (.I0(\Kp[7] ), .I1(n1[16]), .I2(GND_net), 
            .I3(GND_net), .O(n560));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i377_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i743_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n1105_adj_4891));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i743_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i69_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n101));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i69_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i22_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n32));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i22_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i118_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n174));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i118_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i20909_2_lut (.I0(n1[20]), .I1(\PID_CONTROLLER.integral_23__N_3884 ), 
            .I2(GND_net), .I3(GND_net), .O(n4751[20]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i20909_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i3_1_lut (.I0(PWMLimit[2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5235[2]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i167_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n247));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i167_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i20908_2_lut (.I0(n1[21]), .I1(\PID_CONTROLLER.integral_23__N_3884 ), 
            .I2(GND_net), .I3(GND_net), .O(n4751[21]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i20908_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5000_19 (.CI(n39710), .I0(n13104[16]), .I1(GND_net), 
            .CO(n39711));
    SB_LUT4 mult_11_i216_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n320));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i216_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i265_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n393));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i265_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i55_2_lut (.I0(\Kp[1] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n80));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i55_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i4_1_lut (.I0(PWMLimit[3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5235[3]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i8_2_lut (.I0(\Kp[0] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n11_adj_4897));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i8_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i55_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n80_adj_4898));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i55_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i8_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_4899));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i8_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i20907_2_lut (.I0(n1[22]), .I1(\PID_CONTROLLER.integral_23__N_3884 ), 
            .I2(GND_net), .I3(GND_net), .O(n4751[22]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i20907_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i104_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n153));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i104_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i314_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n466));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i314_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i153_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n226));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i153_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i363_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n539));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i363_2_lut.LUT_INIT = 16'h8888;
    SB_DFF result_i0 (.Q(duty[0]), .C(clk32MHz), .D(duty_23__N_3812[0]));   // verilog/motorControl.v(29[14] 48[8])
    SB_LUT4 mult_11_i412_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n612));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i412_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i202_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n299));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i202_2_lut.LUT_INIT = 16'h8888;
    SB_DFF \PID_CONTROLLER.integral_i0  (.Q(\PID_CONTROLLER.integral [0]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3836 [0]));   // verilog/motorControl.v(29[14] 48[8])
    SB_LUT4 unary_minus_16_inv_0_i5_1_lut (.I0(PWMLimit[4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5235[4]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY unary_minus_5_add_3_3 (.CI(n38730), .I0(GND_net), .I1(n1_adj_5234[1]), 
            .CO(n38731));
    SB_LUT4 unary_minus_5_add_3_2_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5234[0]), 
            .I3(VCC_net), .O(\PID_CONTROLLER.integral_23__N_3887 [0])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_5_add_3_2 (.CI(VCC_net), .I0(GND_net), .I1(n1_adj_5234[0]), 
            .CO(n38730));
    SB_LUT4 sub_3_add_2_25_lut (.I0(GND_net), .I1(setpoint[23]), .I2(motor_state[23]), 
            .I3(n38729), .O(n1[23])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_3_add_2_24_lut (.I0(GND_net), .I1(setpoint[22]), .I2(motor_state[22]), 
            .I3(n38728), .O(n1[22])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_3_add_2_24 (.CI(n38728), .I0(setpoint[22]), .I1(motor_state[22]), 
            .CO(n38729));
    SB_LUT4 mult_10_i104_2_lut (.I0(\Kp[2] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n153_adj_4904));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i104_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 IntegralLimit_23__I_0_i17_2_lut (.I0(\PID_CONTROLLER.integral [8]), 
            .I1(IntegralLimit[8]), .I2(GND_net), .I3(GND_net), .O(n17_adj_4905));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 IntegralLimit_23__I_0_i9_2_lut (.I0(\PID_CONTROLLER.integral [4]), 
            .I1(IntegralLimit[4]), .I2(GND_net), .I3(GND_net), .O(n9_adj_4906));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 IntegralLimit_23__I_0_i11_2_lut (.I0(\PID_CONTROLLER.integral [5]), 
            .I1(IntegralLimit[5]), .I2(GND_net), .I3(GND_net), .O(n11_adj_4907));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 sub_3_add_2_23_lut (.I0(GND_net), .I1(setpoint[21]), .I2(motor_state[21]), 
            .I3(n38727), .O(n1[21])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i34066_4_lut (.I0(\PID_CONTROLLER.integral [3]), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(IntegralLimit[3]), .I3(IntegralLimit[2]), .O(n49653));
    defparam i34066_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 i34064_3_lut (.I0(n11_adj_4907), .I1(n9_adj_4906), .I2(n49653), 
            .I3(GND_net), .O(n49651));
    defparam i34064_3_lut.LUT_INIT = 16'habab;
    SB_LUT4 mult_10_i153_2_lut (.I0(\Kp[3] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n226_adj_4908));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i153_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 IntegralLimit_23__I_0_i13_rep_267_2_lut (.I0(\PID_CONTROLLER.integral [6]), 
            .I1(IntegralLimit[6]), .I2(GND_net), .I3(GND_net), .O(n51808));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i13_rep_267_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i34590_4_lut (.I0(\PID_CONTROLLER.integral [7]), .I1(n51808), 
            .I2(IntegralLimit[7]), .I3(n49651), .O(n50178));
    defparam i34590_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 i34371_4_lut (.I0(\PID_CONTROLLER.integral [9]), .I1(n17_adj_4905), 
            .I2(IntegralLimit[9]), .I3(n50178), .O(n49959));
    defparam i34371_4_lut.LUT_INIT = 16'hdeff;
    SB_CARRY sub_3_add_2_23 (.CI(n38727), .I0(setpoint[21]), .I1(motor_state[21]), 
            .CO(n38728));
    SB_LUT4 IntegralLimit_23__I_0_i21_rep_249_2_lut (.I0(\PID_CONTROLLER.integral [10]), 
            .I1(IntegralLimit[10]), .I2(GND_net), .I3(GND_net), .O(n51790));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i21_rep_249_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i34369_4_lut (.I0(\PID_CONTROLLER.integral [9]), .I1(n17_adj_4905), 
            .I2(IntegralLimit[9]), .I3(n9_adj_4906), .O(n49957));
    defparam i34369_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 add_5000_18_lut (.I0(GND_net), .I1(n13104[15]), .I2(GND_net), 
            .I3(n39709), .O(n12180[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5000_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i34367_4_lut (.I0(\PID_CONTROLLER.integral [11]), .I1(n51790), 
            .I2(IntegralLimit[11]), .I3(n49957), .O(n49955));
    defparam i34367_4_lut.LUT_INIT = 16'hdeff;
    SB_LUT4 sub_3_add_2_22_lut (.I0(GND_net), .I1(setpoint[20]), .I2(motor_state[20]), 
            .I3(n38726), .O(n1[20])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 IntegralLimit_23__I_0_i25_rep_243_2_lut (.I0(\PID_CONTROLLER.integral [12]), 
            .I1(IntegralLimit[12]), .I2(GND_net), .I3(GND_net), .O(n51784));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i25_rep_243_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i34013_4_lut (.I0(n27), .I1(n15_adj_4909), .I2(n13_adj_4910), 
            .I3(n11_adj_4911), .O(n49600));
    defparam i34013_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i34019_4_lut (.I0(n21_adj_4912), .I1(n19_adj_4913), .I2(n17_adj_4914), 
            .I3(n9_adj_4915), .O(n49606));
    defparam i34019_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 \PID_CONTROLLER.integral_23__I_0_i16_3_lut  (.I0(\PID_CONTROLLER.integral [9]), 
            .I1(\PID_CONTROLLER.integral [21]), .I2(n43), .I3(GND_net), 
            .O(n16_adj_4916));   // verilog/motorControl.v(31[38:63])
    defparam \PID_CONTROLLER.integral_23__I_0_i16_3_lut .LUT_INIT = 16'hcaca;
    SB_LUT4 i33996_2_lut (.I0(n43), .I1(n19_adj_4913), .I2(GND_net), .I3(GND_net), 
            .O(n49583));
    defparam i33996_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 mult_10_i277_2_lut (.I0(\Kp[5] ), .I1(n1[15]), .I2(GND_net), 
            .I3(GND_net), .O(n411));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i277_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5216_7 (.CI(n39575), .I0(n17024[4]), .I1(n463), .CO(n39576));
    SB_LUT4 \PID_CONTROLLER.integral_23__I_0_i8_3_lut  (.I0(\PID_CONTROLLER.integral [4]), 
            .I1(\PID_CONTROLLER.integral [8]), .I2(n17_adj_4914), .I3(GND_net), 
            .O(n8_adj_4917));   // verilog/motorControl.v(31[38:63])
    defparam \PID_CONTROLLER.integral_23__I_0_i8_3_lut .LUT_INIT = 16'hcaca;
    SB_LUT4 \PID_CONTROLLER.integral_23__I_0_i24_3_lut  (.I0(n16_adj_4916), 
            .I1(\PID_CONTROLLER.integral [22]), .I2(n45), .I3(GND_net), 
            .O(n24_adj_4918));   // verilog/motorControl.v(31[38:63])
    defparam \PID_CONTROLLER.integral_23__I_0_i24_3_lut .LUT_INIT = 16'hcaca;
    SB_CARRY add_5000_18 (.CI(n39709), .I0(n13104[15]), .I1(GND_net), 
            .CO(n39710));
    SB_LUT4 mult_10_i202_2_lut (.I0(\Kp[4] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n299_adj_4919));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i202_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i34032_2_lut (.I0(n7), .I1(n5_adj_4819), .I2(GND_net), .I3(GND_net), 
            .O(n49619));
    defparam i34032_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i34343_4_lut (.I0(n13_adj_4910), .I1(n11_adj_4911), .I2(n9_adj_4915), 
            .I3(n49619), .O(n49931));
    defparam i34343_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i34339_4_lut (.I0(n19_adj_4913), .I1(n17_adj_4914), .I2(n15_adj_4909), 
            .I3(n49931), .O(n49927));
    defparam i34339_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i34766_4_lut (.I0(n25_adj_4920), .I1(n23_adj_4921), .I2(n21_adj_4912), 
            .I3(n49927), .O(n50354));
    defparam i34766_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 unary_minus_16_inv_0_i6_1_lut (.I0(PWMLimit[5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5235[5]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i251_2_lut (.I0(\Kp[5] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n372));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i251_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i34564_4_lut (.I0(n31), .I1(n29), .I2(n27), .I3(n50354), 
            .O(n50152));
    defparam i34564_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i34828_4_lut (.I0(n37), .I1(n35), .I2(n33), .I3(n50152), 
            .O(n50416));
    defparam i34828_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i34373_4_lut (.I0(\PID_CONTROLLER.integral [7]), .I1(n51808), 
            .I2(IntegralLimit[7]), .I3(n11_adj_4907), .O(n49961));
    defparam i34373_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 mult_11_i353_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n524_adj_4923));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i353_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 IntegralLimit_23__I_0_i27_rep_236_2_lut (.I0(\PID_CONTROLLER.integral [13]), 
            .I1(IntegralLimit[13]), .I2(GND_net), .I3(GND_net), .O(n51777));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i27_rep_236_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i34361_4_lut (.I0(\PID_CONTROLLER.integral [14]), .I1(n51777), 
            .I2(IntegralLimit[14]), .I3(n49961), .O(n49949));
    defparam i34361_4_lut.LUT_INIT = 16'hdeff;
    SB_LUT4 IntegralLimit_23__I_0_i31_rep_231_2_lut (.I0(\PID_CONTROLLER.integral [15]), 
            .I1(IntegralLimit[15]), .I2(GND_net), .I3(GND_net), .O(n51772));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i31_rep_231_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 IntegralLimit_23__I_0_i12_3_lut (.I0(IntegralLimit[7]), .I1(IntegralLimit[16]), 
            .I2(\PID_CONTROLLER.integral [16]), .I3(GND_net), .O(n12_adj_4924));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i12_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i34044_4_lut (.I0(\PID_CONTROLLER.integral [16]), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(IntegralLimit[16]), .I3(IntegralLimit[7]), .O(n49631));
    defparam i34044_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 IntegralLimit_23__I_0_i35_rep_254_2_lut (.I0(\PID_CONTROLLER.integral [17]), 
            .I1(IntegralLimit[17]), .I2(GND_net), .I3(GND_net), .O(n51795));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i35_rep_254_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 IntegralLimit_23__I_0_i10_3_lut (.I0(IntegralLimit[5]), .I1(IntegralLimit[6]), 
            .I2(\PID_CONTROLLER.integral [6]), .I3(GND_net), .O(n10_adj_4925));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i10_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 IntegralLimit_23__I_0_i30_3_lut (.I0(n12_adj_4924), .I1(IntegralLimit[17]), 
            .I2(\PID_CONTROLLER.integral [17]), .I3(GND_net), .O(n30));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i30_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i34712_4_lut (.I0(\PID_CONTROLLER.integral [11]), .I1(n51790), 
            .I2(IntegralLimit[11]), .I3(n49959), .O(n50300));
    defparam i34712_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 unary_minus_16_inv_0_i14_1_lut (.I0(PWMLimit[13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5235[13]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i34052_4_lut (.I0(\PID_CONTROLLER.integral [13]), .I1(n51784), 
            .I2(IntegralLimit[13]), .I3(n50300), .O(n49639));
    defparam i34052_4_lut.LUT_INIT = 16'h5a7b;
    SB_LUT4 IntegralLimit_23__I_0_i29_rep_234_2_lut (.I0(\PID_CONTROLLER.integral [14]), 
            .I1(IntegralLimit[14]), .I2(GND_net), .I3(GND_net), .O(n51775));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i29_rep_234_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_10_i300_2_lut (.I0(\Kp[6] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n445));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i300_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i349_2_lut (.I0(\Kp[7] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n518));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i349_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i398_2_lut (.I0(\Kp[8] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n591));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i398_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i447_2_lut (.I0(\Kp[9] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n664));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i447_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i34584_4_lut (.I0(\PID_CONTROLLER.integral [15]), .I1(n51775), 
            .I2(IntegralLimit[15]), .I3(n49639), .O(n50172));
    defparam i34584_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 IntegralLimit_23__I_0_i33_rep_260_2_lut (.I0(\PID_CONTROLLER.integral [16]), 
            .I1(IntegralLimit[16]), .I2(GND_net), .I3(GND_net), .O(n51801));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i33_rep_260_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_5216_6_lut (.I0(GND_net), .I1(n17024[3]), .I2(n390), .I3(n39574), 
            .O(n16544[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5216_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i34772_4_lut (.I0(\PID_CONTROLLER.integral [17]), .I1(n51801), 
            .I2(IntegralLimit[17]), .I3(n50172), .O(n50360));
    defparam i34772_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 IntegralLimit_23__I_0_i37_rep_225_2_lut (.I0(\PID_CONTROLLER.integral [18]), 
            .I1(IntegralLimit[18]), .I2(GND_net), .I3(GND_net), .O(n51766));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i37_rep_225_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_5216_6 (.CI(n39574), .I0(n17024[3]), .I1(n390), .CO(n39575));
    SB_LUT4 add_5216_5_lut (.I0(GND_net), .I1(n17024[2]), .I2(n317), .I3(n39573), 
            .O(n16544[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5216_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5216_5 (.CI(n39573), .I0(n17024[2]), .I1(n317), .CO(n39574));
    SB_LUT4 add_5216_4_lut (.I0(GND_net), .I1(n17024[1]), .I2(n244), .I3(n39572), 
            .O(n16544[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5216_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5216_4 (.CI(n39572), .I0(n17024[1]), .I1(n244), .CO(n39573));
    SB_LUT4 add_5216_3_lut (.I0(GND_net), .I1(n17024[0]), .I2(n171), .I3(n39571), 
            .O(n16544[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5216_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5216_3 (.CI(n39571), .I0(n17024[0]), .I1(n171), .CO(n39572));
    SB_LUT4 add_5216_2_lut (.I0(GND_net), .I1(n29_adj_4927), .I2(n98), 
            .I3(GND_net), .O(n16544[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5216_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i34858_4_lut (.I0(\PID_CONTROLLER.integral [19]), .I1(n51766), 
            .I2(IntegralLimit[19]), .I3(n50360), .O(n50446));
    defparam i34858_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 IntegralLimit_23__I_0_i41_rep_222_2_lut (.I0(\PID_CONTROLLER.integral [20]), 
            .I1(IntegralLimit[20]), .I2(GND_net), .I3(GND_net), .O(n51763));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i41_rep_222_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY sub_3_add_2_22 (.CI(n38726), .I0(setpoint[20]), .I1(motor_state[20]), 
            .CO(n38727));
    SB_CARRY add_5216_2 (.CI(GND_net), .I0(n29_adj_4927), .I1(n98), .CO(n39571));
    SB_LUT4 IntegralLimit_23__I_0_i16_3_lut (.I0(IntegralLimit[9]), .I1(IntegralLimit[21]), 
            .I2(\PID_CONTROLLER.integral [21]), .I3(GND_net), .O(n16_adj_4928));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i16_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 add_5245_15_lut (.I0(GND_net), .I1(n17444[12]), .I2(n1050), 
            .I3(n39570), .O(n17024[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5245_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5000_17_lut (.I0(GND_net), .I1(n13104[14]), .I2(GND_net), 
            .I3(n39708), .O(n12180[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5000_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i34034_4_lut (.I0(\PID_CONTROLLER.integral [21]), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(IntegralLimit[21]), .I3(IntegralLimit[9]), .O(n49621));
    defparam i34034_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 mult_10_i496_2_lut (.I0(\Kp[10] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n737));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i496_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 sub_3_add_2_21_lut (.I0(GND_net), .I1(setpoint[19]), .I2(motor_state[19]), 
            .I3(n38725), .O(n1[19])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i545_2_lut (.I0(\Kp[11] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n810));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i545_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i594_2_lut (.I0(\Kp[12] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n883));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i594_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i643_2_lut (.I0(\Kp[13] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n956));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i643_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i692_2_lut (.I0(\Kp[14] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n1029));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i692_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 IntegralLimit_23__I_0_i24_3_lut (.I0(n16_adj_4928), .I1(IntegralLimit[22]), 
            .I2(\PID_CONTROLLER.integral [22]), .I3(GND_net), .O(n24_adj_4929));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i24_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 IntegralLimit_23__I_0_i6_3_lut (.I0(IntegralLimit[2]), .I1(IntegralLimit[3]), 
            .I2(\PID_CONTROLLER.integral [3]), .I3(GND_net), .O(n6_adj_4930));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i6_3_lut.LUT_INIT = 16'h8e8e;
    SB_CARRY add_5000_17 (.CI(n39708), .I0(n13104[14]), .I1(GND_net), 
            .CO(n39709));
    SB_LUT4 mult_10_i741_2_lut (.I0(\Kp[15] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n1102));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i741_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i34658_3_lut (.I0(n6_adj_4930), .I1(IntegralLimit[10]), .I2(\PID_CONTROLLER.integral [10]), 
            .I3(GND_net), .O(n50246));   // verilog/motorControl.v(31[10:34])
    defparam i34658_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 mult_10_i53_2_lut (.I0(\Kp[1] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n77_adj_4932));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i53_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i6_2_lut (.I0(\Kp[0] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n8_adj_4933));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i6_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i34659_3_lut (.I0(n50246), .I1(IntegralLimit[11]), .I2(\PID_CONTROLLER.integral [11]), 
            .I3(GND_net), .O(n50247));   // verilog/motorControl.v(31[10:34])
    defparam i34659_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 mult_10_i102_2_lut (.I0(\Kp[2] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n150_adj_4934));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i102_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5000_16_lut (.I0(GND_net), .I1(n13104[13]), .I2(n1102_adj_4935), 
            .I3(n39707), .O(n12180[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5000_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5000_16 (.CI(n39707), .I0(n13104[13]), .I1(n1102_adj_4935), 
            .CO(n39708));
    SB_LUT4 add_5000_15_lut (.I0(GND_net), .I1(n13104[12]), .I2(n1029_adj_4936), 
            .I3(n39706), .O(n12180[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5000_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5000_15 (.CI(n39706), .I0(n13104[12]), .I1(n1029_adj_4936), 
            .CO(n39707));
    SB_LUT4 add_5000_14_lut (.I0(GND_net), .I1(n13104[11]), .I2(n956_adj_4937), 
            .I3(n39705), .O(n12180[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5000_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i34036_4_lut (.I0(\PID_CONTROLLER.integral [21]), .I1(n51784), 
            .I2(IntegralLimit[21]), .I3(n49955), .O(n49623));
    defparam i34036_4_lut.LUT_INIT = 16'h5a7b;
    SB_LUT4 mult_10_i151_2_lut (.I0(\Kp[3] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n223_adj_4938));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i151_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5000_14 (.CI(n39705), .I0(n13104[11]), .I1(n956_adj_4937), 
            .CO(n39706));
    SB_LUT4 mult_10_i200_2_lut (.I0(\Kp[4] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n296_adj_4939));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i200_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5245_14_lut (.I0(GND_net), .I1(n17444[11]), .I2(n977), 
            .I3(n39569), .O(n17024[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5245_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5000_13_lut (.I0(GND_net), .I1(n13104[10]), .I2(n883_adj_4940), 
            .I3(n39704), .O(n12180[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5000_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i34660_4_lut (.I0(n24_adj_4929), .I1(n8_adj_4941), .I2(n51761), 
            .I3(n49621), .O(n50248));   // verilog/motorControl.v(31[10:34])
    defparam i34660_4_lut.LUT_INIT = 16'haaac;
    SB_CARRY sub_3_add_2_21 (.CI(n38725), .I0(setpoint[19]), .I1(motor_state[19]), 
            .CO(n38726));
    SB_LUT4 mult_10_i249_2_lut (.I0(\Kp[5] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n369_adj_4942));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i249_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i298_2_lut (.I0(\Kp[6] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n442_adj_4943));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i298_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i34176_3_lut (.I0(n50247), .I1(IntegralLimit[12]), .I2(\PID_CONTROLLER.integral [12]), 
            .I3(GND_net), .O(n49764));   // verilog/motorControl.v(31[10:34])
    defparam i34176_3_lut.LUT_INIT = 16'h8e8e;
    SB_CARRY add_5000_13 (.CI(n39704), .I0(n13104[10]), .I1(n883_adj_4940), 
            .CO(n39705));
    SB_LUT4 mult_10_i347_2_lut (.I0(\Kp[7] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n515_adj_4944));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i347_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 \PID_CONTROLLER.integral_23__I_0_i4_4_lut  (.I0(\PID_CONTROLLER.integral_23__N_3887 [0]), 
            .I1(\PID_CONTROLLER.integral [1]), .I2(n3), .I3(\PID_CONTROLLER.integral [0]), 
            .O(n4_adj_4945));   // verilog/motorControl.v(31[38:63])
    defparam \PID_CONTROLLER.integral_23__I_0_i4_4_lut .LUT_INIT = 16'hc5c0;
    SB_LUT4 mult_10_i396_2_lut (.I0(\Kp[8] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n588_adj_4946));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i396_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i34686_3_lut (.I0(n4_adj_4945), .I1(\PID_CONTROLLER.integral [13]), 
            .I2(n27), .I3(GND_net), .O(n50274));   // verilog/motorControl.v(31[38:63])
    defparam i34686_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34687_3_lut (.I0(n50274), .I1(\PID_CONTROLLER.integral [14]), 
            .I2(n29), .I3(GND_net), .O(n50275));   // verilog/motorControl.v(31[38:63])
    defparam i34687_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_10_i445_2_lut (.I0(\Kp[9] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n661_adj_4947));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i445_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i7_1_lut (.I0(PWMLimit[6]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5235[6]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 \PID_CONTROLLER.integral_23__I_0_i12_3_lut  (.I0(\PID_CONTROLLER.integral [7]), 
            .I1(\PID_CONTROLLER.integral [16]), .I2(n33), .I3(GND_net), 
            .O(n12_adj_4949));   // verilog/motorControl.v(31[38:63])
    defparam \PID_CONTROLLER.integral_23__I_0_i12_3_lut .LUT_INIT = 16'hcaca;
    SB_LUT4 i34007_2_lut (.I0(n33), .I1(n15_adj_4909), .I2(GND_net), .I3(GND_net), 
            .O(n49594));
    defparam i34007_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 \PID_CONTROLLER.integral_23__I_0_i10_3_lut  (.I0(\PID_CONTROLLER.integral [5]), 
            .I1(\PID_CONTROLLER.integral [6]), .I2(n13_adj_4910), .I3(GND_net), 
            .O(n10_adj_4950));   // verilog/motorControl.v(31[38:63])
    defparam \PID_CONTROLLER.integral_23__I_0_i10_3_lut .LUT_INIT = 16'hcaca;
    SB_CARRY add_5245_14 (.CI(n39569), .I0(n17444[11]), .I1(n977), .CO(n39570));
    SB_LUT4 mult_10_i494_2_lut (.I0(\Kp[10] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n734_adj_4951));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i494_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i543_2_lut (.I0(\Kp[11] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n807_adj_4952));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i543_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 \PID_CONTROLLER.integral_23__I_0_i30_3_lut  (.I0(n12_adj_4949), 
            .I1(\PID_CONTROLLER.integral [17]), .I2(n35), .I3(GND_net), 
            .O(n30_adj_4953));   // verilog/motorControl.v(31[38:63])
    defparam \PID_CONTROLLER.integral_23__I_0_i30_3_lut .LUT_INIT = 16'hcaca;
    SB_LUT4 i34009_4_lut (.I0(n33), .I1(n31), .I2(n29), .I3(n49600), 
            .O(n49596));
    defparam i34009_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i34794_4_lut (.I0(n30_adj_4953), .I1(n10_adj_4950), .I2(n35), 
            .I3(n49594), .O(n50382));   // verilog/motorControl.v(31[38:63])
    defparam i34794_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i34188_3_lut (.I0(n50275), .I1(\PID_CONTROLLER.integral [15]), 
            .I2(n31), .I3(GND_net), .O(n49776));   // verilog/motorControl.v(31[38:63])
    defparam i34188_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34872_4_lut (.I0(n49776), .I1(n50382), .I2(n35), .I3(n49596), 
            .O(n50460));   // verilog/motorControl.v(31[38:63])
    defparam i34872_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i34873_3_lut (.I0(n50460), .I1(\PID_CONTROLLER.integral [18]), 
            .I2(n37), .I3(GND_net), .O(n50461));   // verilog/motorControl.v(31[38:63])
    defparam i34873_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_5245_13_lut (.I0(GND_net), .I1(n17444[10]), .I2(n904), 
            .I3(n39568), .O(n17024[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5245_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_3_add_2_20_lut (.I0(GND_net), .I1(setpoint[18]), .I2(motor_state[18]), 
            .I3(n38724), .O(n1[18])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i34851_3_lut (.I0(n50461), .I1(\PID_CONTROLLER.integral [19]), 
            .I2(n39), .I3(GND_net), .O(n50439));   // verilog/motorControl.v(31[38:63])
    defparam i34851_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 \PID_CONTROLLER.integral_23__I_0_i6_3_lut  (.I0(\PID_CONTROLLER.integral [2]), 
            .I1(\PID_CONTROLLER.integral [3]), .I2(n7), .I3(GND_net), 
            .O(n6_adj_4954));   // verilog/motorControl.v(31[38:63])
    defparam \PID_CONTROLLER.integral_23__I_0_i6_3_lut .LUT_INIT = 16'hcaca;
    SB_LUT4 mult_10_i592_2_lut (.I0(\Kp[12] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n880_adj_4955));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i592_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5245_13 (.CI(n39568), .I0(n17444[10]), .I1(n904), .CO(n39569));
    SB_LUT4 unary_minus_16_inv_0_i15_1_lut (.I0(PWMLimit[14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5235[14]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i641_2_lut (.I0(\Kp[13] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n953_adj_4957));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i641_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i690_2_lut (.I0(\Kp[14] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n1026_adj_4958));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i690_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5000_12_lut (.I0(GND_net), .I1(n13104[9]), .I2(n810_adj_4959), 
            .I3(n39703), .O(n12180[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5000_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5000_12 (.CI(n39703), .I0(n13104[9]), .I1(n810_adj_4959), 
            .CO(n39704));
    SB_LUT4 add_5000_11_lut (.I0(GND_net), .I1(n13104[8]), .I2(n737_adj_4960), 
            .I3(n39702), .O(n12180[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5000_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5245_12_lut (.I0(GND_net), .I1(n17444[9]), .I2(n831), 
            .I3(n39567), .O(n17024[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5245_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5245_12 (.CI(n39567), .I0(n17444[9]), .I1(n831), .CO(n39568));
    SB_LUT4 mult_10_i739_2_lut (.I0(\Kp[15] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n1099_adj_4961));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i739_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY sub_3_add_2_20 (.CI(n38724), .I0(setpoint[18]), .I1(motor_state[18]), 
            .CO(n38725));
    SB_LUT4 i34690_3_lut (.I0(n6_adj_4954), .I1(\PID_CONTROLLER.integral [10]), 
            .I2(n21_adj_4912), .I3(GND_net), .O(n50278));   // verilog/motorControl.v(31[38:63])
    defparam i34690_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34691_3_lut (.I0(n50278), .I1(\PID_CONTROLLER.integral [11]), 
            .I2(n23_adj_4921), .I3(GND_net), .O(n50279));   // verilog/motorControl.v(31[38:63])
    defparam i34691_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i33998_4_lut (.I0(n43), .I1(n25_adj_4920), .I2(n23_adj_4921), 
            .I3(n49606), .O(n49585));
    defparam i33998_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i34662_4_lut (.I0(n24_adj_4918), .I1(n8_adj_4917), .I2(n45), 
            .I3(n49583), .O(n50250));   // verilog/motorControl.v(31[38:63])
    defparam i34662_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i34186_3_lut (.I0(n50279), .I1(\PID_CONTROLLER.integral [12]), 
            .I2(n25_adj_4920), .I3(GND_net), .O(n49774));   // verilog/motorControl.v(31[38:63])
    defparam i34186_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34000_4_lut (.I0(n43), .I1(n41_adj_4962), .I2(n39), .I3(n50416), 
            .O(n49587));
    defparam i34000_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 mult_10_i51_2_lut (.I0(\Kp[1] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n74_adj_4964));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i51_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 sub_3_add_2_19_lut (.I0(GND_net), .I1(setpoint[17]), .I2(motor_state[17]), 
            .I3(n38723), .O(n1[17])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i4_2_lut (.I0(\Kp[0] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n5_adj_4965));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i4_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i100_2_lut (.I0(\Kp[2] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n147_adj_4966));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i100_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5000_11 (.CI(n39702), .I0(n13104[8]), .I1(n737_adj_4960), 
            .CO(n39703));
    SB_LUT4 mult_10_i326_2_lut (.I0(\Kp[6] ), .I1(n1[15]), .I2(GND_net), 
            .I3(GND_net), .O(n484));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i326_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i34808_4_lut (.I0(n49774), .I1(n50250), .I2(n45), .I3(n49585), 
            .O(n50396));   // verilog/motorControl.v(31[38:63])
    defparam i34808_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 mult_10_i149_2_lut (.I0(\Kp[3] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n220_adj_4967));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i149_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i198_2_lut (.I0(\Kp[4] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n293_adj_4968));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i198_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5000_10_lut (.I0(GND_net), .I1(n13104[7]), .I2(n664_adj_4969), 
            .I3(n39701), .O(n12180[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5000_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5245_11_lut (.I0(GND_net), .I1(n17444[8]), .I2(n758), 
            .I3(n39566), .O(n17024[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5245_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5245_11 (.CI(n39566), .I0(n17444[8]), .I1(n758), .CO(n39567));
    SB_LUT4 i34194_3_lut (.I0(n50439), .I1(\PID_CONTROLLER.integral [20]), 
            .I2(n41_adj_4962), .I3(GND_net), .O(n49782));   // verilog/motorControl.v(31[38:63])
    defparam i34194_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34810_4_lut (.I0(n49782), .I1(n50396), .I2(n45), .I3(n49587), 
            .O(n50398));   // verilog/motorControl.v(31[38:63])
    defparam i34810_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 IntegralLimit_23__I_0_i4_4_lut (.I0(\PID_CONTROLLER.integral [0]), 
            .I1(IntegralLimit[1]), .I2(\PID_CONTROLLER.integral [1]), .I3(IntegralLimit[0]), 
            .O(n4_adj_4970));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i4_4_lut.LUT_INIT = 16'h4d0c;
    SB_LUT4 i34696_3_lut (.I0(n4_adj_4970), .I1(IntegralLimit[13]), .I2(\PID_CONTROLLER.integral [13]), 
            .I3(GND_net), .O(n50284));   // verilog/motorControl.v(31[10:34])
    defparam i34696_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i34697_3_lut (.I0(n50284), .I1(IntegralLimit[14]), .I2(\PID_CONTROLLER.integral [14]), 
            .I3(GND_net), .O(n50285));   // verilog/motorControl.v(31[10:34])
    defparam i34697_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i34046_4_lut (.I0(\PID_CONTROLLER.integral [16]), .I1(n51772), 
            .I2(IntegralLimit[16]), .I3(n49949), .O(n49633));
    defparam i34046_4_lut.LUT_INIT = 16'h5a7b;
    SB_LUT4 i34792_4_lut (.I0(n30), .I1(n10_adj_4925), .I2(n51795), .I3(n49631), 
            .O(n50380));   // verilog/motorControl.v(31[10:34])
    defparam i34792_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i34178_3_lut (.I0(n50285), .I1(IntegralLimit[15]), .I2(\PID_CONTROLLER.integral [15]), 
            .I3(GND_net), .O(n49766));   // verilog/motorControl.v(31[10:34])
    defparam i34178_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i34870_4_lut (.I0(n49766), .I1(n50380), .I2(n51795), .I3(n49633), 
            .O(n50458));   // verilog/motorControl.v(31[10:34])
    defparam i34870_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 mult_10_i320_2_lut (.I0(\Kp[6] ), .I1(n1[12]), .I2(GND_net), 
            .I3(GND_net), .O(n475_adj_4971));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i320_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i34871_3_lut (.I0(n50458), .I1(IntegralLimit[18]), .I2(\PID_CONTROLLER.integral [18]), 
            .I3(GND_net), .O(n50459));   // verilog/motorControl.v(31[10:34])
    defparam i34871_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i34855_3_lut (.I0(n50459), .I1(IntegralLimit[19]), .I2(\PID_CONTROLLER.integral [19]), 
            .I3(GND_net), .O(n50443));   // verilog/motorControl.v(31[10:34])
    defparam i34855_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 mult_10_i247_2_lut (.I0(\Kp[5] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n366_adj_4972));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i247_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i34038_4_lut (.I0(\PID_CONTROLLER.integral [21]), .I1(n51763), 
            .I2(IntegralLimit[21]), .I3(n50446), .O(n49625));
    defparam i34038_4_lut.LUT_INIT = 16'h5a7b;
    SB_LUT4 mult_10_i296_2_lut (.I0(\Kp[6] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n439_adj_4973));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i296_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 IntegralLimit_23__I_0_i45_rep_220_2_lut (.I0(\PID_CONTROLLER.integral [22]), 
            .I1(IntegralLimit[22]), .I2(GND_net), .I3(GND_net), .O(n51761));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i45_rep_220_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i34804_4_lut (.I0(n49764), .I1(n50248), .I2(n51761), .I3(n49623), 
            .O(n50392));   // verilog/motorControl.v(31[10:34])
    defparam i34804_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i34184_3_lut (.I0(n50443), .I1(IntegralLimit[20]), .I2(\PID_CONTROLLER.integral [20]), 
            .I3(GND_net), .O(n49772));   // verilog/motorControl.v(31[10:34])
    defparam i34184_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 unary_minus_16_inv_0_i8_1_lut (.I0(PWMLimit[7]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5235[7]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_5000_10 (.CI(n39701), .I0(n13104[7]), .I1(n664_adj_4969), 
            .CO(n39702));
    SB_LUT4 mult_10_i369_2_lut (.I0(\Kp[7] ), .I1(n1[12]), .I2(GND_net), 
            .I3(GND_net), .O(n548_adj_4975));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i369_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i345_2_lut (.I0(\Kp[7] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n512_adj_4976));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i345_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i394_2_lut (.I0(\Kp[8] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n585_adj_4977));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i394_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5000_9_lut (.I0(GND_net), .I1(n13104[6]), .I2(n591_adj_4978), 
            .I3(n39700), .O(n12180[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5000_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5245_10_lut (.I0(GND_net), .I1(n17444[7]), .I2(n685), 
            .I3(n39565), .O(n17024[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5245_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i443_2_lut (.I0(\Kp[9] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n658_adj_4979));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i443_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i34811_3_lut (.I0(n50398), .I1(\PID_CONTROLLER.integral_23__N_3887 [23]), 
            .I2(\PID_CONTROLLER.integral [23]), .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3886 ));   // verilog/motorControl.v(31[38:63])
    defparam i34811_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i34806_4_lut (.I0(n49772), .I1(n50392), .I2(n51761), .I3(n49625), 
            .O(n50394));   // verilog/motorControl.v(31[10:34])
    defparam i34806_4_lut.LUT_INIT = 16'hccca;
    SB_CARRY add_5000_9 (.CI(n39700), .I0(n13104[6]), .I1(n591_adj_4978), 
            .CO(n39701));
    SB_LUT4 mult_10_i418_2_lut (.I0(\Kp[8] ), .I1(n1[12]), .I2(GND_net), 
            .I3(GND_net), .O(n621_adj_4980));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i418_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5000_8_lut (.I0(GND_net), .I1(n13104[5]), .I2(n518_adj_4981), 
            .I3(n39699), .O(n12180[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5000_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5000_8 (.CI(n39699), .I0(n13104[5]), .I1(n518_adj_4981), 
            .CO(n39700));
    SB_LUT4 mult_10_i492_2_lut (.I0(\Kp[10] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n731_adj_4982));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i492_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 \PID_CONTROLLER.integral_23__I_936_4_lut  (.I0(n50394), .I1(\PID_CONTROLLER.integral_23__N_3886 ), 
            .I2(\PID_CONTROLLER.integral [23]), .I3(IntegralLimit[23]), 
            .O(\PID_CONTROLLER.integral_23__N_3884 ));   // verilog/motorControl.v(31[10:63])
    defparam \PID_CONTROLLER.integral_23__I_936_4_lut .LUT_INIT = 16'h80c8;
    SB_LUT4 add_5000_7_lut (.I0(GND_net), .I1(n13104[4]), .I2(n445_adj_4983), 
            .I3(n39698), .O(n12180[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5000_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5000_7 (.CI(n39698), .I0(n13104[4]), .I1(n445_adj_4983), 
            .CO(n39699));
    SB_CARRY sub_3_add_2_19 (.CI(n38723), .I0(setpoint[17]), .I1(motor_state[17]), 
            .CO(n38724));
    SB_LUT4 add_5000_6_lut (.I0(GND_net), .I1(n13104[3]), .I2(n372_adj_4984), 
            .I3(n39697), .O(n12180[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5000_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i467_2_lut (.I0(\Kp[9] ), .I1(n1[12]), .I2(GND_net), 
            .I3(GND_net), .O(n694_adj_4985));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i467_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i541_2_lut (.I0(\Kp[11] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n804_adj_4986));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i541_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i590_2_lut (.I0(\Kp[12] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n877_adj_4987));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i590_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i639_2_lut (.I0(\Kp[13] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n950_adj_4988));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i639_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_1008_25_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [23]), 
            .I2(n4751[23]), .I3(n38637), .O(\PID_CONTROLLER.integral_23__N_3836 [23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1008_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_3_add_2_18_lut (.I0(GND_net), .I1(setpoint[16]), .I2(motor_state[16]), 
            .I3(n38722), .O(n1[16])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5000_6 (.CI(n39697), .I0(n13104[3]), .I1(n372_adj_4984), 
            .CO(n39698));
    SB_CARRY add_5245_10 (.CI(n39565), .I0(n17444[7]), .I1(n685), .CO(n39566));
    SB_LUT4 add_5000_5_lut (.I0(GND_net), .I1(n13104[2]), .I2(n299), .I3(n39696), 
            .O(n12180[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5000_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i688_2_lut (.I0(\Kp[14] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n1023_adj_4989));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i688_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i737_2_lut (.I0(\Kp[15] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n1096_adj_4990));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i737_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i375_2_lut (.I0(\Kp[7] ), .I1(n1[15]), .I2(GND_net), 
            .I3(GND_net), .O(n557));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i375_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5245_9_lut (.I0(GND_net), .I1(n17444[6]), .I2(n612), .I3(n39564), 
            .O(n17024[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5245_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5245_9 (.CI(n39564), .I0(n17444[6]), .I1(n612), .CO(n39565));
    SB_CARRY add_5000_5 (.CI(n39696), .I0(n13104[2]), .I1(n299), .CO(n39697));
    SB_LUT4 add_5245_8_lut (.I0(GND_net), .I1(n17444[5]), .I2(n539), .I3(n39563), 
            .O(n17024[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5245_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5245_8 (.CI(n39563), .I0(n17444[5]), .I1(n539), .CO(n39564));
    SB_LUT4 add_5000_4_lut (.I0(GND_net), .I1(n13104[1]), .I2(n226), .I3(n39695), 
            .O(n12180[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5000_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5245_7_lut (.I0(GND_net), .I1(n17444[4]), .I2(n466), .I3(n39562), 
            .O(n17024[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5245_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5000_4 (.CI(n39695), .I0(n13104[1]), .I1(n226), .CO(n39696));
    SB_CARRY add_5245_7 (.CI(n39562), .I0(n17444[4]), .I1(n466), .CO(n39563));
    SB_CARRY sub_3_add_2_18 (.CI(n38722), .I0(setpoint[16]), .I1(motor_state[16]), 
            .CO(n38723));
    SB_LUT4 mult_10_i516_2_lut (.I0(\Kp[10] ), .I1(n1[12]), .I2(GND_net), 
            .I3(GND_net), .O(n767_adj_4991));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i516_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i402_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n597_adj_4992));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i402_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5000_3_lut (.I0(GND_net), .I1(n13104[0]), .I2(n153), .I3(n39694), 
            .O(n12180[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5000_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_1008_24_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [22]), 
            .I2(n4751[22]), .I3(n38636), .O(\PID_CONTROLLER.integral_23__N_3836 [22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1008_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5000_3 (.CI(n39694), .I0(n13104[0]), .I1(n153), .CO(n39695));
    SB_LUT4 add_5000_2_lut (.I0(GND_net), .I1(n11_adj_4899), .I2(n80_adj_4898), 
            .I3(GND_net), .O(n12180[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5000_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_3_add_2_17_lut (.I0(GND_net), .I1(setpoint[15]), .I2(motor_state[15]), 
            .I3(n38721), .O(n1[15])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5000_2 (.CI(GND_net), .I0(n11_adj_4899), .I1(n80_adj_4898), 
            .CO(n39694));
    SB_LUT4 unary_minus_16_inv_0_i9_1_lut (.I0(PWMLimit[8]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5235[8]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_5041_21_lut (.I0(GND_net), .I1(n13944[18]), .I2(GND_net), 
            .I3(n39693), .O(n13104[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5041_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5245_6_lut (.I0(GND_net), .I1(n17444[3]), .I2(n393), .I3(n39561), 
            .O(n17024[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5245_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5041_20_lut (.I0(GND_net), .I1(n13944[17]), .I2(GND_net), 
            .I3(n39692), .O(n13104[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5041_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i424_2_lut (.I0(\Kp[8] ), .I1(n1[15]), .I2(GND_net), 
            .I3(GND_net), .O(n630));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i424_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i565_2_lut (.I0(\Kp[11] ), .I1(n1[12]), .I2(GND_net), 
            .I3(GND_net), .O(n840_adj_4994));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i565_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5041_20 (.CI(n39692), .I0(n13944[17]), .I1(GND_net), 
            .CO(n39693));
    SB_CARRY add_5245_6 (.CI(n39561), .I0(n17444[3]), .I1(n393), .CO(n39562));
    SB_LUT4 add_5041_19_lut (.I0(GND_net), .I1(n13944[16]), .I2(GND_net), 
            .I3(n39691), .O(n13104[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5041_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i73_2_lut (.I0(\Kp[1] ), .I1(n1[11]), .I2(GND_net), 
            .I3(GND_net), .O(n107));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i73_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i26_2_lut (.I0(\Kp[0] ), .I1(n1[12]), .I2(GND_net), 
            .I3(GND_net), .O(n38));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i26_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5245_5_lut (.I0(GND_net), .I1(n17444[2]), .I2(n320), .I3(n39560), 
            .O(n17024[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5245_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1008_24 (.CI(n38636), .I0(\PID_CONTROLLER.integral [22]), 
            .I1(n4751[22]), .CO(n38637));
    SB_CARRY add_5041_19 (.CI(n39691), .I0(n13944[16]), .I1(GND_net), 
            .CO(n39692));
    SB_LUT4 add_5041_18_lut (.I0(GND_net), .I1(n13944[15]), .I2(GND_net), 
            .I3(n39690), .O(n13104[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5041_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_3_add_2_17 (.CI(n38721), .I0(setpoint[15]), .I1(motor_state[15]), 
            .CO(n38722));
    SB_CARRY add_5245_5 (.CI(n39560), .I0(n17444[2]), .I1(n320), .CO(n39561));
    SB_LUT4 add_1008_23_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [21]), 
            .I2(n4751[21]), .I3(n38635), .O(\PID_CONTROLLER.integral_23__N_3836 [21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1008_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5245_4_lut (.I0(GND_net), .I1(n17444[1]), .I2(n247), .I3(n39559), 
            .O(n17024[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5245_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1008_23 (.CI(n38635), .I0(\PID_CONTROLLER.integral [21]), 
            .I1(n4751[21]), .CO(n38636));
    SB_CARRY add_5041_18 (.CI(n39690), .I0(n13944[15]), .I1(GND_net), 
            .CO(n39691));
    SB_LUT4 mult_10_i122_2_lut (.I0(\Kp[2] ), .I1(n1[11]), .I2(GND_net), 
            .I3(GND_net), .O(n180));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i122_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 sub_3_add_2_16_lut (.I0(GND_net), .I1(setpoint[14]), .I2(motor_state[14]), 
            .I3(n38720), .O(n1[14])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5041_17_lut (.I0(GND_net), .I1(n13944[14]), .I2(GND_net), 
            .I3(n39689), .O(n13104[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5041_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_1008_22_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [20]), 
            .I2(n4751[20]), .I3(n38634), .O(\PID_CONTROLLER.integral_23__N_3836 [20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1008_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_3_add_2_16 (.CI(n38720), .I0(setpoint[14]), .I1(motor_state[14]), 
            .CO(n38721));
    SB_CARRY add_5245_4 (.CI(n39559), .I0(n17444[1]), .I1(n247), .CO(n39560));
    SB_LUT4 sub_3_add_2_15_lut (.I0(GND_net), .I1(setpoint[13]), .I2(motor_state[13]), 
            .I3(n38719), .O(n1[13])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5245_3_lut (.I0(GND_net), .I1(n17444[0]), .I2(n174), .I3(n39558), 
            .O(n17024[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5245_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_3_add_2_15 (.CI(n38719), .I0(setpoint[13]), .I1(motor_state[13]), 
            .CO(n38720));
    SB_LUT4 mux_17_i2_3_lut (.I0(duty_23__N_3936[1]), .I1(n257[1]), .I2(n256_adj_4995), 
            .I3(GND_net), .O(duty_23__N_3911[1]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i2_3_lut (.I0(duty_23__N_3911[1]), .I1(PWMLimit[1]), 
            .I2(duty_23__N_3935), .I3(GND_net), .O(duty_23__N_3812[1]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i3_3_lut (.I0(duty_23__N_3936[2]), .I1(n257[2]), .I2(n256_adj_4995), 
            .I3(GND_net), .O(duty_23__N_3911[2]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i3_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 sub_3_add_2_14_lut (.I0(GND_net), .I1(setpoint[12]), .I2(motor_state[12]), 
            .I3(n38718), .O(n1[12])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_3_add_2_14 (.CI(n38718), .I0(setpoint[12]), .I1(motor_state[12]), 
            .CO(n38719));
    SB_CARRY add_5245_3 (.CI(n39558), .I0(n17444[0]), .I1(n174), .CO(n39559));
    SB_CARRY add_5041_17 (.CI(n39689), .I0(n13944[14]), .I1(GND_net), 
            .CO(n39690));
    SB_LUT4 add_5245_2_lut (.I0(GND_net), .I1(n32), .I2(n101), .I3(GND_net), 
            .O(n17024[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5245_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5041_16_lut (.I0(GND_net), .I1(n13944[13]), .I2(n1105_adj_4891), 
            .I3(n39688), .O(n13104[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5041_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5245_2 (.CI(GND_net), .I0(n32), .I1(n101), .CO(n39558));
    SB_LUT4 mult_10_i171_2_lut (.I0(\Kp[3] ), .I1(n1[11]), .I2(GND_net), 
            .I3(GND_net), .O(n253));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i171_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 duty_23__I_0_i3_3_lut (.I0(duty_23__N_3911[2]), .I1(PWMLimit[2]), 
            .I2(duty_23__N_3935), .I3(GND_net), .O(duty_23__N_3812[2]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i3_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_5399_8_lut (.I0(GND_net), .I1(n19088[5]), .I2(n560), .I3(n39557), 
            .O(n18991[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5399_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_17_i4_3_lut (.I0(duty_23__N_3936[3]), .I1(n257[3]), .I2(n256_adj_4995), 
            .I3(GND_net), .O(duty_23__N_3911[3]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i4_3_lut (.I0(duty_23__N_3911[3]), .I1(PWMLimit[3]), 
            .I2(duty_23__N_3935), .I3(GND_net), .O(duty_23__N_3812[3]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i5_3_lut (.I0(duty_23__N_3936[4]), .I1(n257[4]), .I2(n256_adj_4995), 
            .I3(GND_net), .O(duty_23__N_3911[4]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i5_3_lut (.I0(duty_23__N_3911[4]), .I1(PWMLimit[4]), 
            .I2(duty_23__N_3935), .I3(GND_net), .O(duty_23__N_3812[4]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i6_3_lut (.I0(duty_23__N_3936[5]), .I1(n257[5]), .I2(n256_adj_4995), 
            .I3(GND_net), .O(duty_23__N_3911[5]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i6_3_lut (.I0(duty_23__N_3911[5]), .I1(PWMLimit[5]), 
            .I2(duty_23__N_3935), .I3(GND_net), .O(duty_23__N_3812[5]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_10_i220_2_lut (.I0(\Kp[4] ), .I1(n1[11]), .I2(GND_net), 
            .I3(GND_net), .O(n326));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i220_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_17_i7_3_lut (.I0(duty_23__N_3936[6]), .I1(n257[6]), .I2(n256_adj_4995), 
            .I3(GND_net), .O(duty_23__N_3911[6]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i7_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i7_3_lut (.I0(duty_23__N_3911[6]), .I1(PWMLimit[6]), 
            .I2(duty_23__N_3935), .I3(GND_net), .O(duty_23__N_3812[6]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i7_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i8_3_lut (.I0(duty_23__N_3936[7]), .I1(n257[7]), .I2(n256_adj_4995), 
            .I3(GND_net), .O(duty_23__N_3911[7]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i8_3_lut (.I0(duty_23__N_3911[7]), .I1(PWMLimit[7]), 
            .I2(duty_23__N_3935), .I3(GND_net), .O(duty_23__N_3812[7]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_5041_16 (.CI(n39688), .I0(n13944[13]), .I1(n1105_adj_4891), 
            .CO(n39689));
    SB_LUT4 add_5041_15_lut (.I0(GND_net), .I1(n13944[12]), .I2(n1032_adj_4890), 
            .I3(n39687), .O(n13104[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5041_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5041_15 (.CI(n39687), .I0(n13944[12]), .I1(n1032_adj_4890), 
            .CO(n39688));
    SB_LUT4 add_5041_14_lut (.I0(GND_net), .I1(n13944[11]), .I2(n959_adj_4888), 
            .I3(n39686), .O(n13104[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5041_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5041_14 (.CI(n39686), .I0(n13944[11]), .I1(n959_adj_4888), 
            .CO(n39687));
    SB_LUT4 add_5399_7_lut (.I0(GND_net), .I1(n19088[4]), .I2(n487), .I3(n39556), 
            .O(n18991[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5399_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5041_13_lut (.I0(GND_net), .I1(n13944[10]), .I2(n886_adj_4887), 
            .I3(n39685), .O(n13104[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5041_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5399_7 (.CI(n39556), .I0(n19088[4]), .I1(n487), .CO(n39557));
    SB_CARRY add_1008_22 (.CI(n38634), .I0(\PID_CONTROLLER.integral [20]), 
            .I1(n4751[20]), .CO(n38635));
    SB_LUT4 add_5399_6_lut (.I0(GND_net), .I1(n19088[3]), .I2(n414), .I3(n39555), 
            .O(n18991[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5399_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5399_6 (.CI(n39555), .I0(n19088[3]), .I1(n414), .CO(n39556));
    SB_CARRY add_5041_13 (.CI(n39685), .I0(n13944[10]), .I1(n886_adj_4887), 
            .CO(n39686));
    SB_LUT4 add_5399_5_lut (.I0(GND_net), .I1(n19088[2]), .I2(n341), .I3(n39554), 
            .O(n18991[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5399_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_17_i9_3_lut (.I0(duty_23__N_3936[8]), .I1(n257[8]), .I2(n256_adj_4995), 
            .I3(GND_net), .O(duty_23__N_3911[8]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i9_3_lut (.I0(duty_23__N_3911[8]), .I1(PWMLimit[8]), 
            .I2(duty_23__N_3935), .I3(GND_net), .O(duty_23__N_3812[8]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_1008_21_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [19]), 
            .I2(n4751[19]), .I3(n38633), .O(\PID_CONTROLLER.integral_23__N_3836 [19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1008_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1008_21 (.CI(n38633), .I0(\PID_CONTROLLER.integral [19]), 
            .I1(n4751[19]), .CO(n38634));
    SB_LUT4 sub_3_add_2_13_lut (.I0(GND_net), .I1(setpoint[11]), .I2(motor_state[11]), 
            .I3(n38717), .O(n1[11])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5399_5 (.CI(n39554), .I0(n19088[2]), .I1(n341), .CO(n39555));
    SB_LUT4 mux_17_i10_3_lut (.I0(duty_23__N_3936[9]), .I1(n257[9]), .I2(n256_adj_4995), 
            .I3(GND_net), .O(duty_23__N_3911[9]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY sub_3_add_2_13 (.CI(n38717), .I0(setpoint[11]), .I1(motor_state[11]), 
            .CO(n38718));
    SB_LUT4 duty_23__I_0_i10_3_lut (.I0(duty_23__N_3911[9]), .I1(PWMLimit[9]), 
            .I2(duty_23__N_3935), .I3(GND_net), .O(duty_23__N_3812[9]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_5399_4_lut (.I0(GND_net), .I1(n19088[1]), .I2(n268), .I3(n39553), 
            .O(n18991[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5399_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_17_i11_3_lut (.I0(duty_23__N_3936[10]), .I1(n257[10]), .I2(n256_adj_4995), 
            .I3(GND_net), .O(duty_23__N_3911[10]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i11_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 sub_3_add_2_12_lut (.I0(GND_net), .I1(setpoint[10]), .I2(motor_state[10]), 
            .I3(n38716), .O(n1[10])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5041_12_lut (.I0(GND_net), .I1(n13944[9]), .I2(n813_adj_4885), 
            .I3(n39684), .O(n13104[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5041_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5399_4 (.CI(n39553), .I0(n19088[1]), .I1(n268), .CO(n39554));
    SB_CARRY sub_3_add_2_12 (.CI(n38716), .I0(setpoint[10]), .I1(motor_state[10]), 
            .CO(n38717));
    SB_LUT4 duty_23__I_0_i11_3_lut (.I0(duty_23__N_3911[10]), .I1(PWMLimit[10]), 
            .I2(duty_23__N_3935), .I3(GND_net), .O(duty_23__N_3812[10]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i11_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i12_3_lut (.I0(duty_23__N_3936[11]), .I1(n257[11]), .I2(n256_adj_4995), 
            .I3(GND_net), .O(duty_23__N_3911[11]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i12_3_lut (.I0(duty_23__N_3911[11]), .I1(PWMLimit[11]), 
            .I2(duty_23__N_3935), .I3(GND_net), .O(duty_23__N_3812[11]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_10_i269_2_lut (.I0(\Kp[5] ), .I1(n1[11]), .I2(GND_net), 
            .I3(GND_net), .O(n399));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i269_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i20906_2_lut (.I0(n1[23]), .I1(\PID_CONTROLLER.integral_23__N_3884 ), 
            .I2(GND_net), .I3(GND_net), .O(n4751[23]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i20906_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i251_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n372_adj_4984));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i251_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i300_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n445_adj_4983));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i300_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i349_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n518_adj_4981));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i349_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i461_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n685));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i461_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_17_i13_3_lut (.I0(duty_23__N_3936[12]), .I1(n257[12]), .I2(n256_adj_4995), 
            .I3(GND_net), .O(duty_23__N_3911[12]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i13_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i13_3_lut (.I0(duty_23__N_3911[12]), .I1(PWMLimit[12]), 
            .I2(duty_23__N_3935), .I3(GND_net), .O(duty_23__N_3812[12]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i13_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_1008_20_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [18]), 
            .I2(n4751[18]), .I3(n38632), .O(\PID_CONTROLLER.integral_23__N_3836 [18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1008_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_17_i14_3_lut (.I0(duty_23__N_3936[13]), .I1(n257[13]), .I2(n256_adj_4995), 
            .I3(GND_net), .O(duty_23__N_3911[13]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i14_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_1008_20 (.CI(n38632), .I0(\PID_CONTROLLER.integral [18]), 
            .I1(n4751[18]), .CO(n38633));
    SB_LUT4 mult_11_i398_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n591_adj_4978));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i398_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 sub_3_add_2_11_lut (.I0(GND_net), .I1(setpoint[9]), .I2(motor_state[9]), 
            .I3(n38715), .O(n1[9])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_1008_19_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [17]), 
            .I2(n4751[17]), .I3(n38631), .O(\PID_CONTROLLER.integral_23__N_3836 [17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1008_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_3_add_2_11 (.CI(n38715), .I0(setpoint[9]), .I1(motor_state[9]), 
            .CO(n38716));
    SB_LUT4 sub_3_add_2_10_lut (.I0(GND_net), .I1(setpoint[8]), .I2(motor_state[8]), 
            .I3(n38714), .O(n1[8])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 duty_23__I_0_i14_3_lut (.I0(duty_23__N_3911[13]), .I1(PWMLimit[13]), 
            .I2(duty_23__N_3935), .I3(GND_net), .O(duty_23__N_3812[13]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i14_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i15_3_lut (.I0(duty_23__N_3936[14]), .I1(n257[14]), .I2(n256_adj_4995), 
            .I3(GND_net), .O(duty_23__N_3911[14]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i15_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_5399_3_lut (.I0(GND_net), .I1(n19088[0]), .I2(n195), .I3(n39552), 
            .O(n18991[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5399_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5041_12 (.CI(n39684), .I0(n13944[9]), .I1(n813_adj_4885), 
            .CO(n39685));
    SB_LUT4 duty_23__I_0_i15_3_lut (.I0(duty_23__N_3911[14]), .I1(PWMLimit[14]), 
            .I2(duty_23__N_3935), .I3(GND_net), .O(duty_23__N_3812[14]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i15_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i16_3_lut (.I0(duty_23__N_3936[15]), .I1(n257[15]), .I2(n256_adj_4995), 
            .I3(GND_net), .O(duty_23__N_3911[15]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY sub_3_add_2_10 (.CI(n38714), .I0(setpoint[8]), .I1(motor_state[8]), 
            .CO(n38715));
    SB_LUT4 duty_23__I_0_i16_3_lut (.I0(duty_23__N_3911[15]), .I1(PWMLimit[15]), 
            .I2(duty_23__N_3935), .I3(GND_net), .O(duty_23__N_3812[15]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i17_3_lut (.I0(duty_23__N_3936[16]), .I1(n257[16]), .I2(n256_adj_4995), 
            .I3(GND_net), .O(duty_23__N_3911[16]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_11_i510_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n758));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i510_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i447_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n664_adj_4969));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i447_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5041_11_lut (.I0(GND_net), .I1(n13944[8]), .I2(n740_adj_4882), 
            .I3(n39683), .O(n13104[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5041_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_3_add_2_9_lut (.I0(GND_net), .I1(setpoint[7]), .I2(motor_state[7]), 
            .I3(n38713), .O(n1[7])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1008_19 (.CI(n38631), .I0(\PID_CONTROLLER.integral [17]), 
            .I1(n4751[17]), .CO(n38632));
    SB_CARRY add_5399_3 (.CI(n39552), .I0(n19088[0]), .I1(n195), .CO(n39553));
    SB_CARRY add_5041_11 (.CI(n39683), .I0(n13944[8]), .I1(n740_adj_4882), 
            .CO(n39684));
    SB_LUT4 add_5399_2_lut (.I0(GND_net), .I1(n53), .I2(n122), .I3(GND_net), 
            .O(n18991[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5399_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5041_10_lut (.I0(GND_net), .I1(n13944[7]), .I2(n667_adj_4879), 
            .I3(n39682), .O(n13104[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5041_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5399_2 (.CI(GND_net), .I0(n53), .I1(n122), .CO(n39552));
    SB_LUT4 duty_23__I_0_i17_3_lut (.I0(duty_23__N_3911[16]), .I1(PWMLimit[16]), 
            .I2(duty_23__N_3935), .I3(GND_net), .O(duty_23__N_3812[16]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i18_3_lut (.I0(duty_23__N_3936[17]), .I1(n257[17]), .I2(n256_adj_4995), 
            .I3(GND_net), .O(duty_23__N_3911[17]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i18_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i18_3_lut (.I0(duty_23__N_3911[17]), .I1(PWMLimit[17]), 
            .I2(duty_23__N_3935), .I3(GND_net), .O(duty_23__N_3812[17]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i18_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i19_3_lut (.I0(duty_23__N_3936[18]), .I1(n257[18]), .I2(n256_adj_4995), 
            .I3(GND_net), .O(duty_23__N_3911[18]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i19_3_lut (.I0(duty_23__N_3911[18]), .I1(PWMLimit[18]), 
            .I2(duty_23__N_3935), .I3(GND_net), .O(duty_23__N_3812[18]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i20_3_lut (.I0(duty_23__N_3936[19]), .I1(n257[19]), .I2(n256_adj_4995), 
            .I3(GND_net), .O(duty_23__N_3911[19]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i20_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i20_3_lut (.I0(duty_23__N_3911[19]), .I1(PWMLimit[19]), 
            .I2(duty_23__N_3935), .I3(GND_net), .O(duty_23__N_3812[19]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i20_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_11_i559_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n831));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i559_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i496_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n737_adj_4960));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i496_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_17_i21_3_lut (.I0(duty_23__N_3936[20]), .I1(n257[20]), .I2(n256_adj_4995), 
            .I3(GND_net), .O(duty_23__N_3911[20]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i21_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i21_3_lut (.I0(duty_23__N_3911[20]), .I1(PWMLimit[20]), 
            .I2(duty_23__N_3935), .I3(GND_net), .O(duty_23__N_3812[20]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i21_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_11_i545_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n810_adj_4959));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i545_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5272_14_lut (.I0(GND_net), .I1(n17808[11]), .I2(n980), 
            .I3(n39551), .O(n17444[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5272_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_1008_18_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [16]), 
            .I2(n4751[16]), .I3(n38630), .O(\PID_CONTROLLER.integral_23__N_3836 [16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1008_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1008_18 (.CI(n38630), .I0(\PID_CONTROLLER.integral [16]), 
            .I1(n4751[16]), .CO(n38631));
    SB_CARRY sub_3_add_2_9 (.CI(n38713), .I0(setpoint[7]), .I1(motor_state[7]), 
            .CO(n38714));
    SB_LUT4 add_5272_13_lut (.I0(GND_net), .I1(n17808[10]), .I2(n907), 
            .I3(n39550), .O(n17444[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5272_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_1008_17_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [15]), 
            .I2(n4751[15]), .I3(n38629), .O(\PID_CONTROLLER.integral_23__N_3836 [15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1008_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_17_i22_3_lut (.I0(duty_23__N_3936[21]), .I1(n257[21]), .I2(n256_adj_4995), 
            .I3(GND_net), .O(duty_23__N_3911[21]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i22_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i22_3_lut (.I0(duty_23__N_3911[21]), .I1(PWMLimit[21]), 
            .I2(duty_23__N_3935), .I3(GND_net), .O(duty_23__N_3812[21]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i22_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_1008_17 (.CI(n38629), .I0(\PID_CONTROLLER.integral [15]), 
            .I1(n4751[15]), .CO(n38630));
    SB_LUT4 sub_3_add_2_8_lut (.I0(GND_net), .I1(setpoint[6]), .I2(motor_state[6]), 
            .I3(n38712), .O(n1[6])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_3_add_2_8 (.CI(n38712), .I0(setpoint[6]), .I1(motor_state[6]), 
            .CO(n38713));
    SB_LUT4 add_1008_16_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [14]), 
            .I2(n4751[14]), .I3(n38628), .O(\PID_CONTROLLER.integral_23__N_3836 [14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1008_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_3_add_2_7_lut (.I0(GND_net), .I1(setpoint[5]), .I2(motor_state[5]), 
            .I3(n38711), .O(n1[5])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_3_add_2_7 (.CI(n38711), .I0(setpoint[5]), .I1(motor_state[5]), 
            .CO(n38712));
    SB_CARRY add_5272_13 (.CI(n39550), .I0(n17808[10]), .I1(n907), .CO(n39551));
    SB_CARRY add_5041_10 (.CI(n39682), .I0(n13944[7]), .I1(n667_adj_4879), 
            .CO(n39683));
    SB_LUT4 mux_17_i23_3_lut (.I0(duty_23__N_3936[22]), .I1(n257[22]), .I2(n256_adj_4995), 
            .I3(GND_net), .O(duty_23__N_3911[22]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i23_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_5041_9_lut (.I0(GND_net), .I1(n13944[6]), .I2(n594_adj_4874), 
            .I3(n39681), .O(n13104[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5041_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5272_12_lut (.I0(GND_net), .I1(n17808[9]), .I2(n834), 
            .I3(n39549), .O(n17444[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5272_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5272_12 (.CI(n39549), .I0(n17808[9]), .I1(n834), .CO(n39550));
    SB_LUT4 duty_23__I_0_i23_3_lut (.I0(duty_23__N_3911[22]), .I1(PWMLimit[22]), 
            .I2(duty_23__N_3935), .I3(GND_net), .O(duty_23__N_3812[22]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i23_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i24_3_lut (.I0(duty_23__N_3936[23]), .I1(n257[23]), .I2(n256_adj_4995), 
            .I3(GND_net), .O(duty_23__N_3911[23]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i24_3_lut (.I0(duty_23__N_3911[23]), .I1(PWMLimit[23]), 
            .I2(duty_23__N_3935), .I3(GND_net), .O(duty_23__N_3812[23]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 sub_3_add_2_6_lut (.I0(GND_net), .I1(setpoint[4]), .I2(motor_state[4]), 
            .I3(n38710), .O(n1[4])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_3_add_2_6 (.CI(n38710), .I0(setpoint[4]), .I1(motor_state[4]), 
            .CO(n38711));
    SB_CARRY add_5041_9 (.CI(n39681), .I0(n13944[6]), .I1(n594_adj_4874), 
            .CO(n39682));
    SB_LUT4 add_5272_11_lut (.I0(GND_net), .I1(n17808[8]), .I2(n761), 
            .I3(n39548), .O(n17444[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5272_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5272_11 (.CI(n39548), .I0(n17808[8]), .I1(n761), .CO(n39549));
    SB_CARRY add_1008_16 (.CI(n38628), .I0(\PID_CONTROLLER.integral [14]), 
            .I1(n4751[14]), .CO(n38629));
    SB_LUT4 sub_3_add_2_5_lut (.I0(GND_net), .I1(setpoint[3]), .I2(motor_state[3]), 
            .I3(n38709), .O(n1[3])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5272_10_lut (.I0(GND_net), .I1(n17808[7]), .I2(n688), 
            .I3(n39547), .O(n17444[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5272_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_3_add_2_5 (.CI(n38709), .I0(setpoint[3]), .I1(motor_state[3]), 
            .CO(n38710));
    SB_LUT4 add_1008_15_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [13]), 
            .I2(n4751[13]), .I3(n38627), .O(\PID_CONTROLLER.integral_23__N_3836 [13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1008_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_3_add_2_4_lut (.I0(GND_net), .I1(setpoint[2]), .I2(motor_state[2]), 
            .I3(n38708), .O(n1[2])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_3_add_2_4 (.CI(n38708), .I0(setpoint[2]), .I1(motor_state[2]), 
            .CO(n38709));
    SB_LUT4 sub_3_add_2_3_lut (.I0(GND_net), .I1(setpoint[1]), .I2(motor_state[1]), 
            .I3(n38707), .O(n1[1])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_3_add_2_3 (.CI(n38707), .I0(setpoint[1]), .I1(motor_state[1]), 
            .CO(n38708));
    SB_LUT4 add_5041_8_lut (.I0(GND_net), .I1(n13944[5]), .I2(n521_adj_4865), 
            .I3(n39680), .O(n13104[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5041_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i608_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n904));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i608_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_1008_15 (.CI(n38627), .I0(\PID_CONTROLLER.integral [13]), 
            .I1(n4751[13]), .CO(n38628));
    SB_LUT4 mult_11_i594_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n883_adj_4940));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i594_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 sub_3_add_2_2_lut (.I0(GND_net), .I1(setpoint[0]), .I2(motor_state[0]), 
            .I3(VCC_net), .O(n1[0])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_3_add_2_2 (.CI(VCC_net), .I0(setpoint[0]), .I1(motor_state[0]), 
            .CO(n38707));
    SB_CARRY add_5041_8 (.CI(n39680), .I0(n13944[5]), .I1(n521_adj_4865), 
            .CO(n39681));
    SB_CARRY add_5272_10 (.CI(n39547), .I0(n17808[7]), .I1(n688), .CO(n39548));
    SB_LUT4 mult_11_i657_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n977));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i657_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5272_9_lut (.I0(GND_net), .I1(n17808[6]), .I2(n615), .I3(n39546), 
            .O(n17444[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5272_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i643_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n956_adj_4937));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i643_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i692_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n1029_adj_4936));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i692_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_1008_14_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [12]), 
            .I2(n4751[12]), .I3(n38626), .O(\PID_CONTROLLER.integral_23__N_3836 [12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1008_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5041_7_lut (.I0(GND_net), .I1(n13944[4]), .I2(n448_adj_4862), 
            .I3(n39679), .O(n13104[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5041_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1008_14 (.CI(n38626), .I0(\PID_CONTROLLER.integral [12]), 
            .I1(n4751[12]), .CO(n38627));
    SB_CARRY add_5041_7 (.CI(n39679), .I0(n13944[4]), .I1(n448_adj_4862), 
            .CO(n39680));
    SB_LUT4 add_5041_6_lut (.I0(GND_net), .I1(n13944[3]), .I2(n375_adj_4861), 
            .I3(n39678), .O(n13104[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5041_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5272_9 (.CI(n39546), .I0(n17808[6]), .I1(n615), .CO(n39547));
    SB_LUT4 add_5272_8_lut (.I0(GND_net), .I1(n17808[5]), .I2(n542), .I3(n39545), 
            .O(n17444[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5272_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i741_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n1102_adj_4935));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i741_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5041_6 (.CI(n39678), .I0(n13944[3]), .I1(n375_adj_4861), 
            .CO(n39679));
    SB_CARRY add_5272_8 (.CI(n39545), .I0(n17808[5]), .I1(n542), .CO(n39546));
    SB_LUT4 add_5272_7_lut (.I0(GND_net), .I1(n17808[4]), .I2(n469), .I3(n39544), 
            .O(n17444[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5272_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_1008_13_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [11]), 
            .I2(n4751[11]), .I3(n38625), .O(\PID_CONTROLLER.integral_23__N_3836 [11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1008_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5041_5_lut (.I0(GND_net), .I1(n13944[2]), .I2(n302_adj_4859), 
            .I3(n39677), .O(n13104[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5041_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5041_5 (.CI(n39677), .I0(n13944[2]), .I1(n302_adj_4859), 
            .CO(n39678));
    SB_LUT4 mult_10_i318_2_lut (.I0(\Kp[6] ), .I1(n1[11]), .I2(GND_net), 
            .I3(GND_net), .O(n472));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i318_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5272_7 (.CI(n39544), .I0(n17808[4]), .I1(n469), .CO(n39545));
    SB_LUT4 add_5041_4_lut (.I0(GND_net), .I1(n13944[1]), .I2(n229_adj_4858), 
            .I3(n39676), .O(n13104[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5041_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5041_4 (.CI(n39676), .I0(n13944[1]), .I1(n229_adj_4858), 
            .CO(n39677));
    SB_LUT4 add_5272_6_lut (.I0(GND_net), .I1(n17808[3]), .I2(n396), .I3(n39543), 
            .O(n17444[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5272_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5041_3_lut (.I0(GND_net), .I1(n13944[0]), .I2(n156_adj_4857), 
            .I3(n39675), .O(n13104[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5041_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5041_3 (.CI(n39675), .I0(n13944[0]), .I1(n156_adj_4857), 
            .CO(n39676));
    SB_CARRY add_5272_6 (.CI(n39543), .I0(n17808[3]), .I1(n396), .CO(n39544));
    SB_LUT4 add_5041_2_lut (.I0(GND_net), .I1(n14_adj_4856), .I2(n83_adj_4855), 
            .I3(GND_net), .O(n13104[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5041_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5272_5_lut (.I0(GND_net), .I1(n17808[2]), .I2(n323), .I3(n39542), 
            .O(n17444[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5272_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5041_2 (.CI(GND_net), .I0(n14_adj_4856), .I1(n83_adj_4855), 
            .CO(n39675));
    SB_CARRY add_5272_5 (.CI(n39542), .I0(n17808[2]), .I1(n323), .CO(n39543));
    SB_LUT4 mult_11_i706_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n1050));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i706_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5272_4_lut (.I0(GND_net), .I1(n17808[1]), .I2(n250), .I3(n39541), 
            .O(n17444[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5272_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i67_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n98));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i67_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i20_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_4927));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i20_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i367_2_lut (.I0(\Kp[7] ), .I1(n1[11]), .I2(GND_net), 
            .I3(GND_net), .O(n545));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i367_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i416_2_lut (.I0(\Kp[8] ), .I1(n1[11]), .I2(GND_net), 
            .I3(GND_net), .O(n618));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i416_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5351_11_lut (.I0(GND_net), .I1(n18703[8]), .I2(n770), 
            .I3(n39674), .O(n18504[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5351_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5272_4 (.CI(n39541), .I0(n17808[1]), .I1(n250), .CO(n39542));
    SB_LUT4 add_5272_3_lut (.I0(GND_net), .I1(n17808[0]), .I2(n177), .I3(n39540), 
            .O(n17444[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5272_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i116_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n171));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i116_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i465_2_lut (.I0(\Kp[9] ), .I1(n1[11]), .I2(GND_net), 
            .I3(GND_net), .O(n691));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i465_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5351_10_lut (.I0(GND_net), .I1(n18703[7]), .I2(n697), 
            .I3(n39673), .O(n18504[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5351_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i114_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n168));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i114_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5351_10 (.CI(n39673), .I0(n18703[7]), .I1(n697), .CO(n39674));
    SB_CARRY add_5272_3 (.CI(n39540), .I0(n17808[0]), .I1(n177), .CO(n39541));
    SB_LUT4 add_5351_9_lut (.I0(GND_net), .I1(n18703[6]), .I2(n624), .I3(n39672), 
            .O(n18504[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5351_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1008_13 (.CI(n38625), .I0(\PID_CONTROLLER.integral [11]), 
            .I1(n4751[11]), .CO(n38626));
    SB_LUT4 add_1008_12_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [10]), 
            .I2(n4751[10]), .I3(n38624), .O(\PID_CONTROLLER.integral_23__N_3836 [10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1008_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1008_12 (.CI(n38624), .I0(\PID_CONTROLLER.integral [10]), 
            .I1(n4751[10]), .CO(n38625));
    SB_CARRY add_5351_9 (.CI(n39672), .I0(n18703[6]), .I1(n624), .CO(n39673));
    SB_LUT4 unary_minus_16_inv_0_i16_1_lut (.I0(PWMLimit[15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5235[15]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_5272_2_lut (.I0(GND_net), .I1(n35_adj_5004), .I2(n104), 
            .I3(GND_net), .O(n17444[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5272_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5351_8_lut (.I0(GND_net), .I1(n18703[5]), .I2(n551), .I3(n39671), 
            .O(n18504[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5351_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5272_2 (.CI(GND_net), .I0(n35_adj_5004), .I1(n104), .CO(n39540));
    SB_CARRY add_5351_8 (.CI(n39671), .I0(n18703[5]), .I1(n551), .CO(n39672));
    SB_LUT4 add_1008_11_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(n4751[9]), .I3(n38623), .O(\PID_CONTROLLER.integral_23__N_3836 [9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1008_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1008_11 (.CI(n38623), .I0(\PID_CONTROLLER.integral [9]), 
            .I1(n4751[9]), .CO(n38624));
    SB_LUT4 mult_11_i508_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n755));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i508_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5351_7_lut (.I0(GND_net), .I1(n18703[4]), .I2(n478), .I3(n39670), 
            .O(n18504[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5351_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5297_13_lut (.I0(GND_net), .I1(n18120[10]), .I2(n910), 
            .I3(n39539), .O(n17808[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5297_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i163_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n241));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i163_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5297_12_lut (.I0(GND_net), .I1(n18120[9]), .I2(n837), 
            .I3(n39538), .O(n17808[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5297_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5351_7 (.CI(n39670), .I0(n18703[4]), .I1(n478), .CO(n39671));
    SB_LUT4 add_1008_10_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(n4751[8]), .I3(n38622), .O(\PID_CONTROLLER.integral_23__N_3836 [8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1008_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5351_6_lut (.I0(GND_net), .I1(n18703[3]), .I2(n405), .I3(n39669), 
            .O(n18504[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5351_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1008_10 (.CI(n38622), .I0(\PID_CONTROLLER.integral [8]), 
            .I1(n4751[8]), .CO(n38623));
    SB_LUT4 add_1008_9_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(n4751[7]), .I3(n38621), .O(\PID_CONTROLLER.integral_23__N_3836 [7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1008_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1008_9 (.CI(n38621), .I0(\PID_CONTROLLER.integral [7]), 
            .I1(n4751[7]), .CO(n38622));
    SB_LUT4 add_1008_8_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(n4751[6]), .I3(n38620), .O(\PID_CONTROLLER.integral_23__N_3836 [6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1008_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1008_8 (.CI(n38620), .I0(\PID_CONTROLLER.integral [6]), 
            .I1(n4751[6]), .CO(n38621));
    SB_LUT4 add_1008_7_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(n4751[5]), .I3(n38619), .O(\PID_CONTROLLER.integral_23__N_3836 [5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1008_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1008_7 (.CI(n38619), .I0(\PID_CONTROLLER.integral [5]), 
            .I1(n4751[5]), .CO(n38620));
    SB_CARRY add_5297_12 (.CI(n39538), .I0(n18120[9]), .I1(n837), .CO(n39539));
    SB_LUT4 add_1008_6_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(n4751[4]), .I3(n38618), .O(\PID_CONTROLLER.integral_23__N_3836 [4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1008_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5297_11_lut (.I0(GND_net), .I1(n18120[8]), .I2(n764), 
            .I3(n39537), .O(n17808[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5297_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5351_6 (.CI(n39669), .I0(n18703[3]), .I1(n405), .CO(n39670));
    SB_CARRY add_1008_6 (.CI(n38618), .I0(\PID_CONTROLLER.integral [4]), 
            .I1(n4751[4]), .CO(n38619));
    SB_CARRY add_5297_11 (.CI(n39537), .I0(n18120[8]), .I1(n764), .CO(n39538));
    SB_LUT4 add_5351_5_lut (.I0(GND_net), .I1(n18703[2]), .I2(n332), .I3(n39668), 
            .O(n18504[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5351_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_1008_5_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(n4751[3]), .I3(n38617), .O(\PID_CONTROLLER.integral_23__N_3836 [3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1008_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5297_10_lut (.I0(GND_net), .I1(n18120[7]), .I2(n691_adj_5005), 
            .I3(n39536), .O(n17808[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5297_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5351_5 (.CI(n39668), .I0(n18703[2]), .I1(n332), .CO(n39669));
    SB_LUT4 unary_minus_5_inv_0_i4_1_lut (.I0(IntegralLimit[3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5234[3]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_1008_5 (.CI(n38617), .I0(\PID_CONTROLLER.integral [3]), 
            .I1(n4751[3]), .CO(n38618));
    SB_CARRY add_5297_10 (.CI(n39536), .I0(n18120[7]), .I1(n691_adj_5005), 
            .CO(n39537));
    SB_LUT4 add_5351_4_lut (.I0(GND_net), .I1(n18703[1]), .I2(n259_adj_5006), 
            .I3(n39667), .O(n18504[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5351_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_1008_4_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(n4751[2]), .I3(n38616), .O(\PID_CONTROLLER.integral_23__N_3836 [2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1008_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1008_4 (.CI(n38616), .I0(\PID_CONTROLLER.integral [2]), 
            .I1(n4751[2]), .CO(n38617));
    SB_CARRY add_5351_4 (.CI(n39667), .I0(n18703[1]), .I1(n259_adj_5006), 
            .CO(n39668));
    SB_LUT4 add_5351_3_lut (.I0(GND_net), .I1(n18703[0]), .I2(n186), .I3(n39666), 
            .O(n18504[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5351_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5297_9_lut (.I0(GND_net), .I1(n18120[6]), .I2(n618_adj_5007), 
            .I3(n39535), .O(n17808[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5297_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_1008_3_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(n4751[1]), .I3(n38615), .O(\PID_CONTROLLER.integral_23__N_3836 [1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1008_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5351_3 (.CI(n39666), .I0(n18703[0]), .I1(n186), .CO(n39667));
    SB_LUT4 add_5351_2_lut (.I0(GND_net), .I1(n44), .I2(n113), .I3(GND_net), 
            .O(n18504[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5351_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5297_9 (.CI(n39535), .I0(n18120[6]), .I1(n618_adj_5007), 
            .CO(n39536));
    SB_CARRY add_5351_2 (.CI(GND_net), .I0(n44), .I1(n113), .CO(n39666));
    SB_LUT4 add_5297_8_lut (.I0(GND_net), .I1(n18120[5]), .I2(n545_adj_5008), 
            .I3(n39534), .O(n17808[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5297_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5297_8 (.CI(n39534), .I0(n18120[5]), .I1(n545_adj_5008), 
            .CO(n39535));
    SB_LUT4 add_5080_20_lut (.I0(GND_net), .I1(n14704[17]), .I2(GND_net), 
            .I3(n39665), .O(n13944[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5080_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5080_19_lut (.I0(GND_net), .I1(n14704[16]), .I2(GND_net), 
            .I3(n39664), .O(n13944[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5080_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5080_19 (.CI(n39664), .I0(n14704[16]), .I1(GND_net), 
            .CO(n39665));
    SB_LUT4 add_5297_7_lut (.I0(GND_net), .I1(n18120[4]), .I2(n472_adj_5009), 
            .I3(n39533), .O(n17808[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5297_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5297_7 (.CI(n39533), .I0(n18120[4]), .I1(n472_adj_5009), 
            .CO(n39534));
    SB_LUT4 add_5080_18_lut (.I0(GND_net), .I1(n14704[15]), .I2(GND_net), 
            .I3(n39663), .O(n13944[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5080_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5297_6_lut (.I0(GND_net), .I1(n18120[3]), .I2(n399_adj_5010), 
            .I3(n39532), .O(n17808[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5297_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5297_6 (.CI(n39532), .I0(n18120[3]), .I1(n399_adj_5010), 
            .CO(n39533));
    SB_CARRY add_5080_18 (.CI(n39663), .I0(n14704[15]), .I1(GND_net), 
            .CO(n39664));
    SB_LUT4 add_5080_17_lut (.I0(GND_net), .I1(n14704[14]), .I2(GND_net), 
            .I3(n39662), .O(n13944[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5080_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5297_5_lut (.I0(GND_net), .I1(n18120[2]), .I2(n326_adj_5011), 
            .I3(n39531), .O(n17808[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5297_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5297_5 (.CI(n39531), .I0(n18120[2]), .I1(n326_adj_5011), 
            .CO(n39532));
    SB_LUT4 add_5297_4_lut (.I0(GND_net), .I1(n18120[1]), .I2(n253_adj_5012), 
            .I3(n39530), .O(n17808[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5297_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5297_4 (.CI(n39530), .I0(n18120[1]), .I1(n253_adj_5012), 
            .CO(n39531));
    SB_LUT4 mult_11_i212_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n314));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i212_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i451_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n670_adj_5013));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i451_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5297_3_lut (.I0(GND_net), .I1(n18120[0]), .I2(n180_adj_5014), 
            .I3(n39529), .O(n17808[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5297_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5297_3 (.CI(n39529), .I0(n18120[0]), .I1(n180_adj_5014), 
            .CO(n39530));
    SB_LUT4 add_5297_2_lut (.I0(GND_net), .I1(n38_adj_5015), .I2(n107_adj_5016), 
            .I3(GND_net), .O(n17808[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5297_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1008_3 (.CI(n38615), .I0(\PID_CONTROLLER.integral [1]), 
            .I1(n4751[1]), .CO(n38616));
    SB_CARRY add_5080_17 (.CI(n39662), .I0(n14704[14]), .I1(GND_net), 
            .CO(n39663));
    SB_LUT4 unary_minus_5_inv_0_i2_1_lut (.I0(IntegralLimit[1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5234[1]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i514_2_lut (.I0(\Kp[10] ), .I1(n1[11]), .I2(GND_net), 
            .I3(GND_net), .O(n764_adj_5017));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i514_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i563_2_lut (.I0(\Kp[11] ), .I1(n1[11]), .I2(GND_net), 
            .I3(GND_net), .O(n837_adj_5018));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i563_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i612_2_lut (.I0(\Kp[12] ), .I1(n1[11]), .I2(GND_net), 
            .I3(GND_net), .O(n910_adj_5019));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i612_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i261_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n387));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i261_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i310_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n460));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i310_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i85_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [17]), 
            .I2(GND_net), .I3(GND_net), .O(n125));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i85_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i38_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [18]), 
            .I2(GND_net), .I3(GND_net), .O(n56));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i38_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5297_2 (.CI(GND_net), .I0(n38_adj_5015), .I1(n107_adj_5016), 
            .CO(n39529));
    SB_LUT4 add_5411_7_lut (.I0(GND_net), .I1(n45851), .I2(n490), .I3(n39528), 
            .O(n19088[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5411_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5080_16_lut (.I0(GND_net), .I1(n14704[13]), .I2(n1108_adj_5020), 
            .I3(n39661), .O(n13944[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5080_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i134_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [17]), 
            .I2(GND_net), .I3(GND_net), .O(n198));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i134_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i17_1_lut (.I0(PWMLimit[16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5235[16]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i183_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [17]), 
            .I2(GND_net), .I3(GND_net), .O(n271_adj_5022));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i183_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i232_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [17]), 
            .I2(GND_net), .I3(GND_net), .O(n344));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i232_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i281_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [17]), 
            .I2(GND_net), .I3(GND_net), .O(n417));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i281_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_4_lut (.I0(n6_adj_5023), .I1(\Ki[4] ), .I2(n19184[2]), 
            .I3(\PID_CONTROLLER.integral_23__N_3836 [18]), .O(n19124[3]));   // verilog/motorControl.v(34[25:36])
    defparam i2_4_lut.LUT_INIT = 16'h965a;
    SB_LUT4 add_5411_6_lut (.I0(GND_net), .I1(n19159[3]), .I2(n417_adj_5024), 
            .I3(n39527), .O(n19088[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5411_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_1008_2_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [0]), 
            .I2(n4751[0]), .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3836 [0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1008_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5080_16 (.CI(n39661), .I0(n14704[13]), .I1(n1108_adj_5020), 
            .CO(n39662));
    SB_LUT4 add_5080_15_lut (.I0(GND_net), .I1(n14704[12]), .I2(n1035_adj_5025), 
            .I3(n39660), .O(n13944[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5080_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1008_2 (.CI(GND_net), .I0(\PID_CONTROLLER.integral [0]), 
            .I1(n4751[0]), .CO(n38615));
    SB_CARRY add_5080_15 (.CI(n39660), .I0(n14704[12]), .I1(n1035_adj_5025), 
            .CO(n39661));
    SB_LUT4 add_5080_14_lut (.I0(GND_net), .I1(n14704[11]), .I2(n962_adj_5026), 
            .I3(n39659), .O(n13944[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5080_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5411_6 (.CI(n39527), .I0(n19159[3]), .I1(n417_adj_5024), 
            .CO(n39528));
    SB_CARRY add_5080_14 (.CI(n39659), .I0(n14704[11]), .I1(n962_adj_5026), 
            .CO(n39660));
    SB_LUT4 add_5080_13_lut (.I0(GND_net), .I1(n14704[10]), .I2(n889_adj_5027), 
            .I3(n39658), .O(n13944[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5080_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5411_5_lut (.I0(GND_net), .I1(n19159[2]), .I2(n344_adj_5028), 
            .I3(n39526), .O(n19088[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5411_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5411_5 (.CI(n39526), .I0(n19159[2]), .I1(n344_adj_5028), 
            .CO(n39527));
    SB_CARRY add_5080_13 (.CI(n39658), .I0(n14704[10]), .I1(n889_adj_5027), 
            .CO(n39659));
    SB_LUT4 add_5411_4_lut (.I0(GND_net), .I1(n19159[1]), .I2(n271_adj_5029), 
            .I3(n39525), .O(n19088[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5411_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5411_4 (.CI(n39525), .I0(n19159[1]), .I1(n271_adj_5029), 
            .CO(n39526));
    SB_LUT4 add_5411_3_lut (.I0(GND_net), .I1(n19159[0]), .I2(n198_adj_5030), 
            .I3(n39524), .O(n19088[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5411_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5080_12_lut (.I0(GND_net), .I1(n14704[9]), .I2(n816_adj_5031), 
            .I3(n39657), .O(n13944[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5080_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5411_3 (.CI(n39524), .I0(n19159[0]), .I1(n198_adj_5030), 
            .CO(n39525));
    SB_LUT4 add_5411_2_lut (.I0(GND_net), .I1(n56_adj_5032), .I2(n125_adj_5033), 
            .I3(GND_net), .O(n19088[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5411_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5411_2 (.CI(GND_net), .I0(n56_adj_5032), .I1(n125_adj_5033), 
            .CO(n39524));
    SB_CARRY add_5080_12 (.CI(n39657), .I0(n14704[9]), .I1(n816_adj_5031), 
            .CO(n39658));
    SB_LUT4 add_5080_11_lut (.I0(GND_net), .I1(n14704[8]), .I2(n743_adj_5034), 
            .I3(n39656), .O(n13944[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5080_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5080_11 (.CI(n39656), .I0(n14704[8]), .I1(n743_adj_5034), 
            .CO(n39657));
    SB_LUT4 mult_11_i200_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n296));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i200_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_12_25_lut (.I0(GND_net), .I1(n11187[0]), .I2(n10656[0]), 
            .I3(n38614), .O(duty_23__N_3936[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5080_10_lut (.I0(GND_net), .I1(n14704[7]), .I2(n670_adj_5013), 
            .I3(n39655), .O(n13944[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5080_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_12_24_lut (.I0(GND_net), .I1(n106[22]), .I2(n155[22]), 
            .I3(n38613), .O(duty_23__N_3936[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i2_4_lut_adj_1714 (.I0(n4_adj_5035), .I1(\Ki[3] ), .I2(n19224[1]), 
            .I3(\PID_CONTROLLER.integral_23__N_3836 [19]), .O(n19184[2]));   // verilog/motorControl.v(34[25:36])
    defparam i2_4_lut_adj_1714.LUT_INIT = 16'h965a;
    SB_LUT4 i24427_4_lut (.I0(\Ki[0] ), .I1(\Ki[1] ), .I2(\PID_CONTROLLER.integral_23__N_3836 [22]), 
            .I3(\PID_CONTROLLER.integral_23__N_3836 [21]), .O(n19248[0]));   // verilog/motorControl.v(34[25:36])
    defparam i24427_4_lut.LUT_INIT = 16'h6ca0;
    SB_LUT4 mult_11_i330_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [17]), 
            .I2(GND_net), .I3(GND_net), .O(n490_adj_5036));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i330_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_4_lut_adj_1715 (.I0(\Ki[0] ), .I1(\Ki[3] ), .I2(\PID_CONTROLLER.integral_23__N_3836 [23]), 
            .I3(\PID_CONTROLLER.integral_23__N_3836 [20]), .O(n12_adj_5037));   // verilog/motorControl.v(34[25:36])
    defparam i2_4_lut_adj_1715.LUT_INIT = 16'h9c50;
    SB_LUT4 i24349_4_lut (.I0(n19184[2]), .I1(\Ki[4] ), .I2(n6_adj_5023), 
            .I3(\PID_CONTROLLER.integral_23__N_3836 [18]), .O(n8_adj_5038));   // verilog/motorControl.v(34[25:36])
    defparam i24349_4_lut.LUT_INIT = 16'he8a0;
    SB_LUT4 i1_4_lut (.I0(\Ki[4] ), .I1(\Ki[2] ), .I2(\PID_CONTROLLER.integral_23__N_3836 [19]), 
            .I3(\PID_CONTROLLER.integral_23__N_3836 [21]), .O(n11_adj_5039));   // verilog/motorControl.v(34[25:36])
    defparam i1_4_lut.LUT_INIT = 16'h6ca0;
    SB_CARRY add_5080_10 (.CI(n39655), .I0(n14704[7]), .I1(n670_adj_5013), 
            .CO(n39656));
    SB_LUT4 i24303_4_lut (.I0(n19224[1]), .I1(\Ki[3] ), .I2(n4_adj_5035), 
            .I3(\PID_CONTROLLER.integral_23__N_3836 [19]), .O(n6_adj_5040));   // verilog/motorControl.v(34[25:36])
    defparam i24303_4_lut.LUT_INIT = 16'he8a0;
    SB_DFF \PID_CONTROLLER.integral_i23  (.Q(\PID_CONTROLLER.integral [23]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3836 [23]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i22  (.Q(\PID_CONTROLLER.integral [22]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3836 [22]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i21  (.Q(\PID_CONTROLLER.integral [21]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3836 [21]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i20  (.Q(\PID_CONTROLLER.integral [20]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3836 [20]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i19  (.Q(\PID_CONTROLLER.integral [19]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3836 [19]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i18  (.Q(\PID_CONTROLLER.integral [18]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3836 [18]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i17  (.Q(\PID_CONTROLLER.integral [17]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3836 [17]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i16  (.Q(\PID_CONTROLLER.integral [16]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3836 [16]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i15  (.Q(\PID_CONTROLLER.integral [15]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3836 [15]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i14  (.Q(\PID_CONTROLLER.integral [14]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3836 [14]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i13  (.Q(\PID_CONTROLLER.integral [13]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3836 [13]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i12  (.Q(\PID_CONTROLLER.integral [12]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3836 [12]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i11  (.Q(\PID_CONTROLLER.integral [11]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3836 [11]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i10  (.Q(\PID_CONTROLLER.integral [10]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3836 [10]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i9  (.Q(\PID_CONTROLLER.integral [9]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3836 [9]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i8  (.Q(\PID_CONTROLLER.integral [8]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3836 [8]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i7  (.Q(\PID_CONTROLLER.integral [7]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3836 [7]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i6  (.Q(\PID_CONTROLLER.integral [6]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3836 [6]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i5  (.Q(\PID_CONTROLLER.integral [5]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3836 [5]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i4  (.Q(\PID_CONTROLLER.integral [4]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3836 [4]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i3  (.Q(\PID_CONTROLLER.integral [3]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3836 [3]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i2  (.Q(\PID_CONTROLLER.integral [2]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3836 [2]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i1  (.Q(\PID_CONTROLLER.integral [1]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3836 [1]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i23 (.Q(duty[23]), .C(clk32MHz), .D(duty_23__N_3812[23]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i22 (.Q(duty[22]), .C(clk32MHz), .D(duty_23__N_3812[22]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i21 (.Q(duty[21]), .C(clk32MHz), .D(duty_23__N_3812[21]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i20 (.Q(duty[20]), .C(clk32MHz), .D(duty_23__N_3812[20]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i19 (.Q(duty[19]), .C(clk32MHz), .D(duty_23__N_3812[19]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i18 (.Q(duty[18]), .C(clk32MHz), .D(duty_23__N_3812[18]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i17 (.Q(duty[17]), .C(clk32MHz), .D(duty_23__N_3812[17]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i16 (.Q(duty[16]), .C(clk32MHz), .D(duty_23__N_3812[16]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i15 (.Q(duty[15]), .C(clk32MHz), .D(duty_23__N_3812[15]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i14 (.Q(duty[14]), .C(clk32MHz), .D(duty_23__N_3812[14]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i13 (.Q(duty[13]), .C(clk32MHz), .D(duty_23__N_3812[13]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i12 (.Q(duty[12]), .C(clk32MHz), .D(duty_23__N_3812[12]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i11 (.Q(duty[11]), .C(clk32MHz), .D(duty_23__N_3812[11]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i10 (.Q(duty[10]), .C(clk32MHz), .D(duty_23__N_3812[10]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i9 (.Q(duty[9]), .C(clk32MHz), .D(duty_23__N_3812[9]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i8 (.Q(duty[8]), .C(clk32MHz), .D(duty_23__N_3812[8]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i7 (.Q(duty[7]), .C(clk32MHz), .D(duty_23__N_3812[7]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i6 (.Q(duty[6]), .C(clk32MHz), .D(duty_23__N_3812[6]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i5 (.Q(duty[5]), .C(clk32MHz), .D(duty_23__N_3812[5]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i4 (.Q(duty[4]), .C(clk32MHz), .D(duty_23__N_3812[4]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i3 (.Q(duty[3]), .C(clk32MHz), .D(duty_23__N_3812[3]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i2 (.Q(duty[2]), .C(clk32MHz), .D(duty_23__N_3812[2]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i1 (.Q(duty[1]), .C(clk32MHz), .D(duty_23__N_3812[1]));   // verilog/motorControl.v(29[14] 48[8])
    SB_LUT4 i24429_4_lut (.I0(\Ki[0] ), .I1(\Ki[1] ), .I2(\PID_CONTROLLER.integral_23__N_3836 [22]), 
            .I3(\PID_CONTROLLER.integral_23__N_3836 [21]), .O(n38389));   // verilog/motorControl.v(34[25:36])
    defparam i24429_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 add_5080_9_lut (.I0(GND_net), .I1(n14704[6]), .I2(n597_adj_4992), 
            .I3(n39654), .O(n13944[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5080_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i8_4_lut (.I0(n6_adj_5040), .I1(n11_adj_5039), .I2(n8_adj_5038), 
            .I3(n12_adj_5037), .O(n18_adj_5041));   // verilog/motorControl.v(34[25:36])
    defparam i8_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut (.I0(\Ki[5] ), .I1(\Ki[1] ), .I2(\PID_CONTROLLER.integral_23__N_3836 [18]), 
            .I3(\PID_CONTROLLER.integral_23__N_3836 [22]), .O(n13_adj_5042));   // verilog/motorControl.v(34[25:36])
    defparam i3_4_lut.LUT_INIT = 16'h6ca0;
    SB_LUT4 i9_4_lut (.I0(n13_adj_5042), .I1(n18_adj_5041), .I2(n38389), 
            .I3(n4_adj_5043), .O(n46355));   // verilog/motorControl.v(34[25:36])
    defparam i9_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i33898_2_lut_4_lut (.I0(duty_23__N_3936[21]), .I1(n257[21]), 
            .I2(duty_23__N_3936[9]), .I3(n257[9]), .O(n49485));
    defparam i33898_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i33919_2_lut_4_lut (.I0(duty_23__N_3936[16]), .I1(n257[16]), 
            .I2(duty_23__N_3936[7]), .I3(n257[7]), .O(n49506));
    defparam i33919_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 mult_10_add_1225_24_lut (.I0(n1[23]), .I1(n11694[21]), .I2(GND_net), 
            .I3(n39990), .O(n11187[0])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_24_lut.LUT_INIT = 16'h6996;
    SB_LUT4 mult_10_add_1225_23_lut (.I0(GND_net), .I1(n11694[20]), .I2(GND_net), 
            .I3(n39989), .O(n106[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_23 (.CI(n39989), .I0(n11694[20]), .I1(GND_net), 
            .CO(n39990));
    SB_LUT4 mult_10_add_1225_22_lut (.I0(GND_net), .I1(n11694[19]), .I2(GND_net), 
            .I3(n39988), .O(n106[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_22 (.CI(n39988), .I0(n11694[19]), .I1(GND_net), 
            .CO(n39989));
    SB_LUT4 mult_10_add_1225_21_lut (.I0(GND_net), .I1(n11694[18]), .I2(GND_net), 
            .I3(n39987), .O(n106[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_21 (.CI(n39987), .I0(n11694[18]), .I1(GND_net), 
            .CO(n39988));
    SB_LUT4 mult_10_add_1225_20_lut (.I0(GND_net), .I1(n11694[17]), .I2(GND_net), 
            .I3(n39986), .O(n106[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i71_2_lut (.I0(\Kp[1] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n104_adj_5044));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i71_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mult_10_add_1225_20 (.CI(n39986), .I0(n11694[17]), .I1(GND_net), 
            .CO(n39987));
    SB_LUT4 mult_10_add_1225_19_lut (.I0(GND_net), .I1(n11694[16]), .I2(GND_net), 
            .I3(n39985), .O(n106[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_19 (.CI(n39985), .I0(n11694[16]), .I1(GND_net), 
            .CO(n39986));
    SB_LUT4 mult_10_add_1225_18_lut (.I0(GND_net), .I1(n11694[15]), .I2(GND_net), 
            .I3(n39984), .O(n106[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_18 (.CI(n39984), .I0(n11694[15]), .I1(GND_net), 
            .CO(n39985));
    SB_LUT4 mult_10_add_1225_17_lut (.I0(GND_net), .I1(n11694[14]), .I2(GND_net), 
            .I3(n39983), .O(n106[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_17 (.CI(n39983), .I0(n11694[14]), .I1(GND_net), 
            .CO(n39984));
    SB_LUT4 mult_10_add_1225_16_lut (.I0(GND_net), .I1(n11694[13]), .I2(n1096_adj_4990), 
            .I3(n39982), .O(n106[15])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_16 (.CI(n39982), .I0(n11694[13]), .I1(n1096_adj_4990), 
            .CO(n39983));
    SB_LUT4 mult_10_add_1225_15_lut (.I0(GND_net), .I1(n11694[12]), .I2(n1023_adj_4989), 
            .I3(n39981), .O(n106[14])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_15 (.CI(n39981), .I0(n11694[12]), .I1(n1023_adj_4989), 
            .CO(n39982));
    SB_LUT4 mult_10_i24_2_lut (.I0(\Kp[0] ), .I1(n1[11]), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_5045));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i24_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_add_1225_14_lut (.I0(GND_net), .I1(n11694[11]), .I2(n950_adj_4988), 
            .I3(n39980), .O(n106[13])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_14 (.CI(n39980), .I0(n11694[11]), .I1(n950_adj_4988), 
            .CO(n39981));
    SB_LUT4 mult_10_add_1225_13_lut (.I0(GND_net), .I1(n11694[10]), .I2(n877_adj_4987), 
            .I3(n39979), .O(n106[12])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_13 (.CI(n39979), .I0(n11694[10]), .I1(n877_adj_4987), 
            .CO(n39980));
    SB_LUT4 mult_10_i120_2_lut (.I0(\Kp[2] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n177_adj_5046));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i120_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_add_1225_12_lut (.I0(GND_net), .I1(n11694[9]), .I2(n804_adj_4986), 
            .I3(n39978), .O(n106[11])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_12 (.CI(n39978), .I0(n11694[9]), .I1(n804_adj_4986), 
            .CO(n39979));
    SB_LUT4 mult_10_add_1225_11_lut (.I0(GND_net), .I1(n11694[8]), .I2(n731_adj_4982), 
            .I3(n39977), .O(n106[10])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_11 (.CI(n39977), .I0(n11694[8]), .I1(n731_adj_4982), 
            .CO(n39978));
    SB_LUT4 mult_10_add_1225_10_lut (.I0(GND_net), .I1(n11694[7]), .I2(n658_adj_4979), 
            .I3(n39976), .O(n106[9])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_10 (.CI(n39976), .I0(n11694[7]), .I1(n658_adj_4979), 
            .CO(n39977));
    SB_LUT4 mult_10_add_1225_9_lut (.I0(GND_net), .I1(n11694[6]), .I2(n585_adj_4977), 
            .I3(n39975), .O(n106[8])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_9 (.CI(n39975), .I0(n11694[6]), .I1(n585_adj_4977), 
            .CO(n39976));
    SB_LUT4 mult_10_add_1225_8_lut (.I0(GND_net), .I1(n11694[5]), .I2(n512_adj_4976), 
            .I3(n39974), .O(n106[7])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_8 (.CI(n39974), .I0(n11694[5]), .I1(n512_adj_4976), 
            .CO(n39975));
    SB_LUT4 mult_10_add_1225_7_lut (.I0(GND_net), .I1(n11694[4]), .I2(n439_adj_4973), 
            .I3(n39973), .O(n106[6])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_7 (.CI(n39973), .I0(n11694[4]), .I1(n439_adj_4973), 
            .CO(n39974));
    SB_LUT4 mult_10_i169_2_lut (.I0(\Kp[3] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n250_adj_5048));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i169_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i218_2_lut (.I0(\Kp[4] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n323_adj_5049));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i218_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_add_1225_6_lut (.I0(GND_net), .I1(n11694[3]), .I2(n366_adj_4972), 
            .I3(n39972), .O(n106[5])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i33957_2_lut_4_lut (.I0(PWMLimit[21]), .I1(duty_23__N_3936[21]), 
            .I2(PWMLimit[9]), .I3(duty_23__N_3936[9]), .O(n49544));
    defparam i33957_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 mult_10_i267_2_lut (.I0(\Kp[5] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n396_adj_5050));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i267_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i316_2_lut (.I0(\Kp[6] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n469_adj_5051));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i316_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i18_1_lut (.I0(PWMLimit[17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5235[17]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i359_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n533));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i359_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mult_10_add_1225_6 (.CI(n39972), .I0(n11694[3]), .I1(n366_adj_4972), 
            .CO(n39973));
    SB_LUT4 mult_10_add_1225_5_lut (.I0(GND_net), .I1(n11694[2]), .I2(n293_adj_4968), 
            .I3(n39971), .O(n106[4])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_5 (.CI(n39971), .I0(n11694[2]), .I1(n293_adj_4968), 
            .CO(n39972));
    SB_LUT4 mult_10_add_1225_4_lut (.I0(GND_net), .I1(n11694[1]), .I2(n220_adj_4967), 
            .I3(n39970), .O(n106[3])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_4 (.CI(n39970), .I0(n11694[1]), .I1(n220_adj_4967), 
            .CO(n39971));
    SB_LUT4 mult_10_add_1225_3_lut (.I0(GND_net), .I1(n11694[0]), .I2(n147_adj_4966), 
            .I3(n39969), .O(n106[2])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_3 (.CI(n39969), .I0(n11694[0]), .I1(n147_adj_4966), 
            .CO(n39970));
    SB_CARRY add_12_24 (.CI(n38613), .I0(n106[22]), .I1(n155[22]), .CO(n38614));
    SB_LUT4 mult_10_add_1225_2_lut (.I0(GND_net), .I1(n5_adj_4965), .I2(n74_adj_4964), 
            .I3(GND_net), .O(n106[1])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_2 (.CI(GND_net), .I0(n5_adj_4965), .I1(n74_adj_4964), 
            .CO(n39969));
    SB_LUT4 mult_10_i365_2_lut (.I0(\Kp[7] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n542_adj_5055));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i365_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4978_23_lut (.I0(GND_net), .I1(n12663[20]), .I2(GND_net), 
            .I3(n39968), .O(n11694[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4978_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4978_22_lut (.I0(GND_net), .I1(n12663[19]), .I2(GND_net), 
            .I3(n39967), .O(n11694[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4978_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4978_22 (.CI(n39967), .I0(n12663[19]), .I1(GND_net), 
            .CO(n39968));
    SB_LUT4 add_4978_21_lut (.I0(GND_net), .I1(n12663[18]), .I2(GND_net), 
            .I3(n39966), .O(n11694[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4978_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4978_21 (.CI(n39966), .I0(n12663[18]), .I1(GND_net), 
            .CO(n39967));
    SB_LUT4 add_4978_20_lut (.I0(GND_net), .I1(n12663[17]), .I2(GND_net), 
            .I3(n39965), .O(n11694[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4978_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4978_20 (.CI(n39965), .I0(n12663[17]), .I1(GND_net), 
            .CO(n39966));
    SB_LUT4 mult_10_i414_2_lut (.I0(\Kp[8] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n615_adj_5056));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i414_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4978_19_lut (.I0(GND_net), .I1(n12663[16]), .I2(GND_net), 
            .I3(n39964), .O(n11694[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4978_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4978_19 (.CI(n39964), .I0(n12663[16]), .I1(GND_net), 
            .CO(n39965));
    SB_LUT4 add_4978_18_lut (.I0(GND_net), .I1(n12663[15]), .I2(GND_net), 
            .I3(n39963), .O(n11694[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4978_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i463_2_lut (.I0(\Kp[9] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n688_adj_5057));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i463_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4978_18 (.CI(n39963), .I0(n12663[15]), .I1(GND_net), 
            .CO(n39964));
    SB_LUT4 add_4978_17_lut (.I0(GND_net), .I1(n12663[14]), .I2(GND_net), 
            .I3(n39962), .O(n11694[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4978_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i408_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n606));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i408_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4978_17 (.CI(n39962), .I0(n12663[14]), .I1(GND_net), 
            .CO(n39963));
    SB_LUT4 mult_10_i512_2_lut (.I0(\Kp[10] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n761_adj_5058));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i512_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4978_16_lut (.I0(GND_net), .I1(n12663[13]), .I2(n1099_adj_4961), 
            .I3(n39961), .O(n11694[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4978_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4978_16 (.CI(n39961), .I0(n12663[13]), .I1(n1099_adj_4961), 
            .CO(n39962));
    SB_LUT4 add_4978_15_lut (.I0(GND_net), .I1(n12663[12]), .I2(n1026_adj_4958), 
            .I3(n39960), .O(n11694[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4978_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4978_15 (.CI(n39960), .I0(n12663[12]), .I1(n1026_adj_4958), 
            .CO(n39961));
    SB_LUT4 add_4978_14_lut (.I0(GND_net), .I1(n12663[11]), .I2(n953_adj_4957), 
            .I3(n39959), .O(n11694[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4978_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4978_14 (.CI(n39959), .I0(n12663[11]), .I1(n953_adj_4957), 
            .CO(n39960));
    SB_LUT4 add_4978_13_lut (.I0(GND_net), .I1(n12663[10]), .I2(n880_adj_4955), 
            .I3(n39958), .O(n11694[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4978_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i561_2_lut (.I0(\Kp[11] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n834_adj_5059));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i561_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4978_13 (.CI(n39958), .I0(n12663[10]), .I1(n880_adj_4955), 
            .CO(n39959));
    SB_LUT4 add_4978_12_lut (.I0(GND_net), .I1(n12663[9]), .I2(n807_adj_4952), 
            .I3(n39957), .O(n11694[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4978_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4978_12 (.CI(n39957), .I0(n12663[9]), .I1(n807_adj_4952), 
            .CO(n39958));
    SB_LUT4 add_4978_11_lut (.I0(GND_net), .I1(n12663[8]), .I2(n734_adj_4951), 
            .I3(n39956), .O(n11694[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4978_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4978_11 (.CI(n39956), .I0(n12663[8]), .I1(n734_adj_4951), 
            .CO(n39957));
    SB_LUT4 add_4978_10_lut (.I0(GND_net), .I1(n12663[7]), .I2(n661_adj_4947), 
            .I3(n39955), .O(n11694[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4978_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4978_10 (.CI(n39955), .I0(n12663[7]), .I1(n661_adj_4947), 
            .CO(n39956));
    SB_LUT4 add_4978_9_lut (.I0(GND_net), .I1(n12663[6]), .I2(n588_adj_4946), 
            .I3(n39954), .O(n11694[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4978_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4978_9 (.CI(n39954), .I0(n12663[6]), .I1(n588_adj_4946), 
            .CO(n39955));
    SB_LUT4 add_4978_8_lut (.I0(GND_net), .I1(n12663[5]), .I2(n515_adj_4944), 
            .I3(n39953), .O(n11694[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4978_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4978_8 (.CI(n39953), .I0(n12663[5]), .I1(n515_adj_4944), 
            .CO(n39954));
    SB_LUT4 add_4978_7_lut (.I0(GND_net), .I1(n12663[4]), .I2(n442_adj_4943), 
            .I3(n39952), .O(n11694[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4978_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4978_7 (.CI(n39952), .I0(n12663[4]), .I1(n442_adj_4943), 
            .CO(n39953));
    SB_LUT4 add_4978_6_lut (.I0(GND_net), .I1(n12663[3]), .I2(n369_adj_4942), 
            .I3(n39951), .O(n11694[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4978_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4978_6 (.CI(n39951), .I0(n12663[3]), .I1(n369_adj_4942), 
            .CO(n39952));
    SB_LUT4 add_4978_5_lut (.I0(GND_net), .I1(n12663[2]), .I2(n296_adj_4939), 
            .I3(n39950), .O(n11694[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4978_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_inv_0_i19_1_lut (.I0(PWMLimit[18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5235[18]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_4978_5 (.CI(n39950), .I0(n12663[2]), .I1(n296_adj_4939), 
            .CO(n39951));
    SB_LUT4 i33970_2_lut_4_lut (.I0(PWMLimit[16]), .I1(duty_23__N_3936[16]), 
            .I2(PWMLimit[7]), .I3(duty_23__N_3936[7]), .O(n49557));
    defparam i33970_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 mult_10_i610_2_lut (.I0(\Kp[12] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n907_adj_5061));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i610_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4978_4_lut (.I0(GND_net), .I1(n12663[1]), .I2(n223_adj_4938), 
            .I3(n39949), .O(n11694[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4978_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4978_4 (.CI(n39949), .I0(n12663[1]), .I1(n223_adj_4938), 
            .CO(n39950));
    SB_LUT4 add_4978_3_lut (.I0(GND_net), .I1(n12663[0]), .I2(n150_adj_4934), 
            .I3(n39948), .O(n11694[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4978_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4978_3 (.CI(n39948), .I0(n12663[0]), .I1(n150_adj_4934), 
            .CO(n39949));
    SB_LUT4 add_4978_2_lut (.I0(GND_net), .I1(n8_adj_4933), .I2(n77_adj_4932), 
            .I3(GND_net), .O(n11694[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4978_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4978_2 (.CI(GND_net), .I0(n8_adj_4933), .I1(n77_adj_4932), 
            .CO(n39948));
    SB_LUT4 add_5021_22_lut (.I0(GND_net), .I1(n13544[19]), .I2(GND_net), 
            .I3(n39947), .O(n12663[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5021_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_inv_0_i20_1_lut (.I0(PWMLimit[19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5235[19]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_5021_21_lut (.I0(GND_net), .I1(n13544[18]), .I2(GND_net), 
            .I3(n39946), .O(n12663[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5021_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5021_21 (.CI(n39946), .I0(n13544[18]), .I1(GND_net), 
            .CO(n39947));
    SB_LUT4 add_5021_20_lut (.I0(GND_net), .I1(n13544[17]), .I2(GND_net), 
            .I3(n39945), .O(n12663[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5021_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i659_2_lut (.I0(\Kp[13] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n980_adj_5063));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i659_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5021_20 (.CI(n39945), .I0(n13544[17]), .I1(GND_net), 
            .CO(n39946));
    SB_LUT4 add_5021_19_lut (.I0(GND_net), .I1(n13544[16]), .I2(GND_net), 
            .I3(n39944), .O(n12663[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5021_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5021_19 (.CI(n39944), .I0(n13544[16]), .I1(GND_net), 
            .CO(n39945));
    SB_LUT4 add_5021_18_lut (.I0(GND_net), .I1(n13544[15]), .I2(GND_net), 
            .I3(n39943), .O(n12663[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5021_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i165_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n244));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i165_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i214_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n317));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i214_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i69_2_lut (.I0(\Kp[1] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n101_adj_5064));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i69_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i22_2_lut (.I0(\Kp[0] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n32_adj_5065));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i22_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i118_2_lut (.I0(\Kp[2] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n174_adj_5066));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i118_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5021_18 (.CI(n39943), .I0(n13544[15]), .I1(GND_net), 
            .CO(n39944));
    SB_LUT4 add_5021_17_lut (.I0(GND_net), .I1(n13544[14]), .I2(GND_net), 
            .I3(n39942), .O(n12663[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5021_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5021_17 (.CI(n39942), .I0(n13544[14]), .I1(GND_net), 
            .CO(n39943));
    SB_LUT4 add_5021_16_lut (.I0(GND_net), .I1(n13544[13]), .I2(n1102), 
            .I3(n39941), .O(n12663[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5021_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5021_16 (.CI(n39941), .I0(n13544[13]), .I1(n1102), .CO(n39942));
    SB_LUT4 add_5021_15_lut (.I0(GND_net), .I1(n13544[12]), .I2(n1029), 
            .I3(n39940), .O(n12663[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5021_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5021_15 (.CI(n39940), .I0(n13544[12]), .I1(n1029), .CO(n39941));
    SB_LUT4 add_5021_14_lut (.I0(GND_net), .I1(n13544[11]), .I2(n956), 
            .I3(n39939), .O(n12663[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5021_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5021_14 (.CI(n39939), .I0(n13544[11]), .I1(n956), .CO(n39940));
    SB_LUT4 add_5021_13_lut (.I0(GND_net), .I1(n13544[10]), .I2(n883), 
            .I3(n39938), .O(n12663[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5021_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5021_13 (.CI(n39938), .I0(n13544[10]), .I1(n883), .CO(n39939));
    SB_LUT4 add_5021_12_lut (.I0(GND_net), .I1(n13544[9]), .I2(n810), 
            .I3(n39937), .O(n12663[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5021_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i167_2_lut (.I0(\Kp[3] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n247_adj_5067));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i167_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5021_12 (.CI(n39937), .I0(n13544[9]), .I1(n810), .CO(n39938));
    SB_LUT4 add_5021_11_lut (.I0(GND_net), .I1(n13544[8]), .I2(n737), 
            .I3(n39936), .O(n12663[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5021_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5021_11 (.CI(n39936), .I0(n13544[8]), .I1(n737), .CO(n39937));
    SB_LUT4 add_5021_10_lut (.I0(GND_net), .I1(n13544[7]), .I2(n664), 
            .I3(n39935), .O(n12663[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5021_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5021_10 (.CI(n39935), .I0(n13544[7]), .I1(n664), .CO(n39936));
    SB_LUT4 add_5021_9_lut (.I0(GND_net), .I1(n13544[6]), .I2(n591), .I3(n39934), 
            .O(n12663[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5021_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_inv_0_i21_1_lut (.I0(PWMLimit[20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5235[20]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_5021_9 (.CI(n39934), .I0(n13544[6]), .I1(n591), .CO(n39935));
    SB_LUT4 add_5021_8_lut (.I0(GND_net), .I1(n13544[5]), .I2(n518), .I3(n39933), 
            .O(n12663[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5021_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5021_8 (.CI(n39933), .I0(n13544[5]), .I1(n518), .CO(n39934));
    SB_LUT4 add_5021_7_lut (.I0(GND_net), .I1(n13544[4]), .I2(n445), .I3(n39932), 
            .O(n12663[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5021_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i216_2_lut (.I0(\Kp[4] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n320_adj_5069));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i216_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i22_1_lut (.I0(PWMLimit[21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5235[21]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_12_23_lut (.I0(GND_net), .I1(n106[21]), .I2(n155[21]), 
            .I3(n38612), .O(duty_23__N_3936[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_12_23 (.CI(n38612), .I0(n106[21]), .I1(n155[21]), .CO(n38613));
    SB_CARRY add_5080_9 (.CI(n39654), .I0(n14704[6]), .I1(n597_adj_4992), 
            .CO(n39655));
    SB_LUT4 mult_10_i265_2_lut (.I0(\Kp[5] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n393_adj_5071));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i265_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_12_22_lut (.I0(GND_net), .I1(n106[20]), .I2(n155[20]), 
            .I3(n38611), .O(duty_23__N_3936[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_12_22 (.CI(n38611), .I0(n106[20]), .I1(n155[20]), .CO(n38612));
    SB_LUT4 mult_10_i314_2_lut (.I0(\Kp[6] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n466_adj_5073));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i314_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i363_2_lut (.I0(\Kp[7] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n539_adj_5074));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i363_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i457_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n679));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i457_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i412_2_lut (.I0(\Kp[8] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n612_adj_5075));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i412_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5021_7 (.CI(n39932), .I0(n13544[4]), .I1(n445), .CO(n39933));
    SB_LUT4 unary_minus_16_inv_0_i23_1_lut (.I0(PWMLimit[22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5235[22]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i263_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n390));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i263_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5080_8_lut (.I0(GND_net), .I1(n14704[5]), .I2(n524_adj_4923), 
            .I3(n39653), .O(n13944[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5080_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5021_6_lut (.I0(GND_net), .I1(n13544[3]), .I2(n372), .I3(n39931), 
            .O(n12663[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5021_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5021_6 (.CI(n39931), .I0(n13544[3]), .I1(n372), .CO(n39932));
    SB_LUT4 unary_minus_16_inv_0_i24_1_lut (.I0(PWMLimit[23]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5235[23]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_5021_5_lut (.I0(GND_net), .I1(n13544[2]), .I2(n299_adj_4919), 
            .I3(n39930), .O(n12663[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5021_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5021_5 (.CI(n39930), .I0(n13544[2]), .I1(n299_adj_4919), 
            .CO(n39931));
    SB_LUT4 add_5021_4_lut (.I0(GND_net), .I1(n13544[1]), .I2(n226_adj_4908), 
            .I3(n39929), .O(n12663[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5021_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5021_4 (.CI(n39929), .I0(n13544[1]), .I1(n226_adj_4908), 
            .CO(n39930));
    SB_LUT4 add_5021_3_lut (.I0(GND_net), .I1(n13544[0]), .I2(n153_adj_4904), 
            .I3(n39928), .O(n12663[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5021_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5080_8 (.CI(n39653), .I0(n14704[5]), .I1(n524_adj_4923), 
            .CO(n39654));
    SB_CARRY add_5021_3 (.CI(n39928), .I0(n13544[0]), .I1(n153_adj_4904), 
            .CO(n39929));
    SB_LUT4 add_5021_2_lut (.I0(GND_net), .I1(n11_adj_4897), .I2(n80), 
            .I3(GND_net), .O(n12663[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5021_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5021_2 (.CI(GND_net), .I0(n11_adj_4897), .I1(n80), .CO(n39928));
    SB_LUT4 add_5061_21_lut (.I0(GND_net), .I1(n14343[18]), .I2(GND_net), 
            .I3(n39927), .O(n13544[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5061_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i500_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n743_adj_5034));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i500_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i461_2_lut (.I0(\Kp[9] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n685_adj_5078));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i461_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i85_2_lut (.I0(\Kp[1] ), .I1(n1[17]), .I2(GND_net), 
            .I3(GND_net), .O(n125_adj_5033));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i85_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i38_2_lut (.I0(\Kp[0] ), .I1(n1[18]), .I2(GND_net), 
            .I3(GND_net), .O(n56_adj_5032));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i38_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5061_20_lut (.I0(GND_net), .I1(n14343[17]), .I2(GND_net), 
            .I3(n39926), .O(n13544[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5061_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i549_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n816_adj_5031));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i549_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i134_2_lut (.I0(\Kp[2] ), .I1(n1[17]), .I2(GND_net), 
            .I3(GND_net), .O(n198_adj_5030));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i134_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5080_7_lut (.I0(GND_net), .I1(n14704[4]), .I2(n451_adj_4854), 
            .I3(n39652), .O(n13944[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5080_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_12_21_lut (.I0(GND_net), .I1(n106[19]), .I2(n155[19]), 
            .I3(n38610), .O(duty_23__N_3936[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_12_21 (.CI(n38610), .I0(n106[19]), .I1(n155[19]), .CO(n38611));
    SB_LUT4 mult_10_i510_2_lut (.I0(\Kp[10] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n758_adj_5079));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i510_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i183_2_lut (.I0(\Kp[3] ), .I1(n1[17]), .I2(GND_net), 
            .I3(GND_net), .O(n271_adj_5029));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i183_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5061_20 (.CI(n39926), .I0(n14343[17]), .I1(GND_net), 
            .CO(n39927));
    SB_LUT4 add_5061_19_lut (.I0(GND_net), .I1(n14343[16]), .I2(GND_net), 
            .I3(n39925), .O(n13544[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5061_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5061_19 (.CI(n39925), .I0(n14343[16]), .I1(GND_net), 
            .CO(n39926));
    SB_LUT4 add_5061_18_lut (.I0(GND_net), .I1(n14343[15]), .I2(GND_net), 
            .I3(n39924), .O(n13544[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5061_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5061_18 (.CI(n39924), .I0(n14343[15]), .I1(GND_net), 
            .CO(n39925));
    SB_LUT4 mult_10_i232_2_lut (.I0(\Kp[4] ), .I1(n1[17]), .I2(GND_net), 
            .I3(GND_net), .O(n344_adj_5028));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i232_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5061_17_lut (.I0(GND_net), .I1(n14343[14]), .I2(GND_net), 
            .I3(n39923), .O(n13544[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5061_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i598_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n889_adj_5027));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i598_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5061_17 (.CI(n39923), .I0(n14343[14]), .I1(GND_net), 
            .CO(n39924));
    SB_LUT4 add_5061_16_lut (.I0(GND_net), .I1(n14343[13]), .I2(n1105), 
            .I3(n39922), .O(n13544[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5061_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5061_16 (.CI(n39922), .I0(n14343[13]), .I1(n1105), .CO(n39923));
    SB_LUT4 add_5061_15_lut (.I0(GND_net), .I1(n14343[12]), .I2(n1032), 
            .I3(n39921), .O(n13544[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5061_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5061_15 (.CI(n39921), .I0(n14343[12]), .I1(n1032), .CO(n39922));
    SB_LUT4 add_12_20_lut (.I0(GND_net), .I1(n106[18]), .I2(n155[18]), 
            .I3(n38609), .O(duty_23__N_3936[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5061_14_lut (.I0(GND_net), .I1(n14343[11]), .I2(n959), 
            .I3(n39920), .O(n13544[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5061_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5061_14 (.CI(n39920), .I0(n14343[11]), .I1(n959), .CO(n39921));
    SB_LUT4 add_5061_13_lut (.I0(GND_net), .I1(n14343[10]), .I2(n886), 
            .I3(n39919), .O(n13544[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5061_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5061_13 (.CI(n39919), .I0(n14343[10]), .I1(n886), .CO(n39920));
    SB_LUT4 add_5061_12_lut (.I0(GND_net), .I1(n14343[9]), .I2(n813), 
            .I3(n39918), .O(n13544[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5061_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5080_7 (.CI(n39652), .I0(n14704[4]), .I1(n451_adj_4854), 
            .CO(n39653));
    SB_CARRY add_5061_12 (.CI(n39918), .I0(n14343[9]), .I1(n813), .CO(n39919));
    SB_LUT4 add_5061_11_lut (.I0(GND_net), .I1(n14343[8]), .I2(n740), 
            .I3(n39917), .O(n13544[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5061_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5061_11 (.CI(n39917), .I0(n14343[8]), .I1(n740), .CO(n39918));
    SB_LUT4 add_5061_10_lut (.I0(GND_net), .I1(n14343[7]), .I2(n667), 
            .I3(n39916), .O(n13544[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5061_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5061_10 (.CI(n39916), .I0(n14343[7]), .I1(n667), .CO(n39917));
    SB_LUT4 add_5061_9_lut (.I0(GND_net), .I1(n14343[6]), .I2(n594), .I3(n39915), 
            .O(n13544[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5061_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5061_9 (.CI(n39915), .I0(n14343[6]), .I1(n594), .CO(n39916));
    SB_LUT4 add_5080_6_lut (.I0(GND_net), .I1(n14704[3]), .I2(n378_adj_4852), 
            .I3(n39651), .O(n13944[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5080_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5080_6 (.CI(n39651), .I0(n14704[3]), .I1(n378_adj_4852), 
            .CO(n39652));
    SB_LUT4 add_5080_5_lut (.I0(GND_net), .I1(n14704[2]), .I2(n305_adj_4851), 
            .I3(n39650), .O(n13944[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5080_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5080_5 (.CI(n39650), .I0(n14704[2]), .I1(n305_adj_4851), 
            .CO(n39651));
    SB_LUT4 add_5080_4_lut (.I0(GND_net), .I1(n14704[1]), .I2(n232_adj_4849), 
            .I3(n39649), .O(n13944[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5080_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5080_4 (.CI(n39649), .I0(n14704[1]), .I1(n232_adj_4849), 
            .CO(n39650));
    SB_LUT4 add_5080_3_lut (.I0(GND_net), .I1(n14704[0]), .I2(n159_adj_4848), 
            .I3(n39648), .O(n13944[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5080_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5080_3 (.CI(n39648), .I0(n14704[0]), .I1(n159_adj_4848), 
            .CO(n39649));
    SB_LUT4 add_5061_8_lut (.I0(GND_net), .I1(n14343[5]), .I2(n521), .I3(n39914), 
            .O(n13544[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5061_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5080_2_lut (.I0(GND_net), .I1(n17_adj_4847), .I2(n86_adj_4846), 
            .I3(GND_net), .O(n13944[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5080_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5061_8 (.CI(n39914), .I0(n14343[5]), .I1(n521), .CO(n39915));
    SB_LUT4 add_5061_7_lut (.I0(GND_net), .I1(n14343[4]), .I2(n448), .I3(n39913), 
            .O(n13544[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5061_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5061_7 (.CI(n39913), .I0(n14343[4]), .I1(n448), .CO(n39914));
    SB_CARRY add_12_20 (.CI(n38609), .I0(n106[18]), .I1(n155[18]), .CO(n38610));
    SB_LUT4 add_5061_6_lut (.I0(GND_net), .I1(n14343[3]), .I2(n375), .I3(n39912), 
            .O(n13544[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5061_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5061_6 (.CI(n39912), .I0(n14343[3]), .I1(n375), .CO(n39913));
    SB_LUT4 add_5061_5_lut (.I0(GND_net), .I1(n14343[2]), .I2(n302), .I3(n39911), 
            .O(n13544[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5061_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5061_5 (.CI(n39911), .I0(n14343[2]), .I1(n302), .CO(n39912));
    SB_LUT4 add_5061_4_lut (.I0(GND_net), .I1(n14343[1]), .I2(n229), .I3(n39910), 
            .O(n13544[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5061_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5080_2 (.CI(GND_net), .I0(n17_adj_4847), .I1(n86_adj_4846), 
            .CO(n39648));
    SB_LUT4 add_5117_19_lut (.I0(GND_net), .I1(n15388[16]), .I2(GND_net), 
            .I3(n39647), .O(n14704[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5117_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5117_18_lut (.I0(GND_net), .I1(n15388[15]), .I2(GND_net), 
            .I3(n39646), .O(n14704[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5117_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_12_19_lut (.I0(GND_net), .I1(n106[17]), .I2(n155[17]), 
            .I3(n38608), .O(duty_23__N_3936[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5117_18 (.CI(n39646), .I0(n15388[15]), .I1(GND_net), 
            .CO(n39647));
    SB_LUT4 mult_11_i506_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n752));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i506_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5117_17_lut (.I0(GND_net), .I1(n15388[14]), .I2(GND_net), 
            .I3(n39645), .O(n14704[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5117_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_12_19 (.CI(n38608), .I0(n106[17]), .I1(n155[17]), .CO(n38609));
    SB_LUT4 add_12_18_lut (.I0(GND_net), .I1(n106[16]), .I2(n155[16]), 
            .I3(n38607), .O(duty_23__N_3936[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5117_17 (.CI(n39645), .I0(n15388[14]), .I1(GND_net), 
            .CO(n39646));
    SB_LUT4 add_5117_16_lut (.I0(GND_net), .I1(n15388[13]), .I2(n1111_adj_4845), 
            .I3(n39644), .O(n14704[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5117_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5061_4 (.CI(n39910), .I0(n14343[1]), .I1(n229), .CO(n39911));
    SB_LUT4 add_5061_3_lut (.I0(GND_net), .I1(n14343[0]), .I2(n156), .I3(n39909), 
            .O(n13544[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5061_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5061_3 (.CI(n39909), .I0(n14343[0]), .I1(n156), .CO(n39910));
    SB_LUT4 add_5061_2_lut (.I0(GND_net), .I1(n14_adj_4844), .I2(n83), 
            .I3(GND_net), .O(n13544[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5061_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5117_16 (.CI(n39644), .I0(n15388[13]), .I1(n1111_adj_4845), 
            .CO(n39645));
    SB_CARRY add_5061_2 (.CI(GND_net), .I0(n14_adj_4844), .I1(n83), .CO(n39909));
    SB_LUT4 add_5099_20_lut (.I0(GND_net), .I1(n15064[17]), .I2(GND_net), 
            .I3(n39908), .O(n14343[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5099_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5099_19_lut (.I0(GND_net), .I1(n15064[16]), .I2(GND_net), 
            .I3(n39907), .O(n14343[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5099_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5099_19 (.CI(n39907), .I0(n15064[16]), .I1(GND_net), 
            .CO(n39908));
    SB_LUT4 add_5099_18_lut (.I0(GND_net), .I1(n15064[15]), .I2(GND_net), 
            .I3(n39906), .O(n14343[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5099_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_12_18 (.CI(n38607), .I0(n106[16]), .I1(n155[16]), .CO(n38608));
    SB_LUT4 add_12_17_lut (.I0(GND_net), .I1(n106[15]), .I2(n155[15]), 
            .I3(n38606), .O(duty_23__N_3936[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_12_17 (.CI(n38606), .I0(n106[15]), .I1(n155[15]), .CO(n38607));
    SB_LUT4 add_5117_15_lut (.I0(GND_net), .I1(n15388[12]), .I2(n1038_adj_4842), 
            .I3(n39643), .O(n14704[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5117_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_12_16_lut (.I0(GND_net), .I1(n106[14]), .I2(n155[14]), 
            .I3(n38605), .O(duty_23__N_3936[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_12_16 (.CI(n38605), .I0(n106[14]), .I1(n155[14]), .CO(n38606));
    SB_LUT4 add_12_15_lut (.I0(GND_net), .I1(n106[13]), .I2(n155[13]), 
            .I3(n38604), .O(duty_23__N_3936[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5117_15 (.CI(n39643), .I0(n15388[12]), .I1(n1038_adj_4842), 
            .CO(n39644));
    SB_CARRY add_5099_18 (.CI(n39906), .I0(n15064[15]), .I1(GND_net), 
            .CO(n39907));
    SB_CARRY add_12_15 (.CI(n38604), .I0(n106[13]), .I1(n155[13]), .CO(n38605));
    SB_LUT4 add_5099_17_lut (.I0(GND_net), .I1(n15064[14]), .I2(GND_net), 
            .I3(n39905), .O(n14343[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5099_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5099_17 (.CI(n39905), .I0(n15064[14]), .I1(GND_net), 
            .CO(n39906));
    SB_LUT4 add_5099_16_lut (.I0(GND_net), .I1(n15064[13]), .I2(n1108), 
            .I3(n39904), .O(n14343[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5099_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5099_16 (.CI(n39904), .I0(n15064[13]), .I1(n1108), .CO(n39905));
    SB_LUT4 add_5117_14_lut (.I0(GND_net), .I1(n15388[11]), .I2(n965_adj_4841), 
            .I3(n39642), .O(n14704[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5117_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5099_15_lut (.I0(GND_net), .I1(n15064[12]), .I2(n1035), 
            .I3(n39903), .O(n14343[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5099_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5099_15 (.CI(n39903), .I0(n15064[12]), .I1(n1035), .CO(n39904));
    SB_LUT4 add_5099_14_lut (.I0(GND_net), .I1(n15064[11]), .I2(n962), 
            .I3(n39902), .O(n14343[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5099_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5117_14 (.CI(n39642), .I0(n15388[11]), .I1(n965_adj_4841), 
            .CO(n39643));
    SB_LUT4 add_5117_13_lut (.I0(GND_net), .I1(n15388[10]), .I2(n892_adj_4840), 
            .I3(n39641), .O(n14704[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5117_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5117_13 (.CI(n39641), .I0(n15388[10]), .I1(n892_adj_4840), 
            .CO(n39642));
    SB_CARRY add_5099_14 (.CI(n39902), .I0(n15064[11]), .I1(n962), .CO(n39903));
    SB_LUT4 add_5117_12_lut (.I0(GND_net), .I1(n15388[9]), .I2(n819_adj_4839), 
            .I3(n39640), .O(n14704[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5117_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5099_13_lut (.I0(GND_net), .I1(n15064[10]), .I2(n889), 
            .I3(n39901), .O(n14343[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5099_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5117_12 (.CI(n39640), .I0(n15388[9]), .I1(n819_adj_4839), 
            .CO(n39641));
    SB_LUT4 add_5117_11_lut (.I0(GND_net), .I1(n15388[8]), .I2(n746_adj_4838), 
            .I3(n39639), .O(n14704[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5117_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5099_13 (.CI(n39901), .I0(n15064[10]), .I1(n889), .CO(n39902));
    SB_LUT4 add_5099_12_lut (.I0(GND_net), .I1(n15064[9]), .I2(n816), 
            .I3(n39900), .O(n14343[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5099_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5099_12 (.CI(n39900), .I0(n15064[9]), .I1(n816), .CO(n39901));
    SB_LUT4 add_5099_11_lut (.I0(GND_net), .I1(n15064[8]), .I2(n743), 
            .I3(n39899), .O(n14343[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5099_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5099_11 (.CI(n39899), .I0(n15064[8]), .I1(n743), .CO(n39900));
    SB_LUT4 add_12_14_lut (.I0(GND_net), .I1(n106[12]), .I2(n155[12]), 
            .I3(n38603), .O(duty_23__N_3936[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5099_10_lut (.I0(GND_net), .I1(n15064[7]), .I2(n670), 
            .I3(n39898), .O(n14343[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5099_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5099_10 (.CI(n39898), .I0(n15064[7]), .I1(n670), .CO(n39899));
    SB_LUT4 add_5099_9_lut (.I0(GND_net), .I1(n15064[6]), .I2(n597), .I3(n39897), 
            .O(n14343[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5099_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5099_9 (.CI(n39897), .I0(n15064[6]), .I1(n597), .CO(n39898));
    SB_LUT4 add_5099_8_lut (.I0(GND_net), .I1(n15064[5]), .I2(n524), .I3(n39896), 
            .O(n14343[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5099_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5099_8 (.CI(n39896), .I0(n15064[5]), .I1(n524), .CO(n39897));
    SB_LUT4 add_5099_7_lut (.I0(GND_net), .I1(n15064[4]), .I2(n451), .I3(n39895), 
            .O(n14343[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5099_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5099_7 (.CI(n39895), .I0(n15064[4]), .I1(n451), .CO(n39896));
    SB_CARRY add_5117_11 (.CI(n39639), .I0(n15388[8]), .I1(n746_adj_4838), 
            .CO(n39640));
    SB_LUT4 add_5099_6_lut (.I0(GND_net), .I1(n15064[3]), .I2(n378), .I3(n39894), 
            .O(n14343[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5099_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5117_10_lut (.I0(GND_net), .I1(n15388[7]), .I2(n673_adj_4837), 
            .I3(n39638), .O(n14704[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5117_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5117_10 (.CI(n39638), .I0(n15388[7]), .I1(n673_adj_4837), 
            .CO(n39639));
    SB_CARRY add_12_14 (.CI(n38603), .I0(n106[12]), .I1(n155[12]), .CO(n38604));
    SB_LUT4 add_5117_9_lut (.I0(GND_net), .I1(n15388[6]), .I2(n600_adj_4836), 
            .I3(n39637), .O(n14704[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5117_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5117_9 (.CI(n39637), .I0(n15388[6]), .I1(n600_adj_4836), 
            .CO(n39638));
    SB_LUT4 add_12_13_lut (.I0(GND_net), .I1(n106[11]), .I2(n155[11]), 
            .I3(n38602), .O(duty_23__N_3936[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5117_8_lut (.I0(GND_net), .I1(n15388[5]), .I2(n527_adj_4835), 
            .I3(n39636), .O(n14704[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5117_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5117_8 (.CI(n39636), .I0(n15388[5]), .I1(n527_adj_4835), 
            .CO(n39637));
    SB_CARRY add_5099_6 (.CI(n39894), .I0(n15064[3]), .I1(n378), .CO(n39895));
    SB_LUT4 add_5099_5_lut (.I0(GND_net), .I1(n15064[2]), .I2(n305), .I3(n39893), 
            .O(n14343[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5099_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5099_5 (.CI(n39893), .I0(n15064[2]), .I1(n305), .CO(n39894));
    SB_LUT4 add_5099_4_lut (.I0(GND_net), .I1(n15064[1]), .I2(n232), .I3(n39892), 
            .O(n14343[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5099_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5117_7_lut (.I0(GND_net), .I1(n15388[4]), .I2(n454_adj_4834), 
            .I3(n39635), .O(n14704[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5117_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5117_7 (.CI(n39635), .I0(n15388[4]), .I1(n454_adj_4834), 
            .CO(n39636));
    SB_CARRY add_12_13 (.CI(n38602), .I0(n106[11]), .I1(n155[11]), .CO(n38603));
    SB_LUT4 mult_10_i559_2_lut (.I0(\Kp[11] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n831_adj_5083));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i559_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5099_4 (.CI(n39892), .I0(n15064[1]), .I1(n232), .CO(n39893));
    SB_LUT4 mult_10_i608_2_lut (.I0(\Kp[12] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n904_adj_5084));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i608_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5099_3_lut (.I0(GND_net), .I1(n15064[0]), .I2(n159), .I3(n39891), 
            .O(n14343[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5099_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5099_3 (.CI(n39891), .I0(n15064[0]), .I1(n159), .CO(n39892));
    SB_LUT4 add_5099_2_lut (.I0(GND_net), .I1(n17), .I2(n86), .I3(GND_net), 
            .O(n14343[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5099_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5117_6_lut (.I0(GND_net), .I1(n15388[3]), .I2(n381_adj_4832), 
            .I3(n39634), .O(n14704[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5117_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5099_2 (.CI(GND_net), .I0(n17), .I1(n86), .CO(n39891));
    SB_CARRY add_5117_6 (.CI(n39634), .I0(n15388[3]), .I1(n381_adj_4832), 
            .CO(n39635));
    SB_LUT4 add_5360_10_lut (.I0(GND_net), .I1(n18784[7]), .I2(n700_adj_4831), 
            .I3(n39890), .O(n18604[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5360_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5360_9_lut (.I0(GND_net), .I1(n18784[6]), .I2(n627_adj_4830), 
            .I3(n39889), .O(n18604[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5360_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5360_9 (.CI(n39889), .I0(n18784[6]), .I1(n627_adj_4830), 
            .CO(n39890));
    SB_LUT4 add_12_12_lut (.I0(GND_net), .I1(n106[10]), .I2(n155[10]), 
            .I3(n38601), .O(duty_23__N_3936[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_12_12 (.CI(n38601), .I0(n106[10]), .I1(n155[10]), .CO(n38602));
    SB_LUT4 add_12_11_lut (.I0(GND_net), .I1(n106[9]), .I2(n155[9]), .I3(n38600), 
            .O(duty_23__N_3936[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5360_8_lut (.I0(GND_net), .I1(n18784[5]), .I2(n554_adj_4829), 
            .I3(n39888), .O(n18604[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5360_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5360_8 (.CI(n39888), .I0(n18784[5]), .I1(n554_adj_4829), 
            .CO(n39889));
    SB_LUT4 add_5117_5_lut (.I0(GND_net), .I1(n15388[2]), .I2(n308_adj_4828), 
            .I3(n39633), .O(n14704[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5117_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5117_5 (.CI(n39633), .I0(n15388[2]), .I1(n308_adj_4828), 
            .CO(n39634));
    SB_LUT4 add_5360_7_lut (.I0(GND_net), .I1(n18784[4]), .I2(n481_adj_4827), 
            .I3(n39887), .O(n18604[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5360_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5360_7 (.CI(n39887), .I0(n18784[4]), .I1(n481_adj_4827), 
            .CO(n39888));
    SB_CARRY add_12_11 (.CI(n38600), .I0(n106[9]), .I1(n155[9]), .CO(n38601));
    SB_LUT4 add_5360_6_lut (.I0(GND_net), .I1(n18784[3]), .I2(n408_adj_4826), 
            .I3(n39886), .O(n18604[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5360_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5360_6 (.CI(n39886), .I0(n18784[3]), .I1(n408_adj_4826), 
            .CO(n39887));
    SB_LUT4 add_12_10_lut (.I0(GND_net), .I1(n106[8]), .I2(n155[8]), .I3(n38599), 
            .O(duty_23__N_3936[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5117_4_lut (.I0(GND_net), .I1(n15388[1]), .I2(n235_adj_4825), 
            .I3(n39632), .O(n14704[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5117_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5360_5_lut (.I0(GND_net), .I1(n18784[2]), .I2(n335_adj_4824), 
            .I3(n39885), .O(n18604[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5360_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5360_5 (.CI(n39885), .I0(n18784[2]), .I1(n335_adj_4824), 
            .CO(n39886));
    SB_LUT4 add_5360_4_lut (.I0(GND_net), .I1(n18784[1]), .I2(n262_adj_4823), 
            .I3(n39884), .O(n18604[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5360_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5360_4 (.CI(n39884), .I0(n18784[1]), .I1(n262_adj_4823), 
            .CO(n39885));
    SB_LUT4 add_5360_3_lut (.I0(GND_net), .I1(n18784[0]), .I2(n189_adj_4822), 
            .I3(n39883), .O(n18604[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5360_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5360_3 (.CI(n39883), .I0(n18784[0]), .I1(n189_adj_4822), 
            .CO(n39884));
    SB_LUT4 add_5360_2_lut (.I0(GND_net), .I1(n47_adj_4821), .I2(n116_adj_4820), 
            .I3(GND_net), .O(n18604[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5360_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5360_2 (.CI(GND_net), .I0(n47_adj_4821), .I1(n116_adj_4820), 
            .CO(n39883));
    SB_LUT4 add_5135_19_lut (.I0(GND_net), .I1(n15711[16]), .I2(GND_net), 
            .I3(n39882), .O(n15064[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5135_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5135_18_lut (.I0(GND_net), .I1(n15711[15]), .I2(GND_net), 
            .I3(n39881), .O(n15064[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5135_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5135_18 (.CI(n39881), .I0(n15711[15]), .I1(GND_net), 
            .CO(n39882));
    SB_CARRY add_12_10 (.CI(n38599), .I0(n106[8]), .I1(n155[8]), .CO(n38600));
    SB_LUT4 add_5135_17_lut (.I0(GND_net), .I1(n15711[14]), .I2(GND_net), 
            .I3(n39880), .O(n15064[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5135_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5135_17 (.CI(n39880), .I0(n15711[14]), .I1(GND_net), 
            .CO(n39881));
    SB_LUT4 add_5135_16_lut (.I0(GND_net), .I1(n15711[13]), .I2(n1111), 
            .I3(n39879), .O(n15064[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5135_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5117_4 (.CI(n39632), .I0(n15388[1]), .I1(n235_adj_4825), 
            .CO(n39633));
    SB_CARRY add_5135_16 (.CI(n39879), .I0(n15711[13]), .I1(n1111), .CO(n39880));
    SB_LUT4 add_5135_15_lut (.I0(GND_net), .I1(n15711[12]), .I2(n1038), 
            .I3(n39878), .O(n15064[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5135_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5135_15 (.CI(n39878), .I0(n15711[12]), .I1(n1038), .CO(n39879));
    SB_LUT4 add_5135_14_lut (.I0(GND_net), .I1(n15711[11]), .I2(n965), 
            .I3(n39877), .O(n15064[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5135_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_12_9_lut (.I0(GND_net), .I1(n106[7]), .I2(n155[7]), .I3(n38598), 
            .O(duty_23__N_3936[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5135_14 (.CI(n39877), .I0(n15711[11]), .I1(n965), .CO(n39878));
    SB_LUT4 add_5135_13_lut (.I0(GND_net), .I1(n15711[10]), .I2(n892), 
            .I3(n39876), .O(n15064[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5135_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5135_13 (.CI(n39876), .I0(n15711[10]), .I1(n892), .CO(n39877));
    SB_LUT4 add_5135_12_lut (.I0(GND_net), .I1(n15711[9]), .I2(n819), 
            .I3(n39875), .O(n15064[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5135_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5135_12 (.CI(n39875), .I0(n15711[9]), .I1(n819), .CO(n39876));
    SB_LUT4 add_5135_11_lut (.I0(GND_net), .I1(n15711[8]), .I2(n746), 
            .I3(n39874), .O(n15064[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5135_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5135_11 (.CI(n39874), .I0(n15711[8]), .I1(n746), .CO(n39875));
    SB_LUT4 add_5135_10_lut (.I0(GND_net), .I1(n15711[7]), .I2(n673), 
            .I3(n39873), .O(n15064[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5135_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5135_10 (.CI(n39873), .I0(n15711[7]), .I1(n673), .CO(n39874));
    SB_LUT4 add_5135_9_lut (.I0(GND_net), .I1(n15711[6]), .I2(n600), .I3(n39872), 
            .O(n15064[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5135_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5135_9 (.CI(n39872), .I0(n15711[6]), .I1(n600), .CO(n39873));
    SB_LUT4 add_5135_8_lut (.I0(GND_net), .I1(n15711[5]), .I2(n527), .I3(n39871), 
            .O(n15064[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5135_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5117_3_lut (.I0(GND_net), .I1(n15388[0]), .I2(n162_adj_4818), 
            .I3(n39631), .O(n14704[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5117_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5117_3 (.CI(n39631), .I0(n15388[0]), .I1(n162_adj_4818), 
            .CO(n39632));
    SB_CARRY add_5135_8 (.CI(n39871), .I0(n15711[5]), .I1(n527), .CO(n39872));
    SB_LUT4 add_5117_2_lut (.I0(GND_net), .I1(n20_adj_4817), .I2(n89_adj_4816), 
            .I3(GND_net), .O(n14704[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5117_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5135_7_lut (.I0(GND_net), .I1(n15711[4]), .I2(n454), .I3(n39870), 
            .O(n15064[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5135_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5135_7 (.CI(n39870), .I0(n15711[4]), .I1(n454), .CO(n39871));
    SB_LUT4 add_5135_6_lut (.I0(GND_net), .I1(n15711[3]), .I2(n381), .I3(n39869), 
            .O(n15064[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5135_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5135_6 (.CI(n39869), .I0(n15711[3]), .I1(n381), .CO(n39870));
    SB_CARRY add_5117_2 (.CI(GND_net), .I0(n20_adj_4817), .I1(n89_adj_4816), 
            .CO(n39631));
    SB_CARRY add_12_9 (.CI(n38598), .I0(n106[7]), .I1(n155[7]), .CO(n38599));
    SB_LUT4 add_5369_10_lut (.I0(GND_net), .I1(n18864[7]), .I2(n700), 
            .I3(n39630), .O(n18703[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5369_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_12_8_lut (.I0(GND_net), .I1(n106[6]), .I2(n155[6]), .I3(n38597), 
            .O(duty_23__N_3936[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5135_5_lut (.I0(GND_net), .I1(n15711[2]), .I2(n308), .I3(n39868), 
            .O(n15064[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5135_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_12_8 (.CI(n38597), .I0(n106[6]), .I1(n155[6]), .CO(n38598));
    SB_CARRY add_5135_5 (.CI(n39868), .I0(n15711[2]), .I1(n308), .CO(n39869));
    SB_LUT4 add_5135_4_lut (.I0(GND_net), .I1(n15711[1]), .I2(n235), .I3(n39867), 
            .O(n15064[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5135_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i555_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n825));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i555_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5135_4 (.CI(n39867), .I0(n15711[1]), .I1(n235), .CO(n39868));
    SB_LUT4 add_5135_3_lut (.I0(GND_net), .I1(n15711[0]), .I2(n162), .I3(n39866), 
            .O(n15064[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5135_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5369_9_lut (.I0(GND_net), .I1(n18864[6]), .I2(n627), .I3(n39629), 
            .O(n18703[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5369_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5369_9 (.CI(n39629), .I0(n18864[6]), .I1(n627), .CO(n39630));
    SB_LUT4 add_5369_8_lut (.I0(GND_net), .I1(n18864[5]), .I2(n554), .I3(n39628), 
            .O(n18703[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5369_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5320_12_lut (.I0(GND_net), .I1(n18384[9]), .I2(n840), 
            .I3(n39492), .O(n18120[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5320_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5320_11_lut (.I0(GND_net), .I1(n18384[8]), .I2(n767), 
            .I3(n39491), .O(n18120[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5320_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5369_8 (.CI(n39628), .I0(n18864[5]), .I1(n554), .CO(n39629));
    SB_CARRY add_5320_11 (.CI(n39491), .I0(n18384[8]), .I1(n767), .CO(n39492));
    SB_LUT4 add_5320_10_lut (.I0(GND_net), .I1(n18384[7]), .I2(n694), 
            .I3(n39490), .O(n18120[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5320_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5369_7_lut (.I0(GND_net), .I1(n18864[4]), .I2(n481), .I3(n39627), 
            .O(n18703[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5369_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_12_7_lut (.I0(GND_net), .I1(n106[5]), .I2(n155[5]), .I3(n38596), 
            .O(duty_23__N_3936[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5320_10 (.CI(n39490), .I0(n18384[7]), .I1(n694), .CO(n39491));
    SB_CARRY add_5369_7 (.CI(n39627), .I0(n18864[4]), .I1(n481), .CO(n39628));
    SB_LUT4 add_5320_9_lut (.I0(GND_net), .I1(n18384[6]), .I2(n621), .I3(n39489), 
            .O(n18120[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5320_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5320_9 (.CI(n39489), .I0(n18384[6]), .I1(n621), .CO(n39490));
    SB_LUT4 add_5320_8_lut (.I0(GND_net), .I1(n18384[5]), .I2(n548), .I3(n39488), 
            .O(n18120[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5320_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5135_3 (.CI(n39866), .I0(n15711[0]), .I1(n162), .CO(n39867));
    SB_LUT4 add_5369_6_lut (.I0(GND_net), .I1(n18864[3]), .I2(n408), .I3(n39626), 
            .O(n18703[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5369_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5320_8 (.CI(n39488), .I0(n18384[5]), .I1(n548), .CO(n39489));
    SB_CARRY add_5369_6 (.CI(n39626), .I0(n18864[3]), .I1(n408), .CO(n39627));
    SB_LUT4 add_5320_7_lut (.I0(GND_net), .I1(n18384[4]), .I2(n475), .I3(n39487), 
            .O(n18120[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5320_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5369_5_lut (.I0(GND_net), .I1(n18864[2]), .I2(n335), .I3(n39625), 
            .O(n18703[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5369_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5320_7 (.CI(n39487), .I0(n18384[4]), .I1(n475), .CO(n39488));
    SB_CARRY add_12_7 (.CI(n38596), .I0(n106[5]), .I1(n155[5]), .CO(n38597));
    SB_CARRY add_5369_5 (.CI(n39625), .I0(n18864[2]), .I1(n335), .CO(n39626));
    SB_LUT4 add_5320_6_lut (.I0(GND_net), .I1(n18384[3]), .I2(n402), .I3(n39486), 
            .O(n18120[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5320_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5135_2_lut (.I0(GND_net), .I1(n20_adj_4815), .I2(n89), 
            .I3(GND_net), .O(n15064[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5135_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5135_2 (.CI(GND_net), .I0(n20_adj_4815), .I1(n89), .CO(n39866));
    SB_LUT4 add_5169_18_lut (.I0(GND_net), .I1(n16288[15]), .I2(GND_net), 
            .I3(n39865), .O(n15711[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5169_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5169_17_lut (.I0(GND_net), .I1(n16288[14]), .I2(GND_net), 
            .I3(n39864), .O(n15711[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5169_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5169_17 (.CI(n39864), .I0(n16288[14]), .I1(GND_net), 
            .CO(n39865));
    SB_LUT4 add_5369_4_lut (.I0(GND_net), .I1(n18864[1]), .I2(n262), .I3(n39624), 
            .O(n18703[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5369_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5320_6 (.CI(n39486), .I0(n18384[3]), .I1(n402), .CO(n39487));
    SB_CARRY add_5369_4 (.CI(n39624), .I0(n18864[1]), .I1(n262), .CO(n39625));
    SB_LUT4 add_5369_3_lut (.I0(GND_net), .I1(n18864[0]), .I2(n189), .I3(n39623), 
            .O(n18703[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5369_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5320_5_lut (.I0(GND_net), .I1(n18384[2]), .I2(n329), .I3(n39485), 
            .O(n18120[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5320_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5369_3 (.CI(n39623), .I0(n18864[0]), .I1(n189), .CO(n39624));
    SB_CARRY add_5320_5 (.CI(n39485), .I0(n18384[2]), .I1(n329), .CO(n39486));
    SB_LUT4 add_5320_4_lut (.I0(GND_net), .I1(n18384[1]), .I2(n256), .I3(n39484), 
            .O(n18120[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5320_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5169_16_lut (.I0(GND_net), .I1(n16288[13]), .I2(n1114), 
            .I3(n39863), .O(n15711[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5169_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5369_2_lut (.I0(GND_net), .I1(n47), .I2(n116), .I3(GND_net), 
            .O(n18703[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5369_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5169_16 (.CI(n39863), .I0(n16288[13]), .I1(n1114), .CO(n39864));
    SB_LUT4 add_5169_15_lut (.I0(GND_net), .I1(n16288[12]), .I2(n1041), 
            .I3(n39862), .O(n15711[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5169_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5169_15 (.CI(n39862), .I0(n16288[12]), .I1(n1041), .CO(n39863));
    SB_LUT4 add_5169_14_lut (.I0(GND_net), .I1(n16288[11]), .I2(n968), 
            .I3(n39861), .O(n15711[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5169_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5169_14 (.CI(n39861), .I0(n16288[11]), .I1(n968), .CO(n39862));
    SB_LUT4 add_5169_13_lut (.I0(GND_net), .I1(n16288[10]), .I2(n895), 
            .I3(n39860), .O(n15711[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5169_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5169_13 (.CI(n39860), .I0(n16288[10]), .I1(n895), .CO(n39861));
    SB_LUT4 add_5169_12_lut (.I0(GND_net), .I1(n16288[9]), .I2(n822), 
            .I3(n39859), .O(n15711[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5169_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5169_12 (.CI(n39859), .I0(n16288[9]), .I1(n822), .CO(n39860));
    SB_LUT4 add_12_6_lut (.I0(GND_net), .I1(n106[4]), .I2(n155[4]), .I3(n38595), 
            .O(duty_23__N_3936[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5169_11_lut (.I0(GND_net), .I1(n16288[8]), .I2(n749), 
            .I3(n39858), .O(n15711[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5169_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5169_11 (.CI(n39858), .I0(n16288[8]), .I1(n749), .CO(n39859));
    SB_LUT4 add_5169_10_lut (.I0(GND_net), .I1(n16288[7]), .I2(n676), 
            .I3(n39857), .O(n15711[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5169_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5169_10 (.CI(n39857), .I0(n16288[7]), .I1(n676), .CO(n39858));
    SB_LUT4 add_5169_9_lut (.I0(GND_net), .I1(n16288[6]), .I2(n603), .I3(n39856), 
            .O(n15711[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5169_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5169_9 (.CI(n39856), .I0(n16288[6]), .I1(n603), .CO(n39857));
    SB_LUT4 add_5169_8_lut (.I0(GND_net), .I1(n16288[5]), .I2(n530), .I3(n39855), 
            .O(n15711[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5169_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5169_8 (.CI(n39855), .I0(n16288[5]), .I1(n530), .CO(n39856));
    SB_LUT4 add_5169_7_lut (.I0(GND_net), .I1(n16288[4]), .I2(n457), .I3(n39854), 
            .O(n15711[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5169_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5369_2 (.CI(GND_net), .I0(n47), .I1(n116), .CO(n39623));
    SB_CARRY add_5169_7 (.CI(n39854), .I0(n16288[4]), .I1(n457), .CO(n39855));
    SB_CARRY add_5320_4 (.CI(n39484), .I0(n18384[1]), .I1(n256), .CO(n39485));
    SB_LUT4 add_5169_6_lut (.I0(GND_net), .I1(n16288[3]), .I2(n384), .I3(n39853), 
            .O(n15711[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5169_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5169_6 (.CI(n39853), .I0(n16288[3]), .I1(n384), .CO(n39854));
    SB_LUT4 add_5320_3_lut (.I0(GND_net), .I1(n18384[0]), .I2(n183_adj_5087), 
            .I3(n39483), .O(n18120[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5320_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5169_5_lut (.I0(GND_net), .I1(n16288[2]), .I2(n311), .I3(n39852), 
            .O(n15711[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5169_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_12_6 (.CI(n38595), .I0(n106[4]), .I1(n155[4]), .CO(n38596));
    SB_CARRY add_5169_5 (.CI(n39852), .I0(n16288[2]), .I1(n311), .CO(n39853));
    SB_LUT4 add_5169_4_lut (.I0(GND_net), .I1(n16288[1]), .I2(n238), .I3(n39851), 
            .O(n15711[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5169_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5169_4 (.CI(n39851), .I0(n16288[1]), .I1(n238), .CO(n39852));
    SB_LUT4 add_5169_3_lut (.I0(GND_net), .I1(n16288[0]), .I2(n165), .I3(n39850), 
            .O(n15711[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5169_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5169_3 (.CI(n39850), .I0(n16288[0]), .I1(n165), .CO(n39851));
    SB_LUT4 add_5169_2_lut (.I0(GND_net), .I1(n23_adj_5088), .I2(n92), 
            .I3(GND_net), .O(n15711[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5169_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5169_2 (.CI(GND_net), .I0(n23_adj_5088), .I1(n92), .CO(n39850));
    SB_LUT4 add_5377_9_lut (.I0(GND_net), .I1(n18928[6]), .I2(n630_adj_5089), 
            .I3(n39849), .O(n18784[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5377_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_12_5_lut (.I0(GND_net), .I1(n106[3]), .I2(n155[3]), .I3(n38594), 
            .O(duty_23__N_3936[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5152_18_lut (.I0(GND_net), .I1(n16000[15]), .I2(GND_net), 
            .I3(n39622), .O(n15388[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5152_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_12_5 (.CI(n38594), .I0(n106[3]), .I1(n155[3]), .CO(n38595));
    SB_LUT4 add_5377_8_lut (.I0(GND_net), .I1(n18928[5]), .I2(n557_adj_5090), 
            .I3(n39848), .O(n18784[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5377_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5377_8 (.CI(n39848), .I0(n18928[5]), .I1(n557_adj_5090), 
            .CO(n39849));
    SB_LUT4 add_5377_7_lut (.I0(GND_net), .I1(n18928[4]), .I2(n484_adj_5091), 
            .I3(n39847), .O(n18784[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5377_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5377_7 (.CI(n39847), .I0(n18928[4]), .I1(n484_adj_5091), 
            .CO(n39848));
    SB_LUT4 add_5377_6_lut (.I0(GND_net), .I1(n18928[3]), .I2(n411_adj_5092), 
            .I3(n39846), .O(n18784[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5377_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5377_6 (.CI(n39846), .I0(n18928[3]), .I1(n411_adj_5092), 
            .CO(n39847));
    SB_LUT4 add_5377_5_lut (.I0(GND_net), .I1(n18928[2]), .I2(n338_adj_5093), 
            .I3(n39845), .O(n18784[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5377_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5377_5 (.CI(n39845), .I0(n18928[2]), .I1(n338_adj_5093), 
            .CO(n39846));
    SB_LUT4 add_5377_4_lut (.I0(GND_net), .I1(n18928[1]), .I2(n265_adj_5094), 
            .I3(n39844), .O(n18784[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5377_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5377_4 (.CI(n39844), .I0(n18928[1]), .I1(n265_adj_5094), 
            .CO(n39845));
    SB_LUT4 add_5341_11_lut (.I0(GND_net), .I1(n18604[8]), .I2(n770_adj_5095), 
            .I3(n38820), .O(n18384[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5341_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5377_3_lut (.I0(GND_net), .I1(n18928[0]), .I2(n192_adj_5096), 
            .I3(n39843), .O(n18784[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5377_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5377_3 (.CI(n39843), .I0(n18928[0]), .I1(n192_adj_5096), 
            .CO(n39844));
    SB_LUT4 add_12_4_lut (.I0(GND_net), .I1(n106[2]), .I2(n155[2]), .I3(n38593), 
            .O(duty_23__N_3936[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5152_17_lut (.I0(GND_net), .I1(n16000[14]), .I2(GND_net), 
            .I3(n39621), .O(n15388[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5152_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5320_3 (.CI(n39483), .I0(n18384[0]), .I1(n183_adj_5087), 
            .CO(n39484));
    SB_LUT4 add_5320_2_lut (.I0(GND_net), .I1(n41_adj_5097), .I2(n110_adj_5098), 
            .I3(GND_net), .O(n18120[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5320_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_12_4 (.CI(n38593), .I0(n106[2]), .I1(n155[2]), .CO(n38594));
    SB_LUT4 add_5341_10_lut (.I0(GND_net), .I1(n18604[7]), .I2(n697_adj_5099), 
            .I3(n38819), .O(n18384[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5341_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5377_2_lut (.I0(GND_net), .I1(n50_adj_5100), .I2(n119_adj_5101), 
            .I3(GND_net), .O(n18784[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5377_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5320_2 (.CI(GND_net), .I0(n41_adj_5097), .I1(n110_adj_5098), 
            .CO(n39483));
    SB_CARRY add_5152_17 (.CI(n39621), .I0(n16000[14]), .I1(GND_net), 
            .CO(n39622));
    SB_LUT4 add_12_3_lut (.I0(GND_net), .I1(n106[1]), .I2(n155[1]), .I3(n38592), 
            .O(duty_23__N_3936[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5341_10 (.CI(n38819), .I0(n18604[7]), .I1(n697_adj_5099), 
            .CO(n38820));
    SB_CARRY add_12_3 (.CI(n38592), .I0(n106[1]), .I1(n155[1]), .CO(n38593));
    SB_LUT4 add_5152_16_lut (.I0(GND_net), .I1(n16000[13]), .I2(n1114_adj_5102), 
            .I3(n39620), .O(n15388[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5152_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5152_16 (.CI(n39620), .I0(n16000[13]), .I1(n1114_adj_5102), 
            .CO(n39621));
    SB_CARRY add_5377_2 (.CI(GND_net), .I0(n50_adj_5100), .I1(n119_adj_5101), 
            .CO(n39843));
    SB_LUT4 add_5341_9_lut (.I0(GND_net), .I1(n18604[6]), .I2(n624_adj_5103), 
            .I3(n38818), .O(n18384[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5341_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5341_9 (.CI(n38818), .I0(n18604[6]), .I1(n624_adj_5103), 
            .CO(n38819));
    SB_LUT4 add_5152_15_lut (.I0(GND_net), .I1(n16000[12]), .I2(n1041_adj_5104), 
            .I3(n39619), .O(n15388[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5152_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5201_17_lut (.I0(GND_net), .I1(n16799[14]), .I2(GND_net), 
            .I3(n39842), .O(n16288[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5201_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5201_16_lut (.I0(GND_net), .I1(n16799[13]), .I2(n1117), 
            .I3(n39841), .O(n16288[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5201_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5201_16 (.CI(n39841), .I0(n16799[13]), .I1(n1117), .CO(n39842));
    SB_LUT4 add_5201_15_lut (.I0(GND_net), .I1(n16799[12]), .I2(n1044), 
            .I3(n39840), .O(n16288[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5201_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5341_8_lut (.I0(GND_net), .I1(n18604[5]), .I2(n551_adj_5105), 
            .I3(n38817), .O(n18384[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5341_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5341_8 (.CI(n38817), .I0(n18604[5]), .I1(n551_adj_5105), 
            .CO(n38818));
    SB_CARRY add_5152_15 (.CI(n39619), .I0(n16000[12]), .I1(n1041_adj_5104), 
            .CO(n39620));
    SB_CARRY add_5201_15 (.CI(n39840), .I0(n16799[12]), .I1(n1044), .CO(n39841));
    SB_LUT4 add_5341_7_lut (.I0(GND_net), .I1(n18604[4]), .I2(n478_adj_5106), 
            .I3(n38816), .O(n18384[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5341_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5341_7 (.CI(n38816), .I0(n18604[4]), .I1(n478_adj_5106), 
            .CO(n38817));
    SB_LUT4 add_12_2_lut (.I0(GND_net), .I1(n106[0]), .I2(n155[0]), .I3(GND_net), 
            .O(duty_23__N_3936[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5341_6_lut (.I0(GND_net), .I1(n18604[3]), .I2(n405_adj_5107), 
            .I3(n38815), .O(n18384[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5341_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5152_14_lut (.I0(GND_net), .I1(n16000[11]), .I2(n968_adj_5108), 
            .I3(n39618), .O(n15388[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5152_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_12_2 (.CI(GND_net), .I0(n106[0]), .I1(n155[0]), .CO(n38592));
    SB_LUT4 add_5201_14_lut (.I0(GND_net), .I1(n16799[11]), .I2(n971), 
            .I3(n39839), .O(n16288[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5201_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5341_6 (.CI(n38815), .I0(n18604[3]), .I1(n405_adj_5107), 
            .CO(n38816));
    SB_CARRY add_5201_14 (.CI(n39839), .I0(n16799[11]), .I1(n971), .CO(n39840));
    SB_LUT4 add_5341_5_lut (.I0(GND_net), .I1(n18604[2]), .I2(n332_adj_5109), 
            .I3(n38814), .O(n18384[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5341_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5341_5 (.CI(n38814), .I0(n18604[2]), .I1(n332_adj_5109), 
            .CO(n38815));
    SB_LUT4 add_5201_13_lut (.I0(GND_net), .I1(n16799[10]), .I2(n898), 
            .I3(n39838), .O(n16288[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5201_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5341_4_lut (.I0(GND_net), .I1(n18604[1]), .I2(n259_adj_5110), 
            .I3(n38813), .O(n18384[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5341_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5341_4 (.CI(n38813), .I0(n18604[1]), .I1(n259_adj_5110), 
            .CO(n38814));
    SB_CARRY add_5201_13 (.CI(n39838), .I0(n16799[10]), .I1(n898), .CO(n39839));
    SB_LUT4 add_5201_12_lut (.I0(GND_net), .I1(n16799[9]), .I2(n825_adj_5111), 
            .I3(n39837), .O(n16288[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5201_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5201_12 (.CI(n39837), .I0(n16799[9]), .I1(n825_adj_5111), 
            .CO(n39838));
    SB_LUT4 add_5201_11_lut (.I0(GND_net), .I1(n16799[8]), .I2(n752_adj_5112), 
            .I3(n39836), .O(n16288[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5201_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5201_11 (.CI(n39836), .I0(n16799[8]), .I1(n752_adj_5112), 
            .CO(n39837));
    SB_LUT4 add_5341_3_lut (.I0(GND_net), .I1(n18604[0]), .I2(n186_adj_5113), 
            .I3(n38812), .O(n18384[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5341_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5152_14 (.CI(n39618), .I0(n16000[11]), .I1(n968_adj_5108), 
            .CO(n39619));
    SB_CARRY add_5341_3 (.CI(n38812), .I0(n18604[0]), .I1(n186_adj_5113), 
            .CO(n38813));
    SB_LUT4 add_5341_2_lut (.I0(GND_net), .I1(n44_adj_5114), .I2(n113_adj_5115), 
            .I3(GND_net), .O(n18384[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5341_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5152_13_lut (.I0(GND_net), .I1(n16000[10]), .I2(n895_adj_5116), 
            .I3(n39617), .O(n15388[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5152_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5152_13 (.CI(n39617), .I0(n16000[10]), .I1(n895_adj_5116), 
            .CO(n39618));
    SB_LUT4 add_5152_12_lut (.I0(GND_net), .I1(n16000[9]), .I2(n822_adj_5117), 
            .I3(n39616), .O(n15388[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5152_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5201_10_lut (.I0(GND_net), .I1(n16799[7]), .I2(n679_adj_5118), 
            .I3(n39835), .O(n16288[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5201_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5152_12 (.CI(n39616), .I0(n16000[9]), .I1(n822_adj_5117), 
            .CO(n39617));
    SB_LUT4 add_5152_11_lut (.I0(GND_net), .I1(n16000[8]), .I2(n749_adj_5119), 
            .I3(n39615), .O(n15388[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5152_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5152_11 (.CI(n39615), .I0(n16000[8]), .I1(n749_adj_5119), 
            .CO(n39616));
    SB_CARRY add_5341_2 (.CI(GND_net), .I0(n44_adj_5114), .I1(n113_adj_5115), 
            .CO(n38812));
    SB_LUT4 add_5152_10_lut (.I0(GND_net), .I1(n16000[7]), .I2(n676_adj_5120), 
            .I3(n39614), .O(n15388[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5152_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5152_10 (.CI(n39614), .I0(n16000[7]), .I1(n676_adj_5120), 
            .CO(n39615));
    SB_LUT4 add_5152_9_lut (.I0(GND_net), .I1(n16000[6]), .I2(n603_adj_5121), 
            .I3(n39613), .O(n15388[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5152_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5152_9 (.CI(n39613), .I0(n16000[6]), .I1(n603_adj_5121), 
            .CO(n39614));
    SB_LUT4 mult_11_i647_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n962_adj_5026));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i647_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5152_8_lut (.I0(GND_net), .I1(n16000[5]), .I2(n530_adj_5122), 
            .I3(n39612), .O(n15388[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5152_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5201_10 (.CI(n39835), .I0(n16799[7]), .I1(n679_adj_5118), 
            .CO(n39836));
    SB_CARRY add_5152_8 (.CI(n39612), .I0(n16000[5]), .I1(n530_adj_5122), 
            .CO(n39613));
    SB_LUT4 add_5201_9_lut (.I0(GND_net), .I1(n16799[6]), .I2(n606_adj_5123), 
            .I3(n39834), .O(n16288[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5201_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5201_9 (.CI(n39834), .I0(n16799[6]), .I1(n606_adj_5123), 
            .CO(n39835));
    SB_LUT4 add_5201_8_lut (.I0(GND_net), .I1(n16799[5]), .I2(n533_adj_5124), 
            .I3(n39833), .O(n16288[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5201_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5201_8 (.CI(n39833), .I0(n16799[5]), .I1(n533_adj_5124), 
            .CO(n39834));
    SB_LUT4 add_5201_7_lut (.I0(GND_net), .I1(n16799[4]), .I2(n460_adj_5125), 
            .I3(n39832), .O(n16288[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5201_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5201_7 (.CI(n39832), .I0(n16799[4]), .I1(n460_adj_5125), 
            .CO(n39833));
    SB_LUT4 add_5201_6_lut (.I0(GND_net), .I1(n16799[3]), .I2(n387_adj_5126), 
            .I3(n39831), .O(n16288[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5201_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5201_6 (.CI(n39831), .I0(n16799[3]), .I1(n387_adj_5126), 
            .CO(n39832));
    SB_LUT4 add_5201_5_lut (.I0(GND_net), .I1(n16799[2]), .I2(n314_adj_5127), 
            .I3(n39830), .O(n16288[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5201_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5201_5 (.CI(n39830), .I0(n16799[2]), .I1(n314_adj_5127), 
            .CO(n39831));
    SB_LUT4 add_5201_4_lut (.I0(GND_net), .I1(n16799[1]), .I2(n241_adj_5128), 
            .I3(n39829), .O(n16288[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5201_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5201_4 (.CI(n39829), .I0(n16799[1]), .I1(n241_adj_5128), 
            .CO(n39830));
    SB_LUT4 add_5152_7_lut (.I0(GND_net), .I1(n16000[4]), .I2(n457_adj_5129), 
            .I3(n39611), .O(n15388[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5152_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5201_3_lut (.I0(GND_net), .I1(n16799[0]), .I2(n168_adj_5130), 
            .I3(n39828), .O(n16288[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5201_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5152_7 (.CI(n39611), .I0(n16000[4]), .I1(n457_adj_5129), 
            .CO(n39612));
    SB_CARRY add_5201_3 (.CI(n39828), .I0(n16799[0]), .I1(n168_adj_5130), 
            .CO(n39829));
    SB_LUT4 add_5152_6_lut (.I0(GND_net), .I1(n16000[3]), .I2(n384_adj_5131), 
            .I3(n39610), .O(n15388[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5152_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5201_2_lut (.I0(GND_net), .I1(n26_adj_5132), .I2(n95_adj_5133), 
            .I3(GND_net), .O(n16288[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5201_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5201_2 (.CI(GND_net), .I0(n26_adj_5132), .I1(n95_adj_5133), 
            .CO(n39828));
    SB_LUT4 add_5231_16_lut (.I0(GND_net), .I1(n17248[13]), .I2(n1120_adj_5134), 
            .I3(n39827), .O(n16799[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5231_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5231_15_lut (.I0(GND_net), .I1(n17248[12]), .I2(n1047_adj_5135), 
            .I3(n39826), .O(n16799[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5231_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5231_15 (.CI(n39826), .I0(n17248[12]), .I1(n1047_adj_5135), 
            .CO(n39827));
    SB_LUT4 add_5231_14_lut (.I0(GND_net), .I1(n17248[11]), .I2(n974_adj_5136), 
            .I3(n39825), .O(n16799[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5231_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5231_14 (.CI(n39825), .I0(n17248[11]), .I1(n974_adj_5136), 
            .CO(n39826));
    SB_LUT4 add_5231_13_lut (.I0(GND_net), .I1(n17248[10]), .I2(n901_adj_5137), 
            .I3(n39824), .O(n16799[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5231_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5231_13 (.CI(n39824), .I0(n17248[10]), .I1(n901_adj_5137), 
            .CO(n39825));
    SB_LUT4 add_5231_12_lut (.I0(GND_net), .I1(n17248[9]), .I2(n828_adj_5138), 
            .I3(n39823), .O(n16799[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5231_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5231_12 (.CI(n39823), .I0(n17248[9]), .I1(n828_adj_5138), 
            .CO(n39824));
    SB_LUT4 add_5231_11_lut (.I0(GND_net), .I1(n17248[8]), .I2(n755_adj_5139), 
            .I3(n39822), .O(n16799[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5231_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5152_6 (.CI(n39610), .I0(n16000[3]), .I1(n384_adj_5131), 
            .CO(n39611));
    SB_CARRY add_5231_11 (.CI(n39822), .I0(n17248[8]), .I1(n755_adj_5139), 
            .CO(n39823));
    SB_LUT4 add_5231_10_lut (.I0(GND_net), .I1(n17248[7]), .I2(n682_adj_5140), 
            .I3(n39821), .O(n16799[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5231_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5152_5_lut (.I0(GND_net), .I1(n16000[2]), .I2(n311_adj_5141), 
            .I3(n39609), .O(n15388[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5152_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5152_5 (.CI(n39609), .I0(n16000[2]), .I1(n311_adj_5141), 
            .CO(n39610));
    SB_CARRY add_5231_10 (.CI(n39821), .I0(n17248[7]), .I1(n682_adj_5140), 
            .CO(n39822));
    SB_LUT4 add_5231_9_lut (.I0(GND_net), .I1(n17248[6]), .I2(n609_adj_5142), 
            .I3(n39820), .O(n16799[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5231_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5231_9 (.CI(n39820), .I0(n17248[6]), .I1(n609_adj_5142), 
            .CO(n39821));
    SB_LUT4 i33955_3_lut_4_lut (.I0(duty_23__N_3936[3]), .I1(n257[3]), .I2(n257[2]), 
            .I3(duty_23__N_3936[2]), .O(n49542));   // verilog/motorControl.v(38[19:35])
    defparam i33955_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 add_5152_4_lut (.I0(GND_net), .I1(n16000[1]), .I2(n238_adj_5143), 
            .I3(n39608), .O(n15388[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5152_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5231_8_lut (.I0(GND_net), .I1(n17248[5]), .I2(n536_adj_5144), 
            .I3(n39819), .O(n16799[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5231_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5231_8 (.CI(n39819), .I0(n17248[5]), .I1(n536_adj_5144), 
            .CO(n39820));
    SB_LUT4 add_5231_7_lut (.I0(GND_net), .I1(n17248[4]), .I2(n463_adj_5145), 
            .I3(n39818), .O(n16799[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5231_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5231_7 (.CI(n39818), .I0(n17248[4]), .I1(n463_adj_5145), 
            .CO(n39819));
    SB_LUT4 add_5231_6_lut (.I0(GND_net), .I1(n17248[3]), .I2(n390_adj_5146), 
            .I3(n39817), .O(n16799[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5231_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5231_6 (.CI(n39817), .I0(n17248[3]), .I1(n390_adj_5146), 
            .CO(n39818));
    SB_LUT4 add_5231_5_lut (.I0(GND_net), .I1(n17248[2]), .I2(n317_adj_5147), 
            .I3(n39816), .O(n16799[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5231_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5231_5 (.CI(n39816), .I0(n17248[2]), .I1(n317_adj_5147), 
            .CO(n39817));
    SB_LUT4 add_5231_4_lut (.I0(GND_net), .I1(n17248[1]), .I2(n244_adj_5148), 
            .I3(n39815), .O(n16799[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5231_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5231_4 (.CI(n39815), .I0(n17248[1]), .I1(n244_adj_5148), 
            .CO(n39816));
    SB_LUT4 add_5231_3_lut (.I0(GND_net), .I1(n17248[0]), .I2(n171_adj_5149), 
            .I3(n39814), .O(n16799[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5231_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5231_3 (.CI(n39814), .I0(n17248[0]), .I1(n171_adj_5149), 
            .CO(n39815));
    SB_LUT4 add_5231_2_lut (.I0(GND_net), .I1(n29_adj_5150), .I2(n98_adj_5151), 
            .I3(GND_net), .O(n16799[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5231_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5231_2 (.CI(GND_net), .I0(n29_adj_5150), .I1(n98_adj_5151), 
            .CO(n39814));
    SB_LUT4 add_5392_8_lut (.I0(GND_net), .I1(n19040[5]), .I2(n560_adj_5152), 
            .I3(n39813), .O(n18928[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5392_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5392_7_lut (.I0(GND_net), .I1(n19040[4]), .I2(n487_adj_5153), 
            .I3(n39812), .O(n18928[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5392_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5392_7 (.CI(n39812), .I0(n19040[4]), .I1(n487_adj_5153), 
            .CO(n39813));
    SB_LUT4 LessThan_15_i6_3_lut_3_lut (.I0(duty_23__N_3936[3]), .I1(n257[3]), 
            .I2(n257[2]), .I3(GND_net), .O(n6_adj_5154));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 mult_11_i604_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n898_adj_5155));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i604_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5152_4 (.CI(n39608), .I0(n16000[1]), .I1(n238_adj_5143), 
            .CO(n39609));
    SB_LUT4 add_5392_6_lut (.I0(GND_net), .I1(n19040[3]), .I2(n414_adj_5156), 
            .I3(n39811), .O(n18928[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5392_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5392_6 (.CI(n39811), .I0(n19040[3]), .I1(n414_adj_5156), 
            .CO(n39812));
    SB_LUT4 add_5392_5_lut (.I0(GND_net), .I1(n19040[2]), .I2(n341_adj_5157), 
            .I3(n39810), .O(n18928[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5392_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5392_5 (.CI(n39810), .I0(n19040[2]), .I1(n341_adj_5157), 
            .CO(n39811));
    SB_LUT4 add_5392_4_lut (.I0(GND_net), .I1(n19040[1]), .I2(n268_adj_5158), 
            .I3(n39809), .O(n18928[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5392_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5392_4 (.CI(n39809), .I0(n19040[1]), .I1(n268_adj_5158), 
            .CO(n39810));
    SB_LUT4 add_5152_3_lut (.I0(GND_net), .I1(n16000[0]), .I2(n165_adj_5159), 
            .I3(n39607), .O(n15388[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5152_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5392_3_lut (.I0(GND_net), .I1(n19040[0]), .I2(n195_adj_5160), 
            .I3(n39808), .O(n18928[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5392_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5392_3 (.CI(n39808), .I0(n19040[0]), .I1(n195_adj_5160), 
            .CO(n39809));
    SB_LUT4 add_5392_2_lut (.I0(GND_net), .I1(n53_adj_5161), .I2(n122_adj_5162), 
            .I3(GND_net), .O(n18928[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5392_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5392_2 (.CI(GND_net), .I0(n53_adj_5161), .I1(n122_adj_5162), 
            .CO(n39808));
    SB_LUT4 add_5259_15_lut (.I0(GND_net), .I1(n17639[12]), .I2(n1050_adj_5163), 
            .I3(n39807), .O(n17248[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5259_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5259_14_lut (.I0(GND_net), .I1(n17639[11]), .I2(n977_adj_5164), 
            .I3(n39806), .O(n17248[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5259_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i33994_3_lut_4_lut (.I0(PWMLimit[3]), .I1(duty_23__N_3936[3]), 
            .I2(duty_23__N_3936[2]), .I3(PWMLimit[2]), .O(n49581));   // verilog/motorControl.v(36[10:25])
    defparam i33994_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_CARRY add_5152_3 (.CI(n39607), .I0(n16000[0]), .I1(n165_adj_5159), 
            .CO(n39608));
    SB_LUT4 add_5152_2_lut (.I0(GND_net), .I1(n23_adj_5165), .I2(n92_adj_5166), 
            .I3(GND_net), .O(n15388[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5152_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5152_2 (.CI(GND_net), .I0(n23_adj_5165), .I1(n92_adj_5166), 
            .CO(n39607));
    SB_CARRY add_5259_14 (.CI(n39806), .I0(n17639[11]), .I1(n977_adj_5164), 
            .CO(n39807));
    SB_LUT4 add_5185_17_lut (.I0(GND_net), .I1(n16544[14]), .I2(GND_net), 
            .I3(n39606), .O(n16000[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5185_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5185_16_lut (.I0(GND_net), .I1(n16544[13]), .I2(n1117_adj_5167), 
            .I3(n39605), .O(n16000[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5185_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5185_16 (.CI(n39605), .I0(n16544[13]), .I1(n1117_adj_5167), 
            .CO(n39606));
    SB_LUT4 add_5185_15_lut (.I0(GND_net), .I1(n16544[12]), .I2(n1044_adj_5168), 
            .I3(n39604), .O(n16000[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5185_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5185_15 (.CI(n39604), .I0(n16544[12]), .I1(n1044_adj_5168), 
            .CO(n39605));
    SB_LUT4 add_5185_14_lut (.I0(GND_net), .I1(n16544[11]), .I2(n971_adj_5169), 
            .I3(n39603), .O(n16000[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5185_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5185_14 (.CI(n39603), .I0(n16544[11]), .I1(n971_adj_5169), 
            .CO(n39604));
    SB_LUT4 add_5185_13_lut (.I0(GND_net), .I1(n16544[10]), .I2(n898_adj_5155), 
            .I3(n39602), .O(n16000[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5185_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5185_13 (.CI(n39602), .I0(n16544[10]), .I1(n898_adj_5155), 
            .CO(n39603));
    SB_LUT4 add_5185_12_lut (.I0(GND_net), .I1(n16544[9]), .I2(n825), 
            .I3(n39601), .O(n16000[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5185_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5259_13_lut (.I0(GND_net), .I1(n17639[10]), .I2(n904_adj_5084), 
            .I3(n39805), .O(n17248[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5259_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5259_13 (.CI(n39805), .I0(n17639[10]), .I1(n904_adj_5084), 
            .CO(n39806));
    SB_CARRY add_5185_12 (.CI(n39601), .I0(n16544[9]), .I1(n825), .CO(n39602));
    SB_LUT4 add_5259_12_lut (.I0(GND_net), .I1(n17639[9]), .I2(n831_adj_5083), 
            .I3(n39804), .O(n17248[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5259_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5185_11_lut (.I0(GND_net), .I1(n16544[8]), .I2(n752), 
            .I3(n39600), .O(n16000[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5185_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5259_12 (.CI(n39804), .I0(n17639[9]), .I1(n831_adj_5083), 
            .CO(n39805));
    SB_LUT4 add_5259_11_lut (.I0(GND_net), .I1(n17639[8]), .I2(n758_adj_5079), 
            .I3(n39803), .O(n17248[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5259_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5259_11 (.CI(n39803), .I0(n17639[8]), .I1(n758_adj_5079), 
            .CO(n39804));
    SB_LUT4 add_5259_10_lut (.I0(GND_net), .I1(n17639[7]), .I2(n685_adj_5078), 
            .I3(n39802), .O(n17248[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5259_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5185_11 (.CI(n39600), .I0(n16544[8]), .I1(n752), .CO(n39601));
    SB_CARRY add_5259_10 (.CI(n39802), .I0(n17639[7]), .I1(n685_adj_5078), 
            .CO(n39803));
    SB_LUT4 duty_23__I_937_i6_3_lut_3_lut (.I0(PWMLimit[3]), .I1(duty_23__N_3936[3]), 
            .I2(duty_23__N_3936[2]), .I3(GND_net), .O(n6_adj_5170));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_937_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 unary_minus_16_add_3_25_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5235[23]), 
            .I3(n38775), .O(n257[23])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_add_3_24_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5235[22]), 
            .I3(n38774), .O(n257[22])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5259_9_lut (.I0(GND_net), .I1(n17639[6]), .I2(n612_adj_5075), 
            .I3(n39801), .O(n17248[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5259_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5259_9 (.CI(n39801), .I0(n17639[6]), .I1(n612_adj_5075), 
            .CO(n39802));
    SB_LUT4 add_5185_10_lut (.I0(GND_net), .I1(n16544[7]), .I2(n679), 
            .I3(n39599), .O(n16000[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5185_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5259_8_lut (.I0(GND_net), .I1(n17639[5]), .I2(n539_adj_5074), 
            .I3(n39800), .O(n17248[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5259_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5259_8 (.CI(n39800), .I0(n17639[5]), .I1(n539_adj_5074), 
            .CO(n39801));
    SB_LUT4 add_5259_7_lut (.I0(GND_net), .I1(n17639[4]), .I2(n466_adj_5073), 
            .I3(n39799), .O(n17248[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5259_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_24 (.CI(n38774), .I0(GND_net), .I1(n1_adj_5235[22]), 
            .CO(n38775));
    SB_CARRY add_5259_7 (.CI(n39799), .I0(n17639[4]), .I1(n466_adj_5073), 
            .CO(n39800));
    SB_LUT4 add_5259_6_lut (.I0(GND_net), .I1(n17639[3]), .I2(n393_adj_5071), 
            .I3(n39798), .O(n17248[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5259_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_add_3_23_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5235[21]), 
            .I3(n38773), .O(n257[21])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5259_6 (.CI(n39798), .I0(n17639[3]), .I1(n393_adj_5071), 
            .CO(n39799));
    SB_CARRY unary_minus_16_add_3_23 (.CI(n38773), .I0(GND_net), .I1(n1_adj_5235[21]), 
            .CO(n38774));
    SB_LUT4 add_5259_5_lut (.I0(GND_net), .I1(n17639[2]), .I2(n320_adj_5069), 
            .I3(n39797), .O(n17248[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5259_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_add_3_22_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5235[20]), 
            .I3(n38772), .O(n257[20])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5259_5 (.CI(n39797), .I0(n17639[2]), .I1(n320_adj_5069), 
            .CO(n39798));
    SB_LUT4 add_5259_4_lut (.I0(GND_net), .I1(n17639[1]), .I2(n247_adj_5067), 
            .I3(n39796), .O(n17248[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5259_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5259_4 (.CI(n39796), .I0(n17639[1]), .I1(n247_adj_5067), 
            .CO(n39797));
    SB_LUT4 add_5259_3_lut (.I0(GND_net), .I1(n17639[0]), .I2(n174_adj_5066), 
            .I3(n39795), .O(n17248[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5259_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5259_3 (.CI(n39795), .I0(n17639[0]), .I1(n174_adj_5066), 
            .CO(n39796));
    SB_LUT4 add_5259_2_lut (.I0(GND_net), .I1(n32_adj_5065), .I2(n101_adj_5064), 
            .I3(GND_net), .O(n17248[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5259_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5259_2 (.CI(GND_net), .I0(n32_adj_5065), .I1(n101_adj_5064), 
            .CO(n39795));
    SB_CARRY unary_minus_16_add_3_22 (.CI(n38772), .I0(GND_net), .I1(n1_adj_5235[20]), 
            .CO(n38773));
    SB_LUT4 add_5285_14_lut (.I0(GND_net), .I1(n17976[11]), .I2(n980_adj_5063), 
            .I3(n39794), .O(n17639[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5285_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_add_3_21_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5235[19]), 
            .I3(n38771), .O(n257[19])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5285_13_lut (.I0(GND_net), .I1(n17976[10]), .I2(n907_adj_5061), 
            .I3(n39793), .O(n17639[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5285_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_21 (.CI(n38771), .I0(GND_net), .I1(n1_adj_5235[19]), 
            .CO(n38772));
    SB_LUT4 unary_minus_16_add_3_20_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5235[18]), 
            .I3(n38770), .O(n257[18])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5285_13 (.CI(n39793), .I0(n17976[10]), .I1(n907_adj_5061), 
            .CO(n39794));
    SB_LUT4 add_5285_12_lut (.I0(GND_net), .I1(n17976[9]), .I2(n834_adj_5059), 
            .I3(n39792), .O(n17639[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5285_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5285_12 (.CI(n39792), .I0(n17976[9]), .I1(n834_adj_5059), 
            .CO(n39793));
    SB_CARRY add_5185_10 (.CI(n39599), .I0(n16544[7]), .I1(n679), .CO(n39600));
    SB_LUT4 add_5285_11_lut (.I0(GND_net), .I1(n17976[8]), .I2(n761_adj_5058), 
            .I3(n39791), .O(n17639[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5285_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5185_9_lut (.I0(GND_net), .I1(n16544[6]), .I2(n606), .I3(n39598), 
            .O(n16000[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5185_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5285_11 (.CI(n39791), .I0(n17976[8]), .I1(n761_adj_5058), 
            .CO(n39792));
    SB_LUT4 add_5285_10_lut (.I0(GND_net), .I1(n17976[7]), .I2(n688_adj_5057), 
            .I3(n39790), .O(n17639[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5285_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5285_10 (.CI(n39790), .I0(n17976[7]), .I1(n688_adj_5057), 
            .CO(n39791));
    SB_LUT4 add_5285_9_lut (.I0(GND_net), .I1(n17976[6]), .I2(n615_adj_5056), 
            .I3(n39789), .O(n17639[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5285_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_20 (.CI(n38770), .I0(GND_net), .I1(n1_adj_5235[18]), 
            .CO(n38771));
    SB_CARRY add_5185_9 (.CI(n39598), .I0(n16544[6]), .I1(n606), .CO(n39599));
    SB_CARRY add_5285_9 (.CI(n39789), .I0(n17976[6]), .I1(n615_adj_5056), 
            .CO(n39790));
    SB_LUT4 add_5285_8_lut (.I0(GND_net), .I1(n17976[5]), .I2(n542_adj_5055), 
            .I3(n39788), .O(n17639[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5285_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5185_8_lut (.I0(GND_net), .I1(n16544[5]), .I2(n533), .I3(n39597), 
            .O(n16000[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5185_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_add_3_19_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5235[17]), 
            .I3(n38769), .O(n257[17])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5285_8 (.CI(n39788), .I0(n17976[5]), .I1(n542_adj_5055), 
            .CO(n39789));
    SB_LUT4 add_5285_7_lut (.I0(GND_net), .I1(n17976[4]), .I2(n469_adj_5051), 
            .I3(n39787), .O(n17639[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5285_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5285_7 (.CI(n39787), .I0(n17976[4]), .I1(n469_adj_5051), 
            .CO(n39788));
    SB_LUT4 add_5285_6_lut (.I0(GND_net), .I1(n17976[3]), .I2(n396_adj_5050), 
            .I3(n39786), .O(n17639[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5285_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_19 (.CI(n38769), .I0(GND_net), .I1(n1_adj_5235[17]), 
            .CO(n38770));
    SB_CARRY add_5185_8 (.CI(n39597), .I0(n16544[5]), .I1(n533), .CO(n39598));
    SB_CARRY add_5285_6 (.CI(n39786), .I0(n17976[3]), .I1(n396_adj_5050), 
            .CO(n39787));
    SB_LUT4 add_5285_5_lut (.I0(GND_net), .I1(n17976[2]), .I2(n323_adj_5049), 
            .I3(n39785), .O(n17639[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5285_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5285_5 (.CI(n39785), .I0(n17976[2]), .I1(n323_adj_5049), 
            .CO(n39786));
    SB_LUT4 add_5285_4_lut (.I0(GND_net), .I1(n17976[1]), .I2(n250_adj_5048), 
            .I3(n39784), .O(n17639[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5285_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5285_4 (.CI(n39784), .I0(n17976[1]), .I1(n250_adj_5048), 
            .CO(n39785));
    SB_LUT4 add_5285_3_lut (.I0(GND_net), .I1(n17976[0]), .I2(n177_adj_5046), 
            .I3(n39783), .O(n17639[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5285_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5285_3 (.CI(n39783), .I0(n17976[0]), .I1(n177_adj_5046), 
            .CO(n39784));
    SB_LUT4 add_5285_2_lut (.I0(GND_net), .I1(n35_adj_5045), .I2(n104_adj_5044), 
            .I3(GND_net), .O(n17639[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5285_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5285_2 (.CI(GND_net), .I0(n35_adj_5045), .I1(n104_adj_5044), 
            .CO(n39783));
    SB_LUT4 add_5405_7_lut (.I0(GND_net), .I1(n46355), .I2(n490_adj_5036), 
            .I3(n39782), .O(n19040[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5405_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5405_6_lut (.I0(GND_net), .I1(n19124[3]), .I2(n417), .I3(n39781), 
            .O(n19040[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5405_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5405_6 (.CI(n39781), .I0(n19124[3]), .I1(n417), .CO(n39782));
    SB_LUT4 add_5405_5_lut (.I0(GND_net), .I1(n19124[2]), .I2(n344), .I3(n39780), 
            .O(n19040[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5405_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5405_5 (.CI(n39780), .I0(n19124[2]), .I1(n344), .CO(n39781));
    SB_LUT4 add_5405_4_lut (.I0(GND_net), .I1(n19124[1]), .I2(n271_adj_5022), 
            .I3(n39779), .O(n19040[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5405_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_add_3_18_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5235[16]), 
            .I3(n38768), .O(n257[16])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5405_4 (.CI(n39779), .I0(n19124[1]), .I1(n271_adj_5022), 
            .CO(n39780));
    SB_LUT4 add_5405_3_lut (.I0(GND_net), .I1(n19124[0]), .I2(n198), .I3(n39778), 
            .O(n19040[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5405_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5405_3 (.CI(n39778), .I0(n19124[0]), .I1(n198), .CO(n39779));
    SB_LUT4 add_5405_2_lut (.I0(GND_net), .I1(n56), .I2(n125), .I3(GND_net), 
            .O(n19040[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5405_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_18 (.CI(n38768), .I0(GND_net), .I1(n1_adj_5235[16]), 
            .CO(n38769));
    SB_LUT4 add_5185_7_lut (.I0(GND_net), .I1(n16544[4]), .I2(n460), .I3(n39596), 
            .O(n16000[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5185_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5405_2 (.CI(GND_net), .I0(n56), .I1(n125), .CO(n39778));
    SB_CARRY add_5185_7 (.CI(n39596), .I0(n16544[4]), .I1(n460), .CO(n39597));
    SB_LUT4 add_5185_6_lut (.I0(GND_net), .I1(n16544[3]), .I2(n387), .I3(n39595), 
            .O(n16000[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5185_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5309_13_lut (.I0(GND_net), .I1(n18263[10]), .I2(n910_adj_5019), 
            .I3(n39777), .O(n17976[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5309_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5309_12_lut (.I0(GND_net), .I1(n18263[9]), .I2(n837_adj_5018), 
            .I3(n39776), .O(n17976[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5309_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5185_6 (.CI(n39595), .I0(n16544[3]), .I1(n387), .CO(n39596));
    SB_CARRY add_5309_12 (.CI(n39776), .I0(n18263[9]), .I1(n837_adj_5018), 
            .CO(n39777));
    SB_LUT4 add_5309_11_lut (.I0(GND_net), .I1(n18263[8]), .I2(n764_adj_5017), 
            .I3(n39775), .O(n17976[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5309_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5185_5_lut (.I0(GND_net), .I1(n16544[2]), .I2(n314), .I3(n39594), 
            .O(n16000[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5185_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5185_5 (.CI(n39594), .I0(n16544[2]), .I1(n314), .CO(n39595));
    SB_LUT4 add_5185_4_lut (.I0(GND_net), .I1(n16544[1]), .I2(n241), .I3(n39593), 
            .O(n16000[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5185_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_add_3_17_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5235[15]), 
            .I3(n38767), .O(n257[15])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5185_4 (.CI(n39593), .I0(n16544[1]), .I1(n241), .CO(n39594));
    SB_LUT4 add_5185_3_lut (.I0(GND_net), .I1(n16544[0]), .I2(n168), .I3(n39592), 
            .O(n16000[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5185_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5309_11 (.CI(n39775), .I0(n18263[8]), .I1(n764_adj_5017), 
            .CO(n39776));
    SB_LUT4 add_5309_10_lut (.I0(GND_net), .I1(n18263[7]), .I2(n691), 
            .I3(n39774), .O(n17976[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5309_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5309_10 (.CI(n39774), .I0(n18263[7]), .I1(n691), .CO(n39775));
    SB_LUT4 add_5309_9_lut (.I0(GND_net), .I1(n18263[6]), .I2(n618), .I3(n39773), 
            .O(n17976[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5309_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5309_9 (.CI(n39773), .I0(n18263[6]), .I1(n618), .CO(n39774));
    SB_LUT4 add_5309_8_lut (.I0(GND_net), .I1(n18263[5]), .I2(n545), .I3(n39772), 
            .O(n17976[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5309_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5309_8 (.CI(n39772), .I0(n18263[5]), .I1(n545), .CO(n39773));
    SB_LUT4 add_5309_7_lut (.I0(GND_net), .I1(n18263[4]), .I2(n472), .I3(n39771), 
            .O(n17976[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5309_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5185_3 (.CI(n39592), .I0(n16544[0]), .I1(n168), .CO(n39593));
    SB_CARRY add_5309_7 (.CI(n39771), .I0(n18263[4]), .I1(n472), .CO(n39772));
    SB_LUT4 add_5309_6_lut (.I0(GND_net), .I1(n18263[3]), .I2(n399), .I3(n39770), 
            .O(n17976[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5309_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5309_6 (.CI(n39770), .I0(n18263[3]), .I1(n399), .CO(n39771));
    SB_LUT4 add_5309_5_lut (.I0(GND_net), .I1(n18263[2]), .I2(n326), .I3(n39769), 
            .O(n17976[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5309_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5309_5 (.CI(n39769), .I0(n18263[2]), .I1(n326), .CO(n39770));
    SB_LUT4 add_5309_4_lut (.I0(GND_net), .I1(n18263[1]), .I2(n253), .I3(n39768), 
            .O(n17976[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5309_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5309_4 (.CI(n39768), .I0(n18263[1]), .I1(n253), .CO(n39769));
    SB_LUT4 add_5309_3_lut (.I0(GND_net), .I1(n18263[0]), .I2(n180), .I3(n39767), 
            .O(n17976[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5309_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5309_3 (.CI(n39767), .I0(n18263[0]), .I1(n180), .CO(n39768));
    SB_LUT4 add_5309_2_lut (.I0(GND_net), .I1(n38), .I2(n107), .I3(GND_net), 
            .O(n17976[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5309_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5309_2 (.CI(GND_net), .I0(n38), .I1(n107), .CO(n39767));
    SB_LUT4 add_5331_12_lut (.I0(GND_net), .I1(n18504[9]), .I2(n840_adj_4994), 
            .I3(n39766), .O(n18263[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5331_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5331_11_lut (.I0(GND_net), .I1(n18504[8]), .I2(n767_adj_4991), 
            .I3(n39765), .O(n18263[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5331_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5331_11 (.CI(n39765), .I0(n18504[8]), .I1(n767_adj_4991), 
            .CO(n39766));
    SB_LUT4 add_5331_10_lut (.I0(GND_net), .I1(n18504[7]), .I2(n694_adj_4985), 
            .I3(n39764), .O(n18263[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5331_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5331_10 (.CI(n39764), .I0(n18504[7]), .I1(n694_adj_4985), 
            .CO(n39765));
    SB_LUT4 add_5331_9_lut (.I0(GND_net), .I1(n18504[6]), .I2(n621_adj_4980), 
            .I3(n39763), .O(n18263[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5331_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5331_9 (.CI(n39763), .I0(n18504[6]), .I1(n621_adj_4980), 
            .CO(n39764));
    SB_LUT4 add_5331_8_lut (.I0(GND_net), .I1(n18504[5]), .I2(n548_adj_4975), 
            .I3(n39762), .O(n18263[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5331_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5331_8 (.CI(n39762), .I0(n18504[5]), .I1(n548_adj_4975), 
            .CO(n39763));
    SB_LUT4 add_5331_7_lut (.I0(GND_net), .I1(n18504[4]), .I2(n475_adj_4971), 
            .I3(n39761), .O(n18263[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5331_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5331_7 (.CI(n39761), .I0(n18504[4]), .I1(n475_adj_4971), 
            .CO(n39762));
    SB_CARRY unary_minus_16_add_3_17 (.CI(n38767), .I0(GND_net), .I1(n1_adj_5235[15]), 
            .CO(n38768));
    SB_LUT4 unary_minus_16_add_3_16_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5235[14]), 
            .I3(n38766), .O(n257[14])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_16 (.CI(n38766), .I0(GND_net), .I1(n1_adj_5235[14]), 
            .CO(n38767));
    SB_LUT4 unary_minus_16_add_3_15_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5235[13]), 
            .I3(n38765), .O(n257[13])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_15 (.CI(n38765), .I0(GND_net), .I1(n1_adj_5235[13]), 
            .CO(n38766));
    SB_LUT4 unary_minus_16_add_3_14_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5235[12]), 
            .I3(n38764), .O(n257[12])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5331_6_lut (.I0(GND_net), .I1(n18504[3]), .I2(n402_adj_4881), 
            .I3(n39760), .O(n18263[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5331_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5331_6 (.CI(n39760), .I0(n18504[3]), .I1(n402_adj_4881), 
            .CO(n39761));
    SB_LUT4 add_5331_5_lut (.I0(GND_net), .I1(n18504[2]), .I2(n329_adj_4877), 
            .I3(n39759), .O(n18263[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5331_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5331_5 (.CI(n39759), .I0(n18504[2]), .I1(n329_adj_4877), 
            .CO(n39760));
    SB_LUT4 add_5331_4_lut (.I0(GND_net), .I1(n18504[1]), .I2(n256_adj_4873), 
            .I3(n39758), .O(n18263[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5331_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5331_4 (.CI(n39758), .I0(n18504[1]), .I1(n256_adj_4873), 
            .CO(n39759));
    SB_LUT4 add_5331_3_lut (.I0(GND_net), .I1(n18504[0]), .I2(n183), .I3(n39757), 
            .O(n18263[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5331_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5331_3 (.CI(n39757), .I0(n18504[0]), .I1(n183), .CO(n39758));
    SB_LUT4 add_5331_2_lut (.I0(GND_net), .I1(n41), .I2(n110), .I3(GND_net), 
            .O(n18263[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5331_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5331_2 (.CI(GND_net), .I0(n41), .I1(n110), .CO(n39757));
    SB_LUT4 mult_11_add_1225_24_lut (.I0(\PID_CONTROLLER.integral_23__N_3836 [23]), 
            .I1(n11163[21]), .I2(GND_net), .I3(n39756), .O(n10656[0])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_24_lut.LUT_INIT = 16'h6996;
    SB_LUT4 mult_11_add_1225_23_lut (.I0(GND_net), .I1(n11163[20]), .I2(GND_net), 
            .I3(n39755), .O(n155[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_23 (.CI(n39755), .I0(n11163[20]), .I1(GND_net), 
            .CO(n39756));
    SB_LUT4 mult_11_add_1225_22_lut (.I0(GND_net), .I1(n11163[19]), .I2(GND_net), 
            .I3(n39754), .O(n155[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_22 (.CI(n39754), .I0(n11163[19]), .I1(GND_net), 
            .CO(n39755));
    SB_LUT4 mult_11_add_1225_21_lut (.I0(GND_net), .I1(n11163[18]), .I2(GND_net), 
            .I3(n39753), .O(n155[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_21 (.CI(n39753), .I0(n11163[18]), .I1(GND_net), 
            .CO(n39754));
    SB_LUT4 mult_11_add_1225_20_lut (.I0(GND_net), .I1(n11163[17]), .I2(GND_net), 
            .I3(n39752), .O(n155[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_20 (.CI(n39752), .I0(n11163[17]), .I1(GND_net), 
            .CO(n39753));
    SB_LUT4 mult_11_add_1225_19_lut (.I0(GND_net), .I1(n11163[16]), .I2(GND_net), 
            .I3(n39751), .O(n155[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_19 (.CI(n39751), .I0(n11163[16]), .I1(GND_net), 
            .CO(n39752));
    SB_LUT4 mult_11_add_1225_18_lut (.I0(GND_net), .I1(n11163[15]), .I2(GND_net), 
            .I3(n39750), .O(n155[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_18 (.CI(n39750), .I0(n11163[15]), .I1(GND_net), 
            .CO(n39751));
    SB_LUT4 mult_11_add_1225_17_lut (.I0(GND_net), .I1(n11163[14]), .I2(GND_net), 
            .I3(n39749), .O(n155[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_17 (.CI(n39749), .I0(n11163[14]), .I1(GND_net), 
            .CO(n39750));
    SB_LUT4 mult_11_add_1225_16_lut (.I0(GND_net), .I1(n11163[13]), .I2(n1096), 
            .I3(n39748), .O(n155[15])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_16 (.CI(n39748), .I0(n11163[13]), .I1(n1096), 
            .CO(n39749));
    SB_LUT4 mult_11_add_1225_15_lut (.I0(GND_net), .I1(n11163[12]), .I2(n1023), 
            .I3(n39747), .O(n155[14])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_15 (.CI(n39747), .I0(n11163[12]), .I1(n1023), 
            .CO(n39748));
    SB_LUT4 mult_11_add_1225_14_lut (.I0(GND_net), .I1(n11163[11]), .I2(n950), 
            .I3(n39746), .O(n155[13])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i696_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n1035_adj_5025));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i696_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY unary_minus_16_add_3_14 (.CI(n38764), .I0(GND_net), .I1(n1_adj_5235[12]), 
            .CO(n38765));
    SB_CARRY mult_11_add_1225_14 (.CI(n39746), .I0(n11163[11]), .I1(n950), 
            .CO(n39747));
    SB_LUT4 mult_11_add_1225_13_lut (.I0(GND_net), .I1(n11163[10]), .I2(n877), 
            .I3(n39745), .O(n155[12])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_13 (.CI(n39745), .I0(n11163[10]), .I1(n877), 
            .CO(n39746));
    SB_LUT4 mult_11_add_1225_12_lut (.I0(GND_net), .I1(n11163[9]), .I2(n804), 
            .I3(n39744), .O(n155[11])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_12 (.CI(n39744), .I0(n11163[9]), .I1(n804), 
            .CO(n39745));
    SB_LUT4 mult_11_add_1225_11_lut (.I0(GND_net), .I1(n11163[8]), .I2(n731), 
            .I3(n39743), .O(n155[10])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_11 (.CI(n39743), .I0(n11163[8]), .I1(n731), 
            .CO(n39744));
    SB_LUT4 mult_11_add_1225_10_lut (.I0(GND_net), .I1(n11163[7]), .I2(n658), 
            .I3(n39742), .O(n155[9])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_10 (.CI(n39742), .I0(n11163[7]), .I1(n658), 
            .CO(n39743));
    SB_LUT4 mult_11_add_1225_9_lut (.I0(GND_net), .I1(n11163[6]), .I2(n585), 
            .I3(n39741), .O(n155[8])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_9 (.CI(n39741), .I0(n11163[6]), .I1(n585), 
            .CO(n39742));
    SB_LUT4 mult_11_add_1225_8_lut (.I0(GND_net), .I1(n11163[5]), .I2(n512), 
            .I3(n39740), .O(n155[7])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_8 (.CI(n39740), .I0(n11163[5]), .I1(n512), 
            .CO(n39741));
    SB_LUT4 mult_11_add_1225_7_lut (.I0(GND_net), .I1(n11163[4]), .I2(n439), 
            .I3(n39739), .O(n155[6])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_7 (.CI(n39739), .I0(n11163[4]), .I1(n439), 
            .CO(n39740));
    SB_LUT4 mult_11_add_1225_6_lut (.I0(GND_net), .I1(n11163[3]), .I2(n366), 
            .I3(n39738), .O(n155[5])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_6 (.CI(n39738), .I0(n11163[3]), .I1(n366), 
            .CO(n39739));
    SB_LUT4 mult_11_add_1225_5_lut (.I0(GND_net), .I1(n11163[2]), .I2(n293), 
            .I3(n39737), .O(n155[4])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_5 (.CI(n39737), .I0(n11163[2]), .I1(n293), 
            .CO(n39738));
    SB_LUT4 mult_11_add_1225_4_lut (.I0(GND_net), .I1(n11163[1]), .I2(n220), 
            .I3(n39736), .O(n155[3])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_4 (.CI(n39736), .I0(n11163[1]), .I1(n220), 
            .CO(n39737));
    SB_LUT4 mult_11_add_1225_3_lut (.I0(GND_net), .I1(n11163[0]), .I2(n147), 
            .I3(n39735), .O(n155[2])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_3 (.CI(n39735), .I0(n11163[0]), .I1(n147), 
            .CO(n39736));
    SB_LUT4 mult_11_add_1225_2_lut (.I0(GND_net), .I1(n5), .I2(n74), .I3(GND_net), 
            .O(n155[1])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_2 (.CI(GND_net), .I0(n5), .I1(n74), .CO(n39735));
    SB_LUT4 add_4955_23_lut (.I0(GND_net), .I1(n12180[20]), .I2(GND_net), 
            .I3(n39734), .O(n11163[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4955_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_add_3_13_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5235[11]), 
            .I3(n38763), .O(n257[11])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4955_22_lut (.I0(GND_net), .I1(n12180[19]), .I2(GND_net), 
            .I3(n39733), .O(n11163[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4955_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4955_22 (.CI(n39733), .I0(n12180[19]), .I1(GND_net), 
            .CO(n39734));
    SB_LUT4 add_5185_2_lut (.I0(GND_net), .I1(n26), .I2(n95), .I3(GND_net), 
            .O(n16000[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5185_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4955_21_lut (.I0(GND_net), .I1(n12180[18]), .I2(GND_net), 
            .I3(n39732), .O(n11163[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4955_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i557_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n828));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i557_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY unary_minus_16_add_3_13 (.CI(n38763), .I0(GND_net), .I1(n1_adj_5235[11]), 
            .CO(n38764));
    SB_LUT4 unary_minus_16_add_3_12_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5235[10]), 
            .I3(n38762), .O(n257[10])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5185_2 (.CI(GND_net), .I0(n26), .I1(n95), .CO(n39592));
    SB_CARRY add_4955_21 (.CI(n39732), .I0(n12180[18]), .I1(GND_net), 
            .CO(n39733));
    SB_CARRY unary_minus_16_add_3_12 (.CI(n38762), .I0(GND_net), .I1(n1_adj_5235[10]), 
            .CO(n38763));
    SB_LUT4 i20711_2_lut (.I0(n1[0]), .I1(\PID_CONTROLLER.integral_23__N_3884 ), 
            .I2(GND_net), .I3(GND_net), .O(n4751[0]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i20711_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i281_2_lut (.I0(\Kp[5] ), .I1(n1[17]), .I2(GND_net), 
            .I3(GND_net), .O(n417_adj_5024));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i281_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i653_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n971_adj_5169));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i653_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_4_lut_adj_1716 (.I0(n6_adj_5171), .I1(\Kp[4] ), .I2(n19208[2]), 
            .I3(n1[18]), .O(n19159[3]));   // verilog/motorControl.v(34[16:22])
    defparam i2_4_lut_adj_1716.LUT_INIT = 16'h965a;
    SB_LUT4 mult_11_i606_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n901));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i606_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i151_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n223));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i151_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i3_1_lut (.I0(IntegralLimit[2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5234[2]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_16_add_3_11_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5235[9]), 
            .I3(n38761), .O(n257[9])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_11 (.CI(n38761), .I0(GND_net), .I1(n1_adj_5235[9]), 
            .CO(n38762));
    SB_LUT4 add_4955_20_lut (.I0(GND_net), .I1(n12180[17]), .I2(GND_net), 
            .I3(n39731), .O(n11163[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4955_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4955_20 (.CI(n39731), .I0(n12180[17]), .I1(GND_net), 
            .CO(n39732));
    SB_LUT4 add_5385_9_lut (.I0(GND_net), .I1(n18991[6]), .I2(n630), .I3(n39591), 
            .O(n18864[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5385_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_add_3_10_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5235[8]), 
            .I3(n38760), .O(n257[8])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5385_8_lut (.I0(GND_net), .I1(n18991[5]), .I2(n557), .I3(n39590), 
            .O(n18864[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5385_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_10 (.CI(n38760), .I0(GND_net), .I1(n1_adj_5235[8]), 
            .CO(n38761));
    SB_LUT4 unary_minus_16_add_3_9_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5235[7]), 
            .I3(n38759), .O(n257[7])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_9 (.CI(n38759), .I0(GND_net), .I1(n1_adj_5235[7]), 
            .CO(n38760));
    SB_LUT4 add_4955_19_lut (.I0(GND_net), .I1(n12180[16]), .I2(GND_net), 
            .I3(n39730), .O(n11163[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4955_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4955_19 (.CI(n39730), .I0(n12180[16]), .I1(GND_net), 
            .CO(n39731));
    SB_CARRY add_5385_8 (.CI(n39590), .I0(n18991[5]), .I1(n557), .CO(n39591));
    SB_LUT4 add_5385_7_lut (.I0(GND_net), .I1(n18991[4]), .I2(n484), .I3(n39589), 
            .O(n18864[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5385_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_add_3_8_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5235[6]), 
            .I3(n38758), .O(n257[6])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_8 (.CI(n38758), .I0(GND_net), .I1(n1_adj_5235[6]), 
            .CO(n38759));
    SB_LUT4 add_4955_18_lut (.I0(GND_net), .I1(n12180[15]), .I2(GND_net), 
            .I3(n39729), .O(n11163[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4955_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5385_7 (.CI(n39589), .I0(n18991[4]), .I1(n484), .CO(n39590));
    SB_LUT4 unary_minus_16_add_3_7_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5235[5]), 
            .I3(n38757), .O(n257[5])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_7 (.CI(n38757), .I0(GND_net), .I1(n1_adj_5235[5]), 
            .CO(n38758));
    SB_LUT4 add_5385_6_lut (.I0(GND_net), .I1(n18991[3]), .I2(n411), .I3(n39588), 
            .O(n18864[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5385_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_add_3_6_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5235[4]), 
            .I3(n38756), .O(n257[4])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_6 (.CI(n38756), .I0(GND_net), .I1(n1_adj_5235[4]), 
            .CO(n38757));
    SB_LUT4 unary_minus_16_add_3_5_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5235[3]), 
            .I3(n38755), .O(n257[3])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5385_6 (.CI(n39588), .I0(n18991[3]), .I1(n411), .CO(n39589));
    SB_CARRY unary_minus_16_add_3_5 (.CI(n38755), .I0(GND_net), .I1(n1_adj_5235[3]), 
            .CO(n38756));
    SB_LUT4 unary_minus_16_add_3_4_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5235[2]), 
            .I3(n38754), .O(n257[2])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4955_18 (.CI(n39729), .I0(n12180[15]), .I1(GND_net), 
            .CO(n39730));
    SB_LUT4 add_4955_17_lut (.I0(GND_net), .I1(n12180[14]), .I2(GND_net), 
            .I3(n39728), .O(n11163[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4955_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5385_5_lut (.I0(GND_net), .I1(n18991[2]), .I2(n338), .I3(n39587), 
            .O(n18864[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5385_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_4 (.CI(n38754), .I0(GND_net), .I1(n1_adj_5235[2]), 
            .CO(n38755));
    SB_LUT4 unary_minus_16_add_3_3_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5235[1]), 
            .I3(n38753), .O(n257[1])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5385_5 (.CI(n39587), .I0(n18991[2]), .I1(n338), .CO(n39588));
    SB_CARRY unary_minus_16_add_3_3 (.CI(n38753), .I0(GND_net), .I1(n1_adj_5235[1]), 
            .CO(n38754));
    SB_LUT4 unary_minus_16_add_3_2_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5235[0]), 
            .I3(VCC_net), .O(n257[0])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_2 (.CI(VCC_net), .I0(GND_net), .I1(n1_adj_5235[0]), 
            .CO(n38753));
    SB_LUT4 unary_minus_5_add_3_25_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5234[23]), 
            .I3(n38752), .O(\PID_CONTROLLER.integral_23__N_3887 [23])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_24_lut (.I0(\PID_CONTROLLER.integral [22]), 
            .I1(GND_net), .I2(n1_adj_5234[22]), .I3(n38751), .O(n45)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_24_lut.LUT_INIT = 16'h6996;
    SB_CARRY unary_minus_5_add_3_24 (.CI(n38751), .I0(GND_net), .I1(n1_adj_5234[22]), 
            .CO(n38752));
    SB_LUT4 unary_minus_5_add_3_23_lut (.I0(\PID_CONTROLLER.integral [21]), 
            .I1(GND_net), .I2(n1_adj_5234[21]), .I3(n38750), .O(n43)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_23_lut.LUT_INIT = 16'h6996;
    SB_CARRY add_4955_17 (.CI(n39728), .I0(n12180[14]), .I1(GND_net), 
            .CO(n39729));
    SB_CARRY unary_minus_5_add_3_23 (.CI(n38750), .I0(GND_net), .I1(n1_adj_5234[21]), 
            .CO(n38751));
    SB_LUT4 add_5385_4_lut (.I0(GND_net), .I1(n18991[1]), .I2(n265), .I3(n39586), 
            .O(n18864[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5385_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_22_lut (.I0(\PID_CONTROLLER.integral [20]), 
            .I1(GND_net), .I2(n1_adj_5234[20]), .I3(n38749), .O(n41_adj_4962)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_22_lut.LUT_INIT = 16'h6996;
    SB_CARRY unary_minus_5_add_3_22 (.CI(n38749), .I0(GND_net), .I1(n1_adj_5234[20]), 
            .CO(n38750));
    SB_LUT4 unary_minus_5_add_3_21_lut (.I0(\PID_CONTROLLER.integral [19]), 
            .I1(GND_net), .I2(n1_adj_5234[19]), .I3(n38748), .O(n39)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_21_lut.LUT_INIT = 16'h6996;
    SB_CARRY add_5385_4 (.CI(n39586), .I0(n18991[1]), .I1(n265), .CO(n39587));
    SB_CARRY unary_minus_5_add_3_21 (.CI(n38748), .I0(GND_net), .I1(n1_adj_5234[19]), 
            .CO(n38749));
    SB_LUT4 unary_minus_5_add_3_20_lut (.I0(\PID_CONTROLLER.integral [18]), 
            .I1(GND_net), .I2(n1_adj_5234[18]), .I3(n38747), .O(n37)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_20_lut.LUT_INIT = 16'h6996;
    SB_CARRY unary_minus_5_add_3_20 (.CI(n38747), .I0(GND_net), .I1(n1_adj_5234[18]), 
            .CO(n38748));
    SB_LUT4 unary_minus_5_add_3_19_lut (.I0(\PID_CONTROLLER.integral [17]), 
            .I1(GND_net), .I2(n1_adj_5234[17]), .I3(n38746), .O(n35)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_19_lut.LUT_INIT = 16'h6996;
    SB_CARRY unary_minus_5_add_3_19 (.CI(n38746), .I0(GND_net), .I1(n1_adj_5234[17]), 
            .CO(n38747));
    SB_LUT4 unary_minus_5_add_3_18_lut (.I0(\PID_CONTROLLER.integral [16]), 
            .I1(GND_net), .I2(n1_adj_5234[16]), .I3(n38745), .O(n33)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_18_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_4955_16_lut (.I0(GND_net), .I1(n12180[13]), .I2(n1099), 
            .I3(n39727), .O(n11163[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4955_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5385_3_lut (.I0(GND_net), .I1(n18991[0]), .I2(n192), .I3(n39585), 
            .O(n18864[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5385_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_5_add_3_18 (.CI(n38745), .I0(GND_net), .I1(n1_adj_5234[16]), 
            .CO(n38746));
    SB_LUT4 unary_minus_5_add_3_17_lut (.I0(\PID_CONTROLLER.integral [15]), 
            .I1(GND_net), .I2(n1_adj_5234[15]), .I3(n38744), .O(n31)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_17_lut.LUT_INIT = 16'h6996;
    SB_CARRY add_5385_3 (.CI(n39585), .I0(n18991[0]), .I1(n192), .CO(n39586));
    SB_CARRY unary_minus_5_add_3_17 (.CI(n38744), .I0(GND_net), .I1(n1_adj_5234[15]), 
            .CO(n38745));
    SB_LUT4 unary_minus_5_add_3_16_lut (.I0(\PID_CONTROLLER.integral [14]), 
            .I1(GND_net), .I2(n1_adj_5234[14]), .I3(n38743), .O(n29)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_16_lut.LUT_INIT = 16'h6996;
    SB_CARRY unary_minus_5_add_3_16 (.CI(n38743), .I0(GND_net), .I1(n1_adj_5234[14]), 
            .CO(n38744));
    SB_LUT4 unary_minus_5_add_3_15_lut (.I0(\PID_CONTROLLER.integral [13]), 
            .I1(GND_net), .I2(n1_adj_5234[13]), .I3(n38742), .O(n27)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_15_lut.LUT_INIT = 16'h6996;
    SB_CARRY unary_minus_5_add_3_15 (.CI(n38742), .I0(GND_net), .I1(n1_adj_5234[13]), 
            .CO(n38743));
    SB_LUT4 unary_minus_5_add_3_14_lut (.I0(\PID_CONTROLLER.integral [12]), 
            .I1(GND_net), .I2(n1_adj_5234[12]), .I3(n38741), .O(n25_adj_4920)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_14_lut.LUT_INIT = 16'h6996;
    SB_CARRY add_4955_16 (.CI(n39727), .I0(n12180[13]), .I1(n1099), .CO(n39728));
    SB_CARRY unary_minus_5_add_3_14 (.CI(n38741), .I0(GND_net), .I1(n1_adj_5234[12]), 
            .CO(n38742));
    SB_LUT4 add_4955_15_lut (.I0(GND_net), .I1(n12180[12]), .I2(n1026), 
            .I3(n39726), .O(n11163[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4955_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4955_15 (.CI(n39726), .I0(n12180[12]), .I1(n1026), .CO(n39727));
    SB_LUT4 unary_minus_5_add_3_13_lut (.I0(\PID_CONTROLLER.integral [11]), 
            .I1(GND_net), .I2(n1_adj_5234[11]), .I3(n38740), .O(n23_adj_4921)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_13_lut.LUT_INIT = 16'h6996;
    SB_CARRY unary_minus_5_add_3_13 (.CI(n38740), .I0(GND_net), .I1(n1_adj_5234[11]), 
            .CO(n38741));
    SB_LUT4 add_4955_14_lut (.I0(GND_net), .I1(n12180[11]), .I2(n953), 
            .I3(n39725), .O(n11163[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4955_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4955_14 (.CI(n39725), .I0(n12180[11]), .I1(n953), .CO(n39726));
    SB_LUT4 unary_minus_5_add_3_12_lut (.I0(\PID_CONTROLLER.integral [10]), 
            .I1(GND_net), .I2(n1_adj_5234[10]), .I3(n38739), .O(n21_adj_4912)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_12_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_4955_13_lut (.I0(GND_net), .I1(n12180[10]), .I2(n880), 
            .I3(n39724), .O(n11163[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4955_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4955_13 (.CI(n39724), .I0(n12180[10]), .I1(n880), .CO(n39725));
    SB_CARRY unary_minus_5_add_3_12 (.CI(n38739), .I0(GND_net), .I1(n1_adj_5234[10]), 
            .CO(n38740));
    SB_LUT4 add_4955_12_lut (.I0(GND_net), .I1(n12180[9]), .I2(n807), 
            .I3(n39723), .O(n11163[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4955_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4955_12 (.CI(n39723), .I0(n12180[9]), .I1(n807), .CO(n39724));
    SB_LUT4 add_5385_2_lut (.I0(GND_net), .I1(n50), .I2(n119), .I3(GND_net), 
            .O(n18864[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5385_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_11_lut (.I0(\PID_CONTROLLER.integral [9]), 
            .I1(GND_net), .I2(n1_adj_5234[9]), .I3(n38738), .O(n19_adj_4913)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_11_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_4955_11_lut (.I0(GND_net), .I1(n12180[8]), .I2(n734), 
            .I3(n39722), .O(n11163[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4955_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4955_11 (.CI(n39722), .I0(n12180[8]), .I1(n734), .CO(n39723));
    SB_LUT4 add_4955_10_lut (.I0(GND_net), .I1(n12180[7]), .I2(n661), 
            .I3(n39721), .O(n11163[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4955_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4955_10 (.CI(n39721), .I0(n12180[7]), .I1(n661), .CO(n39722));
    SB_LUT4 add_4955_9_lut (.I0(GND_net), .I1(n12180[6]), .I2(n588), .I3(n39720), 
            .O(n11163[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4955_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4955_9 (.CI(n39720), .I0(n12180[6]), .I1(n588), .CO(n39721));
    SB_CARRY unary_minus_5_add_3_11 (.CI(n38738), .I0(GND_net), .I1(n1_adj_5234[9]), 
            .CO(n38739));
    SB_LUT4 unary_minus_5_add_3_10_lut (.I0(\PID_CONTROLLER.integral [8]), 
            .I1(GND_net), .I2(n1_adj_5234[8]), .I3(n38737), .O(n17_adj_4914)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_10_lut.LUT_INIT = 16'h6996;
    SB_CARRY unary_minus_5_add_3_10 (.CI(n38737), .I0(GND_net), .I1(n1_adj_5234[8]), 
            .CO(n38738));
    SB_LUT4 add_4955_8_lut (.I0(GND_net), .I1(n12180[5]), .I2(n515), .I3(n39719), 
            .O(n11163[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4955_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_9_lut (.I0(\PID_CONTROLLER.integral [7]), 
            .I1(GND_net), .I2(n1_adj_5234[7]), .I3(n38736), .O(n15_adj_4909)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_9_lut.LUT_INIT = 16'h6996;
    SB_CARRY unary_minus_5_add_3_9 (.CI(n38736), .I0(GND_net), .I1(n1_adj_5234[7]), 
            .CO(n38737));
    SB_CARRY add_4955_8 (.CI(n39719), .I0(n12180[5]), .I1(n515), .CO(n39720));
    SB_LUT4 add_4955_7_lut (.I0(GND_net), .I1(n12180[4]), .I2(n442), .I3(n39718), 
            .O(n11163[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4955_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_8_lut (.I0(\PID_CONTROLLER.integral [6]), 
            .I1(GND_net), .I2(n1_adj_5234[6]), .I3(n38735), .O(n13_adj_4910)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_8_lut.LUT_INIT = 16'h6996;
    SB_CARRY unary_minus_5_add_3_8 (.CI(n38735), .I0(GND_net), .I1(n1_adj_5234[6]), 
            .CO(n38736));
    SB_CARRY add_5385_2 (.CI(GND_net), .I0(n50), .I1(n119), .CO(n39585));
    SB_LUT4 add_5216_16_lut (.I0(GND_net), .I1(n17024[13]), .I2(n1120), 
            .I3(n39584), .O(n16544[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5216_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_7_lut (.I0(\PID_CONTROLLER.integral [5]), 
            .I1(GND_net), .I2(n1_adj_5234[5]), .I3(n38734), .O(n11_adj_4911)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_7_lut.LUT_INIT = 16'h6996;
    SB_CARRY add_4955_7 (.CI(n39718), .I0(n12180[4]), .I1(n442), .CO(n39719));
    SB_LUT4 add_5216_15_lut (.I0(GND_net), .I1(n17024[12]), .I2(n1047), 
            .I3(n39583), .O(n16544[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5216_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_5_add_3_7 (.CI(n38734), .I0(GND_net), .I1(n1_adj_5234[5]), 
            .CO(n38735));
    SB_LUT4 add_4955_6_lut (.I0(GND_net), .I1(n12180[3]), .I2(n369), .I3(n39717), 
            .O(n11163[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4955_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_6_lut (.I0(\PID_CONTROLLER.integral [4]), 
            .I1(GND_net), .I2(n1_adj_5234[4]), .I3(n38733), .O(n9_adj_4915)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_6_lut.LUT_INIT = 16'h6996;
    SB_CARRY add_4955_6 (.CI(n39717), .I0(n12180[3]), .I1(n369), .CO(n39718));
    SB_LUT4 add_4955_5_lut (.I0(GND_net), .I1(n12180[2]), .I2(n296), .I3(n39716), 
            .O(n11163[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4955_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i702_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n1044_adj_5168));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i702_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5216_15 (.CI(n39583), .I0(n17024[12]), .I1(n1047), .CO(n39584));
    SB_LUT4 mult_11_i751_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n1117_adj_5167));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i751_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i63_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n92_adj_5166));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i63_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i5_1_lut (.I0(IntegralLimit[4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5234[4]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i16_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_5165));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i16_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i745_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n1108_adj_5020));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i745_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i657_2_lut (.I0(\Kp[13] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n977_adj_5164));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i657_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i24267_4_lut (.I0(\Kp[0] ), .I1(\Kp[1] ), .I2(n1[22]), .I3(n1[21]), 
            .O(n19256[0]));   // verilog/motorControl.v(34[16:22])
    defparam i24267_4_lut.LUT_INIT = 16'h6ca0;
    SB_LUT4 mult_10_i706_2_lut (.I0(\Kp[14] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n1050_adj_5163));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i706_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_4_lut_adj_1717 (.I0(n4_adj_5172), .I1(\Kp[3] ), .I2(n19239[1]), 
            .I3(n1[19]), .O(n19208[2]));   // verilog/motorControl.v(34[16:22])
    defparam i2_4_lut_adj_1717.LUT_INIT = 16'h965a;
    SB_LUT4 mult_10_i330_2_lut (.I0(\Kp[6] ), .I1(n1[17]), .I2(GND_net), 
            .I3(GND_net), .O(n490));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i330_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i83_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [16]), 
            .I2(GND_net), .I3(GND_net), .O(n122_adj_5162));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i83_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i36_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [17]), 
            .I2(GND_net), .I3(GND_net), .O(n53_adj_5161));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i36_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i132_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [16]), 
            .I2(GND_net), .I3(GND_net), .O(n195_adj_5160));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i132_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_4_lut_adj_1718 (.I0(\Kp[0] ), .I1(\Kp[3] ), .I2(n1[23]), 
            .I3(n1[20]), .O(n12_adj_5173));   // verilog/motorControl.v(34[16:22])
    defparam i2_4_lut_adj_1718.LUT_INIT = 16'h9c50;
    SB_LUT4 i24471_4_lut (.I0(n19208[2]), .I1(\Kp[4] ), .I2(n6_adj_5171), 
            .I3(n1[18]), .O(n8_adj_5174));   // verilog/motorControl.v(34[16:22])
    defparam i24471_4_lut.LUT_INIT = 16'he8a0;
    SB_LUT4 i1_4_lut_adj_1719 (.I0(\Kp[4] ), .I1(\Kp[2] ), .I2(n1[19]), 
            .I3(n1[21]), .O(n11_adj_5175));   // verilog/motorControl.v(34[16:22])
    defparam i1_4_lut_adj_1719.LUT_INIT = 16'h6ca0;
    SB_LUT4 i24417_4_lut (.I0(n19239[1]), .I1(\Kp[3] ), .I2(n4_adj_5172), 
            .I3(n1[19]), .O(n6_adj_5176));   // verilog/motorControl.v(34[16:22])
    defparam i24417_4_lut.LUT_INIT = 16'he8a0;
    SB_LUT4 i24269_4_lut (.I0(\Kp[0] ), .I1(\Kp[1] ), .I2(n1[22]), .I3(n1[21]), 
            .O(n38216));   // verilog/motorControl.v(34[16:22])
    defparam i24269_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i24463_3_lut_4_lut (.I0(\Kp[3] ), .I1(n1[18]), .I2(n4_adj_5177), 
            .I3(n19208[1]), .O(n6_adj_5171));   // verilog/motorControl.v(34[16:22])
    defparam i24463_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 i8_4_lut_adj_1720 (.I0(n6_adj_5176), .I1(n11_adj_5175), .I2(n8_adj_5174), 
            .I3(n12_adj_5173), .O(n18_adj_5178));   // verilog/motorControl.v(34[16:22])
    defparam i8_4_lut_adj_1720.LUT_INIT = 16'h6996;
    SB_LUT4 mult_11_i655_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n974));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i655_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i112_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n165_adj_5159));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i112_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i181_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [16]), 
            .I2(GND_net), .I3(GND_net), .O(n268_adj_5158));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i181_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i3_4_lut_adj_1721 (.I0(\Kp[5] ), .I1(\Kp[1] ), .I2(n1[18]), 
            .I3(n1[22]), .O(n13_adj_5179));   // verilog/motorControl.v(34[16:22])
    defparam i3_4_lut_adj_1721.LUT_INIT = 16'h6ca0;
    SB_LUT4 i9_4_lut_adj_1722 (.I0(n13_adj_5179), .I1(n18_adj_5178), .I2(n38216), 
            .I3(n4_adj_5180), .O(n45851));   // verilog/motorControl.v(34[16:22])
    defparam i9_4_lut_adj_1722.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut (.I0(\Kp[3] ), .I1(n1[18]), .I2(n19208[1]), 
            .I3(n4_adj_5177), .O(n19159[2]));   // verilog/motorControl.v(34[16:22])
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h8778;
    SB_LUT4 i2_3_lut_4_lut_adj_1723 (.I0(\Kp[2] ), .I1(n1[19]), .I2(n19239[0]), 
            .I3(n38355), .O(n19208[1]));   // verilog/motorControl.v(34[16:22])
    defparam i2_3_lut_4_lut_adj_1723.LUT_INIT = 16'h8778;
    SB_LUT4 i24409_3_lut_4_lut (.I0(\Kp[2] ), .I1(n1[19]), .I2(n38355), 
            .I3(n19239[0]), .O(n4_adj_5172));   // verilog/motorControl.v(34[16:22])
    defparam i24409_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 i24396_2_lut_3_lut_4_lut (.I0(\Kp[0] ), .I1(n1[20]), .I2(n1[19]), 
            .I3(\Kp[1] ), .O(n19208[0]));   // verilog/motorControl.v(34[16:22])
    defparam i24396_2_lut_3_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 i24398_2_lut_3_lut_4_lut (.I0(\Kp[0] ), .I1(n1[20]), .I2(n1[19]), 
            .I3(\Kp[1] ), .O(n38355));   // verilog/motorControl.v(34[16:22])
    defparam i24398_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i24379_3_lut_4_lut (.I0(\Kp[2] ), .I1(n1[20]), .I2(n38323), 
            .I3(n19256[0]), .O(n4_adj_5180));   // verilog/motorControl.v(34[16:22])
    defparam i24379_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 i2_3_lut_4_lut_adj_1724 (.I0(\Kp[2] ), .I1(n1[20]), .I2(n19256[0]), 
            .I3(n38323), .O(n19239[1]));   // verilog/motorControl.v(34[16:22])
    defparam i2_3_lut_4_lut_adj_1724.LUT_INIT = 16'h8778;
    SB_LUT4 i24368_2_lut_3_lut_4_lut (.I0(\Kp[0] ), .I1(n1[21]), .I2(n1[20]), 
            .I3(\Kp[1] ), .O(n38323));   // verilog/motorControl.v(34[16:22])
    defparam i24368_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i24366_2_lut_3_lut_4_lut (.I0(\Kp[0] ), .I1(n1[21]), .I2(n1[20]), 
            .I3(\Kp[1] ), .O(n19239[0]));   // verilog/motorControl.v(34[16:22])
    defparam i24366_2_lut_3_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 i2_3_lut_4_lut_adj_1725 (.I0(\Kp[2] ), .I1(n1[18]), .I2(n19208[0]), 
            .I3(n38405), .O(n19159[1]));   // verilog/motorControl.v(34[16:22])
    defparam i2_3_lut_4_lut_adj_1725.LUT_INIT = 16'h8778;
    SB_LUT4 i24455_3_lut_4_lut (.I0(\Kp[2] ), .I1(n1[18]), .I2(n38405), 
            .I3(n19208[0]), .O(n4_adj_5177));   // verilog/motorControl.v(34[16:22])
    defparam i24455_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 i24442_2_lut_3_lut_4_lut (.I0(\Kp[0] ), .I1(n1[19]), .I2(n1[18]), 
            .I3(\Kp[1] ), .O(n19159[0]));   // verilog/motorControl.v(34[16:22])
    defparam i24442_2_lut_3_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 i24444_2_lut_3_lut_4_lut (.I0(\Kp[0] ), .I1(n1[19]), .I2(n1[18]), 
            .I3(\Kp[1] ), .O(n38405));   // verilog/motorControl.v(34[16:22])
    defparam i24444_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 mult_11_i230_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [16]), 
            .I2(GND_net), .I3(GND_net), .O(n341_adj_5157));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i230_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i279_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [16]), 
            .I2(GND_net), .I3(GND_net), .O(n414_adj_5156));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i279_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i328_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [16]), 
            .I2(GND_net), .I3(GND_net), .O(n487_adj_5153));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i328_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i377_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [16]), 
            .I2(GND_net), .I3(GND_net), .O(n560_adj_5152));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i377_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i67_2_lut (.I0(\Kp[1] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n98_adj_5151));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i67_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i20_2_lut (.I0(\Kp[0] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_5150));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i20_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i116_2_lut (.I0(\Kp[2] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n171_adj_5149));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i116_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i24295_3_lut_4_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [19]), 
            .I2(n38232), .I3(n19224[0]), .O(n4_adj_5035));   // verilog/motorControl.v(34[25:36])
    defparam i24295_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 i2_3_lut_4_lut_adj_1726 (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [19]), 
            .I2(n19224[0]), .I3(n38232), .O(n19184[1]));   // verilog/motorControl.v(34[25:36])
    defparam i2_3_lut_4_lut_adj_1726.LUT_INIT = 16'h8778;
    SB_LUT4 i24257_3_lut_4_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [20]), 
            .I2(n38191), .I3(n19248[0]), .O(n4_adj_5043));   // verilog/motorControl.v(34[25:36])
    defparam i24257_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 i2_3_lut_4_lut_adj_1727 (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [20]), 
            .I2(n19248[0]), .I3(n38191), .O(n19224[1]));   // verilog/motorControl.v(34[25:36])
    defparam i2_3_lut_4_lut_adj_1727.LUT_INIT = 16'h8778;
    SB_LUT4 i24246_2_lut_3_lut_4_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [21]), 
            .I2(\PID_CONTROLLER.integral_23__N_3836 [20]), .I3(\Ki[1] ), 
            .O(n38191));   // verilog/motorControl.v(34[25:36])
    defparam i24246_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i24244_2_lut_3_lut_4_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [21]), 
            .I2(\PID_CONTROLLER.integral_23__N_3836 [20]), .I3(\Ki[1] ), 
            .O(n19224[0]));   // verilog/motorControl.v(34[25:36])
    defparam i24244_2_lut_3_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 i24341_3_lut_4_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [18]), 
            .I2(n4_adj_5181), .I3(n19184[1]), .O(n6_adj_5023));   // verilog/motorControl.v(34[25:36])
    defparam i24341_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 mult_10_i165_2_lut (.I0(\Kp[3] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n244_adj_5148));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i165_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_3_lut_4_lut_adj_1728 (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [18]), 
            .I2(n19184[1]), .I3(n4_adj_5181), .O(n19124[2]));   // verilog/motorControl.v(34[25:36])
    defparam i2_3_lut_4_lut_adj_1728.LUT_INIT = 16'h8778;
    SB_LUT4 mult_11_i73_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n107_adj_5016));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i73_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_3_lut_4_lut_adj_1729 (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [18]), 
            .I2(n19184[0]), .I3(n38273), .O(n19124[1]));   // verilog/motorControl.v(34[25:36])
    defparam i2_3_lut_4_lut_adj_1729.LUT_INIT = 16'h8778;
    SB_LUT4 i24333_3_lut_4_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [18]), 
            .I2(n38273), .I3(n19184[0]), .O(n4_adj_5181));   // verilog/motorControl.v(34[25:36])
    defparam i24333_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 i24320_2_lut_3_lut_4_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [19]), 
            .I2(\PID_CONTROLLER.integral_23__N_3836 [18]), .I3(\Ki[1] ), 
            .O(n19124[0]));   // verilog/motorControl.v(34[25:36])
    defparam i24320_2_lut_3_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 mult_11_i26_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n38_adj_5015));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i26_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i214_2_lut (.I0(\Kp[4] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n317_adj_5147));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i214_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i122_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n180_adj_5014));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i122_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i171_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n253_adj_5012));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i171_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i220_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n326_adj_5011));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i220_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i269_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n399_adj_5010));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i269_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i318_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n472_adj_5009));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i318_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i367_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n545_adj_5008));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i367_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i263_2_lut (.I0(\Kp[5] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n390_adj_5146));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i263_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i77_2_lut (.I0(\Kp[1] ), .I1(n1[13]), .I2(GND_net), 
            .I3(GND_net), .O(n113));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i77_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i30_2_lut (.I0(\Kp[0] ), .I1(n1[14]), .I2(GND_net), 
            .I3(GND_net), .O(n44));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i30_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i20928_2_lut (.I0(n1[1]), .I1(\PID_CONTROLLER.integral_23__N_3884 ), 
            .I2(GND_net), .I3(GND_net), .O(n4751[1]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i20928_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i416_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n618_adj_5007));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i416_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i24322_2_lut_3_lut_4_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [19]), 
            .I2(\PID_CONTROLLER.integral_23__N_3836 [18]), .I3(\Ki[1] ), 
            .O(n38273));   // verilog/motorControl.v(34[25:36])
    defparam i24322_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i24282_2_lut_3_lut_4_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [20]), 
            .I2(\PID_CONTROLLER.integral_23__N_3836 [19]), .I3(\Ki[1] ), 
            .O(n19184[0]));   // verilog/motorControl.v(34[25:36])
    defparam i24282_2_lut_3_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 mult_10_i312_2_lut (.I0(\Kp[6] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n463_adj_5145));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i312_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i24284_2_lut_3_lut_4_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [20]), 
            .I2(\PID_CONTROLLER.integral_23__N_3836 [19]), .I3(\Ki[1] ), 
            .O(n38232));   // verilog/motorControl.v(34[25:36])
    defparam i24284_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 mult_10_i361_2_lut (.I0(\Kp[7] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n536_adj_5144));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i361_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i126_2_lut (.I0(\Kp[2] ), .I1(n1[13]), .I2(GND_net), 
            .I3(GND_net), .O(n186));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i126_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i20927_2_lut (.I0(n1[2]), .I1(\PID_CONTROLLER.integral_23__N_3884 ), 
            .I2(GND_net), .I3(GND_net), .O(n4751[2]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i20927_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i175_2_lut (.I0(\Kp[3] ), .I1(n1[13]), .I2(GND_net), 
            .I3(GND_net), .O(n259_adj_5006));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i175_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i1_1_lut (.I0(IntegralLimit[0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5234[0]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i161_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n238_adj_5143));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i161_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i465_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n691_adj_5005));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i465_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i20926_2_lut (.I0(n1[3]), .I1(\PID_CONTROLLER.integral_23__N_3884 ), 
            .I2(GND_net), .I3(GND_net), .O(n4751[3]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i20926_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i224_2_lut (.I0(\Kp[4] ), .I1(n1[13]), .I2(GND_net), 
            .I3(GND_net), .O(n332));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i224_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i514_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n764));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i514_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i20925_2_lut (.I0(n1[4]), .I1(\PID_CONTROLLER.integral_23__N_3884 ), 
            .I2(GND_net), .I3(GND_net), .O(n4751[4]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i20925_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i20924_2_lut (.I0(n1[5]), .I1(\PID_CONTROLLER.integral_23__N_3884 ), 
            .I2(GND_net), .I3(GND_net), .O(n4751[5]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i20924_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i20923_2_lut (.I0(n1[6]), .I1(\PID_CONTROLLER.integral_23__N_3884 ), 
            .I2(GND_net), .I3(GND_net), .O(n4751[6]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i20923_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i20922_2_lut (.I0(n1[7]), .I1(\PID_CONTROLLER.integral_23__N_3884 ), 
            .I2(GND_net), .I3(GND_net), .O(n4751[7]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i20922_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i410_2_lut (.I0(\Kp[8] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n609_adj_5142));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i410_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i273_2_lut (.I0(\Kp[5] ), .I1(n1[13]), .I2(GND_net), 
            .I3(GND_net), .O(n405));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i273_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i20921_2_lut (.I0(n1[8]), .I1(\PID_CONTROLLER.integral_23__N_3884 ), 
            .I2(GND_net), .I3(GND_net), .O(n4751[8]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i20921_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i563_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n837));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i563_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i210_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n311_adj_5141));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i210_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i612_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n910));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i612_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i322_2_lut (.I0(\Kp[6] ), .I1(n1[13]), .I2(GND_net), 
            .I3(GND_net), .O(n478));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i322_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i20920_2_lut (.I0(n1[9]), .I1(\PID_CONTROLLER.integral_23__N_3884 ), 
            .I2(GND_net), .I3(GND_net), .O(n4751[9]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i20920_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i371_2_lut (.I0(\Kp[7] ), .I1(n1[13]), .I2(GND_net), 
            .I3(GND_net), .O(n551));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i371_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i71_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n104));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i71_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i459_2_lut (.I0(\Kp[9] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n682_adj_5140));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i459_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i24_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_5004));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i24_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i508_2_lut (.I0(\Kp[10] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n755_adj_5139));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i508_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 IntegralLimit_23__I_0_i8_3_lut_3_lut (.I0(IntegralLimit[4]), .I1(IntegralLimit[8]), 
            .I2(\PID_CONTROLLER.integral [8]), .I3(GND_net), .O(n8_adj_4941));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i8_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 mult_10_i557_2_lut (.I0(\Kp[11] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n828_adj_5138));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i557_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 duty_23__I_937_i41_2_lut (.I0(PWMLimit[20]), .I1(duty_23__N_3936[20]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_5182));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_937_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_937_i39_2_lut (.I0(PWMLimit[19]), .I1(duty_23__N_3936[19]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_5183));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_937_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_937_i45_2_lut (.I0(PWMLimit[22]), .I1(duty_23__N_3936[22]), 
            .I2(GND_net), .I3(GND_net), .O(n45_adj_5184));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_937_i45_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_937_i37_2_lut (.I0(PWMLimit[18]), .I1(duty_23__N_3936[18]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_5185));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_937_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_937_i23_2_lut (.I0(PWMLimit[11]), .I1(duty_23__N_3936[11]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_5186));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_937_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_937_i25_2_lut (.I0(PWMLimit[12]), .I1(duty_23__N_3936[12]), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_5187));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_937_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_937_i43_2_lut (.I0(PWMLimit[21]), .I1(duty_23__N_3936[21]), 
            .I2(GND_net), .I3(GND_net), .O(n43_adj_5188));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_937_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_937_i29_2_lut (.I0(PWMLimit[14]), .I1(duty_23__N_3936[14]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_5189));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_937_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_10_i606_2_lut (.I0(\Kp[12] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n901_adj_5137));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i606_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 duty_23__I_937_i31_2_lut (.I0(PWMLimit[15]), .I1(duty_23__N_3936[15]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_5190));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_937_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_10_i655_2_lut (.I0(\Kp[13] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n974_adj_5136));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i655_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 duty_23__I_937_i35_2_lut (.I0(PWMLimit[17]), .I1(duty_23__N_3936[17]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_5191));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_937_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_937_i11_2_lut (.I0(PWMLimit[5]), .I1(duty_23__N_3936[5]), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_5192));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_937_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_937_i13_2_lut (.I0(PWMLimit[6]), .I1(duty_23__N_3936[6]), 
            .I2(GND_net), .I3(GND_net), .O(n13_adj_5193));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_937_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_937_i15_2_lut (.I0(PWMLimit[7]), .I1(duty_23__N_3936[7]), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_5194));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_937_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_937_i27_2_lut (.I0(PWMLimit[13]), .I1(duty_23__N_3936[13]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_5195));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_937_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_937_i33_2_lut (.I0(PWMLimit[16]), .I1(duty_23__N_3936[16]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_5196));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_937_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_937_i9_2_lut (.I0(PWMLimit[4]), .I1(duty_23__N_3936[4]), 
            .I2(GND_net), .I3(GND_net), .O(n9_adj_5197));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_937_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_937_i17_2_lut (.I0(PWMLimit[8]), .I1(duty_23__N_3936[8]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_5198));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_937_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_937_i19_2_lut (.I0(PWMLimit[9]), .I1(duty_23__N_3936[9]), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_5199));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_937_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_937_i21_2_lut (.I0(PWMLimit[10]), .I1(duty_23__N_3936[10]), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_5200));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_937_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i33984_4_lut (.I0(n21_adj_5200), .I1(n19_adj_5199), .I2(n17_adj_5198), 
            .I3(n9_adj_5197), .O(n49571));
    defparam i33984_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 mult_10_i704_2_lut (.I0(\Kp[14] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n1047_adj_5135));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i704_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i33976_4_lut (.I0(n27_adj_5195), .I1(n15_adj_5194), .I2(n13_adj_5193), 
            .I3(n11_adj_5192), .O(n49563));
    defparam i33976_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 duty_23__I_937_i12_3_lut (.I0(duty_23__N_3936[7]), .I1(duty_23__N_3936[16]), 
            .I2(n33_adj_5196), .I3(GND_net), .O(n12_adj_5201));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_937_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_937_i10_3_lut (.I0(duty_23__N_3936[5]), .I1(duty_23__N_3936[6]), 
            .I2(n13_adj_5193), .I3(GND_net), .O(n10_adj_5202));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_937_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_937_i30_3_lut (.I0(n12_adj_5201), .I1(duty_23__N_3936[17]), 
            .I2(n35_adj_5191), .I3(GND_net), .O(n30_adj_5203));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_937_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34309_4_lut (.I0(n13_adj_5193), .I1(n11_adj_5192), .I2(n9_adj_5197), 
            .I3(n49581), .O(n49897));
    defparam i34309_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i34305_4_lut (.I0(n19_adj_5199), .I1(n17_adj_5198), .I2(n15_adj_5194), 
            .I3(n49897), .O(n49893));
    defparam i34305_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i34754_4_lut (.I0(n25_adj_5187), .I1(n23_adj_5186), .I2(n21_adj_5200), 
            .I3(n49893), .O(n50342));
    defparam i34754_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 mult_10_i753_2_lut (.I0(\Kp[15] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n1120_adj_5134));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i753_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i34516_4_lut (.I0(n31_adj_5190), .I1(n29_adj_5189), .I2(n27_adj_5195), 
            .I3(n50342), .O(n50104));
    defparam i34516_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i34822_4_lut (.I0(n37_adj_5185), .I1(n35_adj_5191), .I2(n33_adj_5196), 
            .I3(n50104), .O(n50410));
    defparam i34822_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 duty_23__I_937_i16_3_lut (.I0(duty_23__N_3936[9]), .I1(duty_23__N_3936[21]), 
            .I2(n43_adj_5188), .I3(GND_net), .O(n16_adj_5204));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_937_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34548_3_lut (.I0(n6_adj_5170), .I1(duty_23__N_3936[10]), .I2(n21_adj_5200), 
            .I3(GND_net), .O(n50136));   // verilog/motorControl.v(36[10:25])
    defparam i34548_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34549_3_lut (.I0(n50136), .I1(duty_23__N_3936[11]), .I2(n23_adj_5186), 
            .I3(GND_net), .O(n50137));   // verilog/motorControl.v(36[10:25])
    defparam i34549_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_937_i8_3_lut (.I0(duty_23__N_3936[4]), .I1(duty_23__N_3936[8]), 
            .I2(n17_adj_5198), .I3(GND_net), .O(n8_adj_5205));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_937_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_937_i24_3_lut (.I0(n16_adj_5204), .I1(duty_23__N_3936[22]), 
            .I2(n45_adj_5184), .I3(GND_net), .O(n24_adj_5206));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_937_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i33959_4_lut (.I0(n43_adj_5188), .I1(n25_adj_5187), .I2(n23_adj_5186), 
            .I3(n49571), .O(n49546));
    defparam i33959_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i34664_4_lut (.I0(n24_adj_5206), .I1(n8_adj_5205), .I2(n45_adj_5184), 
            .I3(n49544), .O(n50252));   // verilog/motorControl.v(36[10:25])
    defparam i34664_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 mult_10_i65_2_lut (.I0(\Kp[1] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n95_adj_5133));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i65_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i18_2_lut (.I0(\Kp[0] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n26_adj_5132));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i18_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i34196_3_lut (.I0(n50137), .I1(duty_23__N_3936[12]), .I2(n25_adj_5187), 
            .I3(GND_net), .O(n49784));   // verilog/motorControl.v(36[10:25])
    defparam i34196_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_937_i4_4_lut (.I0(duty_23__N_3936[0]), .I1(duty_23__N_3936[1]), 
            .I2(PWMLimit[1]), .I3(PWMLimit[0]), .O(n4_adj_5207));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_937_i4_4_lut.LUT_INIT = 16'h0c8e;
    SB_LUT4 i34534_3_lut (.I0(n4_adj_5207), .I1(duty_23__N_3936[13]), .I2(n27_adj_5195), 
            .I3(GND_net), .O(n50122));   // verilog/motorControl.v(36[10:25])
    defparam i34534_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34535_3_lut (.I0(n50122), .I1(duty_23__N_3936[14]), .I2(n29_adj_5189), 
            .I3(GND_net), .O(n50123));   // verilog/motorControl.v(36[10:25])
    defparam i34535_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i33972_4_lut (.I0(n33_adj_5196), .I1(n31_adj_5190), .I2(n29_adj_5189), 
            .I3(n49563), .O(n49559));
    defparam i33972_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i20919_2_lut (.I0(n1[10]), .I1(\PID_CONTROLLER.integral_23__N_3884 ), 
            .I2(GND_net), .I3(GND_net), .O(n4751[10]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i20919_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i34742_4_lut (.I0(n30_adj_5203), .I1(n10_adj_5202), .I2(n35_adj_5191), 
            .I3(n49557), .O(n50330));   // verilog/motorControl.v(36[10:25])
    defparam i34742_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i34198_3_lut (.I0(n50123), .I1(duty_23__N_3936[15]), .I2(n31_adj_5190), 
            .I3(GND_net), .O(n49786));   // verilog/motorControl.v(36[10:25])
    defparam i34198_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34848_4_lut (.I0(n49786), .I1(n50330), .I2(n35_adj_5191), 
            .I3(n49559), .O(n50436));   // verilog/motorControl.v(36[10:25])
    defparam i34848_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i34849_3_lut (.I0(n50436), .I1(duty_23__N_3936[18]), .I2(n37_adj_5185), 
            .I3(GND_net), .O(n50437));   // verilog/motorControl.v(36[10:25])
    defparam i34849_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34827_3_lut (.I0(n50437), .I1(duty_23__N_3936[19]), .I2(n39_adj_5183), 
            .I3(GND_net), .O(n50415));   // verilog/motorControl.v(36[10:25])
    defparam i34827_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i33961_4_lut (.I0(n43_adj_5188), .I1(n41_adj_5182), .I2(n39_adj_5183), 
            .I3(n50410), .O(n49548));
    defparam i33961_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i34812_4_lut (.I0(n49784), .I1(n50252), .I2(n45_adj_5184), 
            .I3(n49546), .O(n50400));   // verilog/motorControl.v(36[10:25])
    defparam i34812_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i34204_3_lut (.I0(n50415), .I1(duty_23__N_3936[20]), .I2(n41_adj_5182), 
            .I3(GND_net), .O(n49792));   // verilog/motorControl.v(36[10:25])
    defparam i34204_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34814_4_lut (.I0(n49792), .I1(n50400), .I2(n45_adj_5184), 
            .I3(n49548), .O(n50402));   // verilog/motorControl.v(36[10:25])
    defparam i34814_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 mult_11_i259_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n384_adj_5131));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i259_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i114_2_lut (.I0(\Kp[2] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n168_adj_5130));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i114_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i308_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n457_adj_5129));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i308_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i163_2_lut (.I0(\Kp[3] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n241_adj_5128));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i163_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i34815_3_lut (.I0(n50402), .I1(PWMLimit[23]), .I2(duty_23__N_3936[23]), 
            .I3(GND_net), .O(duty_23__N_3935));   // verilog/motorControl.v(36[10:25])
    defparam i34815_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 LessThan_15_i39_2_lut (.I0(duty_23__N_3936[19]), .I1(n257[19]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_5208));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i41_2_lut (.I0(duty_23__N_3936[20]), .I1(n257[20]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_5209));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i45_2_lut (.I0(duty_23__N_3936[22]), .I1(n257[22]), 
            .I2(GND_net), .I3(GND_net), .O(n45_adj_5210));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i45_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i37_2_lut (.I0(duty_23__N_3936[18]), .I1(n257[18]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_5211));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i29_2_lut (.I0(duty_23__N_3936[14]), .I1(n257[14]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_5212));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i31_2_lut (.I0(duty_23__N_3936[15]), .I1(n257[15]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_5213));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_10_i420_2_lut (.I0(\Kp[8] ), .I1(n1[13]), .I2(GND_net), 
            .I3(GND_net), .O(n624));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i420_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_15_i23_2_lut (.I0(duty_23__N_3936[11]), .I1(n257[11]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_5214));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i25_2_lut (.I0(duty_23__N_3936[12]), .I1(n257[12]), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_5215));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i43_2_lut (.I0(duty_23__N_3936[21]), .I1(n257[21]), 
            .I2(GND_net), .I3(GND_net), .O(n43_adj_5216));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_10_i212_2_lut (.I0(\Kp[4] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n314_adj_5127));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i212_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i261_2_lut (.I0(\Kp[5] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n387_adj_5126));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i261_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_15_i35_2_lut (.I0(duty_23__N_3936[17]), .I1(n257[17]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_5217));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i33_2_lut (.I0(duty_23__N_3936[16]), .I1(n257[16]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_5218));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i11_2_lut (.I0(duty_23__N_3936[5]), .I1(n257[5]), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_5219));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i13_2_lut (.I0(duty_23__N_3936[6]), .I1(n257[6]), 
            .I2(GND_net), .I3(GND_net), .O(n13_adj_5220));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i15_2_lut (.I0(duty_23__N_3936[7]), .I1(n257[7]), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_5221));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i27_2_lut (.I0(duty_23__N_3936[13]), .I1(n257[13]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_5222));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i9_2_lut (.I0(duty_23__N_3936[4]), .I1(n257[4]), 
            .I2(GND_net), .I3(GND_net), .O(n9_adj_5223));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i17_2_lut (.I0(duty_23__N_3936[8]), .I1(n257[8]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_5224));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i19_2_lut (.I0(duty_23__N_3936[9]), .I1(n257[9]), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_5225));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i21_2_lut (.I0(duty_23__N_3936[10]), .I1(n257[10]), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_5226));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i33944_4_lut (.I0(n21_adj_5226), .I1(n19_adj_5225), .I2(n17_adj_5224), 
            .I3(n9_adj_5223), .O(n49531));
    defparam i33944_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i33933_4_lut (.I0(n27_adj_5222), .I1(n15_adj_5221), .I2(n13_adj_5220), 
            .I3(n11_adj_5219), .O(n49520));
    defparam i33933_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 LessThan_15_i12_3_lut (.I0(n257[7]), .I1(n257[16]), .I2(n33_adj_5218), 
            .I3(GND_net), .O(n12_adj_5227));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_15_i10_3_lut (.I0(n257[5]), .I1(n257[6]), .I2(n13_adj_5220), 
            .I3(GND_net), .O(n10_adj_5228));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_15_i30_3_lut (.I0(n12_adj_5227), .I1(n257[17]), .I2(n35_adj_5217), 
            .I3(GND_net), .O(n30_adj_5229));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_10_i310_2_lut (.I0(\Kp[6] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n460_adj_5125));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i310_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i34277_4_lut (.I0(n13_adj_5220), .I1(n11_adj_5219), .I2(n9_adj_5223), 
            .I3(n49542), .O(n49865));
    defparam i34277_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i34273_4_lut (.I0(n19_adj_5225), .I1(n17_adj_5224), .I2(n15_adj_5221), 
            .I3(n49865), .O(n49861));
    defparam i34273_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i34746_4_lut (.I0(n25_adj_5215), .I1(n23_adj_5214), .I2(n21_adj_5226), 
            .I3(n49861), .O(n50334));
    defparam i34746_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 mult_10_i359_2_lut (.I0(\Kp[7] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n533_adj_5124));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i359_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i34500_4_lut (.I0(n31_adj_5213), .I1(n29_adj_5212), .I2(n27_adj_5222), 
            .I3(n50334), .O(n50088));
    defparam i34500_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i34820_4_lut (.I0(n37_adj_5211), .I1(n35_adj_5217), .I2(n33_adj_5218), 
            .I3(n50088), .O(n50408));
    defparam i34820_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 LessThan_15_i16_3_lut (.I0(n257[9]), .I1(n257[21]), .I2(n43_adj_5216), 
            .I3(GND_net), .O(n16_adj_5230));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34524_3_lut (.I0(n6_adj_5154), .I1(n257[10]), .I2(n21_adj_5226), 
            .I3(GND_net), .O(n50112));   // verilog/motorControl.v(38[19:35])
    defparam i34524_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34525_3_lut (.I0(n50112), .I1(n257[11]), .I2(n23_adj_5214), 
            .I3(GND_net), .O(n50113));   // verilog/motorControl.v(38[19:35])
    defparam i34525_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_15_i8_3_lut (.I0(n257[4]), .I1(n257[8]), .I2(n17_adj_5224), 
            .I3(GND_net), .O(n8_adj_5231));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_10_i408_2_lut (.I0(\Kp[8] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n606_adj_5123));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i408_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_15_i24_3_lut (.I0(n16_adj_5230), .I1(n257[22]), .I2(n45_adj_5210), 
            .I3(GND_net), .O(n24_adj_5232));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i33902_4_lut (.I0(n43_adj_5216), .I1(n25_adj_5215), .I2(n23_adj_5214), 
            .I3(n49531), .O(n49489));
    defparam i33902_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i34666_4_lut (.I0(n24_adj_5232), .I1(n8_adj_5231), .I2(n45_adj_5210), 
            .I3(n49485), .O(n50254));   // verilog/motorControl.v(38[19:35])
    defparam i34666_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i34206_3_lut (.I0(n50113), .I1(n257[12]), .I2(n25_adj_5215), 
            .I3(GND_net), .O(n49794));   // verilog/motorControl.v(38[19:35])
    defparam i34206_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_15_i4_4_lut (.I0(duty_23__N_3936[0]), .I1(n257[1]), 
            .I2(duty_23__N_3936[1]), .I3(n257[0]), .O(n4_adj_5233));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i4_4_lut.LUT_INIT = 16'h4d0c;
    SB_LUT4 i34520_3_lut (.I0(n4_adj_5233), .I1(n257[13]), .I2(n27_adj_5222), 
            .I3(GND_net), .O(n50108));   // verilog/motorControl.v(38[19:35])
    defparam i34520_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34521_3_lut (.I0(n50108), .I1(n257[14]), .I2(n29_adj_5212), 
            .I3(GND_net), .O(n50109));   // verilog/motorControl.v(38[19:35])
    defparam i34521_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i33924_4_lut (.I0(n33_adj_5218), .I1(n31_adj_5213), .I2(n29_adj_5212), 
            .I3(n49520), .O(n49511));
    defparam i33924_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 mult_11_i357_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n530_adj_5122));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i357_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i34748_4_lut (.I0(n30_adj_5229), .I1(n10_adj_5228), .I2(n35_adj_5217), 
            .I3(n49506), .O(n50336));   // verilog/motorControl.v(38[19:35])
    defparam i34748_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i34208_3_lut (.I0(n50109), .I1(n257[15]), .I2(n31_adj_5213), 
            .I3(GND_net), .O(n49796));   // verilog/motorControl.v(38[19:35])
    defparam i34208_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34844_4_lut (.I0(n49796), .I1(n50336), .I2(n35_adj_5217), 
            .I3(n49511), .O(n50432));   // verilog/motorControl.v(38[19:35])
    defparam i34844_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i34845_3_lut (.I0(n50432), .I1(n257[18]), .I2(n37_adj_5211), 
            .I3(GND_net), .O(n50433));   // verilog/motorControl.v(38[19:35])
    defparam i34845_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34825_3_lut (.I0(n50433), .I1(n257[19]), .I2(n39_adj_5208), 
            .I3(GND_net), .O(n50413));   // verilog/motorControl.v(38[19:35])
    defparam i34825_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_11_i406_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n603_adj_5121));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i406_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i33904_4_lut (.I0(n43_adj_5216), .I1(n41_adj_5209), .I2(n39_adj_5208), 
            .I3(n50408), .O(n49491));
    defparam i33904_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i34816_4_lut (.I0(n49794), .I1(n50254), .I2(n45_adj_5210), 
            .I3(n49489), .O(n50404));   // verilog/motorControl.v(38[19:35])
    defparam i34816_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i34214_3_lut (.I0(n50413), .I1(n257[20]), .I2(n41_adj_5209), 
            .I3(GND_net), .O(n49802));   // verilog/motorControl.v(38[19:35])
    defparam i34214_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34818_4_lut (.I0(n49802), .I1(n50404), .I2(n45_adj_5210), 
            .I3(n49491), .O(n50406));   // verilog/motorControl.v(38[19:35])
    defparam i34818_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 mult_11_i455_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n676_adj_5120));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i455_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i34819_3_lut (.I0(n50406), .I1(duty_23__N_3936[23]), .I2(n257[23]), 
            .I3(GND_net), .O(n256_adj_4995));   // verilog/motorControl.v(38[19:35])
    defparam i34819_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 mux_17_i1_3_lut (.I0(duty_23__N_3936[0]), .I1(n257[0]), .I2(n256_adj_4995), 
            .I3(GND_net), .O(duty_23__N_3911[0]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i1_3_lut (.I0(duty_23__N_3911[0]), .I1(PWMLimit[0]), 
            .I2(duty_23__N_3935), .I3(GND_net), .O(duty_23__N_3812[0]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_11_i504_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n749_adj_5119));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i504_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i457_2_lut (.I0(\Kp[9] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n679_adj_5118));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i457_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i553_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n822_adj_5117));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i553_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i602_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n895_adj_5116));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i602_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i77_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [13]), 
            .I2(GND_net), .I3(GND_net), .O(n113_adj_5115));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i77_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i30_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [14]), 
            .I2(GND_net), .I3(GND_net), .O(n44_adj_5114));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i30_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i126_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [13]), 
            .I2(GND_net), .I3(GND_net), .O(n186_adj_5113));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i126_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i506_2_lut (.I0(\Kp[10] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n752_adj_5112));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i506_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i555_2_lut (.I0(\Kp[11] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n825_adj_5111));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i555_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i175_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [13]), 
            .I2(GND_net), .I3(GND_net), .O(n259_adj_5110));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i175_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i604_2_lut (.I0(\Kp[12] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n898));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i604_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i224_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [13]), 
            .I2(GND_net), .I3(GND_net), .O(n332_adj_5109));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i224_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i653_2_lut (.I0(\Kp[13] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n971));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i653_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i651_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n968_adj_5108));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i651_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i273_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [13]), 
            .I2(GND_net), .I3(GND_net), .O(n405_adj_5107));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i273_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i2_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n155[0]));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i2_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i2_2_lut (.I0(\Kp[0] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n106[0]));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i2_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i322_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [13]), 
            .I2(GND_net), .I3(GND_net), .O(n478_adj_5106));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i322_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i371_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [13]), 
            .I2(GND_net), .I3(GND_net), .O(n551_adj_5105));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i371_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i702_2_lut (.I0(\Kp[14] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n1044));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i702_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i751_2_lut (.I0(\Kp[15] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n1117));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i751_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i700_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n1041_adj_5104));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i700_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i420_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [13]), 
            .I2(GND_net), .I3(GND_net), .O(n624_adj_5103));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i420_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i749_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n1114_adj_5102));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i749_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i81_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [15]), 
            .I2(GND_net), .I3(GND_net), .O(n119_adj_5101));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i81_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i34_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [16]), 
            .I2(GND_net), .I3(GND_net), .O(n50_adj_5100));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i34_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i469_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [13]), 
            .I2(GND_net), .I3(GND_net), .O(n697_adj_5099));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i469_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i75_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n110_adj_5098));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i75_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i28_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [13]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_5097));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i28_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i130_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [15]), 
            .I2(GND_net), .I3(GND_net), .O(n192_adj_5096));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i130_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i518_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [13]), 
            .I2(GND_net), .I3(GND_net), .O(n770_adj_5095));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i518_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i179_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [15]), 
            .I2(GND_net), .I3(GND_net), .O(n265_adj_5094));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i179_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i228_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [15]), 
            .I2(GND_net), .I3(GND_net), .O(n338_adj_5093));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i228_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i277_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [15]), 
            .I2(GND_net), .I3(GND_net), .O(n411_adj_5092));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i277_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i326_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [15]), 
            .I2(GND_net), .I3(GND_net), .O(n484_adj_5091));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i326_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i375_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [15]), 
            .I2(GND_net), .I3(GND_net), .O(n557_adj_5090));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i375_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i424_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [15]), 
            .I2(GND_net), .I3(GND_net), .O(n630_adj_5089));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i424_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i63_2_lut (.I0(\Kp[1] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n92));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i63_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i16_2_lut (.I0(\Kp[0] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_5088));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i16_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i112_2_lut (.I0(\Kp[2] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n165));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i112_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i161_2_lut (.I0(\Kp[3] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n238));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i161_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i210_2_lut (.I0(\Kp[4] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n311));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i210_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i124_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3836 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n183_adj_5087));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i124_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i259_2_lut (.I0(\Kp[5] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n384));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i259_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i308_2_lut (.I0(\Kp[6] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n457));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i308_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i357_2_lut (.I0(\Kp[7] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n530));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i357_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i406_2_lut (.I0(\Kp[8] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n603));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i406_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i455_2_lut (.I0(\Kp[9] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n676));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i455_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i504_2_lut (.I0(\Kp[10] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n749));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i504_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i553_2_lut (.I0(\Kp[11] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n822));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i553_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i602_2_lut (.I0(\Kp[12] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n895));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i602_2_lut.LUT_INIT = 16'h8888;
    
endmodule
//
// Verilog Description of module pll32MHz
//

module pll32MHz (GND_net, CLK_c, VCC_net, clk32MHz) /* synthesis syn_module_defined=1 */ ;
    input GND_net;
    input CLK_c;
    input VCC_net;
    output clk32MHz;
    
    wire CLK_c /* synthesis SET_AS_NETWORK=CLK_c, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(3[9:12])
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    
    SB_PLL40_CORE pll32MHz_inst (.REFERENCECLK(CLK_c), .PLLOUTGLOBAL(clk32MHz), 
            .BYPASS(GND_net), .RESETB(VCC_net)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=52, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=34, LSE_RLINE=37 */ ;   // verilog/TinyFPGA_B.v(34[10] 37[2])
    defparam pll32MHz_inst.FEEDBACK_PATH = "PHASE_AND_DELAY";
    defparam pll32MHz_inst.DELAY_ADJUSTMENT_MODE_FEEDBACK = "FIXED";
    defparam pll32MHz_inst.DELAY_ADJUSTMENT_MODE_RELATIVE = "FIXED";
    defparam pll32MHz_inst.SHIFTREG_DIV_MODE = 2'b00;
    defparam pll32MHz_inst.FDA_FEEDBACK = 4'b0000;
    defparam pll32MHz_inst.FDA_RELATIVE = 4'b0000;
    defparam pll32MHz_inst.PLLOUT_SELECT = "SHIFTREG_0deg";
    defparam pll32MHz_inst.DIVR = 4'b0000;
    defparam pll32MHz_inst.DIVF = 7'b0000001;
    defparam pll32MHz_inst.DIVQ = 3'b011;
    defparam pll32MHz_inst.FILTER_RANGE = 3'b001;
    defparam pll32MHz_inst.ENABLE_ICEGATE = 1'b0;
    defparam pll32MHz_inst.TEST_MODE = 1'b0;
    defparam pll32MHz_inst.EXTERNAL_DIVIDE_FACTOR = 1;
    
endmodule
//
// Verilog Description of module \quadrature_decoder(1,500000)_U0 
//

module \quadrature_decoder(1,500000)_U0  (b_prev, n1891, encoder0_position, 
            GND_net, a_new, direction_N_4071, ENCODER0_B_N_keep, ENCODER0_A_N_keep, 
            VCC_net, n29249, n1855) /* synthesis lattice_noprune=1 */ ;
    output b_prev;
    input n1891;
    output [31:0]encoder0_position;
    input GND_net;
    output [1:0]a_new;
    output direction_N_4071;
    input ENCODER0_B_N_keep;
    input ENCODER0_A_N_keep;
    input VCC_net;
    input n29249;
    output n1855;
    
    
    wire n29166, n29163, a_prev, n39449, direction_N_4070, n39450;
    wire [31:0]n133;
    
    wire n39448, n39447;
    wire [1:0]b_new;   // vhdl/quadrature_decoder.vhd(41[9:14])
    
    wire direction_N_4074, debounce_cnt, n39446, n39445, n39444;
    wire [1:0]a_new_c;   // vhdl/quadrature_decoder.vhd(40[9:14])
    
    wire n39443, n39442, n39441, n39440, a_prev_N_4077, n39470, 
        n39469, n39468, n39467, n39466, n39465, n39464, n39463, 
        n39462, n39461, n39460, n39459, n39458, n39457, n39456, 
        n39455, n39454, n39453, n39452, n39451;
    
    SB_DFF b_prev_52 (.Q(b_prev), .C(n1891), .D(n29166));   // vhdl/quadrature_decoder.vhd(52[3] 89[10])
    SB_DFF a_prev_51 (.Q(a_prev), .C(n1891), .D(n29163));   // vhdl/quadrature_decoder.vhd(52[3] 89[10])
    SB_CARRY position_2257_add_4_12 (.CI(n39449), .I0(direction_N_4070), 
            .I1(encoder0_position[10]), .CO(n39450));
    SB_LUT4 position_2257_add_4_11_lut (.I0(GND_net), .I1(direction_N_4070), 
            .I2(encoder0_position[9]), .I3(n39448), .O(n133[9])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2257_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2257_add_4_11 (.CI(n39448), .I0(direction_N_4070), 
            .I1(encoder0_position[9]), .CO(n39449));
    SB_LUT4 position_2257_add_4_10_lut (.I0(GND_net), .I1(direction_N_4070), 
            .I2(encoder0_position[8]), .I3(n39447), .O(n133[8])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2257_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2257_add_4_10 (.CI(n39447), .I0(direction_N_4070), 
            .I1(encoder0_position[8]), .CO(n39448));
    SB_LUT4 b_prev_I_0_65_2_lut (.I0(b_prev), .I1(b_new[1]), .I2(GND_net), 
            .I3(GND_net), .O(direction_N_4074));   // vhdl/quadrature_decoder.vhd(80[37:56])
    defparam b_prev_I_0_65_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 debounce_cnt_I_0_4_lut (.I0(debounce_cnt), .I1(a_prev), .I2(direction_N_4074), 
            .I3(a_new[1]), .O(direction_N_4071));   // vhdl/quadrature_decoder.vhd(79[10] 80[64])
    defparam debounce_cnt_I_0_4_lut.LUT_INIT = 16'ha2a8;
    SB_LUT4 position_2257_add_4_9_lut (.I0(GND_net), .I1(direction_N_4070), 
            .I2(encoder0_position[7]), .I3(n39446), .O(n133[7])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2257_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2257_add_4_9 (.CI(n39446), .I0(direction_N_4070), 
            .I1(encoder0_position[7]), .CO(n39447));
    SB_LUT4 position_2257_add_4_8_lut (.I0(GND_net), .I1(direction_N_4070), 
            .I2(encoder0_position[6]), .I3(n39445), .O(n133[6])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2257_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2257_add_4_8 (.CI(n39445), .I0(direction_N_4070), 
            .I1(encoder0_position[6]), .CO(n39446));
    SB_LUT4 position_2257_add_4_7_lut (.I0(GND_net), .I1(direction_N_4070), 
            .I2(encoder0_position[5]), .I3(n39444), .O(n133[5])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2257_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_DFF b_new_i0 (.Q(b_new[0]), .C(n1891), .D(ENCODER0_B_N_keep));   // vhdl/quadrature_decoder.vhd(52[3] 89[10])
    SB_CARRY position_2257_add_4_7 (.CI(n39444), .I0(direction_N_4070), 
            .I1(encoder0_position[5]), .CO(n39445));
    SB_DFF a_new_i0 (.Q(a_new_c[0]), .C(n1891), .D(ENCODER0_A_N_keep));   // vhdl/quadrature_decoder.vhd(52[3] 89[10])
    SB_LUT4 position_2257_add_4_6_lut (.I0(GND_net), .I1(direction_N_4070), 
            .I2(encoder0_position[4]), .I3(n39443), .O(n133[4])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2257_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2257_add_4_6 (.CI(n39443), .I0(direction_N_4070), 
            .I1(encoder0_position[4]), .CO(n39444));
    SB_LUT4 position_2257_add_4_5_lut (.I0(GND_net), .I1(direction_N_4070), 
            .I2(encoder0_position[3]), .I3(n39442), .O(n133[3])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2257_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2257_add_4_5 (.CI(n39442), .I0(direction_N_4070), 
            .I1(encoder0_position[3]), .CO(n39443));
    SB_LUT4 position_2257_add_4_4_lut (.I0(GND_net), .I1(direction_N_4070), 
            .I2(encoder0_position[2]), .I3(n39441), .O(n133[2])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2257_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2257_add_4_4 (.CI(n39441), .I0(direction_N_4070), 
            .I1(encoder0_position[2]), .CO(n39442));
    SB_LUT4 position_2257_add_4_3_lut (.I0(GND_net), .I1(direction_N_4070), 
            .I2(encoder0_position[1]), .I3(n39440), .O(n133[1])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2257_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2257_add_4_3 (.CI(n39440), .I0(direction_N_4070), 
            .I1(encoder0_position[1]), .CO(n39441));
    SB_LUT4 position_2257_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(encoder0_position[0]), 
            .I3(VCC_net), .O(n133[0])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2257_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2257_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(encoder0_position[0]), 
            .CO(n39440));
    SB_DFF debounce_cnt_50 (.Q(debounce_cnt), .C(n1891), .D(a_prev_N_4077));   // vhdl/quadrature_decoder.vhd(52[3] 89[10])
    SB_DFFE position_2257__i31 (.Q(encoder0_position[31]), .C(n1891), .E(direction_N_4071), 
            .D(n133[31]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2257__i30 (.Q(encoder0_position[30]), .C(n1891), .E(direction_N_4071), 
            .D(n133[30]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2257__i29 (.Q(encoder0_position[29]), .C(n1891), .E(direction_N_4071), 
            .D(n133[29]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2257__i28 (.Q(encoder0_position[28]), .C(n1891), .E(direction_N_4071), 
            .D(n133[28]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2257__i27 (.Q(encoder0_position[27]), .C(n1891), .E(direction_N_4071), 
            .D(n133[27]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2257__i26 (.Q(encoder0_position[26]), .C(n1891), .E(direction_N_4071), 
            .D(n133[26]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2257__i25 (.Q(encoder0_position[25]), .C(n1891), .E(direction_N_4071), 
            .D(n133[25]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2257__i24 (.Q(encoder0_position[24]), .C(n1891), .E(direction_N_4071), 
            .D(n133[24]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2257__i23 (.Q(encoder0_position[23]), .C(n1891), .E(direction_N_4071), 
            .D(n133[23]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2257__i22 (.Q(encoder0_position[22]), .C(n1891), .E(direction_N_4071), 
            .D(n133[22]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2257__i21 (.Q(encoder0_position[21]), .C(n1891), .E(direction_N_4071), 
            .D(n133[21]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2257__i20 (.Q(encoder0_position[20]), .C(n1891), .E(direction_N_4071), 
            .D(n133[20]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2257__i19 (.Q(encoder0_position[19]), .C(n1891), .E(direction_N_4071), 
            .D(n133[19]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2257__i18 (.Q(encoder0_position[18]), .C(n1891), .E(direction_N_4071), 
            .D(n133[18]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2257__i17 (.Q(encoder0_position[17]), .C(n1891), .E(direction_N_4071), 
            .D(n133[17]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2257__i16 (.Q(encoder0_position[16]), .C(n1891), .E(direction_N_4071), 
            .D(n133[16]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2257__i15 (.Q(encoder0_position[15]), .C(n1891), .E(direction_N_4071), 
            .D(n133[15]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2257__i14 (.Q(encoder0_position[14]), .C(n1891), .E(direction_N_4071), 
            .D(n133[14]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2257__i13 (.Q(encoder0_position[13]), .C(n1891), .E(direction_N_4071), 
            .D(n133[13]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2257__i12 (.Q(encoder0_position[12]), .C(n1891), .E(direction_N_4071), 
            .D(n133[12]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2257__i11 (.Q(encoder0_position[11]), .C(n1891), .E(direction_N_4071), 
            .D(n133[11]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2257__i10 (.Q(encoder0_position[10]), .C(n1891), .E(direction_N_4071), 
            .D(n133[10]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2257__i9 (.Q(encoder0_position[9]), .C(n1891), .E(direction_N_4071), 
            .D(n133[9]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2257__i8 (.Q(encoder0_position[8]), .C(n1891), .E(direction_N_4071), 
            .D(n133[8]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2257__i7 (.Q(encoder0_position[7]), .C(n1891), .E(direction_N_4071), 
            .D(n133[7]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2257__i6 (.Q(encoder0_position[6]), .C(n1891), .E(direction_N_4071), 
            .D(n133[6]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2257__i5 (.Q(encoder0_position[5]), .C(n1891), .E(direction_N_4071), 
            .D(n133[5]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2257__i4 (.Q(encoder0_position[4]), .C(n1891), .E(direction_N_4071), 
            .D(n133[4]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2257__i3 (.Q(encoder0_position[3]), .C(n1891), .E(direction_N_4071), 
            .D(n133[3]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2257__i2 (.Q(encoder0_position[2]), .C(n1891), .E(direction_N_4071), 
            .D(n133[2]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2257__i1 (.Q(encoder0_position[1]), .C(n1891), .E(direction_N_4071), 
            .D(n133[1]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2257__i0 (.Q(encoder0_position[0]), .C(n1891), .E(direction_N_4071), 
            .D(n133[0]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFF a_new_i1 (.Q(a_new[1]), .C(n1891), .D(a_new_c[0]));   // vhdl/quadrature_decoder.vhd(52[3] 89[10])
    SB_DFF b_new_i1 (.Q(b_new[1]), .C(n1891), .D(b_new[0]));   // vhdl/quadrature_decoder.vhd(52[3] 89[10])
    SB_LUT4 position_2257_add_4_33_lut (.I0(GND_net), .I1(direction_N_4070), 
            .I2(encoder0_position[31]), .I3(n39470), .O(n133[31])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2257_add_4_33_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 position_2257_add_4_32_lut (.I0(GND_net), .I1(direction_N_4070), 
            .I2(encoder0_position[30]), .I3(n39469), .O(n133[30])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2257_add_4_32_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2257_add_4_32 (.CI(n39469), .I0(direction_N_4070), 
            .I1(encoder0_position[30]), .CO(n39470));
    SB_LUT4 position_2257_add_4_31_lut (.I0(GND_net), .I1(direction_N_4070), 
            .I2(encoder0_position[29]), .I3(n39468), .O(n133[29])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2257_add_4_31_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2257_add_4_31 (.CI(n39468), .I0(direction_N_4070), 
            .I1(encoder0_position[29]), .CO(n39469));
    SB_LUT4 position_2257_add_4_30_lut (.I0(GND_net), .I1(direction_N_4070), 
            .I2(encoder0_position[28]), .I3(n39467), .O(n133[28])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2257_add_4_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2257_add_4_30 (.CI(n39467), .I0(direction_N_4070), 
            .I1(encoder0_position[28]), .CO(n39468));
    SB_LUT4 position_2257_add_4_29_lut (.I0(GND_net), .I1(direction_N_4070), 
            .I2(encoder0_position[27]), .I3(n39466), .O(n133[27])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2257_add_4_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2257_add_4_29 (.CI(n39466), .I0(direction_N_4070), 
            .I1(encoder0_position[27]), .CO(n39467));
    SB_LUT4 position_2257_add_4_28_lut (.I0(GND_net), .I1(direction_N_4070), 
            .I2(encoder0_position[26]), .I3(n39465), .O(n133[26])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2257_add_4_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2257_add_4_28 (.CI(n39465), .I0(direction_N_4070), 
            .I1(encoder0_position[26]), .CO(n39466));
    SB_LUT4 position_2257_add_4_27_lut (.I0(GND_net), .I1(direction_N_4070), 
            .I2(encoder0_position[25]), .I3(n39464), .O(n133[25])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2257_add_4_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2257_add_4_27 (.CI(n39464), .I0(direction_N_4070), 
            .I1(encoder0_position[25]), .CO(n39465));
    SB_LUT4 position_2257_add_4_26_lut (.I0(GND_net), .I1(direction_N_4070), 
            .I2(encoder0_position[24]), .I3(n39463), .O(n133[24])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2257_add_4_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2257_add_4_26 (.CI(n39463), .I0(direction_N_4070), 
            .I1(encoder0_position[24]), .CO(n39464));
    SB_LUT4 position_2257_add_4_25_lut (.I0(GND_net), .I1(direction_N_4070), 
            .I2(encoder0_position[23]), .I3(n39462), .O(n133[23])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2257_add_4_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2257_add_4_25 (.CI(n39462), .I0(direction_N_4070), 
            .I1(encoder0_position[23]), .CO(n39463));
    SB_LUT4 position_2257_add_4_24_lut (.I0(GND_net), .I1(direction_N_4070), 
            .I2(encoder0_position[22]), .I3(n39461), .O(n133[22])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2257_add_4_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2257_add_4_24 (.CI(n39461), .I0(direction_N_4070), 
            .I1(encoder0_position[22]), .CO(n39462));
    SB_LUT4 position_2257_add_4_23_lut (.I0(GND_net), .I1(direction_N_4070), 
            .I2(encoder0_position[21]), .I3(n39460), .O(n133[21])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2257_add_4_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2257_add_4_23 (.CI(n39460), .I0(direction_N_4070), 
            .I1(encoder0_position[21]), .CO(n39461));
    SB_LUT4 position_2257_add_4_22_lut (.I0(GND_net), .I1(direction_N_4070), 
            .I2(encoder0_position[20]), .I3(n39459), .O(n133[20])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2257_add_4_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2257_add_4_22 (.CI(n39459), .I0(direction_N_4070), 
            .I1(encoder0_position[20]), .CO(n39460));
    SB_LUT4 position_2257_add_4_21_lut (.I0(GND_net), .I1(direction_N_4070), 
            .I2(encoder0_position[19]), .I3(n39458), .O(n133[19])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2257_add_4_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2257_add_4_21 (.CI(n39458), .I0(direction_N_4070), 
            .I1(encoder0_position[19]), .CO(n39459));
    SB_LUT4 position_2257_add_4_20_lut (.I0(GND_net), .I1(direction_N_4070), 
            .I2(encoder0_position[18]), .I3(n39457), .O(n133[18])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2257_add_4_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2257_add_4_20 (.CI(n39457), .I0(direction_N_4070), 
            .I1(encoder0_position[18]), .CO(n39458));
    SB_LUT4 position_2257_add_4_19_lut (.I0(GND_net), .I1(direction_N_4070), 
            .I2(encoder0_position[17]), .I3(n39456), .O(n133[17])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2257_add_4_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2257_add_4_19 (.CI(n39456), .I0(direction_N_4070), 
            .I1(encoder0_position[17]), .CO(n39457));
    SB_LUT4 b_prev_I_0_63_2_lut (.I0(b_prev), .I1(a_new[1]), .I2(GND_net), 
            .I3(GND_net), .O(direction_N_4070));   // vhdl/quadrature_decoder.vhd(81[18:37])
    defparam b_prev_I_0_63_2_lut.LUT_INIT = 16'h9999;
    SB_DFF direction_57 (.Q(n1855), .C(n1891), .D(n29249));   // vhdl/quadrature_decoder.vhd(52[3] 89[10])
    SB_LUT4 position_2257_add_4_18_lut (.I0(GND_net), .I1(direction_N_4070), 
            .I2(encoder0_position[16]), .I3(n39455), .O(n133[16])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2257_add_4_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2257_add_4_18 (.CI(n39455), .I0(direction_N_4070), 
            .I1(encoder0_position[16]), .CO(n39456));
    SB_LUT4 position_2257_add_4_17_lut (.I0(GND_net), .I1(direction_N_4070), 
            .I2(encoder0_position[15]), .I3(n39454), .O(n133[15])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2257_add_4_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2257_add_4_17 (.CI(n39454), .I0(direction_N_4070), 
            .I1(encoder0_position[15]), .CO(n39455));
    SB_LUT4 position_2257_add_4_16_lut (.I0(GND_net), .I1(direction_N_4070), 
            .I2(encoder0_position[14]), .I3(n39453), .O(n133[14])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2257_add_4_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2257_add_4_16 (.CI(n39453), .I0(direction_N_4070), 
            .I1(encoder0_position[14]), .CO(n39454));
    SB_LUT4 position_2257_add_4_15_lut (.I0(GND_net), .I1(direction_N_4070), 
            .I2(encoder0_position[13]), .I3(n39452), .O(n133[13])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2257_add_4_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2257_add_4_15 (.CI(n39452), .I0(direction_N_4070), 
            .I1(encoder0_position[13]), .CO(n39453));
    SB_LUT4 position_2257_add_4_14_lut (.I0(GND_net), .I1(direction_N_4070), 
            .I2(encoder0_position[12]), .I3(n39451), .O(n133[12])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2257_add_4_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2257_add_4_14 (.CI(n39451), .I0(direction_N_4070), 
            .I1(encoder0_position[12]), .CO(n39452));
    SB_LUT4 position_2257_add_4_13_lut (.I0(GND_net), .I1(direction_N_4070), 
            .I2(encoder0_position[11]), .I3(n39450), .O(n133[11])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2257_add_4_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2257_add_4_13 (.CI(n39450), .I0(direction_N_4070), 
            .I1(encoder0_position[11]), .CO(n39451));
    SB_LUT4 position_2257_add_4_12_lut (.I0(GND_net), .I1(direction_N_4070), 
            .I2(encoder0_position[10]), .I3(n39449), .O(n133[10])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2257_add_4_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15218_3_lut_4_lut (.I0(debounce_cnt), .I1(a_prev_N_4077), .I2(b_new[1]), 
            .I3(b_prev), .O(n29166));   // vhdl/quadrature_decoder.vhd(52[3] 89[10])
    defparam i15218_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i15215_3_lut_4_lut (.I0(debounce_cnt), .I1(a_prev_N_4077), .I2(a_new[1]), 
            .I3(a_prev), .O(n29163));   // vhdl/quadrature_decoder.vhd(52[3] 89[10])
    defparam i15215_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i34896_4_lut (.I0(a_new_c[0]), .I1(b_new[0]), .I2(a_new[1]), 
            .I3(b_new[1]), .O(a_prev_N_4077));   // vhdl/quadrature_decoder.vhd(52[3] 89[10])
    defparam i34896_4_lut.LUT_INIT = 16'h8421;
    
endmodule
//
// Verilog Description of module \grp_debouncer(3,1000) 
//

module \grp_debouncer(3,1000)  (n29162, data_o, CLK_c, n29161, reg_B, 
            n46440, data_i, n29025, GND_net, VCC_net);
    input n29162;
    output [2:0]data_o;
    input CLK_c;
    input n29161;
    output [2:0]reg_B;
    output n46440;
    input [2:0]data_i;
    input n29025;
    input GND_net;
    input VCC_net;
    
    wire CLK_c /* synthesis SET_AS_NETWORK=CLK_c, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(3[9:12])
    wire [2:0]reg_A;   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(142[12:17])
    
    wire n6, cnt_next_9__N_836;
    wire [9:0]n45;
    wire [9:0]cnt_reg;   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(149[12:19])
    
    wire n16, n17, n39376, n39375, n39374, n39373, n39372, n39371, 
        n39370, n39369, n39368;
    
    SB_DFF reg_out_i0_i1 (.Q(data_o[1]), .C(CLK_c), .D(n29162));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    SB_DFF reg_out_i0_i2 (.Q(data_o[2]), .C(CLK_c), .D(n29161));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    SB_DFF reg_B_i0 (.Q(reg_B[0]), .C(CLK_c), .D(reg_A[0]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_LUT4 i2_4_lut (.I0(reg_B[0]), .I1(reg_B[1]), .I2(reg_A[0]), .I3(reg_A[1]), 
            .O(n6));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[40:72])
    defparam i2_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 i3_4_lut (.I0(n46440), .I1(n6), .I2(reg_B[2]), .I3(reg_A[2]), 
            .O(cnt_next_9__N_836));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[40:72])
    defparam i3_4_lut.LUT_INIT = 16'hdffd;
    SB_DFF reg_B_i2 (.Q(reg_B[2]), .C(CLK_c), .D(reg_A[2]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_DFF reg_B_i1 (.Q(reg_B[1]), .C(CLK_c), .D(reg_A[1]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_DFF reg_A_i1 (.Q(reg_A[1]), .C(CLK_c), .D(data_i[1]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_DFF reg_A_i0 (.Q(reg_A[0]), .C(CLK_c), .D(data_i[0]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_DFFSR cnt_reg_2247__i9 (.Q(cnt_reg[9]), .C(CLK_c), .D(n45[9]), 
            .R(cnt_next_9__N_836));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFFSR cnt_reg_2247__i8 (.Q(cnt_reg[8]), .C(CLK_c), .D(n45[8]), 
            .R(cnt_next_9__N_836));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFFSR cnt_reg_2247__i7 (.Q(cnt_reg[7]), .C(CLK_c), .D(n45[7]), 
            .R(cnt_next_9__N_836));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFFSR cnt_reg_2247__i6 (.Q(cnt_reg[6]), .C(CLK_c), .D(n45[6]), 
            .R(cnt_next_9__N_836));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFFSR cnt_reg_2247__i5 (.Q(cnt_reg[5]), .C(CLK_c), .D(n45[5]), 
            .R(cnt_next_9__N_836));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFFSR cnt_reg_2247__i4 (.Q(cnt_reg[4]), .C(CLK_c), .D(n45[4]), 
            .R(cnt_next_9__N_836));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFFSR cnt_reg_2247__i3 (.Q(cnt_reg[3]), .C(CLK_c), .D(n45[3]), 
            .R(cnt_next_9__N_836));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFFSR cnt_reg_2247__i2 (.Q(cnt_reg[2]), .C(CLK_c), .D(n45[2]), 
            .R(cnt_next_9__N_836));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFFSR cnt_reg_2247__i1 (.Q(cnt_reg[1]), .C(CLK_c), .D(n45[1]), 
            .R(cnt_next_9__N_836));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFF reg_out_i0_i0 (.Q(data_o[0]), .C(CLK_c), .D(n29025));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    SB_DFFSR cnt_reg_2247__i0 (.Q(cnt_reg[0]), .C(CLK_c), .D(n45[0]), 
            .R(cnt_next_9__N_836));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_LUT4 i6_4_lut (.I0(cnt_reg[0]), .I1(cnt_reg[1]), .I2(cnt_reg[7]), 
            .I3(cnt_reg[2]), .O(n16));
    defparam i6_4_lut.LUT_INIT = 16'hffef;
    SB_LUT4 i7_4_lut (.I0(cnt_reg[4]), .I1(cnt_reg[9]), .I2(cnt_reg[8]), 
            .I3(cnt_reg[5]), .O(n17));
    defparam i7_4_lut.LUT_INIT = 16'hbfff;
    SB_LUT4 i9_4_lut (.I0(n17), .I1(cnt_reg[6]), .I2(n16), .I3(cnt_reg[3]), 
            .O(n46440));
    defparam i9_4_lut.LUT_INIT = 16'hfbff;
    SB_LUT4 cnt_reg_2247_add_4_11_lut (.I0(GND_net), .I1(GND_net), .I2(cnt_reg[9]), 
            .I3(n39376), .O(n45[9])) /* synthesis syn_instantiated=1 */ ;
    defparam cnt_reg_2247_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 cnt_reg_2247_add_4_10_lut (.I0(GND_net), .I1(GND_net), .I2(cnt_reg[8]), 
            .I3(n39375), .O(n45[8])) /* synthesis syn_instantiated=1 */ ;
    defparam cnt_reg_2247_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY cnt_reg_2247_add_4_10 (.CI(n39375), .I0(GND_net), .I1(cnt_reg[8]), 
            .CO(n39376));
    SB_LUT4 cnt_reg_2247_add_4_9_lut (.I0(GND_net), .I1(GND_net), .I2(cnt_reg[7]), 
            .I3(n39374), .O(n45[7])) /* synthesis syn_instantiated=1 */ ;
    defparam cnt_reg_2247_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY cnt_reg_2247_add_4_9 (.CI(n39374), .I0(GND_net), .I1(cnt_reg[7]), 
            .CO(n39375));
    SB_LUT4 cnt_reg_2247_add_4_8_lut (.I0(GND_net), .I1(GND_net), .I2(cnt_reg[6]), 
            .I3(n39373), .O(n45[6])) /* synthesis syn_instantiated=1 */ ;
    defparam cnt_reg_2247_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY cnt_reg_2247_add_4_8 (.CI(n39373), .I0(GND_net), .I1(cnt_reg[6]), 
            .CO(n39374));
    SB_LUT4 cnt_reg_2247_add_4_7_lut (.I0(GND_net), .I1(GND_net), .I2(cnt_reg[5]), 
            .I3(n39372), .O(n45[5])) /* synthesis syn_instantiated=1 */ ;
    defparam cnt_reg_2247_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY cnt_reg_2247_add_4_7 (.CI(n39372), .I0(GND_net), .I1(cnt_reg[5]), 
            .CO(n39373));
    SB_LUT4 cnt_reg_2247_add_4_6_lut (.I0(GND_net), .I1(GND_net), .I2(cnt_reg[4]), 
            .I3(n39371), .O(n45[4])) /* synthesis syn_instantiated=1 */ ;
    defparam cnt_reg_2247_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY cnt_reg_2247_add_4_6 (.CI(n39371), .I0(GND_net), .I1(cnt_reg[4]), 
            .CO(n39372));
    SB_LUT4 cnt_reg_2247_add_4_5_lut (.I0(GND_net), .I1(GND_net), .I2(cnt_reg[3]), 
            .I3(n39370), .O(n45[3])) /* synthesis syn_instantiated=1 */ ;
    defparam cnt_reg_2247_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY cnt_reg_2247_add_4_5 (.CI(n39370), .I0(GND_net), .I1(cnt_reg[3]), 
            .CO(n39371));
    SB_LUT4 cnt_reg_2247_add_4_4_lut (.I0(GND_net), .I1(GND_net), .I2(cnt_reg[2]), 
            .I3(n39369), .O(n45[2])) /* synthesis syn_instantiated=1 */ ;
    defparam cnt_reg_2247_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY cnt_reg_2247_add_4_4 (.CI(n39369), .I0(GND_net), .I1(cnt_reg[2]), 
            .CO(n39370));
    SB_LUT4 cnt_reg_2247_add_4_3_lut (.I0(GND_net), .I1(GND_net), .I2(cnt_reg[1]), 
            .I3(n39368), .O(n45[1])) /* synthesis syn_instantiated=1 */ ;
    defparam cnt_reg_2247_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY cnt_reg_2247_add_4_3 (.CI(n39368), .I0(GND_net), .I1(cnt_reg[1]), 
            .CO(n39369));
    SB_LUT4 cnt_reg_2247_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(cnt_reg[0]), 
            .I3(VCC_net), .O(n45[0])) /* synthesis syn_instantiated=1 */ ;
    defparam cnt_reg_2247_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY cnt_reg_2247_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(cnt_reg[0]), 
            .CO(n39368));
    SB_DFF reg_A_i2 (.Q(reg_A[2]), .C(CLK_c), .D(data_i[2]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    
endmodule
//
// Verilog Description of module TLI4970
//

module TLI4970 (n29164, \data[8] , n29160, \data[7] , n10, GND_net, 
            n11, n15, \state[1] , \state[0] , n29154, \data[6] , 
            CLK_c, n29152, \data[5] , n29138, \data[4] , n34688, 
            VCC_net, \data[12] , n29103, \data[3] , n29073, \data[2] , 
            n9, clk_out, n29057, CS_c, n29052, \data[1] , n29051, 
            \current[0] , n27177, n28537, \current[15] , \data[15] , 
            n29553, \current[1] , n29552, \current[2] , n29551, \current[3] , 
            n29550, \current[4] , n29549, \current[5] , n29548, \current[6] , 
            n29547, \current[7] , n29546, \current[8] , n29545, \current[9] , 
            n29544, \current[10] , state_7__N_4460, n29543, \current[11] , 
            n27143, n6, n29324, n29323, n29290, \data[11] , n29288, 
            \data[10] , n29238, \data[0] , n29184, \data[9] , n34690, 
            n27167, n27180, n6_adj_14, n27174, CS_CLK_c, n5) /* synthesis syn_noprune=1, syn_module_defined=1 */ ;
    input n29164;
    output \data[8] ;
    input n29160;
    output \data[7] ;
    output n10;
    input GND_net;
    output n11;
    output n15;
    output \state[1] ;
    output \state[0] ;
    input n29154;
    output \data[6] ;
    input CLK_c;
    input n29152;
    output \data[5] ;
    input n29138;
    output \data[4] ;
    output n34688;
    input VCC_net;
    output \data[12] ;
    input n29103;
    output \data[3] ;
    input n29073;
    output \data[2] ;
    input n9;
    output clk_out;
    input n29057;
    output CS_c;
    input n29052;
    output \data[1] ;
    input n29051;
    output \current[0] ;
    output n27177;
    output n28537;
    output \current[15] ;
    output \data[15] ;
    input n29553;
    output \current[1] ;
    input n29552;
    output \current[2] ;
    input n29551;
    output \current[3] ;
    input n29550;
    output \current[4] ;
    input n29549;
    output \current[5] ;
    input n29548;
    output \current[6] ;
    input n29547;
    output \current[7] ;
    input n29546;
    output \current[8] ;
    input n29545;
    output \current[9] ;
    input n29544;
    output \current[10] ;
    output state_7__N_4460;
    input n29543;
    output \current[11] ;
    output n27143;
    output n6;
    input n29324;
    input n29323;
    input n29290;
    output \data[11] ;
    input n29288;
    output \data[10] ;
    input n29238;
    output \data[0] ;
    input n29184;
    output \data[9] ;
    output n34690;
    output n27167;
    output n27180;
    output n6_adj_14;
    output n27174;
    output CS_CLK_c;
    output n5;
    
    wire clk_slow /* synthesis is_clock=1, SET_AS_NETWORK=\tli/clk_slow */ ;   // verilog/tli4970.v(11[7:15])
    wire CLK_c /* synthesis SET_AS_NETWORK=CLK_c, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(3[9:12])
    wire [7:0]bit_counter;   // verilog/tli4970.v(26[13:24])
    
    wire n6_c;
    wire [15:0]delay_counter;   // verilog/tli4970.v(28[14:27])
    
    wire n6_adj_4810, n45207, n45996, n45968, delay_counter_15__N_4455, 
        n10652;
    wire [7:0]n37;
    
    wire n28609, n28867, n28689, n28846, n35257, clk_slow_N_4373;
    wire [4:0]n25;
    wire [7:0]counter;   // verilog/tli4970.v(12[13:20])
    
    wire n39424, n39423, n39422, n39421;
    wire [13:0]n61;
    
    wire n39420, n39419, n39418, n39417, n39416, n39415;
    wire [7:0]n47;
    
    wire clk_slow_N_4374;
    wire [13:0]n241;
    
    wire n39414, n39413, n39412, n39411, n39410, n39409, n39408, 
        n39477, n39476, n39475, n39474, n39473, n39472, n39471, 
        n6_adj_4813;
    
    SB_DFFN data_i8 (.Q(\data[8] ), .C(clk_slow), .D(n29164));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i7 (.Q(\data[7] ), .C(clk_slow), .D(n29160));   // verilog/tli4970.v(35[10] 68[6])
    SB_LUT4 equal_269_i10_2_lut (.I0(bit_counter[2]), .I1(bit_counter[3]), 
            .I2(GND_net), .I3(GND_net), .O(n10));   // verilog/tli4970.v(56[12:26])
    defparam equal_269_i10_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut (.I0(bit_counter[5]), .I1(bit_counter[4]), .I2(GND_net), 
            .I3(GND_net), .O(n6_c));   // verilog/tli4970.v(56[12:26])
    defparam i1_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i4_4_lut (.I0(bit_counter[6]), .I1(bit_counter[7]), .I2(n11), 
            .I3(n6_c), .O(n15));   // verilog/tli4970.v(56[12:26])
    defparam i4_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_2_lut (.I0(delay_counter[5]), .I1(delay_counter[6]), .I2(GND_net), 
            .I3(GND_net), .O(n6_adj_4810));
    defparam i2_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i3_4_lut (.I0(delay_counter[0]), .I1(delay_counter[1]), .I2(delay_counter[3]), 
            .I3(delay_counter[2]), .O(n45207));
    defparam i3_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i3_4_lut_adj_1708 (.I0(n45207), .I1(n6_adj_4810), .I2(delay_counter[7]), 
            .I3(delay_counter[4]), .O(n45996));
    defparam i3_4_lut_adj_1708.LUT_INIT = 16'hfefc;
    SB_LUT4 i3_4_lut_adj_1709 (.I0(n45996), .I1(delay_counter[8]), .I2(delay_counter[10]), 
            .I3(delay_counter[9]), .O(n45968));
    defparam i3_4_lut_adj_1709.LUT_INIT = 16'h8000;
    SB_LUT4 i2360_4_lut (.I0(n45968), .I1(delay_counter[13]), .I2(delay_counter[12]), 
            .I3(delay_counter[11]), .O(delay_counter_15__N_4455));
    defparam i2360_4_lut.LUT_INIT = 16'hccc8;
    SB_LUT4 mux_2351_i2_3_lut (.I0(n15), .I1(\state[1] ), .I2(\state[0] ), 
            .I3(GND_net), .O(n10652));
    defparam mux_2351_i2_3_lut.LUT_INIT = 16'h3535;
    SB_DFFNESR bit_counter_2258__i4 (.Q(bit_counter[4]), .C(clk_slow), .E(n28609), 
            .D(n37[4]), .R(n28867));   // verilog/tli4970.v(55[24:39])
    SB_DFFNESR bit_counter_2258__i5 (.Q(bit_counter[5]), .C(clk_slow), .E(n28609), 
            .D(n37[5]), .R(n28867));   // verilog/tli4970.v(55[24:39])
    SB_DFFNESR bit_counter_2258__i6 (.Q(bit_counter[6]), .C(clk_slow), .E(n28609), 
            .D(n37[6]), .R(n28867));   // verilog/tli4970.v(55[24:39])
    SB_DFFNESR state_i1 (.Q(\state[1] ), .C(clk_slow), .E(n28689), .D(n10652), 
            .R(n28846));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i6 (.Q(\data[6] ), .C(clk_slow), .D(n29154));   // verilog/tli4970.v(35[10] 68[6])
    SB_LUT4 i35019_2_lut (.I0(n15), .I1(\state[0] ), .I2(GND_net), .I3(GND_net), 
            .O(n35257));
    defparam i35019_2_lut.LUT_INIT = 16'h1111;
    SB_DFFNESR bit_counter_2258__i7 (.Q(bit_counter[7]), .C(clk_slow), .E(n28609), 
            .D(n37[7]), .R(n28867));   // verilog/tli4970.v(55[24:39])
    SB_DFF clk_slow_63 (.Q(clk_slow), .C(CLK_c), .D(clk_slow_N_4373));   // verilog/tli4970.v(13[10] 19[6])
    SB_DFFN data_i5 (.Q(\data[5] ), .C(clk_slow), .D(n29152));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i4 (.Q(\data[4] ), .C(clk_slow), .D(n29138));   // verilog/tli4970.v(35[10] 68[6])
    SB_LUT4 i20758_2_lut (.I0(bit_counter[2]), .I1(bit_counter[3]), .I2(GND_net), 
            .I3(GND_net), .O(n34688));
    defparam i20758_2_lut.LUT_INIT = 16'h8888;
    SB_DFFNESS state_i0 (.Q(\state[0] ), .C(clk_slow), .E(n28689), .D(n35257), 
            .S(n28846));   // verilog/tli4970.v(35[10] 68[6])
    SB_LUT4 counter_2251_2252_add_4_6_lut (.I0(GND_net), .I1(GND_net), .I2(counter[4]), 
            .I3(n39424), .O(n25[4])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2251_2252_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 counter_2251_2252_add_4_5_lut (.I0(GND_net), .I1(GND_net), .I2(counter[3]), 
            .I3(n39423), .O(n25[3])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2251_2252_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_2251_2252_add_4_5 (.CI(n39423), .I0(GND_net), .I1(counter[3]), 
            .CO(n39424));
    SB_LUT4 counter_2251_2252_add_4_4_lut (.I0(GND_net), .I1(GND_net), .I2(counter[2]), 
            .I3(n39422), .O(n25[2])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2251_2252_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_2251_2252_add_4_4 (.CI(n39422), .I0(GND_net), .I1(counter[2]), 
            .CO(n39423));
    SB_LUT4 counter_2251_2252_add_4_3_lut (.I0(GND_net), .I1(GND_net), .I2(counter[1]), 
            .I3(n39421), .O(n25[1])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2251_2252_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_2251_2252_add_4_3 (.CI(n39421), .I0(GND_net), .I1(counter[1]), 
            .CO(n39422));
    SB_LUT4 counter_2251_2252_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(counter[0]), 
            .I3(VCC_net), .O(n25[0])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2251_2252_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_2251_2252_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(counter[0]), 
            .CO(n39421));
    SB_LUT4 delay_counter_2249_2250_add_4_15_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[13]), .I3(n39420), .O(n61[13])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_2249_2250_add_4_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 delay_counter_2249_2250_add_4_14_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[12]), .I3(n39419), .O(n61[12])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_2249_2250_add_4_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_2249_2250_add_4_14 (.CI(n39419), .I0(GND_net), 
            .I1(delay_counter[12]), .CO(n39420));
    SB_LUT4 delay_counter_2249_2250_add_4_13_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[11]), .I3(n39418), .O(n61[11])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_2249_2250_add_4_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_2249_2250_add_4_13 (.CI(n39418), .I0(GND_net), 
            .I1(delay_counter[11]), .CO(n39419));
    SB_LUT4 delay_counter_2249_2250_add_4_12_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[10]), .I3(n39417), .O(n61[10])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_2249_2250_add_4_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_2249_2250_add_4_12 (.CI(n39417), .I0(GND_net), 
            .I1(delay_counter[10]), .CO(n39418));
    SB_LUT4 delay_counter_2249_2250_add_4_11_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[9]), .I3(n39416), .O(n61[9])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_2249_2250_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_2249_2250_add_4_11 (.CI(n39416), .I0(GND_net), 
            .I1(delay_counter[9]), .CO(n39417));
    SB_LUT4 delay_counter_2249_2250_add_4_10_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[8]), .I3(n39415), .O(n61[8])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_2249_2250_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_DFFNE bit_counter_2258__i3 (.Q(bit_counter[3]), .C(clk_slow), .E(n28609), 
            .D(n47[3]));   // verilog/tli4970.v(55[24:39])
    SB_DFFNE bit_counter_2258__i2 (.Q(bit_counter[2]), .C(clk_slow), .E(n28609), 
            .D(n47[2]));   // verilog/tli4970.v(55[24:39])
    SB_DFFNE bit_counter_2258__i1 (.Q(bit_counter[1]), .C(clk_slow), .E(n28609), 
            .D(n47[1]));   // verilog/tli4970.v(55[24:39])
    SB_DFFSR counter_2251_2252__i5 (.Q(counter[4]), .C(CLK_c), .D(n25[4]), 
            .R(clk_slow_N_4374));   // verilog/tli4970.v(14[16:27])
    SB_DFFSR counter_2251_2252__i4 (.Q(counter[3]), .C(CLK_c), .D(n25[3]), 
            .R(clk_slow_N_4374));   // verilog/tli4970.v(14[16:27])
    SB_DFFSR counter_2251_2252__i3 (.Q(counter[2]), .C(CLK_c), .D(n25[2]), 
            .R(clk_slow_N_4374));   // verilog/tli4970.v(14[16:27])
    SB_DFFSR counter_2251_2252__i2 (.Q(counter[1]), .C(CLK_c), .D(n25[1]), 
            .R(clk_slow_N_4374));   // verilog/tli4970.v(14[16:27])
    SB_DFFNSR delay_counter_2249_2250__i14 (.Q(delay_counter[13]), .C(clk_slow), 
            .D(n61[13]), .R(delay_counter_15__N_4455));   // verilog/tli4970.v(40[24:39])
    SB_DFFNSR delay_counter_2249_2250__i13 (.Q(delay_counter[12]), .C(clk_slow), 
            .D(n61[12]), .R(delay_counter_15__N_4455));   // verilog/tli4970.v(40[24:39])
    SB_DFFNSR delay_counter_2249_2250__i12 (.Q(delay_counter[11]), .C(clk_slow), 
            .D(n61[11]), .R(delay_counter_15__N_4455));   // verilog/tli4970.v(40[24:39])
    SB_DFFNSR delay_counter_2249_2250__i11 (.Q(delay_counter[10]), .C(clk_slow), 
            .D(n61[10]), .R(delay_counter_15__N_4455));   // verilog/tli4970.v(40[24:39])
    SB_DFFNSR delay_counter_2249_2250__i10 (.Q(delay_counter[9]), .C(clk_slow), 
            .D(n61[9]), .R(delay_counter_15__N_4455));   // verilog/tli4970.v(40[24:39])
    SB_DFFNSR delay_counter_2249_2250__i9 (.Q(delay_counter[8]), .C(clk_slow), 
            .D(n61[8]), .R(delay_counter_15__N_4455));   // verilog/tli4970.v(40[24:39])
    SB_DFFNSR delay_counter_2249_2250__i8 (.Q(delay_counter[7]), .C(clk_slow), 
            .D(n61[7]), .R(delay_counter_15__N_4455));   // verilog/tli4970.v(40[24:39])
    SB_DFFNSR delay_counter_2249_2250__i7 (.Q(delay_counter[6]), .C(clk_slow), 
            .D(n61[6]), .R(delay_counter_15__N_4455));   // verilog/tli4970.v(40[24:39])
    SB_DFFNSR delay_counter_2249_2250__i6 (.Q(delay_counter[5]), .C(clk_slow), 
            .D(n61[5]), .R(delay_counter_15__N_4455));   // verilog/tli4970.v(40[24:39])
    SB_DFFNSR delay_counter_2249_2250__i5 (.Q(delay_counter[4]), .C(clk_slow), 
            .D(n61[4]), .R(delay_counter_15__N_4455));   // verilog/tli4970.v(40[24:39])
    SB_DFFNSR delay_counter_2249_2250__i4 (.Q(delay_counter[3]), .C(clk_slow), 
            .D(n61[3]), .R(delay_counter_15__N_4455));   // verilog/tli4970.v(40[24:39])
    SB_DFFNSR delay_counter_2249_2250__i3 (.Q(delay_counter[2]), .C(clk_slow), 
            .D(n61[2]), .R(delay_counter_15__N_4455));   // verilog/tli4970.v(40[24:39])
    SB_DFFNSR delay_counter_2249_2250__i2 (.Q(delay_counter[1]), .C(clk_slow), 
            .D(n61[1]), .R(delay_counter_15__N_4455));   // verilog/tli4970.v(40[24:39])
    SB_LUT4 i2383_1_lut (.I0(\data[12] ), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n241[13]));
    defparam i2383_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY delay_counter_2249_2250_add_4_10 (.CI(n39415), .I0(GND_net), 
            .I1(delay_counter[8]), .CO(n39416));
    SB_LUT4 delay_counter_2249_2250_add_4_9_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[7]), .I3(n39414), .O(n61[7])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_2249_2250_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_2249_2250_add_4_9 (.CI(n39414), .I0(GND_net), 
            .I1(delay_counter[7]), .CO(n39415));
    SB_LUT4 delay_counter_2249_2250_add_4_8_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[6]), .I3(n39413), .O(n61[6])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_2249_2250_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_2249_2250_add_4_8 (.CI(n39413), .I0(GND_net), 
            .I1(delay_counter[6]), .CO(n39414));
    SB_LUT4 delay_counter_2249_2250_add_4_7_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[5]), .I3(n39412), .O(n61[5])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_2249_2250_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_2249_2250_add_4_7 (.CI(n39412), .I0(GND_net), 
            .I1(delay_counter[5]), .CO(n39413));
    SB_LUT4 i14819_2_lut (.I0(\state[1] ), .I1(\state[0] ), .I2(GND_net), 
            .I3(GND_net), .O(n28609));
    defparam i14819_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 delay_counter_2249_2250_add_4_6_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[4]), .I3(n39411), .O(n61[4])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_2249_2250_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_2249_2250_add_4_6 (.CI(n39411), .I0(GND_net), 
            .I1(delay_counter[4]), .CO(n39412));
    SB_LUT4 delay_counter_2249_2250_add_4_5_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[3]), .I3(n39410), .O(n61[3])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_2249_2250_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_2249_2250_add_4_5 (.CI(n39410), .I0(GND_net), 
            .I1(delay_counter[3]), .CO(n39411));
    SB_LUT4 delay_counter_2249_2250_add_4_4_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[2]), .I3(n39409), .O(n61[2])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_2249_2250_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_2249_2250_add_4_4 (.CI(n39409), .I0(GND_net), 
            .I1(delay_counter[2]), .CO(n39410));
    SB_LUT4 delay_counter_2249_2250_add_4_3_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[1]), .I3(n39408), .O(n61[1])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_2249_2250_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_2249_2250_add_4_3 (.CI(n39408), .I0(GND_net), 
            .I1(delay_counter[1]), .CO(n39409));
    SB_LUT4 delay_counter_2249_2250_add_4_2_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[0]), .I3(VCC_net), .O(n61[0])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_2249_2250_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_2249_2250_add_4_2 (.CI(VCC_net), .I0(GND_net), 
            .I1(delay_counter[0]), .CO(n39408));
    SB_DFFN data_i3 (.Q(\data[3] ), .C(clk_slow), .D(n29103));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i2 (.Q(\data[2] ), .C(clk_slow), .D(n29073));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN clk_out_67 (.Q(clk_out), .C(clk_slow), .D(n9));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN slave_select_66 (.Q(CS_c), .C(clk_slow), .D(n29057));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i1 (.Q(\data[1] ), .C(clk_slow), .D(n29052));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i1 (.Q(\current[0] ), .C(clk_slow), .D(n29051));   // verilog/tli4970.v(35[10] 68[6])
    SB_LUT4 i1_2_lut_4_lut (.I0(\state[0] ), .I1(\state[1] ), .I2(bit_counter[0]), 
            .I3(bit_counter[1]), .O(n27177));   // verilog/tli4970.v(43[5] 67[12])
    defparam i1_2_lut_4_lut.LUT_INIT = 16'hfbff;
    SB_DFFNSR delay_counter_2249_2250__i1 (.Q(delay_counter[0]), .C(clk_slow), 
            .D(n61[0]), .R(delay_counter_15__N_4455));   // verilog/tli4970.v(40[24:39])
    SB_DFFSR counter_2251_2252__i1 (.Q(counter[0]), .C(CLK_c), .D(n25[0]), 
            .R(clk_slow_N_4374));   // verilog/tli4970.v(14[16:27])
    SB_DFFNE bit_counter_2258__i0 (.Q(bit_counter[0]), .C(clk_slow), .E(n28609), 
            .D(n47[0]));   // verilog/tli4970.v(55[24:39])
    SB_DFFNE current__i13 (.Q(\current[15] ), .C(clk_slow), .E(n28537), 
            .D(n241[13]));   // verilog/tli4970.v(35[10] 68[6])
    SB_LUT4 i34912_3_lut (.I0(\data[15] ), .I1(\state[1] ), .I2(\state[0] ), 
            .I3(GND_net), .O(n28537));
    defparam i34912_3_lut.LUT_INIT = 16'h4040;
    SB_DFFN current__i2 (.Q(\current[1] ), .C(clk_slow), .D(n29553));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i3 (.Q(\current[2] ), .C(clk_slow), .D(n29552));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i4 (.Q(\current[3] ), .C(clk_slow), .D(n29551));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i5 (.Q(\current[4] ), .C(clk_slow), .D(n29550));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i6 (.Q(\current[5] ), .C(clk_slow), .D(n29549));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i7 (.Q(\current[6] ), .C(clk_slow), .D(n29548));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i8 (.Q(\current[7] ), .C(clk_slow), .D(n29547));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i9 (.Q(\current[8] ), .C(clk_slow), .D(n29546));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i10 (.Q(\current[9] ), .C(clk_slow), .D(n29545));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i11 (.Q(\current[10] ), .C(clk_slow), .D(n29544));   // verilog/tli4970.v(35[10] 68[6])
    SB_LUT4 state_7__I_0_77_i9_2_lut (.I0(\state[0] ), .I1(\state[1] ), 
            .I2(GND_net), .I3(GND_net), .O(state_7__N_4460));   // verilog/tli4970.v(53[7:17])
    defparam state_7__I_0_77_i9_2_lut.LUT_INIT = 16'hbbbb;
    SB_DFFN current__i12 (.Q(\current[11] ), .C(clk_slow), .D(n29543));   // verilog/tli4970.v(35[10] 68[6])
    SB_LUT4 equal_269_i11_2_lut_3_lut_4_lut (.I0(bit_counter[0]), .I1(bit_counter[1]), 
            .I2(bit_counter[2]), .I3(bit_counter[3]), .O(n11));   // verilog/tli4970.v(56[12:26])
    defparam equal_269_i11_2_lut_3_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 bit_counter_2258_add_4_9_lut (.I0(GND_net), .I1(VCC_net), .I2(bit_counter[7]), 
            .I3(n39477), .O(n37[7])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_counter_2258_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 bit_counter_2258_add_4_8_lut (.I0(GND_net), .I1(VCC_net), .I2(bit_counter[6]), 
            .I3(n39476), .O(n37[6])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_counter_2258_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY bit_counter_2258_add_4_8 (.CI(n39476), .I0(VCC_net), .I1(bit_counter[6]), 
            .CO(n39477));
    SB_LUT4 bit_counter_2258_add_4_7_lut (.I0(GND_net), .I1(VCC_net), .I2(bit_counter[5]), 
            .I3(n39475), .O(n37[5])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_counter_2258_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY bit_counter_2258_add_4_7 (.CI(n39475), .I0(VCC_net), .I1(bit_counter[5]), 
            .CO(n39476));
    SB_LUT4 bit_counter_2258_add_4_6_lut (.I0(GND_net), .I1(VCC_net), .I2(bit_counter[4]), 
            .I3(n39474), .O(n37[4])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_counter_2258_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY bit_counter_2258_add_4_6 (.CI(n39474), .I0(VCC_net), .I1(bit_counter[4]), 
            .CO(n39475));
    SB_LUT4 bit_counter_2258_mux_6_i1_3_lut_4_lut (.I0(\state[1] ), .I1(\state[0] ), 
            .I2(state_7__N_4460), .I3(n37[0]), .O(n47[0]));
    defparam bit_counter_2258_mux_6_i1_3_lut_4_lut.LUT_INIT = 16'h4f40;
    SB_LUT4 bit_counter_2258_add_4_5_lut (.I0(GND_net), .I1(VCC_net), .I2(bit_counter[3]), 
            .I3(n39473), .O(n37[3])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_counter_2258_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY bit_counter_2258_add_4_5 (.CI(n39473), .I0(VCC_net), .I1(bit_counter[3]), 
            .CO(n39474));
    SB_LUT4 bit_counter_2258_mux_6_i2_3_lut_4_lut (.I0(\state[1] ), .I1(\state[0] ), 
            .I2(state_7__N_4460), .I3(n37[1]), .O(n47[1]));
    defparam bit_counter_2258_mux_6_i2_3_lut_4_lut.LUT_INIT = 16'h4f40;
    SB_LUT4 bit_counter_2258_add_4_4_lut (.I0(GND_net), .I1(VCC_net), .I2(bit_counter[2]), 
            .I3(n39472), .O(n37[2])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_counter_2258_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY bit_counter_2258_add_4_4 (.CI(n39472), .I0(VCC_net), .I1(bit_counter[2]), 
            .CO(n39473));
    SB_LUT4 bit_counter_2258_add_4_3_lut (.I0(GND_net), .I1(VCC_net), .I2(bit_counter[1]), 
            .I3(n39471), .O(n37[1])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_counter_2258_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY bit_counter_2258_add_4_3 (.CI(n39471), .I0(VCC_net), .I1(bit_counter[1]), 
            .CO(n39472));
    SB_LUT4 bit_counter_2258_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(bit_counter[0]), 
            .I3(VCC_net), .O(n37[0])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_counter_2258_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY bit_counter_2258_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(bit_counter[0]), 
            .CO(n39471));
    SB_LUT4 i1_2_lut_3_lut_4_lut (.I0(bit_counter[0]), .I1(bit_counter[1]), 
            .I2(\state[0] ), .I3(\state[1] ), .O(n27143));   // verilog/tli4970.v(56[12:26])
    defparam i1_2_lut_3_lut_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 bit_counter_2258_mux_6_i3_3_lut_4_lut (.I0(\state[1] ), .I1(\state[0] ), 
            .I2(state_7__N_4460), .I3(n37[2]), .O(n47[2]));
    defparam bit_counter_2258_mux_6_i3_3_lut_4_lut.LUT_INIT = 16'h4f40;
    SB_LUT4 bit_counter_2258_mux_6_i4_3_lut_4_lut (.I0(\state[1] ), .I1(\state[0] ), 
            .I2(state_7__N_4460), .I3(n37[3]), .O(n47[3]));
    defparam bit_counter_2258_mux_6_i4_3_lut_4_lut.LUT_INIT = 16'h4f40;
    SB_LUT4 equal_329_i6_2_lut (.I0(bit_counter[2]), .I1(bit_counter[3]), 
            .I2(GND_net), .I3(GND_net), .O(n6));   // verilog/tli4970.v(54[9:26])
    defparam equal_329_i6_2_lut.LUT_INIT = 16'hbbbb;
    SB_DFFN data_i15 (.Q(\data[15] ), .C(clk_slow), .D(n29324));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i12 (.Q(\data[12] ), .C(clk_slow), .D(n29323));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i11 (.Q(\data[11] ), .C(clk_slow), .D(n29290));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i10 (.Q(\data[10] ), .C(clk_slow), .D(n29288));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i0 (.Q(\data[0] ), .C(clk_slow), .D(n29238));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i9 (.Q(\data[9] ), .C(clk_slow), .D(n29184));   // verilog/tli4970.v(35[10] 68[6])
    SB_LUT4 i20760_2_lut (.I0(bit_counter[0]), .I1(bit_counter[1]), .I2(GND_net), 
            .I3(GND_net), .O(n34690));
    defparam i20760_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_3_lut_4_lut (.I0(bit_counter[0]), .I1(bit_counter[1]), .I2(\state[0] ), 
            .I3(\state[1] ), .O(n27167));   // verilog/tli4970.v(43[5] 67[12])
    defparam i2_3_lut_4_lut.LUT_INIT = 16'hfdff;
    SB_LUT4 i1_2_lut_4_lut_adj_1710 (.I0(\state[0] ), .I1(\state[1] ), .I2(bit_counter[0]), 
            .I3(bit_counter[1]), .O(n27180));   // verilog/tli4970.v(43[5] 67[12])
    defparam i1_2_lut_4_lut_adj_1710.LUT_INIT = 16'hbfff;
    SB_LUT4 equal_333_i6_2_lut (.I0(bit_counter[2]), .I1(bit_counter[3]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_14));   // verilog/tli4970.v(54[9:26])
    defparam equal_333_i6_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 i14920_2_lut_2_lut (.I0(\state[1] ), .I1(\state[0] ), .I2(GND_net), 
            .I3(GND_net), .O(n28867));   // verilog/tli4970.v(55[24:39])
    defparam i14920_2_lut_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i2_2_lut_adj_1711 (.I0(counter[1]), .I1(counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n6_adj_4813));
    defparam i2_2_lut_adj_1711.LUT_INIT = 16'heeee;
    SB_LUT4 i2355_4_lut (.I0(counter[0]), .I1(counter[4]), .I2(n6_adj_4813), 
            .I3(counter[3]), .O(clk_slow_N_4374));
    defparam i2355_4_lut.LUT_INIT = 16'hccc8;
    SB_LUT4 clk_slow_I_0_72_2_lut (.I0(clk_slow), .I1(clk_slow_N_4374), 
            .I2(GND_net), .I3(GND_net), .O(clk_slow_N_4373));   // verilog/tli4970.v(15[5] 18[8])
    defparam clk_slow_I_0_72_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_4_lut_adj_1712 (.I0(\state[0] ), .I1(\state[1] ), .I2(bit_counter[2]), 
            .I3(bit_counter[3]), .O(n27174));   // verilog/tli4970.v(43[5] 67[12])
    defparam i1_2_lut_4_lut_adj_1712.LUT_INIT = 16'hfbff;
    SB_LUT4 i1_2_lut_4_lut_adj_1713 (.I0(n15), .I1(\state[1] ), .I2(\state[0] ), 
            .I3(delay_counter_15__N_4455), .O(n28689));
    defparam i1_2_lut_4_lut_adj_1713.LUT_INIT = 16'hfff4;
    SB_LUT4 i14898_2_lut_4_lut (.I0(n15), .I1(\state[1] ), .I2(\state[0] ), 
            .I3(delay_counter_15__N_4455), .O(n28846));
    defparam i14898_2_lut_4_lut.LUT_INIT = 16'h0b00;
    SB_LUT4 spi_clk_I_0_i1_3_lut (.I0(clk_slow), .I1(clk_out), .I2(CS_c), 
            .I3(GND_net), .O(CS_CLK_c));   // verilog/tli4970.v(23[20:53])
    defparam spi_clk_I_0_i1_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 equal_326_i5_2_lut (.I0(bit_counter[0]), .I1(bit_counter[1]), 
            .I2(GND_net), .I3(GND_net), .O(n5));   // verilog/tli4970.v(54[9:26])
    defparam equal_326_i5_2_lut.LUT_INIT = 16'hbbbb;
    
endmodule
//
// Verilog Description of module coms
//

module coms (\data_out_frame[13] , GND_net, \data_out_frame[20] , \data_out_frame[23] , 
            CLK_c, \data_in_frame[3] , \data_out_frame[25] , \data_in_frame[5] , 
            rx_data, \data_out_frame[10] , \data_out_frame[6] , \data_out_frame[8] , 
            \data_out_frame[17] , \data_out_frame[15] , \data_out_frame[16] , 
            \data_out_frame[19] , \data_out_frame[21] , \data_out_frame[12] , 
            \data_out_frame[14] , \data_out_frame[5] , \data_out_frame[4] , 
            \data_in_frame[11] , \data_in_frame[14] , \data_in_frame[13] , 
            \data_out_frame[11] , \data_out_frame[9] , \data_out_frame[7] , 
            \data_in_frame[10] , \data_in_frame[12] , \data_out_frame[18] , 
            \data_out_frame[22] , \data_in_frame[1] , n29158, IntegralLimit, 
            \data_in[1] , \data_in[3] , \data_in[0] , \data_in_frame[21] , 
            n29157, n29156, n29155, \data_in_frame[2] , \data_in_frame[20] , 
            \data_in_frame[9] , \data_in_frame[4] , rx_data_ready, setpoint, 
            \data_in_frame[6] , n29153, n29151, n29018, n29150, n29149, 
            n29148, n29147, n29145, n29144, n29143, n29142, n29141, 
            n29140, n29139, n29137, n29136, n29135, n29134, n29133, 
            n29132, n29131, n29130, n29129, ID, n29128, n29127, 
            \data_in_frame[8] , \data_out_frame[24] , n29126, n29125, 
            \data_in_frame[22] , n29124, n29123, n29122, n29121, n29120, 
            n29119, n29118, n29117, n29116, n29115, n29114, n29113, 
            n29112, n29111, n29110, n29109, n29108, n29107, n28521, 
            n29106, n29105, \data_in[2] , n29679, n29678, n29677, 
            n29676, n29675, n29674, n29673, n29672, n29671, n29670, 
            n29669, n29668, n29667, n29666, n29665, n29664, n29663, 
            n29662, n29661, n29660, n29659, n29658, n29657, n29656, 
            n29655, n29654, n29653, n29652, n29651, n29650, n29649, 
            n29648, n29647, n29646, n29645, n29644, n29643, n29642, 
            n29641, n29640, n29639, n29638, n29637, n29636, n29635, 
            n29634, n29633, n29632, n29631, n29630, n29629, n29628, 
            n29104, n29102, n29101, n29100, n29099, n29098, n29097, 
            n29096, n29095, n29094, n29093, n29092, n29091, n29090, 
            n29089, n29088, n29087, n29086, n29085, n29084, n29083, 
            n29082, n29081, n29080, n29079, n29078, n29077, n29076, 
            n29075, n29074, DE_c, n29067, n29065, n29064, n29063, 
            n29062, n29061, n29060, n29056, n29627, LED_c, n29626, 
            n29625, n29624, n29623, n29622, n29621, n29620, n29619, 
            n29618, n29617, n29616, n29615, n29614, n29613, n29612, 
            n29611, n29610, n29609, n29608, n29607, n29606, n29605, 
            n29604, n29602, n29599, control_mode, n29598, n29597, 
            n29596, n29595, n29055, n29050, n29049, n29047, PWMLimit, 
            n29046, current_limit, n29045, n29043, neopxl_color, n29042, 
            \Ki[0] , n29041, \Kp[0] , n29040, n29026, n29594, n29593, 
            n29592, n29591, n29590, n29024, n29589, n29023, n29588, 
            n29587, n29586, n29585, n29584, n29583, n29582, n29581, 
            n29580, n29579, n29578, n29577, n29576, n29575, n29574, 
            n29573, n43838, n29572, n29571, n29570, n29569, n29568, 
            n43847, n43822, n29567, n29566, n29021, n29565, n29564, 
            n29563, n29562, n29561, n29560, n29559, n29558, n29557, 
            n29556, n29555, n24278, n29020, n29542, n29541, n29540, 
            n29539, n29538, n29537, n29529, n29528, n29527, n29526, 
            n29525, n29523, n29522, n29521, n29520, n29519, n29518, 
            n29517, n29506, n29505, n29504, n29503, n29501, n29500, 
            n29499, n29466, n29465, n29464, n29463, n29462, n29461, 
            n29460, n29459, n29458, n29457, n29456, n29455, n29454, 
            n29453, n29452, n29451, n29450, n29449, n29448, n29447, 
            n29446, n29445, n29444, n28522, n29403, n29402, n29401, 
            n29400, n29399, n29398, n29397, n29396, n29395, n29394, 
            n29393, n29392, n29391, n29390, n29389, n29388, n29339, 
            n29338, n29336, n29335, n29334, n29333, n29332, n29331, 
            n29330, n29329, n29328, n29327, n29326, n29325, n29322, 
            n29321, n29270, n29269, n29268, n29267, n29266, n29265, 
            n29264, n29263, n29262, n29261, n29260, n29259, n29258, 
            n29257, n29256, n29255, n29244, n29243, n29242, n29241, 
            n29240, n29239, n29225, n29224, n29223, n29221, n29220, 
            n29219, n29218, n29217, n29216, n29215, n29214, n29213, 
            n29212, n29211, n29210, n29209, n29208, n29207, n29206, 
            n29205, n29204, n29203, n29202, n29201, n29200, n29199, 
            \Kp[1] , n29198, \Kp[2] , n29197, \Kp[3] , n29196, \Kp[4] , 
            n29195, \Kp[5] , n29194, \Kp[6] , n29193, \Kp[7] , n29192, 
            \Kp[8] , n29191, \Kp[9] , n29190, \Kp[10] , n29189, 
            \Kp[11] , n29188, \Kp[12] , n29187, \Kp[13] , n29183, 
            \Kp[14] , n29182, \Kp[15] , n29181, \Ki[1] , n29180, 
            \Ki[2] , n29179, \Ki[3] , n29178, \Ki[4] , n29177, \Ki[5] , 
            n29176, \Ki[6] , n29175, \Ki[7] , n29174, \Ki[8] , n29173, 
            \Ki[9] , n29172, \Ki[10] , n29171, \Ki[11] , n29019, 
            n29170, \Ki[12] , n29169, \Ki[13] , n29168, \Ki[14] , 
            n29167, \Ki[15] , \state[0] , \state[2] , \state[3] , 
            n7754, n43824, n43848, n43839, tx_active, \r_Bit_Index[0] , 
            tx_o, r_SM_Main, VCC_net, \r_SM_Main_2__N_3777[1] , n29230, 
            n51602, n29066, n28662, n28970, n19541, n4, tx_enable, 
            \r_SM_Main_2__N_3706[2] , n4_adj_6, r_SM_Main_adj_13, r_Rx_Data, 
            RX_N_10, \r_Bit_Index[0]_adj_10 , n4_adj_11, n4_adj_12, 
            n34695, n29233, n43326, n28666, n28972, n28562, n29524, 
            n29516, n29510, n29508, n29502, n29467, n29404, n43724, 
            n29237, n27131, n27126) /* synthesis syn_module_defined=1 */ ;
    output [7:0]\data_out_frame[13] ;
    input GND_net;
    output [7:0]\data_out_frame[20] ;
    output [7:0]\data_out_frame[23] ;
    input CLK_c;
    output [7:0]\data_in_frame[3] ;
    output [7:0]\data_out_frame[25] ;
    output [7:0]\data_in_frame[5] ;
    output [7:0]rx_data;
    output [7:0]\data_out_frame[10] ;
    output [7:0]\data_out_frame[6] ;
    output [7:0]\data_out_frame[8] ;
    output [7:0]\data_out_frame[17] ;
    output [7:0]\data_out_frame[15] ;
    output [7:0]\data_out_frame[16] ;
    output [7:0]\data_out_frame[19] ;
    output [7:0]\data_out_frame[21] ;
    output [7:0]\data_out_frame[12] ;
    output [7:0]\data_out_frame[14] ;
    output [7:0]\data_out_frame[5] ;
    output [7:0]\data_out_frame[4] ;
    output [7:0]\data_in_frame[11] ;
    output [7:0]\data_in_frame[14] ;
    output [7:0]\data_in_frame[13] ;
    output [7:0]\data_out_frame[11] ;
    output [7:0]\data_out_frame[9] ;
    output [7:0]\data_out_frame[7] ;
    output [7:0]\data_in_frame[10] ;
    output [7:0]\data_in_frame[12] ;
    output [7:0]\data_out_frame[18] ;
    output [7:0]\data_out_frame[22] ;
    output [7:0]\data_in_frame[1] ;
    input n29158;
    output [23:0]IntegralLimit;
    output [7:0]\data_in[1] ;
    output [7:0]\data_in[3] ;
    output [7:0]\data_in[0] ;
    output [7:0]\data_in_frame[21] ;
    input n29157;
    input n29156;
    input n29155;
    output [7:0]\data_in_frame[2] ;
    output [7:0]\data_in_frame[20] ;
    output [7:0]\data_in_frame[9] ;
    output [7:0]\data_in_frame[4] ;
    output rx_data_ready;
    output [23:0]setpoint;
    output [7:0]\data_in_frame[6] ;
    input n29153;
    input n29151;
    input n29018;
    input n29150;
    input n29149;
    input n29148;
    input n29147;
    input n29145;
    input n29144;
    input n29143;
    input n29142;
    input n29141;
    input n29140;
    input n29139;
    input n29137;
    input n29136;
    input n29135;
    input n29134;
    input n29133;
    input n29132;
    input n29131;
    input n29130;
    input n29129;
    input [7:0]ID;
    input n29128;
    input n29127;
    output [7:0]\data_in_frame[8] ;
    output [7:0]\data_out_frame[24] ;
    input n29126;
    input n29125;
    output [7:0]\data_in_frame[22] ;
    input n29124;
    input n29123;
    input n29122;
    input n29121;
    input n29120;
    input n29119;
    input n29118;
    input n29117;
    input n29116;
    input n29115;
    input n29114;
    input n29113;
    input n29112;
    input n29111;
    input n29110;
    input n29109;
    input n29108;
    input n29107;
    output n28521;
    input n29106;
    input n29105;
    output [7:0]\data_in[2] ;
    input n29679;
    input n29678;
    input n29677;
    input n29676;
    input n29675;
    input n29674;
    input n29673;
    input n29672;
    input n29671;
    input n29670;
    input n29669;
    input n29668;
    input n29667;
    input n29666;
    input n29665;
    input n29664;
    input n29663;
    input n29662;
    input n29661;
    input n29660;
    input n29659;
    input n29658;
    input n29657;
    input n29656;
    input n29655;
    input n29654;
    input n29653;
    input n29652;
    input n29651;
    input n29650;
    input n29649;
    input n29648;
    input n29647;
    input n29646;
    input n29645;
    input n29644;
    input n29643;
    input n29642;
    input n29641;
    input n29640;
    input n29639;
    input n29638;
    input n29637;
    input n29636;
    input n29635;
    input n29634;
    input n29633;
    input n29632;
    input n29631;
    input n29630;
    input n29629;
    input n29628;
    input n29104;
    input n29102;
    input n29101;
    input n29100;
    input n29099;
    input n29098;
    input n29097;
    input n29096;
    input n29095;
    input n29094;
    input n29093;
    input n29092;
    input n29091;
    input n29090;
    input n29089;
    input n29088;
    input n29087;
    input n29086;
    input n29085;
    input n29084;
    input n29083;
    input n29082;
    input n29081;
    input n29080;
    input n29079;
    input n29078;
    input n29077;
    input n29076;
    input n29075;
    input n29074;
    output DE_c;
    input n29067;
    input n29065;
    input n29064;
    input n29063;
    input n29062;
    input n29061;
    input n29060;
    input n29056;
    input n29627;
    output LED_c;
    input n29626;
    input n29625;
    input n29624;
    input n29623;
    input n29622;
    input n29621;
    input n29620;
    input n29619;
    input n29618;
    input n29617;
    input n29616;
    input n29615;
    input n29614;
    input n29613;
    input n29612;
    input n29611;
    input n29610;
    input n29609;
    input n29608;
    input n29607;
    input n29606;
    input n29605;
    input n29604;
    input n29602;
    input n29599;
    output [7:0]control_mode;
    input n29598;
    input n29597;
    input n29596;
    input n29595;
    input n29055;
    input n29050;
    input n29049;
    input n29047;
    output [23:0]PWMLimit;
    input n29046;
    output [15:0]current_limit;
    input n29045;
    input n29043;
    output [23:0]neopxl_color;
    input n29042;
    output \Ki[0] ;
    input n29041;
    output \Kp[0] ;
    input n29040;
    input n29026;
    input n29594;
    input n29593;
    input n29592;
    input n29591;
    input n29590;
    input n29024;
    input n29589;
    input n29023;
    input n29588;
    input n29587;
    input n29586;
    input n29585;
    input n29584;
    input n29583;
    input n29582;
    input n29581;
    input n29580;
    input n29579;
    input n29578;
    input n29577;
    input n29576;
    input n29575;
    input n29574;
    input n29573;
    output n43838;
    input n29572;
    input n29571;
    input n29570;
    input n29569;
    input n29568;
    output n43847;
    output n43822;
    input n29567;
    input n29566;
    input n29021;
    input n29565;
    input n29564;
    input n29563;
    input n29562;
    input n29561;
    input n29560;
    input n29559;
    input n29558;
    input n29557;
    input n29556;
    input n29555;
    output n24278;
    input n29020;
    input n29542;
    input n29541;
    input n29540;
    input n29539;
    input n29538;
    input n29537;
    input n29529;
    input n29528;
    input n29527;
    input n29526;
    input n29525;
    input n29523;
    input n29522;
    input n29521;
    input n29520;
    input n29519;
    input n29518;
    input n29517;
    input n29506;
    input n29505;
    input n29504;
    input n29503;
    input n29501;
    input n29500;
    input n29499;
    input n29466;
    input n29465;
    input n29464;
    input n29463;
    input n29462;
    input n29461;
    input n29460;
    input n29459;
    input n29458;
    input n29457;
    input n29456;
    input n29455;
    input n29454;
    input n29453;
    input n29452;
    input n29451;
    input n29450;
    input n29449;
    input n29448;
    input n29447;
    input n29446;
    input n29445;
    input n29444;
    output n28522;
    input n29403;
    input n29402;
    input n29401;
    input n29400;
    input n29399;
    input n29398;
    input n29397;
    input n29396;
    input n29395;
    input n29394;
    input n29393;
    input n29392;
    input n29391;
    input n29390;
    input n29389;
    input n29388;
    input n29339;
    input n29338;
    input n29336;
    input n29335;
    input n29334;
    input n29333;
    input n29332;
    input n29331;
    input n29330;
    input n29329;
    input n29328;
    input n29327;
    input n29326;
    input n29325;
    input n29322;
    input n29321;
    input n29270;
    input n29269;
    input n29268;
    input n29267;
    input n29266;
    input n29265;
    input n29264;
    input n29263;
    input n29262;
    input n29261;
    input n29260;
    input n29259;
    input n29258;
    input n29257;
    input n29256;
    input n29255;
    input n29244;
    input n29243;
    input n29242;
    input n29241;
    input n29240;
    input n29239;
    input n29225;
    input n29224;
    input n29223;
    input n29221;
    input n29220;
    input n29219;
    input n29218;
    input n29217;
    input n29216;
    input n29215;
    input n29214;
    input n29213;
    input n29212;
    input n29211;
    input n29210;
    input n29209;
    input n29208;
    input n29207;
    input n29206;
    input n29205;
    input n29204;
    input n29203;
    input n29202;
    input n29201;
    input n29200;
    input n29199;
    output \Kp[1] ;
    input n29198;
    output \Kp[2] ;
    input n29197;
    output \Kp[3] ;
    input n29196;
    output \Kp[4] ;
    input n29195;
    output \Kp[5] ;
    input n29194;
    output \Kp[6] ;
    input n29193;
    output \Kp[7] ;
    input n29192;
    output \Kp[8] ;
    input n29191;
    output \Kp[9] ;
    input n29190;
    output \Kp[10] ;
    input n29189;
    output \Kp[11] ;
    input n29188;
    output \Kp[12] ;
    input n29187;
    output \Kp[13] ;
    input n29183;
    output \Kp[14] ;
    input n29182;
    output \Kp[15] ;
    input n29181;
    output \Ki[1] ;
    input n29180;
    output \Ki[2] ;
    input n29179;
    output \Ki[3] ;
    input n29178;
    output \Ki[4] ;
    input n29177;
    output \Ki[5] ;
    input n29176;
    output \Ki[6] ;
    input n29175;
    output \Ki[7] ;
    input n29174;
    output \Ki[8] ;
    input n29173;
    output \Ki[9] ;
    input n29172;
    output \Ki[10] ;
    input n29171;
    output \Ki[11] ;
    input n29019;
    input n29170;
    output \Ki[12] ;
    input n29169;
    output \Ki[13] ;
    input n29168;
    output \Ki[14] ;
    input n29167;
    output \Ki[15] ;
    input \state[0] ;
    input \state[2] ;
    input \state[3] ;
    output n7754;
    output n43824;
    output n43848;
    output n43839;
    output tx_active;
    output \r_Bit_Index[0] ;
    output tx_o;
    output [2:0]r_SM_Main;
    input VCC_net;
    output \r_SM_Main_2__N_3777[1] ;
    input n29230;
    input n51602;
    input n29066;
    output n28662;
    output n28970;
    output n19541;
    output n4;
    output tx_enable;
    output \r_SM_Main_2__N_3706[2] ;
    output n4_adj_6;
    output [2:0]r_SM_Main_adj_13;
    output r_Rx_Data;
    input RX_N_10;
    output \r_Bit_Index[0]_adj_10 ;
    output n4_adj_11;
    output n4_adj_12;
    output n34695;
    input n29233;
    input n43326;
    output n28666;
    output n28972;
    output n28562;
    input n29524;
    input n29516;
    input n29510;
    input n29508;
    input n29502;
    input n29467;
    input n29404;
    input n43724;
    input n29237;
    output n27131;
    output n27126;
    
    wire CLK_c /* synthesis SET_AS_NETWORK=CLK_c, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(3[9:12])
    
    wire n25208, n44553, n44055, n43964, n44409, n27481, n27901, 
        n44504, n2;
    wire [31:0]\FRAME_MATCHER.i ;   // verilog/coms.v(116[11:12])
    
    wire n3, n44251, n44586, n44498, n25338, n27998, n44175, n6, 
        n44000, n28367, n44391, n47817, n47823, n2_adj_4590, n3_adj_4591, 
        n2_adj_4592, n3_adj_4593, n40728, n44335, n40678, n47829, 
        n2_adj_4594, n3_adj_4595, n47339, n41622, n40702, n26774;
    wire [7:0]\data_in_frame[0] ;   // verilog/coms.v(97[12:25])
    
    wire n44223, n41642, n45482, n45944, n27454, n27590, n44052, 
        n8, n43820;
    wire [7:0]\data_in_frame[18] ;   // verilog/coms.v(97[12:25])
    
    wire n29291, n2_adj_4596, n3_adj_4597, n29292, n2_adj_4598, n38576, 
        n3345, n29293, n43920, n43896, n44316, n10, n44438, n28070, 
        n26718, n10_adj_4599, n44262, n43968, n1519, n15, n44296, 
        n14, n44042, n6_adj_4600, n29294, n27820, n27370, n27933, 
        n44012, n27475, n27850, n43971, n27544, n43926, n27756, 
        n44226, n44338, n44302, n28186, n44485, n41677, n27834, 
        n6_adj_4601, n43908, n43874, n44125, n1516, n27261, n28314, 
        n12, n41653, n13, n45244, n29295, n27619, Kp_23__N_1561;
    wire [7:0]\data_in_frame[15] ;   // verilog/coms.v(97[12:25])
    
    wire n14_adj_4602, n28046, n44015, n6_adj_4603, n26888, n1247, 
        n44525, n1191, n44087, n27242, n1168, n44096;
    wire [7:0]byte_transmit_counter;   // verilog/coms.v(103[12:33])
    
    wire n48219, n27248, n44009, n48220, n48218, n44325, n42, 
        n44322, n43889, n46, n44, n45, n27797, n43, n48, n52;
    wire [7:0]\data_in_frame[16] ;   // verilog/coms.v(97[12:25])
    
    wire n10_adj_4604, n41598, n40620, n43974, n47, n10_adj_4605, 
        n43995, n12_adj_4606, n44313, n16, n44577, n44248, n44544, 
        n44026, n12_adj_4607, n44495, n45559, n40631, n27861, n44379, 
        n16_adj_4608, n44441, n44373, n17, n26875, n44596, n28177, 
        n10_adj_4609, n43941, n16_adj_4610, n17_adj_4611, n43980, 
        n4_c, n44233, n44003, n14_adj_4612, n10_adj_4613, n6_adj_4614, 
        n48143, n48144, n48042, n48041, n10_adj_4615, n27265, n44488, 
        n6_adj_4616, n48186, n44358, n8_adj_4617, n48187, n44137, 
        n48185, n44240, n51507, n49351, n10_adj_4618, n40704, n41611, 
        n48055, n48053;
    wire [7:0]n9046;
    
    wire n28546, n28996, n48134, n48135, n48081, n27599, n45499, 
        n46044, n48080, n29296, n27420, n51579, n49353, n51567, 
        n51261, n50124;
    wire [7:0]\data_in_frame[17] ;   // verilog/coms.v(97[12:25])
    
    wire n41760, n4_adj_4619, n44217, n48048, n48049, n51483, n49350, 
        n48047;
    wire [7:0]\data_in_frame[19] ;   // verilog/coms.v(97[12:25])
    
    wire n43957, n44350, n41302, n44592, n44146, n4141, n3_adj_4620, 
        n3_adj_4621, n3_adj_4622, n3_adj_4623, n48306, n48307, n48213, 
        n48305, n48214, n48212, n28011, n41059, n27526, n45643, 
        n3_adj_4624, n33811, n46168;
    wire [31:0]\FRAME_MATCHER.state ;   // verilog/coms.v(113[11:16])
    
    wire n19692;
    wire [31:0]\FRAME_MATCHER.state_31__N_2808 ;
    
    wire n3303, n1, n55, n6_adj_4625, n63, n44726, n51606, n52_adj_4626, 
        n43829, n85, n27227;
    wire [31:0]\FRAME_MATCHER.state_31__N_2872 ;
    
    wire n10_adj_4627, n3_adj_4628, n10_adj_4629, n43026, n3_adj_4630, 
        n3_adj_4631, n3_adj_4632, n51585, n49347, n3_adj_4633, n3_adj_4634, 
        n3_adj_4635, n3_adj_4636, n6_adj_4637, n44065, n43134, Kp_23__N_1059, 
        n44094;
    wire [7:0]\data_in_frame[7] ;   // verilog/coms.v(97[12:25])
    
    wire n44243, n43132, n3_adj_4638, n44361, n27554, n40638, n38577, 
        n43130, n44214, n43128, n3_adj_4639, n3_adj_4640, n3_adj_4641, 
        n43126, n43124, n3_adj_4642, n3_adj_4643, n3_adj_4644, n43122, 
        n43120, n5, n43172, n43118, n8_adj_4645, n43832, n29429, 
        n43178, n43116, n43180, n4452, n27231, n27061, n43114, 
        n43182, n43112, n43110, n43108, n43106, n43104, n44_adj_4646, 
        n4_adj_4647, n43795, n43102, n29430, n10_adj_4648, n43098, 
        n43096, n43094, n40252, n35234, n43092, n48_adj_4649, n24234, 
        n29431, n35236, n29432, n22132, n4120, n43729, n43088, 
        n29433, n41814, n40745, n26199, n27730, n3_adj_4650, n3_adj_4651, 
        n29434, n29435, n48114, n48113;
    wire [0:0]n5403;
    wire [2:0]r_SM_Main_2__N_3780;
    
    wire n44813, n33827, n63_adj_4652, n63_adj_4653;
    wire [31:0]\FRAME_MATCHER.state_31__N_2968 ;
    
    wire n43859, n6_adj_4654, n51605, n26673, n41715, n44367, n47429, 
        n44479, n47433, n29436, n43954, n44507, n47439, n44403, 
        n47445, n41651, n41606, n41725, n47451, Kp_23__N_1811, n44599, 
        n44465, n41058, n44129, n44370, n43992, n40684, n40734, 
        n47315, n44284, n46393, n44534, n47211, n47223, n47225, 
        n43923, n47233, n44614, n44122, n47237, n47235, n44376, 
        n43951, n47243, n44038, n44347, n44574, n47249, n44161, 
        n44620, n47257, n48119, n44341, n44237, n46024, n46118, 
        n47263, n44462, n44331, n47285, n44272, n44450, n47291, 
        n48120, n44199, n47269, n44196, n41769, n47295, n45675, 
        n45694, n44531, n40653, n40755, n44155, n27668, n45887, 
        n48147, n48146, n43899, \FRAME_MATCHER.rx_data_ready_prev , 
        n41618, n47851, n27536, n45300, n47611, n8_adj_4655, n43841, 
        n29355, n48092, Kp_23__N_1465, Kp_23__N_1468, n27513, n29279, 
        n7570, n28531, n2_adj_4656, n38575, n28033, n48093, n51489, 
        n49352, n28288, n44006, n27457, n48183, n4_adj_4657, n48182, 
        n6_adj_4658, n41303, n47459, n48089, n48090, n48096;
    wire [7:0]\data_out_frame[26] ;   // verilog/coms.v(98[12:26])
    wire [7:0]\data_out_frame[27] ;   // verilog/coms.v(98[12:26])
    
    wire n51480, n27976, n44245, n48095, n47621, n29280, Kp_23__N_1027, 
        n27506, n44397, n47297, n47303, n44602, n44538, n47417, 
        n44023, n4_adj_4659, n47309, n48230, n48231, n47423, n48069, 
        n48068, n48086, n48087, n48198, n48197, n41793, n10_adj_4660, 
        n47509, n2_adj_4661, n38574, n27520, Kp_23__N_1531, n44290, 
        n14_adj_4662, n44491, n44183, n41679, n6_adj_4663, n41644, 
        n2_adj_4664, n38573, n43948, n41184, n43877, n10_adj_4665, 
        n29281, n41762, n29282, n10_adj_4666, n48083, n12_adj_4667, 
        n48084, n2_adj_4668, n38572, n8_adj_4669, n44168, n10_adj_4670, 
        n43871, n12_adj_4671, n44293, n29283, n44179, n51477, n49349, 
        n41688, n27335, n11, n44425, n48205, n48203, n44562, Kp_23__N_1253, 
        n8_adj_4672, n27979, n9, n44513, n6_adj_4673, n27574, n27873, 
        n47743, n47519, n40688, n6_adj_4674, n29284, n47523, n44035, 
        n24450, n29285, n2_adj_4675, n38571, n44205, n44528, n44611, 
        n48192, n48191, n44299, n47467, n47473, n44565, n44617, 
        n47483, n47485, n44516, n47491, n44072, n44589, n44547, 
        n47497, n12_adj_4676, n33840, n62, n2_adj_4677, n38570, 
        n40972, Kp_23__N_1327, n47503, n771, n4_adj_4678, n27230, 
        n12_adj_4679, n43086, n29286, n2_adj_4680, n38569, n8_adj_4681, 
        n29271, n29272, n44105, n47759, n2_adj_4682, n29273, n29274, 
        n2_adj_4683, n27350, n2_adj_4684, n38568, n28228, n44432, 
        n44116, n27461, n47589, n29275, n6_adj_4685, n44020, n51474, 
        n29276, n44355, n29277, n44102, Kp_23__N_1103, n7569, n7571, 
        n7572, n7573, n47781, n7574, n44344, n27817, n29278;
    wire [7:0]\data_in_frame[23] ;   // verilog/coms.v(97[12:25])
    
    wire n45738, n2_adj_4686, n38567, n7575, n7576, n2_adj_4687, 
        n38566, n7577, n7578, n47867, n2_adj_4688, n2_adj_4689, 
        n2_adj_4690, n2_adj_4691, n2_adj_4692, n2_adj_4693, n7579, 
        n7580, n44308, n43885, n7581, n7582, n47773, n7583, n43932, 
        n7584, n41751, n47863, n7585, n7586, n2_adj_4694, n38565, 
        n47857, n47629, n7587, n7588, n2_adj_4695, n38564, n47635, 
        n44559, n47601, n51647, n29421, n7589, n7590, n7591, n46369, 
        n7592, n7593, n27488, n29422, n8_adj_4696, n47373, n45168, 
        n44453, n45428, n29423, n10_adj_4697, n47379, n6_adj_4698, 
        n47381, n28621, n47879, n47383, n47871, n44728, n47385, 
        n43902, n43986, Kp_23__N_1135, Kp_23__N_1132, n27469, n47389, 
        n47407, n26693, n51495, n49354, n27411, n27495, n47391, 
        n40706, n44556, n27235, n47641, n47607, n47727, n44305, 
        n44459, n47535, n48196, n48194, n44446, n46011, n45375, 
        n29424, n2_adj_4699, n38563, n45888, n47395, n51501, n49345, 
        n45371, n45804, n46382, n46335, n41755, n31, n29425, n47575, 
        n29426, n45796, n45385, n3_adj_4700, n44267, n51573, n51321, 
        n50140, n45560, n2_adj_4701, n38562, n28009, n47837, n47843, 
        n44419, n7, n29427, n2_adj_4702, n38561, n3_adj_4703, n51582, 
        n2_adj_4704, n38560, n3_adj_4705, n29428, n2_adj_4706, n38559, 
        n2_adj_4707, n38558, n28357, n41171, n43960, n41701, n47351, 
        n3_adj_4708, n3_adj_4709, n44142, n47349, n51576, n47359, 
        n38557, n47361, n47357, n47367, n44364, n44394, n27948, 
        n43989, n27952, n43914, n43944, n47801, n47805, n47811, 
        n51570, n45472, n46198, n45477, n27189, n53, n65, n16_adj_4710, 
        n17_adj_4711, n51564, n27136, n38556, n27186, n18, n38555, 
        n19, n12_adj_4712, n16_adj_4713, n17_adj_4714, n10_adj_4715, 
        n14_adj_4716, n10_adj_4717, n6_adj_4718, n12_adj_4719, n18_adj_4720, 
        n29413, n7477, n44841, n45285, n47977, n29414, n29415, 
        n44_adj_4721, n28824, n43762, n45257, n29416, n29417, n51318, 
        n48221, n48222, n51312, n48228, n48227, n51315, n48062, 
        n48063, n51306, n48138, n48137, n51309, n48101, n48102, 
        n51300, n48129, n48128, n51303, n48131, n48132, n51294, 
        n29603, n48123, n48122, n51297, n29601, n29600, n48110, 
        n48111, n51288, n48105, n48104, n51291, n43142, n29044, 
        n42_adj_4722, n51552, n43_adj_4723, n41, n40, n39, n50, 
        n41682, n45_adj_4724, n27025, n11_adj_4725, n44275, n44254, 
        n44583, n27745, n29418, n8_adj_4726, n57, n29419, n5_adj_4727, 
        n29420, n41472, n41816, n44571, n43861, n10_adj_4728, n44287, 
        n2263, n43850, n44084, n27232, n8_adj_4729, n44435, n51267, 
        n7_adj_4730;
    wire [7:0]tx_data;   // verilog/coms.v(106[13:20])
    
    wire n4_adj_4731, n51213, n51546, n17_adj_4732, n41801, n40636, 
        n44257, n29405, n29406, n43905, n43210, n29407, n29408, 
        n51276, n29409, n29410, n41615, n29411, n29412, n161, 
        n27885, n10_adj_4733, n35014, n10_adj_4734, n7_adj_4735, n27406, 
        n30, n27004, n51279, n27809, n40665, n10_adj_4736, n40836, 
        n45489, n44029, n41633, n27612, n35382, n27157, n44724, 
        n44829, n41829, n41809, n38554, n23931, n46039, n47279, 
        n29340, n51270, n51273, n51264, n51258, n41805, n51252, 
        n44140, n51255, n51246, n51231, n51540, n47567, n51249, 
        n51240, n51243, n51234, n43208, n43206, n43202, n34596, 
        n43200, n43198, n43196, n34594, n35232, n43194, n43192, 
        n43190, n43188, n43186, n43184, n43166, n43164, n43162, 
        n43160, n43158, n43156, n43154, n43150, n35228, n43146, 
        n43036, n43032, n7_adj_4737, n29341, n44230, n35263, n29380, 
        n6_adj_4738, Kp_23__N_1008, n45873, n26, n30_adj_4739, n23, 
        n22, n47901, n32, n29381, n27, n43727, n29382, n51237, 
        n51534, n47565, n23975, n43719, n29383, n29384, n7_adj_4740, 
        n29385, n29386, n46020, n41637, n43714, n55_adj_4741, n63_adj_4742, 
        n45_adj_4743, n29342, n10_adj_4744, n44388, n48126, n48125, 
        n10_adj_4745, n40821, n44202, n44172, n44456, n46018, n38591, 
        n38590, n44319, n44482, n40764, n19_adj_4746, n41723, n10_adj_4747, 
        n44134, n41718, n38589, n29387, n29343, n44187, n46161, 
        n29344, n38588, n45721, n38587, n38586, n2326, n38585, 
        tx_transmit_N_3677, n51528, n29443, n29442, n29441, n29440, 
        n29439, n29438, n29437, n31_adj_4748, n7_adj_4749, n29379, 
        n29378, n29377, n29376, n29375, n29374, n29373, n29372, 
        n29371, n29370, n29369, n29368, n29367, n29366, n29365, 
        n29364, n29363, n29362, n29361, n29360, n29359, n29358, 
        n29357, n29356, n29354, n29353, n29352, n29351, n29350, 
        n29349, n38584, n27123, n29348, n29347, n29346, n29345, 
        n38583, n29320, n29319, n29318, n29317, n29316, n38582, 
        n29315, n29314, n29313, n29312, n29311, n29310, n29309, 
        n29308, n29307, n29306, n29305, n38581, n29304, n29303, 
        n29302, n29301, n29300, n29299, n29298, n29297, n29289, 
        n29287, n38580, n29254, n29253, n38579, n29252, n29251, 
        n29250, n38578, n51522, n7_adj_4750, n51516, n34607, n43817, 
        n18_adj_4751, n24, n22_adj_4752, n26_adj_4753, n43938, n41807, 
        n43716, n4_adj_4754, n27279, n45977, n51228, n7_adj_4755, 
        n44580, n37, n44049, n44400, n6_adj_4756, n40779, n12_adj_4757, 
        n40676, n14_adj_4758, n45753, n41711, n28, n26_adj_4759, 
        n44193, n44263, n12_adj_4760, n44472, n27_adj_4761, n25, 
        n45503, n43929, n51510, n7_adj_4762, n44211, n10_adj_4763, 
        n44468, n4_adj_4764, n44522, n44281, n2520, n44149, n51504, 
        n44476, n44406, n44032, n10_adj_4765, n27326, n14_adj_4766, 
        n44119, n51498, n45596, n6_adj_4767, n44208, n50_adj_4768, 
        n48_adj_4769, n41661, n49, n47_adj_4770, n44541, n46_adj_4771, 
        n44605, n45_adj_4772, n56, n51, n44447, n44152, n44143, 
        n44444, n10_adj_4773, n41693, n14_adj_4774, n44416, n28221, 
        n14_adj_4775, n44568, n43917, n44519, n44190, n23_adj_4776, 
        n28400, n22_adj_4777, n44278, n26_adj_4778, n41596, n12_adj_4779, 
        n27771, n44501, n14_adj_4780, n43911, n15_adj_4781, n1130, 
        n51210, n16_adj_4782, n44328, n17_adj_4783, n28_adj_4784, 
        n31_adj_4785, n30_adj_4786, n34, n29, n7_adj_4787, n12_adj_4788, 
        n45747, n45357, n28_adj_4789, n26_adj_4790, n27_adj_4791, 
        n25_adj_4792, n4_adj_4793, n4_adj_4794, n51492, n41609, n16_adj_4795, 
        n44268, n17_adj_4796, n28049, n8_adj_4797, n10_adj_4798, n13_adj_4799, 
        n12_adj_4800, n51486;
    
    SB_LUT4 i2_3_lut (.I0(n25208), .I1(n44553), .I2(\data_out_frame[13] [6]), 
            .I3(GND_net), .O(n44055));
    defparam i2_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i2_4_lut (.I0(n44055), .I1(n43964), .I2(n44409), .I3(n27481), 
            .O(n27901));
    defparam i2_4_lut.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut (.I0(\data_out_frame[20] [6]), .I1(\data_out_frame[23] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n44504));
    defparam i1_2_lut.LUT_INIT = 16'h6666;
    SB_DFFSS \FRAME_MATCHER.i_i3  (.Q(\FRAME_MATCHER.i [3]), .C(CLK_c), 
            .D(n2), .S(n3));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i3_4_lut (.I0(n44251), .I1(n44586), .I2(n44504), .I3(n44498), 
            .O(n25338));
    defparam i3_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_957 (.I0(n27998), .I1(n44175), .I2(GND_net), 
            .I3(GND_net), .O(n6));
    defparam i1_2_lut_adj_957.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut (.I0(n44000), .I1(n28367), .I2(n44391), .I3(n47817), 
            .O(n47823));
    defparam i1_4_lut.LUT_INIT = 16'h6996;
    SB_DFFSS \FRAME_MATCHER.i_i4  (.Q(\FRAME_MATCHER.i [4]), .C(CLK_c), 
            .D(n2_adj_4590), .S(n3_adj_4591));   // verilog/coms.v(128[12] 303[6])
    SB_DFFSS \FRAME_MATCHER.i_i2  (.Q(\FRAME_MATCHER.i [2]), .C(CLK_c), 
            .D(n2_adj_4592), .S(n3_adj_4593));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i1_4_lut_adj_958 (.I0(n40728), .I1(n47823), .I2(n44335), .I3(n40678), 
            .O(n47829));
    defparam i1_4_lut_adj_958.LUT_INIT = 16'h6996;
    SB_DFFSS \FRAME_MATCHER.i_i1  (.Q(\FRAME_MATCHER.i [1]), .C(CLK_c), 
            .D(n2_adj_4594), .S(n3_adj_4595));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i1_4_lut_adj_959 (.I0(n47339), .I1(n41622), .I2(n40702), .I3(n47829), 
            .O(n26774));
    defparam i1_4_lut_adj_959.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_960 (.I0(\data_in_frame[0] [7]), .I1(\data_in_frame[3] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n44223));
    defparam i1_2_lut_adj_960.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut (.I0(\data_out_frame[23] [4]), .I1(n41642), .I2(\data_out_frame[23] [3]), 
            .I3(n6), .O(n45482));
    defparam i4_4_lut.LUT_INIT = 16'h9669;
    SB_LUT4 i3_4_lut_adj_961 (.I0(\data_out_frame[25] [4]), .I1(n25338), 
            .I2(n45482), .I3(\data_out_frame[25] [5]), .O(n45944));
    defparam i3_4_lut_adj_961.LUT_INIT = 16'h9669;
    SB_LUT4 i1_4_lut_adj_962 (.I0(n27454), .I1(n27590), .I2(n44223), .I3(\data_in_frame[5] [5]), 
            .O(n44052));
    defparam i1_4_lut_adj_962.LUT_INIT = 16'h6996;
    SB_LUT4 i15343_3_lut_4_lut (.I0(n8), .I1(n43820), .I2(rx_data[5]), 
            .I3(\data_in_frame[18] [5]), .O(n29291));
    defparam i15343_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFFSS \FRAME_MATCHER.i_i0  (.Q(\FRAME_MATCHER.i [0]), .C(CLK_c), 
            .D(n2_adj_4596), .S(n3_adj_4597));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i15344_3_lut_4_lut (.I0(n8), .I1(n43820), .I2(rx_data[4]), 
            .I3(\data_in_frame[18] [4]), .O(n29292));
    defparam i15344_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 add_43_25_lut (.I0(n3345), .I1(\FRAME_MATCHER.i [23]), .I2(GND_net), 
            .I3(n38576), .O(n2_adj_4598)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_25_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i15345_3_lut_4_lut (.I0(n8), .I1(n43820), .I2(rx_data[3]), 
            .I3(\data_in_frame[18] [3]), .O(n29293));
    defparam i15345_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_adj_963 (.I0(\data_out_frame[10] [4]), .I1(n43920), 
            .I2(\data_out_frame[6] [0]), .I3(GND_net), .O(n43896));   // verilog/coms.v(76[16:27])
    defparam i2_3_lut_adj_963.LUT_INIT = 16'h9696;
    SB_LUT4 i4_4_lut_adj_964 (.I0(n43896), .I1(\data_out_frame[8] [2]), 
            .I2(\data_out_frame[8] [3]), .I3(n44316), .O(n10));   // verilog/coms.v(76[16:27])
    defparam i4_4_lut_adj_964.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_965 (.I0(\data_out_frame[17] [2]), .I1(\data_out_frame[17] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n44438));
    defparam i1_2_lut_adj_965.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_966 (.I0(\data_out_frame[15] [0]), .I1(\data_out_frame[15] [1]), 
            .I2(\data_out_frame[13] [0]), .I3(GND_net), .O(n28070));
    defparam i2_3_lut_adj_966.LUT_INIT = 16'h9696;
    SB_LUT4 i4_4_lut_adj_967 (.I0(\data_out_frame[16] [7]), .I1(n28070), 
            .I2(n44438), .I3(n26718), .O(n10_adj_4599));
    defparam i4_4_lut_adj_967.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut (.I0(\data_out_frame[19] [3]), .I1(n10_adj_4599), .I2(\data_out_frame[21] [4]), 
            .I3(GND_net), .O(n44262));
    defparam i5_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_968 (.I0(\data_out_frame[12] [5]), .I1(\data_out_frame[14] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n43968));
    defparam i1_2_lut_adj_968.LUT_INIT = 16'h6666;
    SB_LUT4 i6_4_lut (.I0(\data_out_frame[5] [6]), .I1(n1519), .I2(\data_out_frame[12] [6]), 
            .I3(\data_out_frame[4] [2]), .O(n15));   // verilog/coms.v(73[16:27])
    defparam i6_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut (.I0(n15), .I1(n44296), .I2(n14), .I3(\data_out_frame[10] [5]), 
            .O(n44042));   // verilog/coms.v(73[16:27])
    defparam i8_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_969 (.I0(\data_out_frame[17] [1]), .I1(\data_out_frame[15] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_4600));
    defparam i1_2_lut_adj_969.LUT_INIT = 16'h6666;
    SB_LUT4 i15346_3_lut_4_lut (.I0(n8), .I1(n43820), .I2(rx_data[2]), 
            .I3(\data_in_frame[18] [2]), .O(n29294));
    defparam i15346_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i3_4_lut_adj_970 (.I0(\data_in_frame[11] [2]), .I1(n27820), 
            .I2(n27370), .I3(n27933), .O(n44012));   // verilog/coms.v(72[16:27])
    defparam i3_4_lut_adj_970.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_971 (.I0(\data_in_frame[3] [5]), .I1(\data_in_frame[5] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n27475));   // verilog/coms.v(79[16:27])
    defparam i1_2_lut_adj_971.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_972 (.I0(\data_in_frame[14] [0]), .I1(n27850), 
            .I2(n43971), .I3(n27544), .O(n43926));
    defparam i3_4_lut_adj_972.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_973 (.I0(n27756), .I1(\data_out_frame[16] [7]), 
            .I2(n44042), .I3(n6_adj_4600), .O(n44226));
    defparam i4_4_lut_adj_973.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_974 (.I0(\data_in_frame[13] [6]), .I1(\data_in_frame[13] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n44338));
    defparam i1_2_lut_adj_974.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_975 (.I0(\data_out_frame[19] [2]), .I1(n44302), 
            .I2(GND_net), .I3(GND_net), .O(n28186));   // verilog/coms.v(77[16:43])
    defparam i1_2_lut_adj_975.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_976 (.I0(\data_out_frame[21] [3]), .I1(n44226), 
            .I2(GND_net), .I3(GND_net), .O(n44485));
    defparam i1_2_lut_adj_976.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_977 (.I0(n41677), .I1(n28186), .I2(n27834), .I3(n6_adj_4601), 
            .O(n27998));
    defparam i4_4_lut_adj_977.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_978 (.I0(\data_out_frame[4] [1]), .I1(n43908), 
            .I2(n43874), .I3(\data_out_frame[10] [3]), .O(n1519));   // verilog/coms.v(73[16:27])
    defparam i3_4_lut_adj_978.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_979 (.I0(\data_out_frame[19] [0]), .I1(\data_out_frame[19] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n44125));
    defparam i1_2_lut_adj_979.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_980 (.I0(\data_out_frame[14] [6]), .I1(n1519), 
            .I2(n1516), .I3(n27261), .O(n28314));
    defparam i3_4_lut_adj_980.LUT_INIT = 16'h6996;
    SB_LUT4 i4_2_lut (.I0(\data_out_frame[16] [7]), .I1(n27834), .I2(GND_net), 
            .I3(GND_net), .O(n12));   // verilog/coms.v(86[17:28])
    defparam i4_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i5_4_lut (.I0(\data_out_frame[21] [2]), .I1(n28314), .I2(n41653), 
            .I3(n44125), .O(n13));   // verilog/coms.v(86[17:28])
    defparam i5_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut (.I0(n13), .I1(\data_out_frame[17] [0]), .I2(n12), 
            .I3(n41677), .O(n45244));   // verilog/coms.v(86[17:28])
    defparam i7_4_lut.LUT_INIT = 16'h9669;
    SB_LUT4 i15347_3_lut_4_lut (.I0(n8), .I1(n43820), .I2(rx_data[1]), 
            .I3(\data_in_frame[18] [1]), .O(n29295));
    defparam i15347_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_981 (.I0(\data_out_frame[11] [5]), .I1(\data_out_frame[11] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n27619));
    defparam i1_2_lut_adj_981.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_982 (.I0(\data_out_frame[12] [5]), .I1(\data_out_frame[12] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n27261));   // verilog/coms.v(86[17:63])
    defparam i1_2_lut_adj_982.LUT_INIT = 16'h6666;
    SB_LUT4 i6_4_lut_adj_983 (.I0(n44338), .I1(Kp_23__N_1561), .I2(n43926), 
            .I3(\data_in_frame[15] [6]), .O(n14_adj_4602));
    defparam i6_4_lut_adj_983.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_984 (.I0(n28046), .I1(\data_out_frame[9] [3]), 
            .I2(n44015), .I3(n6_adj_4603), .O(n26888));
    defparam i4_4_lut_adj_984.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_985 (.I0(\data_out_frame[8] [5]), .I1(\data_out_frame[10] [6]), 
            .I2(n1247), .I3(GND_net), .O(n44316));   // verilog/coms.v(76[16:27])
    defparam i2_3_lut_adj_985.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_986 (.I0(\data_out_frame[8] [1]), .I1(\data_out_frame[7] [7]), 
            .I2(\data_out_frame[5] [5]), .I3(GND_net), .O(n44525));
    defparam i2_3_lut_adj_986.LUT_INIT = 16'h9696;
    SB_LUT4 i375_2_lut (.I0(\data_out_frame[5] [7]), .I1(\data_out_frame[5] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n1191));   // verilog/coms.v(72[16:27])
    defparam i375_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_987 (.I0(\data_out_frame[5] [4]), .I1(\data_out_frame[5] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n44087));   // verilog/coms.v(72[16:62])
    defparam i1_2_lut_adj_987.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_988 (.I0(\data_out_frame[5] [5]), .I1(n44087), 
            .I2(n27242), .I3(n1191), .O(n1168));   // verilog/coms.v(72[16:62])
    defparam i3_4_lut_adj_988.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_989 (.I0(\data_out_frame[6] [7]), .I1(\data_out_frame[4] [5]), 
            .I2(n1168), .I3(\data_out_frame[5] [0]), .O(n44015));   // verilog/coms.v(86[17:70])
    defparam i3_4_lut_adj_989.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_990 (.I0(\data_out_frame[9] [5]), .I1(\data_out_frame[9] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n44096));
    defparam i1_2_lut_adj_990.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_991 (.I0(\data_out_frame[8] [4]), .I1(\data_out_frame[8] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n44296));   // verilog/coms.v(73[16:27])
    defparam i1_2_lut_adj_991.LUT_INIT = 16'h6666;
    SB_LUT4 i32632_3_lut (.I0(\data_out_frame[6] [4]), .I1(\data_out_frame[7] [4]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n48219));
    defparam i32632_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2_3_lut_adj_992 (.I0(\data_out_frame[4] [1]), .I1(\data_out_frame[4] [0]), 
            .I2(\data_out_frame[6] [2]), .I3(GND_net), .O(n27248));   // verilog/coms.v(75[16:43])
    defparam i2_3_lut_adj_992.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_993 (.I0(\data_out_frame[4] [4]), .I1(\data_out_frame[6] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n44009));
    defparam i1_2_lut_adj_993.LUT_INIT = 16'h6666;
    SB_LUT4 i32633_4_lut (.I0(n48219), .I1(byte_transmit_counter[1]), .I2(byte_transmit_counter[2]), 
            .I3(byte_transmit_counter[0]), .O(n48220));
    defparam i32633_4_lut.LUT_INIT = 16'haca3;
    SB_LUT4 i32631_3_lut (.I0(\data_out_frame[4] [4]), .I1(\data_out_frame[5] [4]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n48218));
    defparam i32631_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_994 (.I0(\data_out_frame[9] [0]), .I1(\data_out_frame[9] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n44325));
    defparam i1_2_lut_adj_994.LUT_INIT = 16'h6666;
    SB_LUT4 i15_4_lut (.I0(n43908), .I1(\data_out_frame[9] [1]), .I2(\data_out_frame[9] [6]), 
            .I3(n44325), .O(n42));
    defparam i15_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i19_4_lut (.I0(\data_out_frame[7] [6]), .I1(n44322), .I2(n44009), 
            .I3(n43889), .O(n46));
    defparam i19_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i17_4_lut (.I0(\data_out_frame[8] [7]), .I1(\data_out_frame[7] [2]), 
            .I2(\data_out_frame[7] [1]), .I3(n44296), .O(n44));
    defparam i17_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i18_4_lut (.I0(\data_out_frame[8] [6]), .I1(\data_out_frame[7] [3]), 
            .I2(\data_out_frame[7] [0]), .I3(\data_out_frame[8] [0]), .O(n45));
    defparam i18_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i16_4_lut (.I0(n1247), .I1(n27797), .I2(\data_out_frame[9] [3]), 
            .I3(\data_out_frame[6] [3]), .O(n43));
    defparam i16_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i21_4_lut (.I0(\data_out_frame[4] [7]), .I1(n42), .I2(\data_out_frame[9] [7]), 
            .I3(n44096), .O(n48));
    defparam i21_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i25_4_lut (.I0(n43), .I1(n45), .I2(n44), .I3(n46), .O(n52));
    defparam i25_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_995 (.I0(\data_in_frame[16] [0]), .I1(n14_adj_4602), 
            .I2(n10_adj_4604), .I3(n41598), .O(n40620));
    defparam i7_4_lut_adj_995.LUT_INIT = 16'h6996;
    SB_LUT4 i20_4_lut (.I0(\data_out_frame[5] [5]), .I1(n43974), .I2(n44015), 
            .I3(\data_out_frame[4] [6]), .O(n47));
    defparam i20_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_996 (.I0(\data_out_frame[11] [1]), .I1(\data_out_frame[11] [0]), 
            .I2(\data_out_frame[11] [3]), .I3(\data_out_frame[11] [2]), 
            .O(n10_adj_4605));
    defparam i1_4_lut_adj_996.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_997 (.I0(n43995), .I1(n47), .I2(n52), .I3(n48), 
            .O(n12_adj_4606));
    defparam i3_4_lut_adj_997.LUT_INIT = 16'h9669;
    SB_LUT4 i7_4_lut_adj_998 (.I0(n44313), .I1(\data_out_frame[10] [5]), 
            .I2(\data_out_frame[10] [4]), .I3(n10_adj_4605), .O(n16));
    defparam i7_4_lut_adj_998.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut_adj_999 (.I0(n44316), .I1(n16), .I2(n12_adj_4606), 
            .I3(\data_out_frame[10] [7]), .O(n44577));
    defparam i8_4_lut_adj_999.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1000 (.I0(\data_out_frame[11] [6]), .I1(\data_out_frame[11] [7]), 
            .I2(n44577), .I3(GND_net), .O(n44248));   // verilog/coms.v(72[16:27])
    defparam i2_3_lut_adj_1000.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1001 (.I0(\data_out_frame[14] [1]), .I1(n44544), 
            .I2(GND_net), .I3(GND_net), .O(n44026));
    defparam i1_2_lut_adj_1001.LUT_INIT = 16'h6666;
    SB_LUT4 i5_4_lut_adj_1002 (.I0(\data_out_frame[12] [1]), .I1(n44248), 
            .I2(\data_out_frame[12] [2]), .I3(\data_out_frame[12] [0]), 
            .O(n12_adj_4607));
    defparam i5_4_lut_adj_1002.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1003 (.I0(\data_out_frame[11] [4]), .I1(n12_adj_4607), 
            .I2(n44495), .I3(n26888), .O(n45559));
    defparam i6_4_lut_adj_1003.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1004 (.I0(n40631), .I1(n40620), .I2(GND_net), 
            .I3(GND_net), .O(n27861));
    defparam i1_2_lut_adj_1004.LUT_INIT = 16'h6666;
    SB_LUT4 i6_4_lut_adj_1005 (.I0(n44087), .I1(\data_out_frame[13] [7]), 
            .I2(n44495), .I3(n44379), .O(n16_adj_4608));
    defparam i6_4_lut_adj_1005.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1006 (.I0(n45559), .I1(n44441), .I2(n44577), 
            .I3(n44373), .O(n17));
    defparam i7_4_lut_adj_1006.LUT_INIT = 16'h9669;
    SB_LUT4 i9_4_lut (.I0(n17), .I1(\data_out_frame[9] [5]), .I2(n16_adj_4608), 
            .I3(n27619), .O(n26875));
    defparam i9_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1007 (.I0(\data_in_frame[14] [7]), .I1(\data_in_frame[15] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n44596));
    defparam i1_2_lut_adj_1007.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1008 (.I0(\data_out_frame[10] [3]), .I1(\data_out_frame[10] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n44313));   // verilog/coms.v(76[16:27])
    defparam i1_2_lut_adj_1008.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1009 (.I0(\data_out_frame[6] [0]), .I1(\data_out_frame[6] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n43889));
    defparam i1_2_lut_adj_1009.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1010 (.I0(n43889), .I1(\data_out_frame[5] [4]), 
            .I2(n28177), .I3(n44313), .O(n10_adj_4609));   // verilog/coms.v(76[16:27])
    defparam i4_4_lut_adj_1010.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_1011 (.I0(\data_out_frame[8] [2]), .I1(n10_adj_4609), 
            .I2(\data_out_frame[4] [0]), .I3(GND_net), .O(n1516));   // verilog/coms.v(76[16:27])
    defparam i5_3_lut_adj_1011.LUT_INIT = 16'h9696;
    SB_LUT4 i6_4_lut_adj_1012 (.I0(\data_out_frame[12] [3]), .I1(\data_out_frame[9] [7]), 
            .I2(\data_out_frame[8] [1]), .I3(n43941), .O(n16_adj_4610));   // verilog/coms.v(76[16:27])
    defparam i6_4_lut_adj_1012.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1013 (.I0(\data_out_frame[5] [7]), .I1(\data_out_frame[10] [2]), 
            .I2(\data_out_frame[5] [3]), .I3(\data_out_frame[10] [1]), .O(n17_adj_4611));   // verilog/coms.v(76[16:27])
    defparam i7_4_lut_adj_1013.LUT_INIT = 16'h6996;
    SB_LUT4 i9_4_lut_adj_1014 (.I0(n17_adj_4611), .I1(\data_out_frame[6] [0]), 
            .I2(n16_adj_4610), .I3(\data_out_frame[7] [5]), .O(n43980));   // verilog/coms.v(76[16:27])
    defparam i9_4_lut_adj_1014.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1015 (.I0(\data_out_frame[14] [5]), .I1(n43980), 
            .I2(\data_out_frame[12] [4]), .I3(n1516), .O(n27756));   // verilog/coms.v(76[16:43])
    defparam i3_4_lut_adj_1015.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1016 (.I0(\data_out_frame[7] [2]), .I1(\data_out_frame[5] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n4_c));   // verilog/coms.v(86[17:28])
    defparam i1_2_lut_adj_1016.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1017 (.I0(\data_in_frame[10] [5]), .I1(\data_in_frame[12] [6]), 
            .I2(\data_in_frame[12] [4]), .I3(\data_in_frame[12] [5]), .O(n44233));
    defparam i3_4_lut_adj_1017.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1018 (.I0(\data_out_frame[12] [1]), .I1(\data_out_frame[11] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n44379));   // verilog/coms.v(72[16:27])
    defparam i1_2_lut_adj_1018.LUT_INIT = 16'h6666;
    SB_LUT4 i6_4_lut_adj_1019 (.I0(\data_out_frame[9] [4]), .I1(\data_out_frame[12] [0]), 
            .I2(n44003), .I3(\data_out_frame[9] [6]), .O(n14_adj_4612));   // verilog/coms.v(72[16:27])
    defparam i6_4_lut_adj_1019.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1020 (.I0(\data_out_frame[14] [2]), .I1(n14_adj_4612), 
            .I2(n10_adj_4613), .I3(n44379), .O(n44544));   // verilog/coms.v(72[16:27])
    defparam i7_4_lut_adj_1020.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1021 (.I0(n44302), .I1(n44544), .I2(GND_net), 
            .I3(GND_net), .O(n6_adj_4614));
    defparam i1_2_lut_adj_1021.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1022 (.I0(\data_out_frame[16] [4]), .I1(\data_out_frame[18] [6]), 
            .I2(n41677), .I3(n6_adj_4614), .O(n41653));
    defparam i4_4_lut_adj_1022.LUT_INIT = 16'h6996;
    SB_LUT4 i32556_3_lut (.I0(\data_out_frame[16] [6]), .I1(\data_out_frame[17] [6]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n48143));
    defparam i32556_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i32557_3_lut (.I0(\data_out_frame[18] [6]), .I1(\data_out_frame[19] [6]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n48144));
    defparam i32557_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_1023 (.I0(\data_out_frame[7] [7]), .I1(\data_out_frame[7] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n43941));   // verilog/coms.v(76[16:27])
    defparam i1_2_lut_adj_1023.LUT_INIT = 16'h6666;
    SB_LUT4 i32455_3_lut (.I0(\data_out_frame[22] [6]), .I1(\data_out_frame[23] [6]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n48042));
    defparam i32455_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i32454_3_lut (.I0(\data_out_frame[20] [6]), .I1(\data_out_frame[21] [6]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n48041));
    defparam i32454_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_1024 (.I0(\data_out_frame[9] [6]), .I1(\data_out_frame[12] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n44373));   // verilog/coms.v(75[16:27])
    defparam i1_2_lut_adj_1024.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1025 (.I0(\data_out_frame[7] [5]), .I1(\data_out_frame[7] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n27797));   // verilog/coms.v(75[16:27])
    defparam i1_2_lut_adj_1025.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1026 (.I0(\data_out_frame[10] [1]), .I1(\data_out_frame[10] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n43995));   // verilog/coms.v(75[16:27])
    defparam i1_2_lut_adj_1026.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1027 (.I0(n43995), .I1(\data_out_frame[5] [6]), 
            .I2(n27797), .I3(n44373), .O(n10_adj_4615));   // verilog/coms.v(75[16:27])
    defparam i4_4_lut_adj_1027.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_1028 (.I0(\data_out_frame[5] [2]), .I1(n10_adj_4615), 
            .I2(n28177), .I3(GND_net), .O(n27265));   // verilog/coms.v(75[16:27])
    defparam i5_3_lut_adj_1028.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1029 (.I0(\data_out_frame[5] [2]), .I1(\data_out_frame[5] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n27242));   // verilog/coms.v(74[16:34])
    defparam i1_2_lut_adj_1029.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1030 (.I0(n44233), .I1(n44596), .I2(\data_in_frame[16] [7]), 
            .I3(GND_net), .O(n44488));
    defparam i2_3_lut_adj_1030.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1031 (.I0(\data_out_frame[9] [5]), .I1(\data_out_frame[9] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_4616));
    defparam i1_2_lut_adj_1031.LUT_INIT = 16'h6666;
    SB_LUT4 i32599_3_lut (.I0(\data_out_frame[6] [0]), .I1(\data_out_frame[7] [0]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n48186));
    defparam i32599_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3_3_lut (.I0(\data_in_frame[14] [5]), .I1(n44358), .I2(n44488), 
            .I3(GND_net), .O(n8_adj_4617));
    defparam i3_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i32600_4_lut (.I0(n48186), .I1(byte_transmit_counter[1]), .I2(byte_transmit_counter[2]), 
            .I3(byte_transmit_counter[0]), .O(n48187));
    defparam i32600_4_lut.LUT_INIT = 16'ha3a0;
    SB_LUT4 i4_4_lut_adj_1032 (.I0(\data_out_frame[5] [5]), .I1(\data_out_frame[7] [6]), 
            .I2(\data_out_frame[10] [0]), .I3(n6_adj_4616), .O(n44003));
    defparam i4_4_lut_adj_1032.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1033 (.I0(\data_out_frame[7] [5]), .I1(n28046), 
            .I2(GND_net), .I3(GND_net), .O(n44441));
    defparam i1_2_lut_adj_1033.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1034 (.I0(\data_out_frame[5] [2]), .I1(\data_out_frame[7] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n44137));
    defparam i1_2_lut_adj_1034.LUT_INIT = 16'h6666;
    SB_LUT4 i32598_3_lut (.I0(\data_out_frame[4] [0]), .I1(\data_out_frame[5] [0]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n48185));
    defparam i32598_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_1035 (.I0(n27265), .I1(\data_out_frame[14] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n44240));
    defparam i1_2_lut_adj_1035.LUT_INIT = 16'h6666;
    SB_LUT4 i33821_2_lut (.I0(n51507), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n49351));
    defparam i33821_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i4_4_lut_adj_1036 (.I0(n44240), .I1(\data_out_frame[12] [1]), 
            .I2(\data_out_frame[11] [7]), .I3(n44137), .O(n10_adj_4618));
    defparam i4_4_lut_adj_1036.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1037 (.I0(\data_out_frame[16] [3]), .I1(n40704), 
            .I2(GND_net), .I3(GND_net), .O(n41611));
    defparam i1_2_lut_adj_1037.LUT_INIT = 16'h6666;
    SB_LUT4 i32468_4_lut (.I0(\data_out_frame[6] [1]), .I1(byte_transmit_counter[0]), 
            .I2(byte_transmit_counter[2]), .I3(\data_out_frame[7] [1]), 
            .O(n48055));
    defparam i32468_4_lut.LUT_INIT = 16'hec2c;
    SB_LUT4 i32466_3_lut (.I0(\data_out_frame[4] [1]), .I1(\data_out_frame[5] [1]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n48053));
    defparam i32466_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFESR byte_transmit_counter_i0_i1 (.Q(byte_transmit_counter[1]), .C(CLK_c), 
            .E(n28546), .D(n9046[1]), .R(n28996));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i1_2_lut_adj_1038 (.I0(n45244), .I1(\data_out_frame[23] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n44251));
    defparam i1_2_lut_adj_1038.LUT_INIT = 16'h9999;
    SB_LUT4 i32547_3_lut (.I0(\data_out_frame[16] [5]), .I1(\data_out_frame[17] [5]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n48134));
    defparam i32547_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFESR byte_transmit_counter_i0_i2 (.Q(byte_transmit_counter[2]), .C(CLK_c), 
            .E(n28546), .D(n9046[2]), .R(n28996));   // verilog/coms.v(128[12] 303[6])
    SB_DFFESR byte_transmit_counter_i0_i3 (.Q(byte_transmit_counter[3]), .C(CLK_c), 
            .E(n28546), .D(n9046[3]), .R(n28996));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i32548_3_lut (.I0(\data_out_frame[18] [5]), .I1(\data_out_frame[19] [5]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n48135));
    defparam i32548_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i32494_3_lut (.I0(\data_out_frame[22] [5]), .I1(\data_out_frame[23] [5]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n48081));
    defparam i32494_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3_4_lut_adj_1039 (.I0(n27599), .I1(n44251), .I2(n44175), 
            .I3(n41642), .O(n45499));
    defparam i3_4_lut_adj_1039.LUT_INIT = 16'h6996;
    SB_DFFESR byte_transmit_counter_i0_i4 (.Q(byte_transmit_counter[4]), .C(CLK_c), 
            .E(n28546), .D(n9046[4]), .R(n28996));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i2_3_lut_adj_1040 (.I0(n45499), .I1(\data_out_frame[25] [5]), 
            .I2(\data_out_frame[25] [6]), .I3(GND_net), .O(n46044));
    defparam i2_3_lut_adj_1040.LUT_INIT = 16'h6969;
    SB_DFFESR byte_transmit_counter_i0_i5 (.Q(byte_transmit_counter[5]), .C(CLK_c), 
            .E(n28546), .D(n9046[5]), .R(n28996));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i32493_3_lut (.I0(\data_out_frame[20] [5]), .I1(\data_out_frame[21] [5]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n48080));
    defparam i32493_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFESR byte_transmit_counter_i0_i6 (.Q(byte_transmit_counter[6]), .C(CLK_c), 
            .E(n28546), .D(n9046[6]), .R(n28996));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i15348_3_lut_4_lut (.I0(n8), .I1(n43820), .I2(rx_data[0]), 
            .I3(\data_in_frame[18] [0]), .O(n29296));
    defparam i15348_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i26_2_lut (.I0(\data_in_frame[1] [3]), .I1(\data_in_frame[1] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n27420));   // verilog/coms.v(97[12:25])
    defparam i26_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i33820_2_lut (.I0(n51579), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n49353));
    defparam i33820_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i34536_3_lut (.I0(n51567), .I1(n51261), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n50124));
    defparam i34536_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFESR byte_transmit_counter_i0_i7 (.Q(byte_transmit_counter[7]), .C(CLK_c), 
            .E(n28546), .D(n9046[7]), .R(n28996));   // verilog/coms.v(128[12] 303[6])
    SB_DFF IntegralLimit_i0_i1 (.Q(IntegralLimit[1]), .C(CLK_c), .D(n29158));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i1_4_lut_adj_1041 (.I0(\data_in_frame[17] [1]), .I1(n41760), 
            .I2(n8_adj_4617), .I3(n4_adj_4619), .O(n44217));
    defparam i1_4_lut_adj_1041.LUT_INIT = 16'h9669;
    SB_LUT4 i32461_3_lut (.I0(\data_out_frame[6] [2]), .I1(\data_out_frame[7] [2]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n48048));
    defparam i32461_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i32462_4_lut (.I0(n48048), .I1(byte_transmit_counter[0]), .I2(byte_transmit_counter[2]), 
            .I3(byte_transmit_counter[1]), .O(n48049));
    defparam i32462_4_lut.LUT_INIT = 16'ha0a3;
    SB_LUT4 i33822_2_lut (.I0(n51483), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n49350));
    defparam i33822_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i32460_3_lut (.I0(\data_out_frame[4] [2]), .I1(\data_out_frame[5] [2]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n48047));
    defparam i32460_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1042 (.I0(\data_in_frame[19] [0]), .I1(n43957), 
            .I2(n44350), .I3(n41302), .O(n44592));
    defparam i1_4_lut_adj_1042.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1043 (.I0(\data_in_frame[18] [6]), .I1(n44592), 
            .I2(GND_net), .I3(GND_net), .O(n44146));
    defparam i1_2_lut_adj_1043.LUT_INIT = 16'h6666;
    SB_LUT4 select_686_Select_5_i3_2_lut (.I0(\FRAME_MATCHER.i [5]), .I1(n4141), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4620));
    defparam select_686_Select_5_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_686_Select_6_i3_2_lut (.I0(\FRAME_MATCHER.i [6]), .I1(n4141), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4621));
    defparam select_686_Select_6_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_686_Select_7_i3_2_lut (.I0(\FRAME_MATCHER.i [7]), .I1(n4141), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4622));
    defparam select_686_Select_7_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_686_Select_8_i3_2_lut (.I0(\FRAME_MATCHER.i [8]), .I1(n4141), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4623));
    defparam select_686_Select_8_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i32719_3_lut (.I0(\data_out_frame[6] [3]), .I1(\data_out_frame[7] [3]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n48306));
    defparam i32719_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i32720_4_lut (.I0(n48306), .I1(byte_transmit_counter[1]), .I2(byte_transmit_counter[2]), 
            .I3(byte_transmit_counter[0]), .O(n48307));
    defparam i32720_4_lut.LUT_INIT = 16'hafa3;
    SB_LUT4 i32626_3_lut (.I0(\data_out_frame[6] [5]), .I1(\data_out_frame[7] [5]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n48213));
    defparam i32626_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i32718_3_lut (.I0(\data_out_frame[4] [3]), .I1(\data_out_frame[5] [3]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n48305));
    defparam i32718_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i32627_4_lut (.I0(n48213), .I1(byte_transmit_counter[1]), .I2(byte_transmit_counter[2]), 
            .I3(byte_transmit_counter[0]), .O(n48214));
    defparam i32627_4_lut.LUT_INIT = 16'ha3a0;
    SB_LUT4 i32625_3_lut (.I0(\data_out_frame[4] [5]), .I1(\data_out_frame[5] [5]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n48212));
    defparam i32625_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut_4_lut (.I0(n28011), .I1(n41059), .I2(\data_in_frame[14] [7]), 
            .I3(n27526), .O(n45643));
    defparam i1_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 select_686_Select_9_i3_2_lut (.I0(\FRAME_MATCHER.i [9]), .I1(n4141), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4624));
    defparam select_686_Select_9_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i3_4_lut_adj_1044 (.I0(\data_in[1] [0]), .I1(n33811), .I2(\data_in[3] [0]), 
            .I3(\data_in[0] [6]), .O(n46168));   // verilog/coms.v(96[12:19])
    defparam i3_4_lut_adj_1044.LUT_INIT = 16'h0080;
    SB_LUT4 i1_3_lut (.I0(n46168), .I1(\FRAME_MATCHER.state [1]), .I2(n19692), 
            .I3(GND_net), .O(\FRAME_MATCHER.state_31__N_2808 [1]));   // verilog/coms.v(96[12:19])
    defparam i1_3_lut.LUT_INIT = 16'heaea;
    SB_LUT4 i2_4_lut_adj_1045 (.I0(n3303), .I1(n1), .I2(n55), .I3(\FRAME_MATCHER.state_31__N_2808 [1]), 
            .O(n6_adj_4625));   // verilog/coms.v(116[11:12])
    defparam i2_4_lut_adj_1045.LUT_INIT = 16'hcfce;
    SB_LUT4 i3_4_lut_adj_1046 (.I0(n63), .I1(n6_adj_4625), .I2(\FRAME_MATCHER.state_31__N_2808 [1]), 
            .I3(n44726), .O(n51606));   // verilog/coms.v(116[11:12])
    defparam i3_4_lut_adj_1046.LUT_INIT = 16'hddfd;
    SB_LUT4 i1_3_lut_adj_1047 (.I0(\FRAME_MATCHER.state [3]), .I1(n52_adj_4626), 
            .I2(n43829), .I3(GND_net), .O(n85));
    defparam i1_3_lut_adj_1047.LUT_INIT = 16'ha8a8;
    SB_LUT4 i1_4_lut_adj_1048 (.I0(\FRAME_MATCHER.state [2]), .I1(n85), 
            .I2(n27227), .I3(\FRAME_MATCHER.state_31__N_2872 [3]), .O(n10_adj_4627));   // verilog/coms.v(116[11:12])
    defparam i1_4_lut_adj_1048.LUT_INIT = 16'hcdcc;
    SB_LUT4 select_686_Select_15_i3_2_lut (.I0(\FRAME_MATCHER.i [15]), .I1(n4141), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4628));
    defparam select_686_Select_15_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1049 (.I0(\FRAME_MATCHER.state [4]), .I1(n10_adj_4629), 
            .I2(GND_net), .I3(GND_net), .O(n43026));
    defparam i1_2_lut_adj_1049.LUT_INIT = 16'h8888;
    SB_LUT4 select_686_Select_16_i3_2_lut (.I0(\FRAME_MATCHER.i [16]), .I1(n4141), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4630));
    defparam select_686_Select_16_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_686_Select_17_i3_2_lut (.I0(\FRAME_MATCHER.i [17]), .I1(n4141), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4631));
    defparam select_686_Select_17_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_686_Select_18_i3_2_lut (.I0(\FRAME_MATCHER.i [18]), .I1(n4141), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4632));
    defparam select_686_Select_18_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i33789_2_lut (.I0(n51585), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n49347));
    defparam i33789_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 select_686_Select_19_i3_2_lut (.I0(\FRAME_MATCHER.i [19]), .I1(n4141), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4633));
    defparam select_686_Select_19_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_686_Select_20_i3_2_lut (.I0(\FRAME_MATCHER.i [20]), .I1(n4141), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4634));
    defparam select_686_Select_20_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_686_Select_21_i3_2_lut (.I0(\FRAME_MATCHER.i [21]), .I1(n4141), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4635));
    defparam select_686_Select_21_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_686_Select_22_i3_2_lut (.I0(\FRAME_MATCHER.i [22]), .I1(n4141), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4636));
    defparam select_686_Select_22_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut_adj_1050 (.I0(\data_in_frame[21] [2]), .I1(\data_in_frame[19] [2]), 
            .I2(n6_adj_4637), .I3(n44146), .O(n44065));
    defparam i1_4_lut_adj_1050.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1051 (.I0(\FRAME_MATCHER.state [6]), .I1(n10_adj_4629), 
            .I2(GND_net), .I3(GND_net), .O(n43134));
    defparam i1_2_lut_adj_1051.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut_adj_1052 (.I0(Kp_23__N_1059), .I1(n44094), .I2(n44052), 
            .I3(\data_in_frame[7] [7]), .O(n44243));   // verilog/coms.v(79[16:27])
    defparam i1_4_lut_adj_1052.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1053 (.I0(\FRAME_MATCHER.state [7]), .I1(n10_adj_4629), 
            .I2(GND_net), .I3(GND_net), .O(n43132));
    defparam i1_2_lut_adj_1053.LUT_INIT = 16'h8888;
    SB_LUT4 select_686_Select_23_i3_2_lut (.I0(\FRAME_MATCHER.i [23]), .I1(n4141), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4638));
    defparam select_686_Select_23_i3_2_lut.LUT_INIT = 16'h8888;
    SB_DFF IntegralLimit_i0_i2 (.Q(IntegralLimit[2]), .C(CLK_c), .D(n29157));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i1_4_lut_adj_1054 (.I0(n44243), .I1(n44361), .I2(n27554), 
            .I3(\data_in_frame[10] [2]), .O(n40638));
    defparam i1_4_lut_adj_1054.LUT_INIT = 16'h6996;
    SB_CARRY add_43_25 (.CI(n38576), .I0(\FRAME_MATCHER.i [23]), .I1(GND_net), 
            .CO(n38577));
    SB_LUT4 i1_2_lut_adj_1055 (.I0(\FRAME_MATCHER.state [8]), .I1(n10_adj_4629), 
            .I2(GND_net), .I3(GND_net), .O(n43130));
    defparam i1_2_lut_adj_1055.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1056 (.I0(\data_in_frame[12] [2]), .I1(\data_in_frame[12] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n44214));
    defparam i1_2_lut_adj_1056.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1057 (.I0(\FRAME_MATCHER.state [9]), .I1(n10_adj_4629), 
            .I2(GND_net), .I3(GND_net), .O(n43128));
    defparam i1_2_lut_adj_1057.LUT_INIT = 16'h8888;
    SB_LUT4 select_686_Select_24_i3_2_lut (.I0(\FRAME_MATCHER.i [24]), .I1(n4141), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4639));
    defparam select_686_Select_24_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_686_Select_25_i3_2_lut (.I0(\FRAME_MATCHER.i [25]), .I1(n4141), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4640));
    defparam select_686_Select_25_i3_2_lut.LUT_INIT = 16'h8888;
    SB_DFF IntegralLimit_i0_i3 (.Q(IntegralLimit[3]), .C(CLK_c), .D(n29156));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 select_686_Select_26_i3_2_lut (.I0(\FRAME_MATCHER.i [26]), .I1(n4141), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4641));
    defparam select_686_Select_26_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1058 (.I0(\FRAME_MATCHER.state [10]), .I1(n10_adj_4629), 
            .I2(GND_net), .I3(GND_net), .O(n43126));
    defparam i1_2_lut_adj_1058.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1059 (.I0(\FRAME_MATCHER.state [11]), .I1(n10_adj_4629), 
            .I2(GND_net), .I3(GND_net), .O(n43124));
    defparam i1_2_lut_adj_1059.LUT_INIT = 16'h8888;
    SB_LUT4 select_686_Select_27_i3_2_lut (.I0(\FRAME_MATCHER.i [27]), .I1(n4141), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4642));
    defparam select_686_Select_27_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_686_Select_28_i3_2_lut (.I0(\FRAME_MATCHER.i [28]), .I1(n4141), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4643));
    defparam select_686_Select_28_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_686_Select_29_i3_2_lut (.I0(\FRAME_MATCHER.i [29]), .I1(n4141), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4644));
    defparam select_686_Select_29_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1060 (.I0(\FRAME_MATCHER.state [12]), .I1(n10_adj_4629), 
            .I2(GND_net), .I3(GND_net), .O(n43122));
    defparam i1_2_lut_adj_1060.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1061 (.I0(\FRAME_MATCHER.state [13]), .I1(n10_adj_4629), 
            .I2(GND_net), .I3(GND_net), .O(n43120));
    defparam i1_2_lut_adj_1061.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1062 (.I0(\FRAME_MATCHER.state [13]), .I1(n5), 
            .I2(GND_net), .I3(GND_net), .O(n43172));
    defparam i1_2_lut_adj_1062.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1063 (.I0(\FRAME_MATCHER.state [14]), .I1(n10_adj_4629), 
            .I2(GND_net), .I3(GND_net), .O(n43118));
    defparam i1_2_lut_adj_1063.LUT_INIT = 16'h8888;
    SB_LUT4 i15481_3_lut_4_lut (.I0(n8_adj_4645), .I1(n43832), .I2(rx_data[7]), 
            .I3(\data_in_frame[1] [7]), .O(n29429));
    defparam i15481_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1064 (.I0(\FRAME_MATCHER.state [14]), .I1(n5), 
            .I2(GND_net), .I3(GND_net), .O(n43178));
    defparam i1_2_lut_adj_1064.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1065 (.I0(\FRAME_MATCHER.state [15]), .I1(n10_adj_4629), 
            .I2(GND_net), .I3(GND_net), .O(n43116));
    defparam i1_2_lut_adj_1065.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1066 (.I0(\FRAME_MATCHER.state [15]), .I1(n5), 
            .I2(GND_net), .I3(GND_net), .O(n43180));
    defparam i1_2_lut_adj_1066.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut_adj_1067 (.I0(n52_adj_4626), .I1(n4452), .I2(n27231), 
            .I3(n27061), .O(n5));
    defparam i1_4_lut_adj_1067.LUT_INIT = 16'habaa;
    SB_LUT4 i1_2_lut_adj_1068 (.I0(\FRAME_MATCHER.state [16]), .I1(n10_adj_4629), 
            .I2(GND_net), .I3(GND_net), .O(n43114));
    defparam i1_2_lut_adj_1068.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1069 (.I0(\FRAME_MATCHER.state [16]), .I1(n5), 
            .I2(GND_net), .I3(GND_net), .O(n43182));
    defparam i1_2_lut_adj_1069.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1070 (.I0(\FRAME_MATCHER.state [17]), .I1(n10_adj_4629), 
            .I2(GND_net), .I3(GND_net), .O(n43112));
    defparam i1_2_lut_adj_1070.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1071 (.I0(\FRAME_MATCHER.state [18]), .I1(n10_adj_4629), 
            .I2(GND_net), .I3(GND_net), .O(n43110));
    defparam i1_2_lut_adj_1071.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1072 (.I0(\FRAME_MATCHER.state [19]), .I1(n10_adj_4629), 
            .I2(GND_net), .I3(GND_net), .O(n43108));
    defparam i1_2_lut_adj_1072.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1073 (.I0(\FRAME_MATCHER.state [20]), .I1(n10_adj_4629), 
            .I2(GND_net), .I3(GND_net), .O(n43106));
    defparam i1_2_lut_adj_1073.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1074 (.I0(\FRAME_MATCHER.state [21]), .I1(n10_adj_4629), 
            .I2(GND_net), .I3(GND_net), .O(n43104));
    defparam i1_2_lut_adj_1074.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut_adj_1075 (.I0(n44_adj_4646), .I1(\FRAME_MATCHER.state [1]), 
            .I2(n4_adj_4647), .I3(n43795), .O(n10_adj_4629));
    defparam i1_4_lut_adj_1075.LUT_INIT = 16'hbbba;
    SB_LUT4 i1_2_lut_adj_1076 (.I0(\FRAME_MATCHER.state [22]), .I1(n10_adj_4629), 
            .I2(GND_net), .I3(GND_net), .O(n43102));
    defparam i1_2_lut_adj_1076.LUT_INIT = 16'h8888;
    SB_LUT4 i15482_3_lut_4_lut (.I0(n8_adj_4645), .I1(n43832), .I2(rx_data[6]), 
            .I3(\data_in_frame[1] [6]), .O(n29430));
    defparam i15482_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1077 (.I0(\FRAME_MATCHER.state [24]), .I1(n10_adj_4648), 
            .I2(GND_net), .I3(GND_net), .O(n43098));
    defparam i1_2_lut_adj_1077.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1078 (.I0(\FRAME_MATCHER.state [25]), .I1(n10_adj_4648), 
            .I2(GND_net), .I3(GND_net), .O(n43096));
    defparam i1_2_lut_adj_1078.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1079 (.I0(\FRAME_MATCHER.state [26]), .I1(n10_adj_4648), 
            .I2(GND_net), .I3(GND_net), .O(n43094));
    defparam i1_2_lut_adj_1079.LUT_INIT = 16'h8888;
    SB_LUT4 i21294_2_lut (.I0(\FRAME_MATCHER.state [27]), .I1(n40252), .I2(GND_net), 
            .I3(GND_net), .O(n35234));
    defparam i21294_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1080 (.I0(\FRAME_MATCHER.state [28]), .I1(n10_adj_4648), 
            .I2(GND_net), .I3(GND_net), .O(n43092));
    defparam i1_2_lut_adj_1080.LUT_INIT = 16'h8888;
    SB_DFF IntegralLimit_i0_i4 (.Q(IntegralLimit[4]), .C(CLK_c), .D(n29155));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i2_4_lut_adj_1081 (.I0(n48_adj_4649), .I1(n24234), .I2(n44_adj_4646), 
            .I3(n55), .O(n40252));
    defparam i2_4_lut_adj_1081.LUT_INIT = 16'hfafe;
    SB_LUT4 i15483_3_lut_4_lut (.I0(n8_adj_4645), .I1(n43832), .I2(rx_data[5]), 
            .I3(\data_in_frame[1] [5]), .O(n29431));
    defparam i15483_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1082 (.I0(\data_in_frame[1] [2]), .I1(\data_in_frame[1] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n27454));   // verilog/coms.v(74[16:34])
    defparam i1_2_lut_adj_1082.LUT_INIT = 16'h6666;
    SB_LUT4 i21295_2_lut (.I0(\FRAME_MATCHER.state [29]), .I1(n40252), .I2(GND_net), 
            .I3(GND_net), .O(n35236));
    defparam i21295_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i15484_3_lut_4_lut (.I0(n8_adj_4645), .I1(n43832), .I2(rx_data[4]), 
            .I3(\data_in_frame[1] [4]), .O(n29432));
    defparam i15484_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1083 (.I0(n22132), .I1(n4120), .I2(GND_net), 
            .I3(GND_net), .O(n44_adj_4646));   // verilog/coms.v(260[6] 262[9])
    defparam i1_2_lut_adj_1083.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut_adj_1084 (.I0(n44_adj_4646), .I1(\FRAME_MATCHER.state [1]), 
            .I2(n43729), .I3(n4_adj_4647), .O(n10_adj_4648));
    defparam i1_4_lut_adj_1084.LUT_INIT = 16'hbbba;
    SB_LUT4 i1_2_lut_adj_1085 (.I0(\FRAME_MATCHER.state [30]), .I1(n10_adj_4648), 
            .I2(GND_net), .I3(GND_net), .O(n43088));
    defparam i1_2_lut_adj_1085.LUT_INIT = 16'h8888;
    SB_LUT4 i15485_3_lut_4_lut (.I0(n8_adj_4645), .I1(n43832), .I2(rx_data[3]), 
            .I3(\data_in_frame[1] [3]), .O(n29433));
    defparam i15485_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_adj_1086 (.I0(n41814), .I1(n44214), .I2(\data_in_frame[14] [4]), 
            .I3(GND_net), .O(n40745));
    defparam i2_3_lut_adj_1086.LUT_INIT = 16'h6969;
    SB_LUT4 i1_2_lut_adj_1087 (.I0(n26199), .I1(\data_in_frame[2] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n27730));
    defparam i1_2_lut_adj_1087.LUT_INIT = 16'h6666;
    SB_LUT4 select_686_Select_30_i3_2_lut (.I0(\FRAME_MATCHER.i [30]), .I1(n4141), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4650));
    defparam select_686_Select_30_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_686_Select_31_i3_2_lut (.I0(\FRAME_MATCHER.i [31]), .I1(n4141), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4651));
    defparam select_686_Select_31_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i15486_3_lut_4_lut (.I0(n8_adj_4645), .I1(n43832), .I2(rx_data[2]), 
            .I3(\data_in_frame[1] [2]), .O(n29434));
    defparam i15486_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15487_3_lut_4_lut (.I0(n8_adj_4645), .I1(n43832), .I2(rx_data[1]), 
            .I3(\data_in_frame[1] [1]), .O(n29435));
    defparam i15487_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i32527_3_lut (.I0(\data_out_frame[22] [4]), .I1(\data_out_frame[23] [4]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n48114));
    defparam i32527_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i32526_3_lut (.I0(\data_out_frame[20] [4]), .I1(\data_out_frame[21] [4]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n48113));
    defparam i32526_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFSR tx_transmit_4011 (.Q(r_SM_Main_2__N_3780[0]), .C(CLK_c), .D(n5403[0]), 
            .R(n44813));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i1_4_lut_adj_1088 (.I0(n33827), .I1(\FRAME_MATCHER.state [2]), 
            .I2(n63_adj_4652), .I3(n63_adj_4653), .O(\FRAME_MATCHER.state_31__N_2808 [2]));   // verilog/coms.v(96[12:19])
    defparam i1_4_lut_adj_1088.LUT_INIT = 16'h8a0a;
    SB_LUT4 i20710_2_lut (.I0(\FRAME_MATCHER.state_31__N_2808 [2]), .I1(n4452), 
            .I2(GND_net), .I3(GND_net), .O(\FRAME_MATCHER.state_31__N_2968 [2]));   // verilog/coms.v(260[6] 262[9])
    defparam i20710_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i2_4_lut_adj_1089 (.I0(\FRAME_MATCHER.state_31__N_2808 [2]), .I1(n3303), 
            .I2(n43859), .I3(n55), .O(n6_adj_4654));   // verilog/coms.v(202[5:24])
    defparam i2_4_lut_adj_1089.LUT_INIT = 16'ha0ee;
    SB_LUT4 i3_4_lut_adj_1090 (.I0(n63), .I1(n6_adj_4654), .I2(n27231), 
            .I3(\FRAME_MATCHER.state_31__N_2968 [2]), .O(n51605));   // verilog/coms.v(202[5:24])
    defparam i3_4_lut_adj_1090.LUT_INIT = 16'hdfdd;
    SB_LUT4 i1_2_lut_adj_1091 (.I0(n26673), .I1(n41715), .I2(GND_net), 
            .I3(GND_net), .O(n44367));   // verilog/coms.v(79[16:27])
    defparam i1_2_lut_adj_1091.LUT_INIT = 16'h9999;
    SB_LUT4 i1_3_lut_adj_1092 (.I0(\data_in_frame[16] [1]), .I1(\data_in_frame[13] [6]), 
            .I2(\data_in_frame[16] [4]), .I3(GND_net), .O(n47429));
    defparam i1_3_lut_adj_1092.LUT_INIT = 16'h9696;
    SB_LUT4 i1_4_lut_adj_1093 (.I0(n47429), .I1(n44479), .I2(\data_in_frame[17] [1]), 
            .I3(\data_in_frame[14] [5]), .O(n47433));
    defparam i1_4_lut_adj_1093.LUT_INIT = 16'h6996;
    SB_LUT4 i15488_3_lut_4_lut (.I0(n8_adj_4645), .I1(n43832), .I2(rx_data[0]), 
            .I3(\data_in_frame[1] [0]), .O(n29436));
    defparam i15488_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_4_lut_adj_1094 (.I0(n41760), .I1(n43954), .I2(n44507), 
            .I3(n47433), .O(n47439));
    defparam i1_4_lut_adj_1094.LUT_INIT = 16'h9669;
    SB_LUT4 i1_4_lut_adj_1095 (.I0(n40745), .I1(n44403), .I2(n47439), 
            .I3(n28011), .O(n47445));
    defparam i1_4_lut_adj_1095.LUT_INIT = 16'h9669;
    SB_LUT4 i1_4_lut_adj_1096 (.I0(n41651), .I1(n41606), .I2(n41725), 
            .I3(n47445), .O(n47451));
    defparam i1_4_lut_adj_1096.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1097 (.I0(Kp_23__N_1811), .I1(n44599), .I2(n45643), 
            .I3(n47451), .O(n26673));
    defparam i1_4_lut_adj_1097.LUT_INIT = 16'h9669;
    SB_LUT4 i1_3_lut_adj_1098 (.I0(\data_in_frame[16] [5]), .I1(n40745), 
            .I2(n44465), .I3(GND_net), .O(n41058));
    defparam i1_3_lut_adj_1098.LUT_INIT = 16'h9696;
    SB_LUT4 i1_4_lut_adj_1099 (.I0(n44129), .I1(n44370), .I2(n41058), 
            .I3(n43992), .O(n41715));
    defparam i1_4_lut_adj_1099.LUT_INIT = 16'h9669;
    SB_LUT4 i1_4_lut_adj_1100 (.I0(n40684), .I1(n26673), .I2(n40734), 
            .I3(\data_in_frame[18] [0]), .O(n44370));
    defparam i1_4_lut_adj_1100.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1101 (.I0(\data_in_frame[17] [3]), .I1(\data_in_frame[15] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n47315));
    defparam i1_2_lut_adj_1101.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1102 (.I0(n44284), .I1(n46393), .I2(n44534), 
            .I3(n47315), .O(n44599));
    defparam i1_4_lut_adj_1102.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1103 (.I0(\data_in_frame[20] [6]), .I1(\data_in_frame[20] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n47211));
    defparam i1_2_lut_adj_1103.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1104 (.I0(\data_in_frame[13] [0]), .I1(\data_in_frame[10] [6]), 
            .I2(\data_in_frame[21] [7]), .I3(\data_in_frame[21] [1]), .O(n47223));
    defparam i1_4_lut_adj_1104.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1105 (.I0(\data_in_frame[9] [0]), .I1(\data_in_frame[11] [1]), 
            .I2(\data_in_frame[20] [5]), .I3(\data_in_frame[19] [2]), .O(n47225));
    defparam i1_4_lut_adj_1105.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1106 (.I0(\data_in_frame[21] [4]), .I1(\data_in_frame[21] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n43923));
    defparam i1_2_lut_adj_1106.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1107 (.I0(\data_in_frame[21] [6]), .I1(\data_in_frame[20] [3]), 
            .I2(\data_in_frame[21] [5]), .I3(\data_in_frame[20] [4]), .O(n47233));
    defparam i1_4_lut_adj_1107.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1108 (.I0(n44614), .I1(n44122), .I2(n43923), 
            .I3(n47225), .O(n47237));
    defparam i1_4_lut_adj_1108.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1109 (.I0(n47223), .I1(n44338), .I2(n47211), 
            .I3(\data_in_frame[13] [7]), .O(n47235));
    defparam i1_4_lut_adj_1109.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1110 (.I0(\data_in_frame[4] [7]), .I1(n44376), 
            .I2(GND_net), .I3(GND_net), .O(n43951));   // verilog/coms.v(86[17:70])
    defparam i1_2_lut_adj_1110.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1111 (.I0(n44488), .I1(n47235), .I2(n47237), 
            .I3(n47233), .O(n47243));
    defparam i1_4_lut_adj_1111.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1112 (.I0(n44038), .I1(n44347), .I2(n44574), 
            .I3(n47243), .O(n47249));
    defparam i1_4_lut_adj_1112.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1113 (.I0(\data_in_frame[16] [5]), .I1(n44161), 
            .I2(n44620), .I3(n47249), .O(n47257));
    defparam i1_4_lut_adj_1113.LUT_INIT = 16'h6996;
    SB_LUT4 i32532_3_lut (.I0(\data_out_frame[16] [3]), .I1(\data_out_frame[17] [3]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n48119));
    defparam i32532_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_1114 (.I0(\data_in_frame[3] [1]), .I1(\data_in_frame[5] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n44341));   // verilog/coms.v(86[17:70])
    defparam i1_2_lut_adj_1114.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1115 (.I0(n44237), .I1(n47257), .I2(n46024), 
            .I3(n46118), .O(n47263));
    defparam i1_4_lut_adj_1115.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1116 (.I0(n44462), .I1(n44331), .I2(\data_in_frame[19] [7]), 
            .I3(\data_in_frame[19] [6]), .O(n47285));
    defparam i1_4_lut_adj_1116.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1117 (.I0(Kp_23__N_1811), .I1(n44272), .I2(n44450), 
            .I3(n47285), .O(n47291));
    defparam i1_4_lut_adj_1117.LUT_INIT = 16'h6996;
    SB_LUT4 i32533_3_lut (.I0(\data_out_frame[18] [3]), .I1(\data_out_frame[19] [3]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n48120));
    defparam i32533_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1118 (.I0(n44599), .I1(n44199), .I2(n44065), 
            .I3(n47263), .O(n47269));
    defparam i1_4_lut_adj_1118.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1119 (.I0(n44196), .I1(\data_in_frame[19] [3]), 
            .I2(n47291), .I3(n41769), .O(n47295));
    defparam i1_4_lut_adj_1119.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1120 (.I0(n44370), .I1(n47295), .I2(n47269), 
            .I3(n41715), .O(n45675));
    defparam i1_4_lut_adj_1120.LUT_INIT = 16'h9669;
    SB_LUT4 i3_4_lut_adj_1121 (.I0(\data_in_frame[18] [5]), .I1(\data_in_frame[20] [1]), 
            .I2(n27861), .I3(\data_in_frame[20] [2]), .O(n44199));
    defparam i3_4_lut_adj_1121.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1122 (.I0(\data_in_frame[18] [3]), .I1(n45694), 
            .I2(GND_net), .I3(GND_net), .O(n44531));
    defparam i1_2_lut_adj_1122.LUT_INIT = 16'h9999;
    SB_LUT4 i1_2_lut_adj_1123 (.I0(\data_in_frame[15] [5]), .I1(\data_in_frame[20] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n44122));
    defparam i1_2_lut_adj_1123.LUT_INIT = 16'h6666;
    SB_LUT4 i2_4_lut_adj_1124 (.I0(n40653), .I1(n40755), .I2(n44122), 
            .I3(\data_in_frame[17] [6]), .O(n44155));
    defparam i2_4_lut_adj_1124.LUT_INIT = 16'h6996;
    SB_LUT4 i1_3_lut_adj_1125 (.I0(n27668), .I1(n46393), .I2(\data_in_frame[19] [4]), 
            .I3(GND_net), .O(n45887));
    defparam i1_3_lut_adj_1125.LUT_INIT = 16'h6969;
    SB_LUT4 i32560_3_lut (.I0(\data_out_frame[22] [3]), .I1(\data_out_frame[23] [3]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n48147));
    defparam i32560_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i32559_3_lut (.I0(\data_out_frame[20] [3]), .I1(\data_out_frame[21] [3]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n48146));
    defparam i32559_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut_adj_1126 (.I0(\data_in_frame[5] [7]), .I1(\data_in_frame[1] [4]), 
            .I2(\data_in_frame[5] [6]), .I3(GND_net), .O(n43899));   // verilog/coms.v(74[16:42])
    defparam i1_3_lut_adj_1126.LUT_INIT = 16'h9696;
    SB_DFF \FRAME_MATCHER.rx_data_ready_prev_4012  (.Q(\FRAME_MATCHER.rx_data_ready_prev ), 
           .C(CLK_c), .D(rx_data_ready));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i1_3_lut_adj_1127 (.I0(n46024), .I1(n27668), .I2(\data_in_frame[19] [5]), 
            .I3(GND_net), .O(n44272));
    defparam i1_3_lut_adj_1127.LUT_INIT = 16'h6969;
    SB_LUT4 i1_4_lut_adj_1128 (.I0(n41618), .I1(n47851), .I2(n27536), 
            .I3(n45300), .O(n47611));
    defparam i1_4_lut_adj_1128.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1129 (.I0(\data_in_frame[17] [3]), .I1(n45643), 
            .I2(n40653), .I3(n47611), .O(n27668));
    defparam i1_4_lut_adj_1129.LUT_INIT = 16'h6996;
    SB_LUT4 i15407_3_lut_4_lut (.I0(n8_adj_4655), .I1(n43841), .I2(rx_data[0]), 
            .I3(\data_in_frame[11] [0]), .O(n29355));
    defparam i15407_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i32505_3_lut (.I0(\data_out_frame[16] [2]), .I1(\data_out_frame[17] [2]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n48092));
    defparam i32505_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_1130 (.I0(\data_in_frame[17] [7]), .I1(\data_in_frame[17] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n44614));
    defparam i1_2_lut_adj_1130.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1131 (.I0(\data_in_frame[13] [5]), .I1(Kp_23__N_1465), 
            .I2(Kp_23__N_1468), .I3(n27513), .O(n27536));   // verilog/coms.v(76[16:43])
    defparam i3_4_lut_adj_1131.LUT_INIT = 16'h6996;
    SB_LUT4 i15331_3_lut_4_lut (.I0(n8_adj_4655), .I1(n43820), .I2(rx_data[7]), 
            .I3(\data_in_frame[19] [7]), .O(n29279));
    defparam i15331_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFFE setpoint__i0 (.Q(setpoint[0]), .C(CLK_c), .E(n28531), .D(n7570));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 add_43_24_lut (.I0(n3345), .I1(\FRAME_MATCHER.i [22]), .I2(GND_net), 
            .I3(n38575), .O(n2_adj_4656)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_24_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_2_lut_adj_1132 (.I0(\data_in_frame[18] [0]), .I1(n27536), 
            .I2(GND_net), .I3(GND_net), .O(n44347));   // verilog/coms.v(71[16:27])
    defparam i1_2_lut_adj_1132.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1133 (.I0(\data_in_frame[3] [6]), .I1(\data_in_frame[6] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n28033));   // verilog/coms.v(77[16:43])
    defparam i1_2_lut_adj_1133.LUT_INIT = 16'h6666;
    SB_LUT4 i32506_3_lut (.I0(\data_out_frame[18] [2]), .I1(\data_out_frame[19] [2]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n48093));
    defparam i32506_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i33827_2_lut (.I0(n51489), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n49352));
    defparam i33827_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1_4_lut_adj_1134 (.I0(n28033), .I1(n27590), .I2(n43899), 
            .I3(\data_in_frame[1] [5]), .O(n28288));
    defparam i1_4_lut_adj_1134.LUT_INIT = 16'h6996;
    SB_DFF IntegralLimit_i0_i5 (.Q(IntegralLimit[5]), .C(CLK_c), .D(n29153));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i1_4_lut_adj_1135 (.I0(n27475), .I1(n44006), .I2(n27420), 
            .I3(n28033), .O(n27457));   // verilog/coms.v(76[16:27])
    defparam i1_4_lut_adj_1135.LUT_INIT = 16'h6996;
    SB_LUT4 i32596_3_lut (.I0(\data_out_frame[22] [2]), .I1(\data_out_frame[23] [2]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n48183));
    defparam i32596_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_43_24 (.CI(n38575), .I0(\FRAME_MATCHER.i [22]), .I1(GND_net), 
            .CO(n38576));
    SB_LUT4 i2_4_lut_adj_1136 (.I0(\data_in_frame[16] [7]), .I1(n40638), 
            .I2(\data_in_frame[14] [6]), .I3(n4_adj_4657), .O(n43957));   // verilog/coms.v(79[16:27])
    defparam i2_4_lut_adj_1136.LUT_INIT = 16'h9669;
    SB_LUT4 i32595_3_lut (.I0(\data_out_frame[20] [2]), .I1(\data_out_frame[21] [2]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n48182));
    defparam i32595_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4_4_lut_adj_1137 (.I0(n40755), .I1(Kp_23__N_1561), .I2(n43954), 
            .I3(n6_adj_4658), .O(n41303));   // verilog/coms.v(71[16:27])
    defparam i4_4_lut_adj_1137.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1138 (.I0(\data_in_frame[14] [6]), .I1(n40638), 
            .I2(GND_net), .I3(GND_net), .O(n44534));
    defparam i1_2_lut_adj_1138.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1139 (.I0(\data_in_frame[11] [2]), .I1(\data_in_frame[11] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n47459));
    defparam i1_2_lut_adj_1139.LUT_INIT = 16'h6666;
    SB_LUT4 i32502_3_lut (.I0(\data_out_frame[16] [0]), .I1(\data_out_frame[17] [0]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n48089));
    defparam i32502_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i32503_3_lut (.I0(\data_out_frame[18] [0]), .I1(\data_out_frame[19] [0]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n48090));
    defparam i32503_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i32509_3_lut (.I0(\data_out_frame[22] [0]), .I1(\data_out_frame[23] [0]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n48096));
    defparam i32509_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_35849 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [4]), .I2(\data_out_frame[27] [4]), 
            .I3(byte_transmit_counter[1]), .O(n51480));
    defparam byte_transmit_counter_0__bdd_4_lut_35849.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_4_lut_adj_1140 (.I0(n27976), .I1(n45643), .I2(n27820), 
            .I3(n47459), .O(n44237));
    defparam i1_4_lut_adj_1140.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1141 (.I0(n27457), .I1(n28288), .I2(GND_net), 
            .I3(GND_net), .O(n44245));
    defparam i1_2_lut_adj_1141.LUT_INIT = 16'h6666;
    SB_LUT4 i32508_3_lut (.I0(\data_out_frame[20] [0]), .I1(\data_out_frame[21] [0]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n48095));
    defparam i32508_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1142 (.I0(n44341), .I1(\data_in_frame[5] [2]), 
            .I2(\data_in_frame[0] [7]), .I3(\data_in_frame[7] [3]), .O(n47621));   // verilog/coms.v(72[16:69])
    defparam i1_4_lut_adj_1142.LUT_INIT = 16'h6996;
    SB_LUT4 i15332_3_lut_4_lut (.I0(n8_adj_4655), .I1(n43820), .I2(rx_data[6]), 
            .I3(\data_in_frame[19] [6]), .O(n29280));
    defparam i15332_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_4_lut_adj_1143 (.I0(n43951), .I1(n27730), .I2(Kp_23__N_1027), 
            .I3(n47621), .O(n40728));   // verilog/coms.v(72[16:69])
    defparam i1_4_lut_adj_1143.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1144 (.I0(\data_in_frame[10] [5]), .I1(n27506), 
            .I2(GND_net), .I3(GND_net), .O(n44397));
    defparam i1_2_lut_adj_1144.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1145 (.I0(\data_in_frame[17] [2]), .I1(\data_in_frame[15] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n47297));
    defparam i1_2_lut_adj_1145.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1146 (.I0(n44596), .I1(\data_in_frame[10] [4]), 
            .I2(n47297), .I3(\data_in_frame[12] [6]), .O(n47303));
    defparam i1_4_lut_adj_1146.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1147 (.I0(n44397), .I1(n44602), .I2(n44538), 
            .I3(\data_in_frame[11] [4]), .O(n47417));
    defparam i1_4_lut_adj_1147.LUT_INIT = 16'h6996;
    SB_DFF IntegralLimit_i0_i6 (.Q(IntegralLimit[6]), .C(CLK_c), .D(n29151));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i1_4_lut_adj_1148 (.I0(n44023), .I1(n44397), .I2(n4_adj_4659), 
            .I3(n47303), .O(n47309));
    defparam i1_4_lut_adj_1148.LUT_INIT = 16'h6996;
    SB_DFF data_out_frame_0___i106 (.Q(\data_out_frame[13] [1]), .C(CLK_c), 
           .D(n29018));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i32643_3_lut (.I0(\data_out_frame[8] [7]), .I1(\data_out_frame[9] [7]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n48230));
    defparam i32643_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i32644_3_lut (.I0(\data_out_frame[10] [7]), .I1(\data_out_frame[11] [7]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n48231));
    defparam i32644_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF IntegralLimit_i0_i7 (.Q(IntegralLimit[7]), .C(CLK_c), .D(n29150));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i1_4_lut_adj_1149 (.I0(n44237), .I1(n41059), .I2(Kp_23__N_1468), 
            .I3(n47417), .O(n47423));
    defparam i1_4_lut_adj_1149.LUT_INIT = 16'h6996;
    SB_LUT4 i32482_3_lut (.I0(\data_out_frame[14] [7]), .I1(\data_out_frame[15] [7]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n48069));
    defparam i32482_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i32481_3_lut (.I0(\data_out_frame[12] [7]), .I1(\data_out_frame[13] [7]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n48068));
    defparam i32481_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i32499_3_lut (.I0(\data_out_frame[8] [0]), .I1(\data_out_frame[9] [0]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n48086));
    defparam i32499_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i32500_3_lut (.I0(\data_out_frame[10] [0]), .I1(\data_out_frame[11] [0]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n48087));
    defparam i32500_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i32611_3_lut (.I0(\data_out_frame[14] [0]), .I1(\data_out_frame[15] [0]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n48198));
    defparam i32611_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i32610_3_lut (.I0(\data_out_frame[12] [0]), .I1(\data_out_frame[13] [0]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n48197));
    defparam i32610_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF IntegralLimit_i0_i8 (.Q(IntegralLimit[8]), .C(CLK_c), .D(n29149));   // verilog/coms.v(128[12] 303[6])
    SB_DFF IntegralLimit_i0_i9 (.Q(IntegralLimit[9]), .C(CLK_c), .D(n29148));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i1_4_lut_adj_1150 (.I0(n44534), .I1(n47423), .I2(n47309), 
            .I3(n41793), .O(n46393));
    defparam i1_4_lut_adj_1150.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1151 (.I0(n46393), .I1(n44217), .I2(GND_net), 
            .I3(GND_net), .O(n41769));
    defparam i1_2_lut_adj_1151.LUT_INIT = 16'h9999;
    SB_DFF IntegralLimit_i0_i10 (.Q(IntegralLimit[10]), .C(CLK_c), .D(n29147));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i2_2_lut (.I0(\data_in_frame[12] [2]), .I1(\data_in_frame[11] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n10_adj_4660));
    defparam i2_2_lut.LUT_INIT = 16'h6666;
    SB_DFF IntegralLimit_i0_i11 (.Q(IntegralLimit[11]), .C(CLK_c), .D(n29145));   // verilog/coms.v(128[12] 303[6])
    SB_DFF IntegralLimit_i0_i12 (.Q(IntegralLimit[12]), .C(CLK_c), .D(n29144));   // verilog/coms.v(128[12] 303[6])
    SB_DFF IntegralLimit_i0_i13 (.Q(IntegralLimit[13]), .C(CLK_c), .D(n29143));   // verilog/coms.v(128[12] 303[6])
    SB_DFF IntegralLimit_i0_i14 (.Q(IntegralLimit[14]), .C(CLK_c), .D(n29142));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i1_2_lut_adj_1152 (.I0(\data_in_frame[13] [2]), .I1(\data_in_frame[13] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n47509));
    defparam i1_2_lut_adj_1152.LUT_INIT = 16'h6666;
    SB_LUT4 add_43_23_lut (.I0(n3345), .I1(\FRAME_MATCHER.i [21]), .I2(GND_net), 
            .I3(n38574), .O(n2_adj_4661)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_23_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_4_lut_adj_1153 (.I0(n27520), .I1(n44161), .I2(Kp_23__N_1531), 
            .I3(n47509), .O(n41059));
    defparam i1_4_lut_adj_1153.LUT_INIT = 16'h6996;
    SB_DFF IntegralLimit_i0_i15 (.Q(IntegralLimit[15]), .C(CLK_c), .D(n29141));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i1_2_lut_adj_1154 (.I0(\data_in_frame[13] [0]), .I1(n44290), 
            .I2(GND_net), .I3(GND_net), .O(n28011));
    defparam i1_2_lut_adj_1154.LUT_INIT = 16'h6666;
    SB_DFF IntegralLimit_i0_i16 (.Q(IntegralLimit[16]), .C(CLK_c), .D(n29140));   // verilog/coms.v(128[12] 303[6])
    SB_CARRY add_43_23 (.CI(n38574), .I0(\FRAME_MATCHER.i [21]), .I1(GND_net), 
            .CO(n38575));
    SB_DFF IntegralLimit_i0_i17 (.Q(IntegralLimit[17]), .C(CLK_c), .D(n29139));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i6_4_lut_adj_1155 (.I0(n40728), .I1(\data_in_frame[12] [1]), 
            .I2(n44245), .I3(\data_in_frame[10] [1]), .O(n14_adj_4662));
    defparam i6_4_lut_adj_1155.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1156 (.I0(\data_in_frame[14] [3]), .I1(n14_adj_4662), 
            .I2(n10_adj_4660), .I3(n44491), .O(n44183));
    defparam i7_4_lut_adj_1156.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1157 (.I0(\data_in_frame[11] [5]), .I1(n41679), 
            .I2(\data_in_frame[9] [3]), .I3(n6_adj_4663), .O(n41644));
    defparam i4_4_lut_adj_1157.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1158 (.I0(\data_in_frame[15] [5]), .I1(\data_in_frame[16] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n44479));
    defparam i1_2_lut_adj_1158.LUT_INIT = 16'h6666;
    SB_LUT4 add_43_22_lut (.I0(n3345), .I1(\FRAME_MATCHER.i [20]), .I2(GND_net), 
            .I3(n38573), .O(n2_adj_4664)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_22_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i3_4_lut_adj_1159 (.I0(n41644), .I1(n43948), .I2(\data_in_frame[16] [2]), 
            .I3(n41184), .O(n45694));
    defparam i3_4_lut_adj_1159.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1160 (.I0(n45694), .I1(n44479), .I2(n43877), 
            .I3(\data_in_frame[17] [7]), .O(n10_adj_4665));
    defparam i4_4_lut_adj_1160.LUT_INIT = 16'h9669;
    SB_DFF IntegralLimit_i0_i18 (.Q(IntegralLimit[18]), .C(CLK_c), .D(n29137));   // verilog/coms.v(128[12] 303[6])
    SB_DFF IntegralLimit_i0_i19 (.Q(IntegralLimit[19]), .C(CLK_c), .D(n29136));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i15333_3_lut_4_lut (.I0(n8_adj_4655), .I1(n43820), .I2(rx_data[5]), 
            .I3(\data_in_frame[19] [5]), .O(n29281));
    defparam i15333_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF IntegralLimit_i0_i20 (.Q(IntegralLimit[20]), .C(CLK_c), .D(n29135));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i1_2_lut_adj_1161 (.I0(n44183), .I1(n44465), .I2(GND_net), 
            .I3(GND_net), .O(n41762));
    defparam i1_2_lut_adj_1161.LUT_INIT = 16'h6666;
    SB_DFF IntegralLimit_i0_i21 (.Q(IntegralLimit[21]), .C(CLK_c), .D(n29134));   // verilog/coms.v(128[12] 303[6])
    SB_DFF IntegralLimit_i0_i22 (.Q(IntegralLimit[22]), .C(CLK_c), .D(n29133));   // verilog/coms.v(128[12] 303[6])
    SB_DFF IntegralLimit_i0_i23 (.Q(IntegralLimit[23]), .C(CLK_c), .D(n29132));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i33 (.Q(\data_out_frame[4] [0]), .C(CLK_c), 
           .D(n29131));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i34 (.Q(\data_out_frame[4] [1]), .C(CLK_c), 
           .D(n29130));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i15334_3_lut_4_lut (.I0(n8_adj_4655), .I1(n43820), .I2(rx_data[4]), 
            .I3(\data_in_frame[19] [4]), .O(n29282));
    defparam i15334_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i4_4_lut_adj_1162 (.I0(\data_in_frame[19] [1]), .I1(n44350), 
            .I2(\data_in_frame[16] [6]), .I3(n41725), .O(n10_adj_4666));
    defparam i4_4_lut_adj_1162.LUT_INIT = 16'h6996;
    SB_CARRY add_43_22 (.CI(n38573), .I0(\FRAME_MATCHER.i [20]), .I1(GND_net), 
            .CO(n38574));
    SB_LUT4 i32496_3_lut (.I0(\data_out_frame[8] [2]), .I1(\data_out_frame[9] [2]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n48083));
    defparam i32496_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5_3_lut_adj_1163 (.I0(n44183), .I1(n10_adj_4666), .I2(\data_in_frame[16] [5]), 
            .I3(GND_net), .O(n44331));
    defparam i5_3_lut_adj_1163.LUT_INIT = 16'h9696;
    SB_DFF data_out_frame_0___i35 (.Q(\data_out_frame[4] [2]), .C(CLK_c), 
           .D(n29129));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i4_4_lut_adj_1164 (.I0(\data_in_frame[0] [4]), .I1(\data_in_frame[0] [6]), 
            .I2(ID[4]), .I3(ID[6]), .O(n12_adj_4667));   // verilog/coms.v(239[12:32])
    defparam i4_4_lut_adj_1164.LUT_INIT = 16'h7bde;
    SB_LUT4 i32497_3_lut (.I0(\data_out_frame[10] [2]), .I1(\data_out_frame[11] [2]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n48084));
    defparam i32497_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF data_out_frame_0___i36 (.Q(\data_out_frame[4] [3]), .C(CLK_c), 
           .D(n29128));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 add_43_21_lut (.I0(n3345), .I1(\FRAME_MATCHER.i [19]), .I2(GND_net), 
            .I3(n38572), .O(n2_adj_4668)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_21_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_43_21 (.CI(n38572), .I0(\FRAME_MATCHER.i [19]), .I1(GND_net), 
            .CO(n38573));
    SB_LUT4 i1_4_lut_adj_1165 (.I0(\data_in_frame[21] [0]), .I1(n41762), 
            .I2(n8_adj_4669), .I3(n40631), .O(n44168));
    defparam i1_4_lut_adj_1165.LUT_INIT = 16'h6996;
    SB_LUT4 i2_4_lut_adj_1166 (.I0(\data_in_frame[0] [1]), .I1(\data_in_frame[0] [2]), 
            .I2(ID[1]), .I3(ID[2]), .O(n10_adj_4670));   // verilog/coms.v(239[12:32])
    defparam i2_4_lut_adj_1166.LUT_INIT = 16'h7bde;
    SB_LUT4 i2_3_lut_adj_1167 (.I0(n44183), .I1(\data_in_frame[16] [5]), 
            .I2(n40745), .I3(GND_net), .O(n40734));
    defparam i2_3_lut_adj_1167.LUT_INIT = 16'h9696;
    SB_LUT4 i5_4_lut_adj_1168 (.I0(n40728), .I1(n43871), .I2(\data_in_frame[14] [1]), 
            .I3(n41622), .O(n12_adj_4671));
    defparam i5_4_lut_adj_1168.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1169 (.I0(\data_in_frame[13] [7]), .I1(n12_adj_4671), 
            .I2(n44293), .I3(\data_in_frame[11] [5]), .O(n41184));
    defparam i6_4_lut_adj_1169.LUT_INIT = 16'h6996;
    SB_DFF data_out_frame_0___i37 (.Q(\data_out_frame[4] [4]), .C(CLK_c), 
           .D(n29127));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i1_3_lut_adj_1170 (.I0(n41651), .I1(n41762), .I2(\data_in_frame[16] [3]), 
            .I3(GND_net), .O(n44129));
    defparam i1_3_lut_adj_1170.LUT_INIT = 16'h6969;
    SB_LUT4 i15335_3_lut_4_lut (.I0(n8_adj_4655), .I1(n43820), .I2(rx_data[3]), 
            .I3(\data_in_frame[19] [3]), .O(n29283));
    defparam i15335_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1171 (.I0(\data_in_frame[18] [5]), .I1(n44592), 
            .I2(GND_net), .I3(GND_net), .O(n44462));
    defparam i1_2_lut_adj_1171.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1172 (.I0(\data_in_frame[20] [7]), .I1(n40734), 
            .I2(\data_in_frame[18] [7]), .I3(GND_net), .O(n44179));
    defparam i2_3_lut_adj_1172.LUT_INIT = 16'h9696;
    SB_LUT4 i33825_2_lut (.I0(n51477), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n49349));
    defparam i33825_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i2_3_lut_adj_1173 (.I0(n44179), .I1(n44462), .I2(n44129), 
            .I3(GND_net), .O(n41688));
    defparam i2_3_lut_adj_1173.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1174 (.I0(\data_in_frame[18] [2]), .I1(\data_in_frame[18] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n27335));
    defparam i1_2_lut_adj_1174.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1175 (.I0(\data_in_frame[0] [7]), .I1(\data_in_frame[0] [5]), 
            .I2(ID[7]), .I3(ID[5]), .O(n11));   // verilog/coms.v(239[12:32])
    defparam i3_4_lut_adj_1175.LUT_INIT = 16'h7bde;
    SB_LUT4 i1_2_lut_adj_1176 (.I0(\data_in_frame[18] [3]), .I1(\data_in_frame[18] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n44425));
    defparam i1_2_lut_adj_1176.LUT_INIT = 16'h6666;
    SB_LUT4 i32618_4_lut (.I0(\data_out_frame[6] [6]), .I1(byte_transmit_counter[0]), 
            .I2(byte_transmit_counter[2]), .I3(\data_out_frame[7] [6]), 
            .O(n48205));
    defparam i32618_4_lut.LUT_INIT = 16'hec2c;
    SB_LUT4 i32616_3_lut (.I0(\data_out_frame[4] [6]), .I1(\data_out_frame[5] [6]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n48203));
    defparam i32616_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut_adj_1177 (.I0(n27506), .I1(n44562), .I2(\data_in_frame[10] [6]), 
            .I3(GND_net), .O(n41606));
    defparam i1_3_lut_adj_1177.LUT_INIT = 16'h9696;
    SB_LUT4 i1_4_lut_adj_1178 (.I0(\data_in_frame[15] [4]), .I1(\data_in_frame[13] [2]), 
            .I2(n41793), .I3(\data_in_frame[13] [3]), .O(n40755));
    defparam i1_4_lut_adj_1178.LUT_INIT = 16'h9669;
    SB_LUT4 equal_2242_i8_2_lut (.I0(Kp_23__N_1253), .I1(\data_in_frame[8] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n8_adj_4672));   // verilog/coms.v(237[9:81])
    defparam equal_2242_i8_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1179 (.I0(\data_in_frame[12] [7]), .I1(n27979), 
            .I2(GND_net), .I3(GND_net), .O(n44602));
    defparam i1_2_lut_adj_1179.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1180 (.I0(\data_in_frame[0] [0]), .I1(\data_in_frame[0] [3]), 
            .I2(ID[0]), .I3(ID[3]), .O(n9));   // verilog/coms.v(239[12:32])
    defparam i1_4_lut_adj_1180.LUT_INIT = 16'h7bde;
    SB_LUT4 i4_4_lut_adj_1181 (.I0(\data_in_frame[8] [1]), .I1(\data_in_frame[8] [2]), 
            .I2(n44513), .I3(n6_adj_4673), .O(n27574));   // verilog/coms.v(97[12:25])
    defparam i4_4_lut_adj_1181.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1182 (.I0(n27873), .I1(n44562), .I2(n44602), 
            .I3(n47743), .O(n41618));
    defparam i1_4_lut_adj_1182.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1183 (.I0(\data_in_frame[13] [2]), .I1(\data_in_frame[13] [1]), 
            .I2(\data_in_frame[10] [5]), .I3(\data_in_frame[15] [3]), .O(n47519));   // verilog/coms.v(72[16:27])
    defparam i1_4_lut_adj_1183.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1184 (.I0(\data_in_frame[9] [7]), .I1(\data_in_frame[10] [1]), 
            .I2(n40688), .I3(n6_adj_4674), .O(n41760));
    defparam i4_4_lut_adj_1184.LUT_INIT = 16'h6996;
    SB_LUT4 i15336_3_lut_4_lut (.I0(n8_adj_4655), .I1(n43820), .I2(rx_data[2]), 
            .I3(\data_in_frame[19] [2]), .O(n29284));
    defparam i15336_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1185 (.I0(\data_in_frame[12] [4]), .I1(n27574), 
            .I2(GND_net), .I3(GND_net), .O(n44023));
    defparam i1_2_lut_adj_1185.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1186 (.I0(n43877), .I1(n40755), .I2(n27976), 
            .I3(n47523), .O(n44284));   // verilog/coms.v(72[16:27])
    defparam i1_4_lut_adj_1186.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1187 (.I0(\data_in_frame[17] [5]), .I1(n44284), 
            .I2(GND_net), .I3(GND_net), .O(n40684));
    defparam i1_2_lut_adj_1187.LUT_INIT = 16'h6666;
    SB_LUT4 i1_3_lut_adj_1188 (.I0(\data_in_frame[15] [3]), .I1(n41618), 
            .I2(\data_in_frame[17] [4]), .I3(GND_net), .O(n46024));
    defparam i1_3_lut_adj_1188.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1189 (.I0(\data_in_frame[21] [7]), .I1(Kp_23__N_1811), 
            .I2(GND_net), .I3(GND_net), .O(n44035));   // verilog/coms.v(86[17:28])
    defparam i1_2_lut_adj_1189.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1190 (.I0(\data_in_frame[11] [4]), .I1(Kp_23__N_1468), 
            .I2(GND_net), .I3(GND_net), .O(n27526));   // verilog/coms.v(77[16:43])
    defparam i1_2_lut_adj_1190.LUT_INIT = 16'h6666;
    SB_LUT4 data_in_frame_13__7__I_0_2_lut (.I0(\data_in_frame[13] [7]), .I1(\data_in_frame[13] [6]), 
            .I2(GND_net), .I3(GND_net), .O(Kp_23__N_1531));   // verilog/coms.v(86[17:28])
    defparam data_in_frame_13__7__I_0_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1191 (.I0(\data_in_frame[16] [3]), .I1(Kp_23__N_1531), 
            .I2(n43926), .I3(n27526), .O(n44038));   // verilog/coms.v(77[16:43])
    defparam i3_4_lut_adj_1191.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1192 (.I0(n44038), .I1(\data_in_frame[16] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n44403));
    defparam i1_2_lut_adj_1192.LUT_INIT = 16'h6666;
    SB_LUT4 i7_4_lut_adj_1193 (.I0(n9), .I1(n11), .I2(n10_adj_4670), .I3(n12_adj_4667), 
            .O(n24450));   // verilog/coms.v(239[12:32])
    defparam i7_4_lut_adj_1193.LUT_INIT = 16'hfffe;
    SB_LUT4 i15337_3_lut_4_lut (.I0(n8_adj_4655), .I1(n43820), .I2(rx_data[1]), 
            .I3(\data_in_frame[19] [1]), .O(n29285));
    defparam i15337_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 add_43_20_lut (.I0(n3345), .I1(\FRAME_MATCHER.i [18]), .I2(GND_net), 
            .I3(n38571), .O(n2_adj_4675)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_20_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_2_lut_adj_1194 (.I0(\data_in_frame[13] [3]), .I1(\data_in_frame[13] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n27520));   // verilog/coms.v(86[17:63])
    defparam i1_2_lut_adj_1194.LUT_INIT = 16'h6666;
    SB_LUT4 n51480_bdd_4_lut (.I0(n51480), .I1(\data_out_frame[25] [4]), 
            .I2(\data_out_frame[24] [4]), .I3(byte_transmit_counter[1]), 
            .O(n51483));
    defparam n51480_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_adj_1195 (.I0(\data_in_frame[13] [7]), .I1(n41598), 
            .I2(GND_net), .I3(GND_net), .O(n44205));
    defparam i1_2_lut_adj_1195.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1196 (.I0(n46118), .I1(\data_in_frame[16] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n43948));
    defparam i1_2_lut_adj_1196.LUT_INIT = 16'h9999;
    SB_LUT4 i1_3_lut_adj_1197 (.I0(\data_in_frame[12] [0]), .I1(n44528), 
            .I2(\data_in_frame[11] [7]), .I3(GND_net), .O(n43871));
    defparam i1_3_lut_adj_1197.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1198 (.I0(\data_in_frame[11] [1]), .I1(\data_in_frame[11] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n44611));
    defparam i1_2_lut_adj_1198.LUT_INIT = 16'h6666;
    SB_CARRY add_43_20 (.CI(n38571), .I0(\FRAME_MATCHER.i [18]), .I1(GND_net), 
            .CO(n38572));
    SB_LUT4 i32605_3_lut (.I0(\data_out_frame[14] [2]), .I1(\data_out_frame[15] [2]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n48192));
    defparam i32605_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_1199 (.I0(\data_in_frame[11] [3]), .I1(\data_in_frame[11] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n27513));   // verilog/coms.v(76[16:43])
    defparam i1_2_lut_adj_1199.LUT_INIT = 16'h6666;
    SB_LUT4 i32604_3_lut (.I0(\data_out_frame[12] [2]), .I1(\data_out_frame[13] [2]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n48191));
    defparam i32604_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_1200 (.I0(\data_in_frame[10] [6]), .I1(\data_in_frame[12] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n44299));   // verilog/coms.v(72[16:27])
    defparam i1_2_lut_adj_1200.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1201 (.I0(\data_in_frame[6] [2]), .I1(\data_in_frame[7] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n47467));
    defparam i1_2_lut_adj_1201.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1202 (.I0(\data_in_frame[11] [2]), .I1(n47467), 
            .I2(\data_in_frame[10] [4]), .I3(\data_in_frame[10] [1]), .O(n47473));
    defparam i1_4_lut_adj_1202.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1203 (.I0(n44565), .I1(n44617), .I2(n44611), 
            .I3(n44214), .O(n47483));
    defparam i1_4_lut_adj_1203.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1204 (.I0(n44233), .I1(n44299), .I2(n47473), 
            .I3(n27513), .O(n47485));
    defparam i1_4_lut_adj_1204.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1205 (.I0(n47485), .I1(n44516), .I2(n44538), 
            .I3(n47483), .O(n47491));
    defparam i1_4_lut_adj_1205.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1206 (.I0(n44072), .I1(n44589), .I2(n44547), 
            .I3(n47491), .O(n47497));
    defparam i1_4_lut_adj_1206.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1207 (.I0(\data_in_frame[16] [6]), .I1(n43957), 
            .I2(n40745), .I3(GND_net), .O(n41302));   // verilog/coms.v(79[16:27])
    defparam i2_3_lut_adj_1207.LUT_INIT = 16'h9696;
    SB_DFF data_out_frame_0___i38 (.Q(\data_out_frame[4] [5]), .C(CLK_c), 
           .D(n29126));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i1_2_lut_adj_1208 (.I0(n27061), .I1(n3303), .I2(GND_net), 
            .I3(GND_net), .O(n24234));   // verilog/coms.v(96[12:19])
    defparam i1_2_lut_adj_1208.LUT_INIT = 16'h2222;
    SB_LUT4 i5_4_lut_adj_1209 (.I0(\data_in_frame[21] [2]), .I1(n44331), 
            .I2(\data_in_frame[21] [1]), .I3(n41762), .O(n12_adj_4676));
    defparam i5_4_lut_adj_1209.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1210 (.I0(n41302), .I1(\data_in_frame[17] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n41725));
    defparam i1_2_lut_adj_1210.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1211 (.I0(n33840), .I1(n19692), .I2(n62), .I3(GND_net), 
            .O(n22132));   // verilog/coms.v(260[6] 262[9])
    defparam i2_3_lut_adj_1211.LUT_INIT = 16'hc8c8;
    SB_LUT4 add_43_19_lut (.I0(n3345), .I1(\FRAME_MATCHER.i [17]), .I2(GND_net), 
            .I3(n38570), .O(n2_adj_4677)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_19_lut.LUT_INIT = 16'h8228;
    SB_DFF data_out_frame_0___i39 (.Q(\data_out_frame[4] [6]), .C(CLK_c), 
           .D(n29125));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i1_4_lut_adj_1212 (.I0(n40972), .I1(n43871), .I2(Kp_23__N_1327), 
            .I3(n47497), .O(n47503));
    defparam i1_4_lut_adj_1212.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1213 (.I0(n771), .I1(\FRAME_MATCHER.state [1]), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_4678));
    defparam i1_2_lut_adj_1213.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_1214 (.I0(n22132), .I1(n27230), .I2(n4120), .I3(n4_adj_4678), 
            .O(n12_adj_4679));
    defparam i1_4_lut_adj_1214.LUT_INIT = 16'ha0a2;
    SB_LUT4 i1_4_lut_adj_1215 (.I0(\FRAME_MATCHER.state [31]), .I1(\FRAME_MATCHER.state [1]), 
            .I2(n12_adj_4679), .I3(n43729), .O(n43086));
    defparam i1_4_lut_adj_1215.LUT_INIT = 16'ha2a0;
    SB_LUT4 i15338_3_lut_4_lut (.I0(n8_adj_4655), .I1(n43820), .I2(rx_data[0]), 
            .I3(\data_in_frame[19] [0]), .O(n29286));
    defparam i15338_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_CARRY add_43_19 (.CI(n38570), .I0(\FRAME_MATCHER.i [17]), .I1(GND_net), 
            .CO(n38571));
    SB_LUT4 add_43_18_lut (.I0(n3345), .I1(\FRAME_MATCHER.i [16]), .I2(GND_net), 
            .I3(n38569), .O(n2_adj_4680)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_18_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i15323_3_lut_4_lut (.I0(n8_adj_4681), .I1(n43820), .I2(rx_data[7]), 
            .I3(\data_in_frame[20] [7]), .O(n29271));
    defparam i15323_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15324_3_lut_4_lut (.I0(n8_adj_4681), .I1(n43820), .I2(rx_data[6]), 
            .I3(\data_in_frame[20] [6]), .O(n29272));
    defparam i15324_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1216 (.I0(\data_in_frame[9] [1]), .I1(n44574), 
            .I2(GND_net), .I3(GND_net), .O(n44105));   // verilog/coms.v(86[17:63])
    defparam i1_2_lut_adj_1216.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1217 (.I0(\data_in_frame[3] [1]), .I1(\data_in_frame[3] [3]), 
            .I2(\data_in_frame[5] [4]), .I3(\data_in_frame[7] [5]), .O(n47759));   // verilog/coms.v(86[17:63])
    defparam i1_4_lut_adj_1217.LUT_INIT = 16'h6996;
    SB_DFFESR byte_transmit_counter_i0_i0 (.Q(byte_transmit_counter[0]), .C(CLK_c), 
            .E(n28546), .D(n9046[0]), .R(n28996));   // verilog/coms.v(128[12] 303[6])
    SB_CARRY add_43_18 (.CI(n38569), .I0(\FRAME_MATCHER.i [16]), .I1(GND_net), 
            .CO(n38570));
    SB_DFFSS \FRAME_MATCHER.i_i31  (.Q(\FRAME_MATCHER.i [31]), .C(CLK_c), 
            .D(n2_adj_4682), .S(n3_adj_4651));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i15325_3_lut_4_lut (.I0(n8_adj_4681), .I1(n43820), .I2(rx_data[5]), 
            .I3(\data_in_frame[20] [5]), .O(n29273));
    defparam i15325_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15326_3_lut_4_lut (.I0(n8_adj_4681), .I1(n43820), .I2(rx_data[4]), 
            .I3(\data_in_frame[20] [4]), .O(n29274));
    defparam i15326_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_4_lut (.I0(\data_in_frame[11] [3]), .I1(Kp_23__N_1465), 
            .I2(n27520), .I3(n44205), .O(n46118));   // verilog/coms.v(72[16:27])
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_DFFSS \FRAME_MATCHER.i_i30  (.Q(\FRAME_MATCHER.i [30]), .C(CLK_c), 
            .D(n2_adj_4683), .S(n3_adj_4650));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i1_3_lut_adj_1218 (.I0(n27590), .I1(n27350), .I2(\data_in_frame[7] [6]), 
            .I3(GND_net), .O(n27554));
    defparam i1_3_lut_adj_1218.LUT_INIT = 16'h9696;
    SB_LUT4 add_43_17_lut (.I0(n3345), .I1(\FRAME_MATCHER.i [15]), .I2(GND_net), 
            .I3(n38568), .O(n2_adj_4684)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_17_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_43_17 (.CI(n38568), .I0(\FRAME_MATCHER.i [15]), .I1(GND_net), 
            .CO(n38569));
    SB_LUT4 i1_4_lut_adj_1219 (.I0(n28228), .I1(n27730), .I2(n44432), 
            .I3(n44116), .O(n27544));
    defparam i1_4_lut_adj_1219.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1220 (.I0(n27461), .I1(\data_in_frame[5] [1]), 
            .I2(\data_in_frame[2] [7]), .I3(\data_in_frame[7] [2]), .O(n47589));
    defparam i1_4_lut_adj_1220.LUT_INIT = 16'h6996;
    SB_LUT4 i15327_3_lut_4_lut (.I0(n8_adj_4681), .I1(n43820), .I2(rx_data[3]), 
            .I3(\data_in_frame[20] [3]), .O(n29275));
    defparam i15327_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_4_lut_adj_1221 (.I0(n26199), .I1(n44000), .I2(n47589), 
            .I3(n44376), .O(n27850));
    defparam i1_4_lut_adj_1221.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1222 (.I0(n6_adj_4685), .I1(n44391), .I2(n44020), 
            .I3(\data_in_frame[4] [6]), .O(n27820));   // verilog/coms.v(75[16:43])
    defparam i1_4_lut_adj_1222.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_35844 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [3]), .I2(\data_out_frame[27] [3]), 
            .I3(byte_transmit_counter[1]), .O(n51474));
    defparam byte_transmit_counter_0__bdd_4_lut_35844.LUT_INIT = 16'he4aa;
    SB_LUT4 i15328_3_lut_4_lut (.I0(n8_adj_4681), .I1(n43820), .I2(rx_data[2]), 
            .I3(\data_in_frame[20] [2]), .O(n29276));
    defparam i15328_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1223 (.I0(\data_in_frame[6] [7]), .I1(\data_in_frame[6] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n44020));   // verilog/coms.v(75[16:43])
    defparam i1_2_lut_adj_1223.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1224 (.I0(\data_in_frame[4] [5]), .I1(n40678), 
            .I2(GND_net), .I3(GND_net), .O(n44355));   // verilog/coms.v(76[16:43])
    defparam i1_2_lut_adj_1224.LUT_INIT = 16'h6666;
    SB_LUT4 i15329_3_lut_4_lut (.I0(n8_adj_4681), .I1(n43820), .I2(rx_data[1]), 
            .I3(\data_in_frame[20] [1]), .O(n29277));
    defparam i15329_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1225 (.I0(Kp_23__N_1059), .I1(n44094), .I2(GND_net), 
            .I3(GND_net), .O(n44293));
    defparam i1_2_lut_adj_1225.LUT_INIT = 16'h9999;
    SB_LUT4 i1_2_lut_adj_1226 (.I0(n27590), .I1(\data_in_frame[5] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n44102));   // verilog/coms.v(79[16:27])
    defparam i1_2_lut_adj_1226.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1227 (.I0(n44102), .I1(n44293), .I2(Kp_23__N_1103), 
            .I3(\data_in_frame[3] [5]), .O(n40972));   // verilog/coms.v(79[16:27])
    defparam i1_4_lut_adj_1227.LUT_INIT = 16'h6996;
    SB_LUT4 mux_2094_i2_3_lut (.I0(\data_in_frame[19] [1]), .I1(\data_in_frame[3] [1]), 
            .I2(n7569), .I3(GND_net), .O(n7571));
    defparam mux_2094_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_2094_i3_3_lut (.I0(\data_in_frame[19] [2]), .I1(\data_in_frame[3] [2]), 
            .I2(n7569), .I3(GND_net), .O(n7572));
    defparam mux_2094_i3_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_2094_i4_3_lut (.I0(\data_in_frame[19] [3]), .I1(\data_in_frame[3] [3]), 
            .I2(n7569), .I3(GND_net), .O(n7573));
    defparam mux_2094_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_1228 (.I0(\data_in_frame[4] [5]), .I1(\data_in_frame[5] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n47781));   // verilog/coms.v(71[16:27])
    defparam i1_2_lut_adj_1228.LUT_INIT = 16'h6666;
    SB_LUT4 mux_2094_i5_3_lut (.I0(\data_in_frame[19] [4]), .I1(\data_in_frame[3] [4]), 
            .I2(n7569), .I3(GND_net), .O(n7574));
    defparam mux_2094_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1229 (.I0(n43951), .I1(Kp_23__N_1059), .I2(n44344), 
            .I3(n47781), .O(n27817));   // verilog/coms.v(71[16:27])
    defparam i1_4_lut_adj_1229.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1230 (.I0(n27817), .I1(n40728), .I2(GND_net), 
            .I3(GND_net), .O(n41679));
    defparam i1_2_lut_adj_1230.LUT_INIT = 16'h6666;
    SB_LUT4 i1_3_lut_adj_1231 (.I0(n27457), .I1(n40972), .I2(\data_in_frame[8] [1]), 
            .I3(GND_net), .O(n44361));
    defparam i1_3_lut_adj_1231.LUT_INIT = 16'h9696;
    SB_LUT4 i15330_3_lut_4_lut (.I0(n8_adj_4681), .I1(n43820), .I2(rx_data[0]), 
            .I3(\data_in_frame[20] [0]), .O(n29278));
    defparam i15330_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_adj_1232 (.I0(\data_in_frame[21] [3]), .I1(n44065), 
            .I2(\data_in_frame[23] [4]), .I3(GND_net), .O(n45738));
    defparam i2_3_lut_adj_1232.LUT_INIT = 16'h9696;
    SB_LUT4 add_43_16_lut (.I0(n3345), .I1(\FRAME_MATCHER.i [14]), .I2(GND_net), 
            .I3(n38567), .O(n2_adj_4686)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_16_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mux_2094_i6_3_lut (.I0(\data_in_frame[19] [5]), .I1(\data_in_frame[3] [5]), 
            .I2(n7569), .I3(GND_net), .O(n7575));
    defparam mux_2094_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_43_16 (.CI(n38567), .I0(\FRAME_MATCHER.i [14]), .I1(GND_net), 
            .CO(n38568));
    SB_LUT4 mux_2094_i7_3_lut (.I0(\data_in_frame[19] [6]), .I1(\data_in_frame[3] [6]), 
            .I2(n7569), .I3(GND_net), .O(n7576));
    defparam mux_2094_i7_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_43_15_lut (.I0(n3345), .I1(\FRAME_MATCHER.i [13]), .I2(GND_net), 
            .I3(n38566), .O(n2_adj_4687)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_15_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_2_lut_3_lut (.I0(\data_in_frame[14] [2]), .I1(n26774), .I2(n41184), 
            .I3(GND_net), .O(n41651));
    defparam i1_2_lut_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 data_in_frame_1__4__I_0_2_lut (.I0(\data_in_frame[1] [4]), .I1(\data_in_frame[1] [3]), 
            .I2(GND_net), .I3(GND_net), .O(Kp_23__N_1103));   // verilog/coms.v(76[16:27])
    defparam data_in_frame_1__4__I_0_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mux_2094_i8_3_lut (.I0(\data_in_frame[19] [7]), .I1(\data_in_frame[3] [7]), 
            .I2(n7569), .I3(GND_net), .O(n7577));
    defparam mux_2094_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_2094_i9_3_lut (.I0(\data_in_frame[18] [0]), .I1(\data_in_frame[2] [0]), 
            .I2(n7569), .I3(GND_net), .O(n7578));
    defparam mux_2094_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut_adj_1233 (.I0(\data_in_frame[19] [3]), .I1(\data_in_frame[18] [7]), 
            .I2(\data_in_frame[23] [5]), .I3(GND_net), .O(n47867));
    defparam i1_3_lut_adj_1233.LUT_INIT = 16'h9696;
    SB_DFFSS \FRAME_MATCHER.i_i29  (.Q(\FRAME_MATCHER.i [29]), .C(CLK_c), 
            .D(n2_adj_4688), .S(n3_adj_4644));   // verilog/coms.v(128[12] 303[6])
    SB_DFFSS \FRAME_MATCHER.i_i28  (.Q(\FRAME_MATCHER.i [28]), .C(CLK_c), 
            .D(n2_adj_4689), .S(n3_adj_4643));   // verilog/coms.v(128[12] 303[6])
    SB_DFFSS \FRAME_MATCHER.i_i27  (.Q(\FRAME_MATCHER.i [27]), .C(CLK_c), 
            .D(n2_adj_4690), .S(n3_adj_4642));   // verilog/coms.v(128[12] 303[6])
    SB_DFFSS \FRAME_MATCHER.i_i26  (.Q(\FRAME_MATCHER.i [26]), .C(CLK_c), 
            .D(n2_adj_4691), .S(n3_adj_4641));   // verilog/coms.v(128[12] 303[6])
    SB_DFFSS \FRAME_MATCHER.i_i25  (.Q(\FRAME_MATCHER.i [25]), .C(CLK_c), 
            .D(n2_adj_4692), .S(n3_adj_4640));   // verilog/coms.v(128[12] 303[6])
    SB_DFFSS \FRAME_MATCHER.i_i24  (.Q(\FRAME_MATCHER.i [24]), .C(CLK_c), 
            .D(n2_adj_4693), .S(n3_adj_4639));   // verilog/coms.v(128[12] 303[6])
    SB_DFFSS \FRAME_MATCHER.i_i23  (.Q(\FRAME_MATCHER.i [23]), .C(CLK_c), 
            .D(n2_adj_4598), .S(n3_adj_4638));   // verilog/coms.v(128[12] 303[6])
    SB_DFFSS \FRAME_MATCHER.i_i22  (.Q(\FRAME_MATCHER.i [22]), .C(CLK_c), 
            .D(n2_adj_4656), .S(n3_adj_4636));   // verilog/coms.v(128[12] 303[6])
    SB_DFFSS \FRAME_MATCHER.i_i21  (.Q(\FRAME_MATCHER.i [21]), .C(CLK_c), 
            .D(n2_adj_4661), .S(n3_adj_4635));   // verilog/coms.v(128[12] 303[6])
    SB_DFFSS \FRAME_MATCHER.i_i20  (.Q(\FRAME_MATCHER.i [20]), .C(CLK_c), 
            .D(n2_adj_4664), .S(n3_adj_4634));   // verilog/coms.v(128[12] 303[6])
    SB_DFFSS \FRAME_MATCHER.i_i19  (.Q(\FRAME_MATCHER.i [19]), .C(CLK_c), 
            .D(n2_adj_4668), .S(n3_adj_4633));   // verilog/coms.v(128[12] 303[6])
    SB_DFFSS \FRAME_MATCHER.i_i18  (.Q(\FRAME_MATCHER.i [18]), .C(CLK_c), 
            .D(n2_adj_4675), .S(n3_adj_4632));   // verilog/coms.v(128[12] 303[6])
    SB_DFFSS \FRAME_MATCHER.i_i17  (.Q(\FRAME_MATCHER.i [17]), .C(CLK_c), 
            .D(n2_adj_4677), .S(n3_adj_4631));   // verilog/coms.v(128[12] 303[6])
    SB_DFFSS \FRAME_MATCHER.i_i16  (.Q(\FRAME_MATCHER.i [16]), .C(CLK_c), 
            .D(n2_adj_4680), .S(n3_adj_4630));   // verilog/coms.v(128[12] 303[6])
    SB_DFFSS \FRAME_MATCHER.i_i15  (.Q(\FRAME_MATCHER.i [15]), .C(CLK_c), 
            .D(n2_adj_4684), .S(n3_adj_4628));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 mux_2094_i10_3_lut (.I0(\data_in_frame[18] [1]), .I1(\data_in_frame[2] [1]), 
            .I2(n7569), .I3(GND_net), .O(n7579));
    defparam mux_2094_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_2094_i11_3_lut (.I0(\data_in_frame[18] [2]), .I1(\data_in_frame[2] [2]), 
            .I2(n7569), .I3(GND_net), .O(n7580));
    defparam mux_2094_i11_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut_adj_1234 (.I0(n44308), .I1(n43885), .I2(\data_in_frame[6] [1]), 
            .I3(GND_net), .O(n44513));   // verilog/coms.v(79[16:27])
    defparam i1_3_lut_adj_1234.LUT_INIT = 16'h9696;
    SB_LUT4 mux_2094_i12_3_lut (.I0(\data_in_frame[18] [3]), .I1(\data_in_frame[2] [3]), 
            .I2(n7569), .I3(GND_net), .O(n7581));
    defparam mux_2094_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_2094_i13_3_lut (.I0(\data_in_frame[18] [4]), .I1(\data_in_frame[2] [4]), 
            .I2(n7569), .I3(GND_net), .O(n7582));
    defparam mux_2094_i13_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_1235 (.I0(\data_in_frame[4] [0]), .I1(\data_in_frame[1] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n44308));   // verilog/coms.v(79[16:27])
    defparam i1_2_lut_adj_1235.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1236 (.I0(\data_in_frame[2] [0]), .I1(\data_in_frame[4] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n47773));   // verilog/coms.v(79[16:27])
    defparam i1_2_lut_adj_1236.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1237 (.I0(\data_in_frame[1] [4]), .I1(n44308), 
            .I2(n47773), .I3(\data_in_frame[1] [7]), .O(n44516));   // verilog/coms.v(79[16:27])
    defparam i1_4_lut_adj_1237.LUT_INIT = 16'h6996;
    SB_LUT4 mux_2094_i14_3_lut (.I0(\data_in_frame[18] [5]), .I1(\data_in_frame[2] [5]), 
            .I2(n7569), .I3(GND_net), .O(n7583));
    defparam mux_2094_i14_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_adj_1238 (.I0(\data_in_frame[14] [2]), .I1(n26774), 
            .I2(\data_in_frame[16] [4]), .I3(GND_net), .O(n44465));
    defparam i1_2_lut_3_lut_adj_1238.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1239 (.I0(\data_in_frame[1] [5]), .I1(\data_in_frame[3] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n43932));   // verilog/coms.v(79[16:27])
    defparam i1_2_lut_adj_1239.LUT_INIT = 16'h6666;
    SB_LUT4 mux_2094_i15_3_lut (.I0(\data_in_frame[18] [6]), .I1(\data_in_frame[2] [6]), 
            .I2(n7569), .I3(GND_net), .O(n7584));
    defparam mux_2094_i15_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1240 (.I0(n41751), .I1(\data_in_frame[21] [5]), 
            .I2(\data_in_frame[21] [4]), .I3(\data_in_frame[23] [6]), .O(n47863));
    defparam i1_4_lut_adj_1240.LUT_INIT = 16'h9669;
    SB_CARRY add_43_15 (.CI(n38566), .I0(\FRAME_MATCHER.i [13]), .I1(GND_net), 
            .CO(n38567));
    SB_LUT4 mux_2094_i16_3_lut (.I0(\data_in_frame[18] [7]), .I1(\data_in_frame[2] [7]), 
            .I2(n7569), .I3(GND_net), .O(n7585));
    defparam mux_2094_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_2094_i17_3_lut (.I0(\data_in_frame[17] [0]), .I1(\data_in_frame[1] [0]), 
            .I2(n7569), .I3(GND_net), .O(n7586));
    defparam mux_2094_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_43_14_lut (.I0(n3345), .I1(\FRAME_MATCHER.i [12]), .I2(GND_net), 
            .I3(n38565), .O(n2_adj_4694)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_14_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_43_14 (.CI(n38565), .I0(\FRAME_MATCHER.i [12]), .I1(GND_net), 
            .CO(n38566));
    SB_LUT4 i1_4_lut_adj_1241 (.I0(n44035), .I1(\data_in_frame[21] [6]), 
            .I2(\data_in_frame[19] [6]), .I3(\data_in_frame[22] [0]), .O(n47857));   // verilog/coms.v(86[17:28])
    defparam i1_4_lut_adj_1241.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1242 (.I0(\data_in_frame[20] [1]), .I1(\data_in_frame[22] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n47629));   // verilog/coms.v(79[16:27])
    defparam i1_2_lut_adj_1242.LUT_INIT = 16'h6666;
    SB_LUT4 mux_2094_i18_3_lut (.I0(\data_in_frame[17] [1]), .I1(\data_in_frame[1] [1]), 
            .I2(n7569), .I3(GND_net), .O(n7587));
    defparam mux_2094_i18_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_2094_i19_3_lut (.I0(\data_in_frame[17] [2]), .I1(\data_in_frame[1] [2]), 
            .I2(n7569), .I3(GND_net), .O(n7588));
    defparam mux_2094_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_43_13_lut (.I0(n3345), .I1(\FRAME_MATCHER.i [11]), .I2(GND_net), 
            .I3(n38564), .O(n2_adj_4695)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_13_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_4_lut_adj_1243 (.I0(n46024), .I1(n43992), .I2(n47629), 
            .I3(\data_in_frame[19] [6]), .O(n47635));   // verilog/coms.v(79[16:27])
    defparam i1_4_lut_adj_1243.LUT_INIT = 16'h9669;
    SB_LUT4 i1_3_lut_adj_1244 (.I0(n44559), .I1(\data_in_frame[19] [7]), 
            .I2(\data_in_frame[22] [3]), .I3(GND_net), .O(n47601));
    defparam i1_3_lut_adj_1244.LUT_INIT = 16'h9696;
    SB_CARRY add_43_13 (.CI(n38564), .I0(\FRAME_MATCHER.i [11]), .I1(GND_net), 
            .CO(n38565));
    SB_DFF data_out_frame_0___i40 (.Q(\data_out_frame[4] [7]), .C(CLK_c), 
           .D(n29124));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i1_rep_106_2_lut (.I0(\data_in_frame[20] [3]), .I1(\data_in_frame[20] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n51647));
    defparam i1_rep_106_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i15473_3_lut_4_lut (.I0(n8), .I1(n43832), .I2(rx_data[7]), 
            .I3(\data_in_frame[2] [7]), .O(n29421));
    defparam i15473_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 mux_2094_i20_3_lut (.I0(\data_in_frame[17] [3]), .I1(\data_in_frame[1] [3]), 
            .I2(n7569), .I3(GND_net), .O(n7589));
    defparam mux_2094_i20_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF data_out_frame_0___i41 (.Q(\data_out_frame[5] [0]), .C(CLK_c), 
           .D(n29123));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i42 (.Q(\data_out_frame[5] [1]), .C(CLK_c), 
           .D(n29122));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 mux_2094_i21_3_lut (.I0(\data_in_frame[17] [4]), .I1(\data_in_frame[1] [4]), 
            .I2(n7569), .I3(GND_net), .O(n7590));
    defparam mux_2094_i21_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF data_out_frame_0___i43 (.Q(\data_out_frame[5] [2]), .C(CLK_c), 
           .D(n29121));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 mux_2094_i22_3_lut (.I0(\data_in_frame[17] [5]), .I1(\data_in_frame[1] [5]), 
            .I2(n7569), .I3(GND_net), .O(n7591));
    defparam mux_2094_i22_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i6_4_lut_adj_1245 (.I0(n44146), .I1(n12_adj_4676), .I2(\data_in_frame[23] [3]), 
            .I3(n41688), .O(n46369));
    defparam i6_4_lut_adj_1245.LUT_INIT = 16'h6996;
    SB_LUT4 mux_2094_i23_3_lut (.I0(\data_in_frame[17] [6]), .I1(\data_in_frame[1] [6]), 
            .I2(n7569), .I3(GND_net), .O(n7592));
    defparam mux_2094_i23_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_2094_i24_3_lut (.I0(\data_in_frame[17] [7]), .I1(\data_in_frame[1] [7]), 
            .I2(n7569), .I3(GND_net), .O(n7593));
    defparam mux_2094_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut_adj_1246 (.I0(n28288), .I1(n27488), .I2(\data_in_frame[8] [2]), 
            .I3(GND_net), .O(n4_adj_4659));   // verilog/coms.v(77[16:43])
    defparam i1_3_lut_adj_1246.LUT_INIT = 16'h9696;
    SB_LUT4 i15474_3_lut_4_lut (.I0(n8), .I1(n43832), .I2(rx_data[6]), 
            .I3(\data_in_frame[2] [6]), .O(n29422));
    defparam i15474_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_out_frame_0___i44 (.Q(\data_out_frame[5] [3]), .C(CLK_c), 
           .D(n29120));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i45 (.Q(\data_out_frame[5] [4]), .C(CLK_c), 
           .D(n29119));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i1_4_lut_adj_1247 (.I0(\data_in_frame[20] [5]), .I1(n45738), 
            .I2(n8_adj_4696), .I3(n27335), .O(n47373));
    defparam i1_4_lut_adj_1247.LUT_INIT = 16'hedde;
    SB_DFF data_out_frame_0___i46 (.Q(\data_out_frame[5] [5]), .C(CLK_c), 
           .D(n29118));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i47 (.Q(\data_out_frame[5] [6]), .C(CLK_c), 
           .D(n29117));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i48 (.Q(\data_out_frame[5] [7]), .C(CLK_c), 
           .D(n29116));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i49 (.Q(\data_out_frame[6] [0]), .C(CLK_c), 
           .D(n29115));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i50 (.Q(\data_out_frame[6] [1]), .C(CLK_c), 
           .D(n29114));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i51 (.Q(\data_out_frame[6] [2]), .C(CLK_c), 
           .D(n29113));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i52 (.Q(\data_out_frame[6] [3]), .C(CLK_c), 
           .D(n29112));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i53 (.Q(\data_out_frame[6] [4]), .C(CLK_c), 
           .D(n29111));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i54 (.Q(\data_out_frame[6] [5]), .C(CLK_c), 
           .D(n29110));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i55 (.Q(\data_out_frame[6] [6]), .C(CLK_c), 
           .D(n29109));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i56 (.Q(\data_out_frame[6] [7]), .C(CLK_c), 
           .D(n29108));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i57 (.Q(\data_out_frame[7] [0]), .C(CLK_c), 
           .D(n29107));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i3_4_lut_adj_1248 (.I0(\data_in_frame[23] [2]), .I1(n44168), 
            .I2(n41688), .I3(\data_in_frame[21] [1]), .O(n45168));
    defparam i3_4_lut_adj_1248.LUT_INIT = 16'h9669;
    SB_LUT4 i3_4_lut_adj_1249 (.I0(\data_in_frame[22] [5]), .I1(n44453), 
            .I2(n44425), .I3(n51647), .O(n45428));
    defparam i3_4_lut_adj_1249.LUT_INIT = 16'h6996;
    SB_LUT4 i15475_3_lut_4_lut (.I0(n8), .I1(n43832), .I2(rx_data[5]), 
            .I3(\data_in_frame[2] [5]), .O(n29423));
    defparam i15475_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i4_4_lut_adj_1250 (.I0(\data_in_frame[22] [4]), .I1(n41303), 
            .I2(n40620), .I3(\data_in_frame[20] [2]), .O(n10_adj_4697));
    defparam i4_4_lut_adj_1250.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1251 (.I0(n45428), .I1(n45168), .I2(n47373), 
            .I3(n46369), .O(n47379));
    defparam i1_4_lut_adj_1251.LUT_INIT = 16'hfbff;
    SB_LUT4 i2_4_lut_adj_1252 (.I0(\data_in_frame[19] [3]), .I1(\data_in_frame[21] [6]), 
            .I2(n41769), .I3(\data_in_frame[21] [5]), .O(n6_adj_4698));
    defparam i2_4_lut_adj_1252.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1253 (.I0(\data_in_frame[18] [2]), .I1(n47379), 
            .I2(n10_adj_4697), .I3(\data_in_frame[20] [3]), .O(n47381));
    defparam i1_4_lut_adj_1253.LUT_INIT = 16'hdeed;
    SB_DFFE data_out_frame_0___i224 (.Q(\data_out_frame[27] [7]), .C(CLK_c), 
            .E(n28621), .D(n46044));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i1_4_lut_adj_1254 (.I0(n27668), .I1(\data_in_frame[19] [5]), 
            .I2(\data_in_frame[19] [7]), .I3(\data_in_frame[22] [1]), .O(n47879));
    defparam i1_4_lut_adj_1254.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1255 (.I0(n44272), .I1(n47381), .I2(n6_adj_4698), 
            .I3(\data_in_frame[23] [7]), .O(n47383));
    defparam i1_4_lut_adj_1255.LUT_INIT = 16'hedde;
    SB_LUT4 i1_4_lut_adj_1256 (.I0(n44331), .I1(\data_in_frame[21] [4]), 
            .I2(n47867), .I3(\data_in_frame[21] [3]), .O(n47871));
    defparam i1_4_lut_adj_1256.LUT_INIT = 16'h6996;
    SB_LUT4 i3_3_lut_adj_1257 (.I0(\FRAME_MATCHER.state [2]), .I1(n44728), 
            .I2(\FRAME_MATCHER.state [3]), .I3(GND_net), .O(n63));   // verilog/coms.v(202[5:24])
    defparam i3_3_lut_adj_1257.LUT_INIT = 16'hefef;
    SB_LUT4 i1_4_lut_adj_1258 (.I0(n44155), .I1(n47383), .I2(n44035), 
            .I3(n47879), .O(n47385));
    defparam i1_4_lut_adj_1258.LUT_INIT = 16'hdeed;
    SB_LUT4 i1_2_lut_adj_1259 (.I0(n27506), .I1(n27979), .I2(GND_net), 
            .I3(GND_net), .O(Kp_23__N_1327));   // verilog/coms.v(77[16:43])
    defparam i1_2_lut_adj_1259.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1260 (.I0(n27976), .I1(n4_adj_4659), .I2(GND_net), 
            .I3(GND_net), .O(n43902));   // verilog/coms.v(75[16:43])
    defparam i1_2_lut_adj_1260.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1261 (.I0(n27544), .I1(n27554), .I2(GND_net), 
            .I3(GND_net), .O(n43986));
    defparam i1_2_lut_adj_1261.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1262 (.I0(Kp_23__N_1135), .I1(Kp_23__N_1132), .I2(n27469), 
            .I3(\data_in_frame[8] [5]), .O(n27979));
    defparam i1_4_lut_adj_1262.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1263 (.I0(n47857), .I1(n47863), .I2(n45887), 
            .I3(n44196), .O(n47389));
    defparam i1_4_lut_adj_1263.LUT_INIT = 16'h7bde;
    SB_LUT4 i1_4_lut_adj_1264 (.I0(n43986), .I1(n43902), .I2(Kp_23__N_1327), 
            .I3(Kp_23__N_1253), .O(n47407));
    defparam i1_4_lut_adj_1264.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1265 (.I0(n44528), .I1(n44361), .I2(n47407), 
            .I3(n41679), .O(n26693));
    defparam i1_4_lut_adj_1265.LUT_INIT = 16'h6996;
    SB_LUT4 i33824_2_lut (.I0(n51495), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n49354));
    defparam i33824_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1_4_lut_adj_1266 (.I0(n27411), .I1(n27495), .I2(\data_in_frame[4] [5]), 
            .I3(\data_in_frame[6] [6]), .O(Kp_23__N_1253));   // verilog/coms.v(76[16:43])
    defparam i1_4_lut_adj_1266.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1267 (.I0(\data_in_frame[9] [2]), .I1(Kp_23__N_1253), 
            .I2(GND_net), .I3(GND_net), .O(n44072));   // verilog/coms.v(73[16:41])
    defparam i1_2_lut_adj_1267.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1268 (.I0(n47389), .I1(n47385), .I2(n47871), 
            .I3(n41769), .O(n47391));
    defparam i1_4_lut_adj_1268.LUT_INIT = 16'heffe;
    SB_LUT4 i1_3_lut_adj_1269 (.I0(n47339), .I1(n26693), .I2(n27979), 
            .I3(GND_net), .O(n40706));   // verilog/coms.v(86[17:63])
    defparam i1_3_lut_adj_1269.LUT_INIT = 16'h9696;
    SB_LUT4 i1_3_lut_adj_1270 (.I0(\data_in_frame[8] [2]), .I1(n40706), 
            .I2(\data_in_frame[8] [3]), .I3(GND_net), .O(n44556));
    defparam i1_3_lut_adj_1270.LUT_INIT = 16'h9696;
    SB_LUT4 i15053_2_lut (.I0(n63), .I1(n27235), .I2(GND_net), .I3(GND_net), 
            .O(n28996));   // verilog/coms.v(128[12] 303[6])
    defparam i15053_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i1_2_lut_adj_1271 (.I0(\data_in_frame[1] [5]), .I1(\data_in_frame[3] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n43885));   // verilog/coms.v(79[16:27])
    defparam i1_2_lut_adj_1271.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1272 (.I0(n44155), .I1(n44453), .I2(n27861), 
            .I3(n47635), .O(n47641));   // verilog/coms.v(79[16:27])
    defparam i1_4_lut_adj_1272.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1273 (.I0(n41303), .I1(n44531), .I2(n44199), 
            .I3(n47601), .O(n47607));
    defparam i1_4_lut_adj_1273.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1274 (.I0(\data_in_frame[4] [1]), .I1(\data_in_frame[2] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n47727));   // verilog/coms.v(79[16:27])
    defparam i1_2_lut_adj_1274.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1275 (.I0(n43885), .I1(n44305), .I2(n47727), 
            .I3(\data_in_frame[0] [0]), .O(Kp_23__N_1132));   // verilog/coms.v(79[16:27])
    defparam i1_4_lut_adj_1275.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1276 (.I0(n44592), .I1(n44459), .I2(\data_in_frame[20] [5]), 
            .I3(\data_in_frame[22] [7]), .O(n47535));
    defparam i1_4_lut_adj_1276.LUT_INIT = 16'h6996;
    SB_LUT4 i32609_4_lut (.I0(\data_out_frame[6] [7]), .I1(byte_transmit_counter[0]), 
            .I2(byte_transmit_counter[2]), .I3(\data_out_frame[7] [7]), 
            .O(n48196));
    defparam i32609_4_lut.LUT_INIT = 16'hec2c;
    SB_LUT4 i32607_3_lut (.I0(\data_out_frame[4] [7]), .I1(\data_out_frame[5] [7]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n48194));
    defparam i32607_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFE data_out_frame_0___i223 (.Q(\data_out_frame[27] [6]), .C(CLK_c), 
            .E(n28621), .D(n45944));   // verilog/coms.v(128[12] 303[6])
    SB_DFFE data_out_frame_0___i222 (.Q(\data_out_frame[27] [5]), .C(CLK_c), 
            .E(n28621), .D(n44446));   // verilog/coms.v(128[12] 303[6])
    SB_DFFE data_out_frame_0___i221 (.Q(\data_out_frame[27] [4]), .C(CLK_c), 
            .E(n28621), .D(n46011));   // verilog/coms.v(128[12] 303[6])
    SB_DFFE data_out_frame_0___i220 (.Q(\data_out_frame[27] [3]), .C(CLK_c), 
            .E(n28621), .D(n45375));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i15476_3_lut_4_lut (.I0(n8), .I1(n43832), .I2(rx_data[4]), 
            .I3(\data_in_frame[2] [4]), .O(n29424));
    defparam i15476_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 add_43_12_lut (.I0(n3345), .I1(\FRAME_MATCHER.i [10]), .I2(GND_net), 
            .I3(n38563), .O(n2_adj_4699)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_12_lut.LUT_INIT = 16'h8228;
    SB_DFFE data_out_frame_0___i219 (.Q(\data_out_frame[27] [2]), .C(CLK_c), 
            .E(n28621), .D(n45888));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i1_4_lut_adj_1277 (.I0(n47607), .I1(n47641), .I2(n44367), 
            .I3(n47391), .O(n47395));
    defparam i1_4_lut_adj_1277.LUT_INIT = 16'hffbd;
    SB_LUT4 i33819_2_lut (.I0(n51501), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n49345));
    defparam i33819_2_lut.LUT_INIT = 16'h2222;
    SB_CARRY add_43_12 (.CI(n38563), .I0(\FRAME_MATCHER.i [10]), .I1(GND_net), 
            .CO(n38564));
    SB_DFFE data_out_frame_0___i218 (.Q(\data_out_frame[27] [1]), .C(CLK_c), 
            .E(n28621), .D(n45371));   // verilog/coms.v(128[12] 303[6])
    SB_DFFE data_out_frame_0___i217 (.Q(\data_out_frame[27] [0]), .C(CLK_c), 
            .E(n28621), .D(n45804));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i1_4_lut_adj_1278 (.I0(n44531), .I1(n45675), .I2(n44168), 
            .I3(n47535), .O(n46382));
    defparam i1_4_lut_adj_1278.LUT_INIT = 16'h9669;
    SB_LUT4 i1_4_lut_adj_1279 (.I0(n44168), .I1(n41688), .I2(\data_in_frame[23] [0]), 
            .I3(n45675), .O(n46335));
    defparam i1_4_lut_adj_1279.LUT_INIT = 16'h6996;
    SB_LUT4 i1_3_lut_adj_1280 (.I0(\data_in_frame[23] [1]), .I1(n41688), 
            .I2(n45675), .I3(GND_net), .O(n41755));
    defparam i1_3_lut_adj_1280.LUT_INIT = 16'h9696;
    SB_LUT4 i1_4_lut_adj_1281 (.I0(n41755), .I1(n46335), .I2(n46382), 
            .I3(n47395), .O(n31));
    defparam i1_4_lut_adj_1281.LUT_INIT = 16'hff7f;
    SB_LUT4 i15477_3_lut_4_lut (.I0(n8), .I1(n43832), .I2(rx_data[3]), 
            .I3(\data_in_frame[2] [3]), .O(n29425));
    defparam i15477_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1282 (.I0(\FRAME_MATCHER.state [3]), .I1(\FRAME_MATCHER.state [2]), 
            .I2(GND_net), .I3(GND_net), .O(n47575));
    defparam i1_2_lut_adj_1282.LUT_INIT = 16'h4444;
    SB_LUT4 i1_4_lut_adj_1283 (.I0(n44728), .I1(n31), .I2(n24450), .I3(n47575), 
            .O(n28521));
    defparam i1_4_lut_adj_1283.LUT_INIT = 16'h0100;
    SB_LUT4 i15478_3_lut_4_lut (.I0(n8), .I1(n43832), .I2(rx_data[2]), 
            .I3(\data_in_frame[2] [2]), .O(n29426));
    defparam i15478_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_3_lut_adj_1284 (.I0(\data_in_frame[6] [3]), .I1(Kp_23__N_1132), 
            .I2(\data_in_frame[8] [4]), .I3(GND_net), .O(n44358));   // verilog/coms.v(75[16:43])
    defparam i1_3_lut_adj_1284.LUT_INIT = 16'h9696;
    SB_DFFE data_out_frame_0___i216 (.Q(\data_out_frame[26] [7]), .C(CLK_c), 
            .E(n28621), .D(n45796));   // verilog/coms.v(128[12] 303[6])
    SB_DFFE data_out_frame_0___i215 (.Q(\data_out_frame[26] [6]), .C(CLK_c), 
            .E(n28621), .D(n45385));   // verilog/coms.v(128[12] 303[6])
    SB_DFFSS \FRAME_MATCHER.i_i14  (.Q(\FRAME_MATCHER.i [14]), .C(CLK_c), 
            .D(n2_adj_4686), .S(n3_adj_4700));   // verilog/coms.v(128[12] 303[6])
    SB_DFFE data_out_frame_0___i214 (.Q(\data_out_frame[26] [5]), .C(CLK_c), 
            .E(n28621), .D(n44267));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i34552_3_lut (.I0(n51573), .I1(n51321), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n50140));
    defparam i34552_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFE data_out_frame_0___i213 (.Q(\data_out_frame[26] [4]), .C(CLK_c), 
            .E(n28621), .D(n45560));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 add_43_11_lut (.I0(n3345), .I1(\FRAME_MATCHER.i [9]), .I2(GND_net), 
            .I3(n38562), .O(n2_adj_4701)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_11_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_43_11 (.CI(n38562), .I0(\FRAME_MATCHER.i [9]), .I1(GND_net), 
            .CO(n38563));
    SB_LUT4 i1_2_lut_adj_1285 (.I0(n28009), .I1(\data_in_frame[10] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n40702));
    defparam i1_2_lut_adj_1285.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1286 (.I0(\data_in_frame[9] [0]), .I1(\data_in_frame[9] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n47837));
    defparam i1_2_lut_adj_1286.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1287 (.I0(n44006), .I1(n44358), .I2(n47837), 
            .I3(\data_in_frame[8] [1]), .O(n47843));
    defparam i1_4_lut_adj_1287.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1288 (.I0(n28009), .I1(n44556), .I2(n44419), 
            .I3(n47843), .O(n41622));
    defparam i1_4_lut_adj_1288.LUT_INIT = 16'h6996;
    SB_LUT4 i1_3_lut_adj_1289 (.I0(\data_in_frame[0] [4]), .I1(\data_in_frame[0] [5]), 
            .I2(\data_in_frame[2] [6]), .I3(GND_net), .O(n7));   // verilog/coms.v(77[16:27])
    defparam i1_3_lut_adj_1289.LUT_INIT = 16'h9696;
    SB_LUT4 i1_3_lut_adj_1290 (.I0(\data_in_frame[5] [2]), .I1(n7), .I2(\data_in_frame[5] [3]), 
            .I3(GND_net), .O(n44116));
    defparam i1_3_lut_adj_1290.LUT_INIT = 16'h9696;
    SB_LUT4 i15479_3_lut_4_lut (.I0(n8), .I1(n43832), .I2(rx_data[1]), 
            .I3(\data_in_frame[2] [1]), .O(n29427));
    defparam i15479_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1291 (.I0(\data_in_frame[11] [3]), .I1(Kp_23__N_1465), 
            .I2(n44012), .I3(GND_net), .O(Kp_23__N_1561));   // verilog/coms.v(72[16:27])
    defparam i1_2_lut_3_lut_adj_1291.LUT_INIT = 16'h9696;
    SB_LUT4 add_43_10_lut (.I0(n3345), .I1(\FRAME_MATCHER.i [8]), .I2(GND_net), 
            .I3(n38561), .O(n2_adj_4702)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_10_lut.LUT_INIT = 16'h8228;
    SB_DFFSS \FRAME_MATCHER.i_i13  (.Q(\FRAME_MATCHER.i [13]), .C(CLK_c), 
            .D(n2_adj_4687), .S(n3_adj_4703));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [2]), .I2(\data_out_frame[27] [2]), 
            .I3(byte_transmit_counter[1]), .O(n51582));
    defparam byte_transmit_counter_0__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n51582_bdd_4_lut (.I0(n51582), .I1(\data_out_frame[25] [2]), 
            .I2(\data_out_frame[24] [2]), .I3(byte_transmit_counter[1]), 
            .O(n51585));
    defparam n51582_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_CARRY add_43_10 (.CI(n38561), .I0(\FRAME_MATCHER.i [8]), .I1(GND_net), 
            .CO(n38562));
    SB_LUT4 add_43_9_lut (.I0(n3345), .I1(\FRAME_MATCHER.i [7]), .I2(GND_net), 
            .I3(n38560), .O(n2_adj_4704)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_9_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_43_9 (.CI(n38560), .I0(\FRAME_MATCHER.i [7]), .I1(GND_net), 
            .CO(n38561));
    SB_DFFSS \FRAME_MATCHER.i_i12  (.Q(\FRAME_MATCHER.i [12]), .C(CLK_c), 
            .D(n2_adj_4694), .S(n3_adj_4705));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i15480_3_lut_4_lut (.I0(n8), .I1(n43832), .I2(rx_data[0]), 
            .I3(\data_in_frame[2] [0]), .O(n29428));
    defparam i15480_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 add_43_8_lut (.I0(n3345), .I1(\FRAME_MATCHER.i [6]), .I2(GND_net), 
            .I3(n38559), .O(n2_adj_4706)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_8_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_43_8 (.CI(n38559), .I0(\FRAME_MATCHER.i [6]), .I1(GND_net), 
            .CO(n38560));
    SB_LUT4 add_43_7_lut (.I0(n3345), .I1(\FRAME_MATCHER.i [5]), .I2(GND_net), 
            .I3(n38558), .O(n2_adj_4707)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_7_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_43_7 (.CI(n38558), .I0(\FRAME_MATCHER.i [5]), .I1(GND_net), 
            .CO(n38559));
    SB_LUT4 i1_3_lut_adj_1292 (.I0(\data_in_frame[5] [4]), .I1(n28357), 
            .I2(\data_in_frame[5] [5]), .I3(GND_net), .O(n27350));
    defparam i1_3_lut_adj_1292.LUT_INIT = 16'h9696;
    SB_LUT4 equal_306_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8));   // verilog/coms.v(155[7:23])
    defparam equal_306_i8_2_lut_3_lut.LUT_INIT = 16'hfdfd;
    SB_LUT4 i2_3_lut_4_lut_adj_1293 (.I0(\data_out_frame[20] [2]), .I1(n41171), 
            .I2(n43960), .I3(\data_out_frame[22] [4]), .O(n41701));
    defparam i2_3_lut_4_lut_adj_1293.LUT_INIT = 16'h9669;
    SB_LUT4 i1_4_lut_adj_1294 (.I0(\data_in_frame[4] [1]), .I1(\data_in_frame[3] [7]), 
            .I2(\data_in_frame[4] [7]), .I3(\data_in_frame[2] [5]), .O(n47351));   // verilog/coms.v(74[16:42])
    defparam i1_4_lut_adj_1294.LUT_INIT = 16'h6996;
    SB_DFFSS \FRAME_MATCHER.i_i11  (.Q(\FRAME_MATCHER.i [11]), .C(CLK_c), 
            .D(n2_adj_4695), .S(n3_adj_4708));   // verilog/coms.v(128[12] 303[6])
    SB_DFFSS \FRAME_MATCHER.i_i10  (.Q(\FRAME_MATCHER.i [10]), .C(CLK_c), 
            .D(n2_adj_4699), .S(n3_adj_4709));   // verilog/coms.v(128[12] 303[6])
    SB_DFFE data_out_frame_0___i212 (.Q(\data_out_frame[26] [3]), .C(CLK_c), 
            .E(n28621), .D(n44142));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i1_3_lut_adj_1295 (.I0(\data_in_frame[2] [3]), .I1(\data_in_frame[2] [7]), 
            .I2(\data_in_frame[3] [0]), .I3(GND_net), .O(n47349));   // verilog/coms.v(74[16:42])
    defparam i1_3_lut_adj_1295.LUT_INIT = 16'h9696;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_35928 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [1]), .I2(\data_out_frame[27] [1]), 
            .I3(byte_transmit_counter[1]), .O(n51576));
    defparam byte_transmit_counter_0__bdd_4_lut_35928.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_4_lut_adj_1296 (.I0(n27420), .I1(n47349), .I2(\data_in_frame[3] [6]), 
            .I3(\data_in_frame[4] [0]), .O(n47359));   // verilog/coms.v(74[16:42])
    defparam i1_4_lut_adj_1296.LUT_INIT = 16'h6996;
    SB_LUT4 add_43_6_lut (.I0(n3345), .I1(\FRAME_MATCHER.i [4]), .I2(GND_net), 
            .I3(n38557), .O(n2_adj_4590)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_6_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_4_lut_adj_1297 (.I0(n44116), .I1(n47359), .I2(n47361), 
            .I3(n47357), .O(n47367));   // verilog/coms.v(74[16:42])
    defparam i1_4_lut_adj_1297.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1298 (.I0(Kp_23__N_1135), .I1(n44547), .I2(n47367), 
            .I3(n44364), .O(n40678));   // verilog/coms.v(74[16:42])
    defparam i1_4_lut_adj_1298.LUT_INIT = 16'h6996;
    SB_LUT4 equal_297_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8_adj_4655));   // verilog/coms.v(155[7:23])
    defparam equal_297_i8_2_lut_3_lut.LUT_INIT = 16'hdfdf;
    SB_LUT4 n51576_bdd_4_lut (.I0(n51576), .I1(\data_out_frame[25] [1]), 
            .I2(\data_out_frame[24] [1]), .I3(byte_transmit_counter[1]), 
            .O(n51579));
    defparam n51576_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_adj_1299 (.I0(\data_in_frame[9] [5]), .I1(\data_in_frame[11] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n44617));
    defparam i1_2_lut_adj_1299.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1300 (.I0(\data_in_frame[6] [3]), .I1(\data_in_frame[6] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n27469));   // verilog/coms.v(86[17:28])
    defparam i1_2_lut_adj_1300.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1301 (.I0(\data_in_frame[6] [5]), .I1(n27469), 
            .I2(\data_in_frame[6] [2]), .I3(\data_in_frame[6] [1]), .O(n44394));   // verilog/coms.v(86[17:28])
    defparam i1_4_lut_adj_1301.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1302 (.I0(n28357), .I1(\data_in_frame[7] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n44432));
    defparam i1_2_lut_adj_1302.LUT_INIT = 16'h6666;
    SB_LUT4 i1_3_lut_adj_1303 (.I0(\data_in_frame[2] [1]), .I1(n27948), 
            .I2(\data_in_frame[4] [4]), .I3(GND_net), .O(n44364));   // verilog/coms.v(75[16:43])
    defparam i1_3_lut_adj_1303.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1304 (.I0(\data_in_frame[1] [7]), .I1(\data_in_frame[0] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n43989));   // verilog/coms.v(71[16:69])
    defparam i1_2_lut_adj_1304.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1305 (.I0(n43989), .I1(n44364), .I2(\data_in_frame[4] [3]), 
            .I3(\data_in_frame[6] [5]), .O(n27495));   // verilog/coms.v(75[16:43])
    defparam i1_4_lut_adj_1305.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1306 (.I0(n27952), .I1(n44305), .I2(\data_in_frame[2] [0]), 
            .I3(\data_in_frame[4] [3]), .O(Kp_23__N_1135));   // verilog/coms.v(74[16:42])
    defparam i1_4_lut_adj_1306.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1307 (.I0(\data_in_frame[0] [3]), .I1(\data_in_frame[0] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n43914));   // verilog/coms.v(167[9:87])
    defparam i1_2_lut_adj_1307.LUT_INIT = 16'h6666;
    SB_LUT4 i1_3_lut_adj_1308 (.I0(\data_in_frame[0] [1]), .I1(\data_in_frame[0] [0]), 
            .I2(\data_in_frame[2] [2]), .I3(GND_net), .O(n27952));   // verilog/coms.v(76[16:43])
    defparam i1_3_lut_adj_1308.LUT_INIT = 16'h9696;
    SB_LUT4 i1_3_lut_adj_1309 (.I0(n27952), .I1(n27461), .I2(\data_in_frame[4] [4]), 
            .I3(GND_net), .O(n27411));   // verilog/coms.v(76[16:43])
    defparam i1_3_lut_adj_1309.LUT_INIT = 16'h9696;
    SB_LUT4 i1_3_lut_adj_1310 (.I0(\data_in_frame[2] [3]), .I1(\data_in_frame[0] [1]), 
            .I2(\data_in_frame[0] [2]), .I3(GND_net), .O(n27948));   // verilog/coms.v(76[16:43])
    defparam i1_3_lut_adj_1310.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1311 (.I0(\data_in_frame[0] [6]), .I1(\data_in_frame[1] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n43944));
    defparam i1_2_lut_adj_1311.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1312 (.I0(Kp_23__N_1135), .I1(n27495), .I2(\data_in_frame[6] [4]), 
            .I3(\data_in_frame[8] [6]), .O(n27933));   // verilog/coms.v(77[16:43])
    defparam i1_4_lut_adj_1312.LUT_INIT = 16'h6996;
    SB_LUT4 i1_3_lut_adj_1313 (.I0(n27948), .I1(n27411), .I2(\data_in_frame[7] [0]), 
            .I3(GND_net), .O(n44391));   // verilog/coms.v(75[16:43])
    defparam i1_3_lut_adj_1313.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1314 (.I0(\data_in_frame[8] [7]), .I1(n27933), 
            .I2(GND_net), .I3(GND_net), .O(n28367));   // verilog/coms.v(77[16:43])
    defparam i1_2_lut_adj_1314.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1315 (.I0(\data_in_frame[6] [7]), .I1(\data_in_frame[7] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n44344));   // verilog/coms.v(71[16:27])
    defparam i1_2_lut_adj_1315.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1316 (.I0(\data_in_frame[9] [1]), .I1(\data_in_frame[9] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n27370));   // verilog/coms.v(72[16:27])
    defparam i1_2_lut_adj_1316.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1317 (.I0(\data_in_frame[12] [1]), .I1(\data_in_frame[6] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n44565));
    defparam i1_2_lut_adj_1317.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1318 (.I0(\data_in_frame[4] [7]), .I1(\data_in_frame[9] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n47801));
    defparam i1_2_lut_adj_1318.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1319 (.I0(\data_in_frame[9] [7]), .I1(n47801), 
            .I2(\data_in_frame[5] [2]), .I3(\data_in_frame[12] [0]), .O(n47805));
    defparam i1_4_lut_adj_1319.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1320 (.I0(n47805), .I1(n44565), .I2(n27370), 
            .I3(n44344), .O(n47811));
    defparam i1_4_lut_adj_1320.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1321 (.I0(n44432), .I1(n43971), .I2(n44394), 
            .I3(n47811), .O(n47817));
    defparam i1_4_lut_adj_1321.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_35923 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[18] [7]), .I2(\data_out_frame[19] [7]), 
            .I3(byte_transmit_counter[1]), .O(n51570));
    defparam byte_transmit_counter_0__bdd_4_lut_35923.LUT_INIT = 16'he4aa;
    SB_DFF data_out_frame_0___i58 (.Q(\data_out_frame[7] [1]), .C(CLK_c), 
           .D(n29106));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 n51570_bdd_4_lut (.I0(n51570), .I1(\data_out_frame[17] [7]), 
            .I2(\data_out_frame[16] [7]), .I3(byte_transmit_counter[1]), 
            .O(n51573));
    defparam n51570_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFFE data_out_frame_0___i211 (.Q(\data_out_frame[26] [2]), .C(CLK_c), 
            .E(n28621), .D(n45472));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i59 (.Q(\data_out_frame[7] [2]), .C(CLK_c), 
           .D(n29105));   // verilog/coms.v(128[12] 303[6])
    SB_DFFE data_out_frame_0___i210 (.Q(\data_out_frame[26] [1]), .C(CLK_c), 
            .E(n28621), .D(n46198));   // verilog/coms.v(128[12] 303[6])
    SB_DFFE data_out_frame_0___i209 (.Q(\data_out_frame[26] [0]), .C(CLK_c), 
            .E(n28621), .D(n45477));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i20869_4_lut (.I0(\FRAME_MATCHER.i [3]), .I1(\FRAME_MATCHER.i [31]), 
            .I2(n27189), .I3(\FRAME_MATCHER.i [4]), .O(n4452));   // verilog/coms.v(260[9:58])
    defparam i20869_4_lut.LUT_INIT = 16'h3230;
    SB_LUT4 i1_2_lut_adj_1322 (.I0(\FRAME_MATCHER.state [1]), .I1(n27230), 
            .I2(GND_net), .I3(GND_net), .O(n27231));   // verilog/coms.v(255[5:25])
    defparam i1_2_lut_adj_1322.LUT_INIT = 16'hdddd;
    SB_LUT4 i1_2_lut_adj_1323 (.I0(n53), .I1(n65), .I2(GND_net), .I3(GND_net), 
            .O(n33840));   // verilog/coms.v(128[12] 303[6])
    defparam i1_2_lut_adj_1323.LUT_INIT = 16'heeee;
    SB_LUT4 i6_4_lut_adj_1324 (.I0(\data_in[1] [3]), .I1(\data_in[0] [1]), 
            .I2(\data_in[3] [2]), .I3(\data_in[0] [5]), .O(n16_adj_4710));
    defparam i6_4_lut_adj_1324.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_4_lut_adj_1325 (.I0(\data_in[2] [6]), .I1(\data_in[2] [5]), 
            .I2(\data_in[2] [0]), .I3(\data_in[1] [2]), .O(n17_adj_4711));
    defparam i7_4_lut_adj_1325.LUT_INIT = 16'hfffd;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_35918 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[18] [1]), .I2(\data_out_frame[19] [1]), 
            .I3(byte_transmit_counter[1]), .O(n51564));
    defparam byte_transmit_counter_0__bdd_4_lut_35918.LUT_INIT = 16'he4aa;
    SB_LUT4 i9_4_lut_adj_1326 (.I0(n17_adj_4711), .I1(\data_in[1] [6]), 
            .I2(n16_adj_4710), .I3(\data_in[3] [7]), .O(n27136));
    defparam i9_4_lut_adj_1326.LUT_INIT = 16'hfbff;
    SB_LUT4 n51564_bdd_4_lut (.I0(n51564), .I1(\data_out_frame[17] [1]), 
            .I2(\data_out_frame[16] [1]), .I3(byte_transmit_counter[1]), 
            .O(n51567));
    defparam n51564_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF data_out_frame_0___i107 (.Q(\data_out_frame[13] [2]), .C(CLK_c), 
           .D(n29679));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i108 (.Q(\data_out_frame[13] [3]), .C(CLK_c), 
           .D(n29678));   // verilog/coms.v(128[12] 303[6])
    SB_CARRY add_43_6 (.CI(n38557), .I0(\FRAME_MATCHER.i [4]), .I1(GND_net), 
            .CO(n38558));
    SB_DFF data_out_frame_0___i109 (.Q(\data_out_frame[13] [4]), .C(CLK_c), 
           .D(n29677));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 add_43_5_lut (.I0(n3345), .I1(\FRAME_MATCHER.i [3]), .I2(GND_net), 
            .I3(n38556), .O(n2)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_5_lut.LUT_INIT = 16'h8228;
    SB_DFF data_out_frame_0___i110 (.Q(\data_out_frame[13] [5]), .C(CLK_c), 
           .D(n29676));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i111 (.Q(\data_out_frame[13] [6]), .C(CLK_c), 
           .D(n29675));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i112 (.Q(\data_out_frame[13] [7]), .C(CLK_c), 
           .D(n29674));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i113 (.Q(\data_out_frame[14] [0]), .C(CLK_c), 
           .D(n29673));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i114 (.Q(\data_out_frame[14] [1]), .C(CLK_c), 
           .D(n29672));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i115 (.Q(\data_out_frame[14] [2]), .C(CLK_c), 
           .D(n29671));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i116 (.Q(\data_out_frame[14] [3]), .C(CLK_c), 
           .D(n29670));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i117 (.Q(\data_out_frame[14] [4]), .C(CLK_c), 
           .D(n29669));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i118 (.Q(\data_out_frame[14] [5]), .C(CLK_c), 
           .D(n29668));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i119 (.Q(\data_out_frame[14] [6]), .C(CLK_c), 
           .D(n29667));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i120 (.Q(\data_out_frame[14] [7]), .C(CLK_c), 
           .D(n29666));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i121 (.Q(\data_out_frame[15] [0]), .C(CLK_c), 
           .D(n29665));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i122 (.Q(\data_out_frame[15] [1]), .C(CLK_c), 
           .D(n29664));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i123 (.Q(\data_out_frame[15] [2]), .C(CLK_c), 
           .D(n29663));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i1_3_lut_4_lut_adj_1327 (.I0(\data_in_frame[1] [2]), .I1(\data_in_frame[3] [4]), 
            .I2(\data_in_frame[3] [5]), .I3(n27350), .O(n44547));
    defparam i1_3_lut_4_lut_adj_1327.LUT_INIT = 16'h6996;
    SB_DFF data_out_frame_0___i124 (.Q(\data_out_frame[15] [3]), .C(CLK_c), 
           .D(n29662));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i125 (.Q(\data_out_frame[15] [4]), .C(CLK_c), 
           .D(n29661));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i126 (.Q(\data_out_frame[15] [5]), .C(CLK_c), 
           .D(n29660));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i127 (.Q(\data_out_frame[15] [6]), .C(CLK_c), 
           .D(n29659));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i128 (.Q(\data_out_frame[15] [7]), .C(CLK_c), 
           .D(n29658));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i129 (.Q(\data_out_frame[16] [0]), .C(CLK_c), 
           .D(n29657));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i130 (.Q(\data_out_frame[16] [1]), .C(CLK_c), 
           .D(n29656));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i131 (.Q(\data_out_frame[16] [2]), .C(CLK_c), 
           .D(n29655));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i132 (.Q(\data_out_frame[16] [3]), .C(CLK_c), 
           .D(n29654));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i133 (.Q(\data_out_frame[16] [4]), .C(CLK_c), 
           .D(n29653));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i134 (.Q(\data_out_frame[16] [5]), .C(CLK_c), 
           .D(n29652));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i135 (.Q(\data_out_frame[16] [6]), .C(CLK_c), 
           .D(n29651));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i7_4_lut_adj_1328 (.I0(n27186), .I1(\data_in[1] [0]), .I2(\data_in[0] [6]), 
            .I3(\data_in[1] [4]), .O(n18));
    defparam i7_4_lut_adj_1328.LUT_INIT = 16'hefff;
    SB_DFF data_out_frame_0___i136 (.Q(\data_out_frame[16] [7]), .C(CLK_c), 
           .D(n29650));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i137 (.Q(\data_out_frame[17] [0]), .C(CLK_c), 
           .D(n29649));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i138 (.Q(\data_out_frame[17] [1]), .C(CLK_c), 
           .D(n29648));   // verilog/coms.v(128[12] 303[6])
    SB_CARRY add_43_5 (.CI(n38556), .I0(\FRAME_MATCHER.i [3]), .I1(GND_net), 
            .CO(n38557));
    SB_LUT4 add_43_4_lut (.I0(n3345), .I1(\FRAME_MATCHER.i [2]), .I2(GND_net), 
            .I3(n38555), .O(n2_adj_4592)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_4_lut.LUT_INIT = 16'h8228;
    SB_DFF data_out_frame_0___i139 (.Q(\data_out_frame[17] [2]), .C(CLK_c), 
           .D(n29647));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i140 (.Q(\data_out_frame[17] [3]), .C(CLK_c), 
           .D(n29646));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i141 (.Q(\data_out_frame[17] [4]), .C(CLK_c), 
           .D(n29645));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i142 (.Q(\data_out_frame[17] [5]), .C(CLK_c), 
           .D(n29644));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i143 (.Q(\data_out_frame[17] [6]), .C(CLK_c), 
           .D(n29643));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i144 (.Q(\data_out_frame[17] [7]), .C(CLK_c), 
           .D(n29642));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i145 (.Q(\data_out_frame[18] [0]), .C(CLK_c), 
           .D(n29641));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i146 (.Q(\data_out_frame[18] [1]), .C(CLK_c), 
           .D(n29640));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i8_4_lut_adj_1329 (.I0(n27136), .I1(\data_in[0] [3]), .I2(\data_in[3] [0]), 
            .I3(\data_in[2] [2]), .O(n19));
    defparam i8_4_lut_adj_1329.LUT_INIT = 16'hfffe;
    SB_DFF data_out_frame_0___i147 (.Q(\data_out_frame[18] [2]), .C(CLK_c), 
           .D(n29639));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i148 (.Q(\data_out_frame[18] [3]), .C(CLK_c), 
           .D(n29638));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i149 (.Q(\data_out_frame[18] [4]), .C(CLK_c), 
           .D(n29637));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i150 (.Q(\data_out_frame[18] [5]), .C(CLK_c), 
           .D(n29636));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i151 (.Q(\data_out_frame[18] [6]), .C(CLK_c), 
           .D(n29635));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i152 (.Q(\data_out_frame[18] [7]), .C(CLK_c), 
           .D(n29634));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i153 (.Q(\data_out_frame[19] [0]), .C(CLK_c), 
           .D(n29633));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i154 (.Q(\data_out_frame[19] [1]), .C(CLK_c), 
           .D(n29632));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i155 (.Q(\data_out_frame[19] [2]), .C(CLK_c), 
           .D(n29631));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i156 (.Q(\data_out_frame[19] [3]), .C(CLK_c), 
           .D(n29630));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i157 (.Q(\data_out_frame[19] [4]), .C(CLK_c), 
           .D(n29629));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i158 (.Q(\data_out_frame[19] [5]), .C(CLK_c), 
           .D(n29628));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i60 (.Q(\data_out_frame[7] [3]), .C(CLK_c), 
           .D(n29104));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i10_4_lut (.I0(n19), .I1(\data_in[2] [4]), .I2(n18), .I3(n12_adj_4712), 
            .O(n63_adj_4652));
    defparam i10_4_lut.LUT_INIT = 16'hfffb;
    SB_LUT4 i6_4_lut_adj_1330 (.I0(\data_in[3] [6]), .I1(\data_in[0] [7]), 
            .I2(\data_in[2] [1]), .I3(n33840), .O(n16_adj_4713));
    defparam i6_4_lut_adj_1330.LUT_INIT = 16'hffef;
    SB_LUT4 i7_4_lut_adj_1331 (.I0(n27136), .I1(\data_in[3] [3]), .I2(\data_in[0] [2]), 
            .I3(\data_in[2] [3]), .O(n17_adj_4714));
    defparam i7_4_lut_adj_1331.LUT_INIT = 16'hbfff;
    SB_LUT4 i9_4_lut_adj_1332 (.I0(n17_adj_4714), .I1(\data_in[3] [1]), 
            .I2(n16_adj_4713), .I3(\data_in[3] [5]), .O(n63_adj_4653));
    defparam i9_4_lut_adj_1332.LUT_INIT = 16'hfbff;
    SB_LUT4 i2_2_lut_adj_1333 (.I0(\data_in[2] [3]), .I1(\data_in[3] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n10_adj_4715));
    defparam i2_2_lut_adj_1333.LUT_INIT = 16'heeee;
    SB_LUT4 i6_4_lut_adj_1334 (.I0(\data_in[0] [2]), .I1(\data_in[3] [3]), 
            .I2(\data_in[3] [1]), .I3(\data_in[0] [7]), .O(n14_adj_4716));
    defparam i6_4_lut_adj_1334.LUT_INIT = 16'hfeff;
    SB_LUT4 i7_4_lut_adj_1335 (.I0(\data_in[3] [6]), .I1(n14_adj_4716), 
            .I2(n10_adj_4715), .I3(\data_in[2] [1]), .O(n27186));
    defparam i7_4_lut_adj_1335.LUT_INIT = 16'hfffd;
    SB_LUT4 i4_4_lut_adj_1336 (.I0(\data_in[1] [7]), .I1(\data_in[0] [0]), 
            .I2(\data_in[1] [1]), .I3(\data_in[0] [4]), .O(n10_adj_4717));
    defparam i4_4_lut_adj_1336.LUT_INIT = 16'hfdff;
    SB_LUT4 i4_4_lut_adj_1337 (.I0(\data_in[2] [2]), .I1(\data_in[1] [5]), 
            .I2(\data_in[1] [4]), .I3(n6_adj_4718), .O(n65));
    defparam i4_4_lut_adj_1337.LUT_INIT = 16'hfff7;
    SB_LUT4 i1_2_lut_adj_1338 (.I0(\data_in[1] [6]), .I1(\data_in[0] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n12_adj_4719));
    defparam i1_2_lut_adj_1338.LUT_INIT = 16'hbbbb;
    SB_LUT4 i7_4_lut_adj_1339 (.I0(n27186), .I1(\data_in[3] [7]), .I2(\data_in[2] [6]), 
            .I3(\data_in[1] [3]), .O(n18_adj_4720));
    defparam i7_4_lut_adj_1339.LUT_INIT = 16'hfeff;
    SB_LUT4 i1_2_lut_3_lut_adj_1340 (.I0(\data_in_frame[1] [2]), .I1(\data_in_frame[3] [4]), 
            .I2(\data_in_frame[1] [3]), .I3(GND_net), .O(n27590));
    defparam i1_2_lut_3_lut_adj_1340.LUT_INIT = 16'h9696;
    SB_DFF data_out_frame_0___i61 (.Q(\data_out_frame[7] [4]), .C(CLK_c), 
           .D(n29102));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i62 (.Q(\data_out_frame[7] [5]), .C(CLK_c), 
           .D(n29101));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i63 (.Q(\data_out_frame[7] [6]), .C(CLK_c), 
           .D(n29100));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i64 (.Q(\data_out_frame[7] [7]), .C(CLK_c), 
           .D(n29099));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i65 (.Q(\data_out_frame[8] [0]), .C(CLK_c), 
           .D(n29098));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i66 (.Q(\data_out_frame[8] [1]), .C(CLK_c), 
           .D(n29097));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i67 (.Q(\data_out_frame[8] [2]), .C(CLK_c), 
           .D(n29096));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i68 (.Q(\data_out_frame[8] [3]), .C(CLK_c), 
           .D(n29095));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i69 (.Q(\data_out_frame[8] [4]), .C(CLK_c), 
           .D(n29094));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i70 (.Q(\data_out_frame[8] [5]), .C(CLK_c), 
           .D(n29093));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i71 (.Q(\data_out_frame[8] [6]), .C(CLK_c), 
           .D(n29092));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i72 (.Q(\data_out_frame[8] [7]), .C(CLK_c), 
           .D(n29091));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i73 (.Q(\data_out_frame[9] [0]), .C(CLK_c), 
           .D(n29090));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i74 (.Q(\data_out_frame[9] [1]), .C(CLK_c), 
           .D(n29089));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i75 (.Q(\data_out_frame[9] [2]), .C(CLK_c), 
           .D(n29088));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i76 (.Q(\data_out_frame[9] [3]), .C(CLK_c), 
           .D(n29087));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i77 (.Q(\data_out_frame[9] [4]), .C(CLK_c), 
           .D(n29086));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i78 (.Q(\data_out_frame[9] [5]), .C(CLK_c), 
           .D(n29085));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i79 (.Q(\data_out_frame[9] [6]), .C(CLK_c), 
           .D(n29084));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i80 (.Q(\data_out_frame[9] [7]), .C(CLK_c), 
           .D(n29083));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i81 (.Q(\data_out_frame[10] [0]), .C(CLK_c), 
           .D(n29082));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i82 (.Q(\data_out_frame[10] [1]), .C(CLK_c), 
           .D(n29081));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i83 (.Q(\data_out_frame[10] [2]), .C(CLK_c), 
           .D(n29080));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i84 (.Q(\data_out_frame[10] [3]), .C(CLK_c), 
           .D(n29079));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i85 (.Q(\data_out_frame[10] [4]), .C(CLK_c), 
           .D(n29078));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i86 (.Q(\data_out_frame[10] [5]), .C(CLK_c), 
           .D(n29077));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i87 (.Q(\data_out_frame[10] [6]), .C(CLK_c), 
           .D(n29076));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i88 (.Q(\data_out_frame[10] [7]), .C(CLK_c), 
           .D(n29075));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i89 (.Q(\data_out_frame[11] [0]), .C(CLK_c), 
           .D(n29074));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i15465_3_lut_4_lut (.I0(n8_adj_4655), .I1(n43832), .I2(rx_data[7]), 
            .I3(\data_in_frame[3] [7]), .O(n29413));
    defparam i15465_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFFESR driver_enable_4015 (.Q(DE_c), .C(CLK_c), .E(n44841), .D(n7477), 
            .R(n45285));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i32452_4_lut (.I0(\data_in[2] [0]), .I1(\data_in[2] [5]), .I2(\data_in[1] [2]), 
            .I3(\data_in[3] [2]), .O(n47977));
    defparam i32452_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i10_4_lut_adj_1341 (.I0(n47977), .I1(\data_in[0] [5]), .I2(n18_adj_4720), 
            .I3(n12_adj_4719), .O(n62));
    defparam i10_4_lut_adj_1341.LUT_INIT = 16'hfff7;
    SB_LUT4 i5777_2_lut (.I0(n63_adj_4653), .I1(n63_adj_4652), .I2(GND_net), 
            .I3(GND_net), .O(n19692));   // verilog/coms.v(140[4] 142[7])
    defparam i5777_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i15466_3_lut_4_lut (.I0(n8_adj_4655), .I1(n43832), .I2(rx_data[6]), 
            .I3(\data_in_frame[3] [6]), .O(n29414));
    defparam i15466_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15467_3_lut_4_lut (.I0(n8_adj_4655), .I1(n43832), .I2(rx_data[5]), 
            .I3(\data_in_frame[3] [5]), .O(n29415));
    defparam i15467_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_out_frame_0___i90 (.Q(\data_out_frame[11] [1]), .C(CLK_c), 
           .D(n29067));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i91 (.Q(\data_out_frame[11] [2]), .C(CLK_c), 
           .D(n29065));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i92 (.Q(\data_out_frame[11] [3]), .C(CLK_c), 
           .D(n29064));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i93 (.Q(\data_out_frame[11] [4]), .C(CLK_c), 
           .D(n29063));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i94 (.Q(\data_out_frame[11] [5]), .C(CLK_c), 
           .D(n29062));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i95 (.Q(\data_out_frame[11] [6]), .C(CLK_c), 
           .D(n29061));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i96 (.Q(\data_out_frame[11] [7]), .C(CLK_c), 
           .D(n29060));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i97 (.Q(\data_out_frame[12] [0]), .C(CLK_c), 
           .D(n29056));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i159 (.Q(\data_out_frame[19] [6]), .C(CLK_c), 
           .D(n29627));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i18_4_lut_adj_1342 (.I0(\FRAME_MATCHER.i [24]), .I1(\FRAME_MATCHER.i [11]), 
            .I2(\FRAME_MATCHER.i [28]), .I3(\FRAME_MATCHER.i [16]), .O(n44_adj_4721));
    defparam i18_4_lut_adj_1342.LUT_INIT = 16'hfffe;
    SB_DFFESR LED_4014 (.Q(LED_c), .C(CLK_c), .E(n43762), .D(n28824), 
            .R(n45257));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i160 (.Q(\data_out_frame[19] [7]), .C(CLK_c), 
           .D(n29626));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i15468_3_lut_4_lut (.I0(n8_adj_4655), .I1(n43832), .I2(rx_data[4]), 
            .I3(\data_in_frame[3] [4]), .O(n29416));
    defparam i15468_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15469_3_lut_4_lut (.I0(n8_adj_4655), .I1(n43832), .I2(rx_data[3]), 
            .I3(\data_in_frame[3] [3]), .O(n29417));
    defparam i15469_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 select_686_Select_1_i3_2_lut (.I0(\FRAME_MATCHER.i [1]), .I1(n4141), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4595));
    defparam select_686_Select_1_i3_2_lut.LUT_INIT = 16'h8888;
    SB_DFF data_out_frame_0___i161 (.Q(\data_out_frame[20] [0]), .C(CLK_c), 
           .D(n29625));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i162 (.Q(\data_out_frame[20] [1]), .C(CLK_c), 
           .D(n29624));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i163 (.Q(\data_out_frame[20] [2]), .C(CLK_c), 
           .D(n29623));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i164 (.Q(\data_out_frame[20] [3]), .C(CLK_c), 
           .D(n29622));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i165 (.Q(\data_out_frame[20] [4]), .C(CLK_c), 
           .D(n29621));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i166 (.Q(\data_out_frame[20] [5]), .C(CLK_c), 
           .D(n29620));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i167 (.Q(\data_out_frame[20] [6]), .C(CLK_c), 
           .D(n29619));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_35839 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[22] [7]), .I2(\data_out_frame[23] [7]), 
            .I3(byte_transmit_counter[1]), .O(n51318));
    defparam byte_transmit_counter_0__bdd_4_lut_35839.LUT_INIT = 16'he4aa;
    SB_DFF data_out_frame_0___i168 (.Q(\data_out_frame[20] [7]), .C(CLK_c), 
           .D(n29618));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 n51318_bdd_4_lut (.I0(n51318), .I1(\data_out_frame[21] [7]), 
            .I2(\data_out_frame[20] [7]), .I3(byte_transmit_counter[1]), 
            .O(n51321));
    defparam n51318_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF data_out_frame_0___i169 (.Q(\data_out_frame[21] [0]), .C(CLK_c), 
           .D(n29617));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i170 (.Q(\data_out_frame[21] [1]), .C(CLK_c), 
           .D(n29616));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut (.I0(byte_transmit_counter[1]), 
            .I1(n48221), .I2(n48222), .I3(byte_transmit_counter[2]), .O(n51312));
    defparam byte_transmit_counter_1__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_DFF data_out_frame_0___i171 (.Q(\data_out_frame[21] [2]), .C(CLK_c), 
           .D(n29615));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 n51312_bdd_4_lut (.I0(n51312), .I1(n48228), .I2(n48227), .I3(byte_transmit_counter[2]), 
            .O(n51315));
    defparam n51312_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF data_out_frame_0___i172 (.Q(\data_out_frame[21] [3]), .C(CLK_c), 
           .D(n29614));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i173 (.Q(\data_out_frame[21] [4]), .C(CLK_c), 
           .D(n29613));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_35706 (.I0(byte_transmit_counter[1]), 
            .I1(n48062), .I2(n48063), .I3(byte_transmit_counter[2]), .O(n51306));
    defparam byte_transmit_counter_1__bdd_4_lut_35706.LUT_INIT = 16'he4aa;
    SB_DFF data_out_frame_0___i174 (.Q(\data_out_frame[21] [5]), .C(CLK_c), 
           .D(n29612));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 n51306_bdd_4_lut (.I0(n51306), .I1(n48138), .I2(n48137), .I3(byte_transmit_counter[2]), 
            .O(n51309));
    defparam n51306_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF data_out_frame_0___i175 (.Q(\data_out_frame[21] [6]), .C(CLK_c), 
           .D(n29611));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i176 (.Q(\data_out_frame[21] [7]), .C(CLK_c), 
           .D(n29610));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_35701 (.I0(byte_transmit_counter[1]), 
            .I1(n48101), .I2(n48102), .I3(byte_transmit_counter[2]), .O(n51300));
    defparam byte_transmit_counter_1__bdd_4_lut_35701.LUT_INIT = 16'he4aa;
    SB_DFF data_out_frame_0___i177 (.Q(\data_out_frame[22] [0]), .C(CLK_c), 
           .D(n29609));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 n51300_bdd_4_lut (.I0(n51300), .I1(n48129), .I2(n48128), .I3(byte_transmit_counter[2]), 
            .O(n51303));
    defparam n51300_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF data_out_frame_0___i178 (.Q(\data_out_frame[22] [1]), .C(CLK_c), 
           .D(n29608));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i179 (.Q(\data_out_frame[22] [2]), .C(CLK_c), 
           .D(n29607));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_35696 (.I0(byte_transmit_counter[1]), 
            .I1(n48131), .I2(n48132), .I3(byte_transmit_counter[2]), .O(n51294));
    defparam byte_transmit_counter_1__bdd_4_lut_35696.LUT_INIT = 16'he4aa;
    SB_DFF data_out_frame_0___i180 (.Q(\data_out_frame[22] [3]), .C(CLK_c), 
           .D(n29606));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i181 (.Q(\data_out_frame[22] [4]), .C(CLK_c), 
           .D(n29605));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i182 (.Q(\data_out_frame[22] [5]), .C(CLK_c), 
           .D(n29604));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i190 (.Q(\data_in_frame[23] [5]), .C(CLK_c), 
           .D(n29603));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i183 (.Q(\data_out_frame[22] [6]), .C(CLK_c), 
           .D(n29602));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 n51294_bdd_4_lut (.I0(n51294), .I1(n48123), .I2(n48122), .I3(byte_transmit_counter[2]), 
            .O(n51297));
    defparam n51294_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF data_in_frame_0__i192 (.Q(\data_in_frame[23] [7]), .C(CLK_c), 
           .D(n29601));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i191 (.Q(\data_in_frame[23] [6]), .C(CLK_c), 
           .D(n29600));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_35691 (.I0(byte_transmit_counter[1]), 
            .I1(n48110), .I2(n48111), .I3(byte_transmit_counter[2]), .O(n51288));
    defparam byte_transmit_counter_1__bdd_4_lut_35691.LUT_INIT = 16'he4aa;
    SB_DFF control_mode_i0_i1 (.Q(control_mode[1]), .C(CLK_c), .D(n29599));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 n51288_bdd_4_lut (.I0(n51288), .I1(n48105), .I2(n48104), .I3(byte_transmit_counter[2]), 
            .O(n51291));
    defparam n51288_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF control_mode_i0_i2 (.Q(control_mode[2]), .C(CLK_c), .D(n29598));   // verilog/coms.v(128[12] 303[6])
    SB_DFF control_mode_i0_i3 (.Q(control_mode[3]), .C(CLK_c), .D(n29597));   // verilog/coms.v(128[12] 303[6])
    SB_DFF control_mode_i0_i4 (.Q(control_mode[4]), .C(CLK_c), .D(n29596));   // verilog/coms.v(128[12] 303[6])
    SB_DFF control_mode_i0_i5 (.Q(control_mode[5]), .C(CLK_c), .D(n29595));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i98 (.Q(\data_out_frame[12] [1]), .C(CLK_c), 
           .D(n29055));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i99 (.Q(\data_out_frame[12] [2]), .C(CLK_c), 
           .D(n29050));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i100 (.Q(\data_out_frame[12] [3]), .C(CLK_c), 
           .D(n29049));   // verilog/coms.v(128[12] 303[6])
    SB_DFF \FRAME_MATCHER.state_i0  (.Q(\FRAME_MATCHER.state [0]), .C(CLK_c), 
           .D(n43142));   // verilog/coms.v(128[12] 303[6])
    SB_DFF PWMLimit_i0_i0 (.Q(PWMLimit[0]), .C(CLK_c), .D(n29047));   // verilog/coms.v(128[12] 303[6])
    SB_DFF current_limit_i0_i0 (.Q(current_limit[0]), .C(CLK_c), .D(n29046));   // verilog/coms.v(128[12] 303[6])
    SB_DFF control_mode_i0_i0 (.Q(control_mode[0]), .C(CLK_c), .D(n29045));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i1 (.Q(\data_in_frame[0] [0]), .C(CLK_c), .D(n29044));   // verilog/coms.v(128[12] 303[6])
    SB_DFF neopxl_color_i0_i0 (.Q(neopxl_color[0]), .C(CLK_c), .D(n29043));   // verilog/coms.v(128[12] 303[6])
    SB_DFF Ki_i0 (.Q(\Ki[0] ), .C(CLK_c), .D(n29042));   // verilog/coms.v(128[12] 303[6])
    SB_DFF Kp_i0 (.Q(\Kp[0] ), .C(CLK_c), .D(n29041));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_0___i1 (.Q(\data_in[0] [0]), .C(CLK_c), .D(n29040));   // verilog/coms.v(128[12] 303[6])
    SB_DFF IntegralLimit_i0_i0 (.Q(IntegralLimit[0]), .C(CLK_c), .D(n29026));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i16_4_lut_adj_1343 (.I0(\FRAME_MATCHER.i [19]), .I1(\FRAME_MATCHER.i [22]), 
            .I2(\FRAME_MATCHER.i [25]), .I3(\FRAME_MATCHER.i [18]), .O(n42_adj_4722));
    defparam i16_4_lut_adj_1343.LUT_INIT = 16'hfffe;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut (.I0(byte_transmit_counter[3]), 
            .I1(n50140), .I2(n49345), .I3(byte_transmit_counter[4]), .O(n51552));
    defparam byte_transmit_counter_3__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_DFF control_mode_i0_i6 (.Q(control_mode[6]), .C(CLK_c), .D(n29594));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i17_4_lut_adj_1344 (.I0(\FRAME_MATCHER.i [29]), .I1(\FRAME_MATCHER.i [17]), 
            .I2(\FRAME_MATCHER.i [30]), .I3(\FRAME_MATCHER.i [21]), .O(n43_adj_4723));
    defparam i17_4_lut_adj_1344.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut_adj_1345 (.I0(\FRAME_MATCHER.i [6]), .I1(\FRAME_MATCHER.i [8]), 
            .I2(\FRAME_MATCHER.i [23]), .I3(\FRAME_MATCHER.i [5]), .O(n41));
    defparam i15_4_lut_adj_1345.LUT_INIT = 16'hfffe;
    SB_LUT4 i14_4_lut (.I0(\FRAME_MATCHER.i [13]), .I1(\FRAME_MATCHER.i [15]), 
            .I2(\FRAME_MATCHER.i [10]), .I3(\FRAME_MATCHER.i [26]), .O(n40));
    defparam i14_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_2_lut (.I0(\FRAME_MATCHER.i [9]), .I1(\FRAME_MATCHER.i [27]), 
            .I2(GND_net), .I3(GND_net), .O(n39));
    defparam i13_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i24_4_lut (.I0(n41), .I1(n43_adj_4723), .I2(n42_adj_4722), 
            .I3(n44_adj_4721), .O(n50));
    defparam i24_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_4_lut (.I0(\data_out_frame[25] [3]), .I1(\data_out_frame[25] [4]), 
            .I2(n41682), .I3(n25338), .O(n44446));
    defparam i1_2_lut_4_lut.LUT_INIT = 16'h9669;
    SB_LUT4 i19_4_lut_adj_1346 (.I0(\FRAME_MATCHER.i [14]), .I1(\FRAME_MATCHER.i [12]), 
            .I2(\FRAME_MATCHER.i [20]), .I3(\FRAME_MATCHER.i [7]), .O(n45_adj_4724));
    defparam i19_4_lut_adj_1346.LUT_INIT = 16'hfffe;
    SB_LUT4 i25_4_lut_adj_1347 (.I0(n45_adj_4724), .I1(n50), .I2(n39), 
            .I3(n40), .O(n27189));
    defparam i25_4_lut_adj_1347.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_adj_1348 (.I0(\FRAME_MATCHER.i [4]), .I1(n27189), .I2(GND_net), 
            .I3(GND_net), .O(n27025));   // verilog/coms.v(155[7:23])
    defparam i1_2_lut_adj_1348.LUT_INIT = 16'heeee;
    SB_LUT4 i3_2_lut_3_lut (.I0(\data_out_frame[20] [6]), .I1(\data_out_frame[23] [2]), 
            .I2(n44175), .I3(GND_net), .O(n11_adj_4725));
    defparam i3_2_lut_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_4_lut_adj_1349 (.I0(n26888), .I1(\data_out_frame[11] [5]), 
            .I2(\data_out_frame[15] [7]), .I3(n44275), .O(n44254));
    defparam i1_2_lut_4_lut_adj_1349.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1350 (.I0(\data_out_frame[13] [6]), .I1(n44583), 
            .I2(\data_out_frame[11] [4]), .I3(n25208), .O(n44275));
    defparam i1_2_lut_4_lut_adj_1350.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1351 (.I0(\data_out_frame[4] [3]), .I1(\data_out_frame[4] [4]), 
            .I2(\data_out_frame[6] [5]), .I3(GND_net), .O(n27745));
    defparam i1_2_lut_3_lut_adj_1351.LUT_INIT = 16'h9696;
    SB_LUT4 i15470_3_lut_4_lut (.I0(n8_adj_4655), .I1(n43832), .I2(rx_data[2]), 
            .I3(\data_in_frame[3] [2]), .O(n29418));
    defparam i15470_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_4_lut (.I0(\data_in_frame[18] [7]), .I1(\data_in_frame[18] [6]), 
            .I2(\data_in_frame[18] [2]), .I3(\data_in_frame[18] [4]), .O(n44559));   // verilog/coms.v(79[16:27])
    defparam i1_2_lut_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_DFF control_mode_i0_i7 (.Q(control_mode[7]), .C(CLK_c), .D(n29593));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i4_4_lut_adj_1352 (.I0(n27227), .I1(n8_adj_4726), .I2(\FRAME_MATCHER.state [2]), 
            .I3(n57), .O(n4120));
    defparam i4_4_lut_adj_1352.LUT_INIT = 16'h8808;
    SB_LUT4 i15471_3_lut_4_lut (.I0(n8_adj_4655), .I1(n43832), .I2(rx_data[1]), 
            .I3(\data_in_frame[3] [1]), .O(n29419));
    defparam i15471_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF current_limit_i0_i1 (.Q(current_limit[1]), .C(CLK_c), .D(n29592));   // verilog/coms.v(128[12] 303[6])
    SB_DFF current_limit_i0_i2 (.Q(current_limit[2]), .C(CLK_c), .D(n29591));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i20865_4_lut (.I0(n5_adj_4727), .I1(\FRAME_MATCHER.i [31]), 
            .I2(\FRAME_MATCHER.i [2]), .I3(\FRAME_MATCHER.i [3]), .O(n771));   // verilog/coms.v(158[9:60])
    defparam i20865_4_lut.LUT_INIT = 16'h3332;
    SB_DFF current_limit_i0_i3 (.Q(current_limit[3]), .C(CLK_c), .D(n29590));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i101 (.Q(\data_out_frame[12] [4]), .C(CLK_c), 
           .D(n29024));   // verilog/coms.v(128[12] 303[6])
    SB_DFF current_limit_i0_i4 (.Q(current_limit[4]), .C(CLK_c), .D(n29589));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i102 (.Q(\data_out_frame[12] [5]), .C(CLK_c), 
           .D(n29023));   // verilog/coms.v(128[12] 303[6])
    SB_DFF current_limit_i0_i5 (.Q(current_limit[5]), .C(CLK_c), .D(n29588));   // verilog/coms.v(128[12] 303[6])
    SB_DFF current_limit_i0_i6 (.Q(current_limit[6]), .C(CLK_c), .D(n29587));   // verilog/coms.v(128[12] 303[6])
    SB_DFF current_limit_i0_i7 (.Q(current_limit[7]), .C(CLK_c), .D(n29586));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i15472_3_lut_4_lut (.I0(n8_adj_4655), .I1(n43832), .I2(rx_data[0]), 
            .I3(\data_in_frame[3] [0]), .O(n29420));
    defparam i15472_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF current_limit_i0_i8 (.Q(current_limit[8]), .C(CLK_c), .D(n29585));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i1_2_lut_3_lut_adj_1353 (.I0(\data_out_frame[19] [5]), .I1(n41472), 
            .I2(n41816), .I3(GND_net), .O(n44571));
    defparam i1_2_lut_3_lut_adj_1353.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_4_lut_adj_1354 (.I0(n43861), .I1(n44015), .I2(n10_adj_4728), 
            .I3(\data_out_frame[9] [1]), .O(n44287));
    defparam i1_2_lut_4_lut_adj_1354.LUT_INIT = 16'h6996;
    SB_LUT4 i1_3_lut_adj_1355 (.I0(n4120), .I1(n27235), .I2(n2263), .I3(GND_net), 
            .O(n43850));
    defparam i1_3_lut_adj_1355.LUT_INIT = 16'hbaba;
    SB_LUT4 i1_2_lut_3_lut_adj_1356 (.I0(\data_out_frame[15] [6]), .I1(\data_out_frame[15] [4]), 
            .I2(\data_out_frame[15] [3]), .I3(GND_net), .O(n44084));
    defparam i1_2_lut_3_lut_adj_1356.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1357 (.I0(\FRAME_MATCHER.state [1]), .I1(n27230), 
            .I2(GND_net), .I3(GND_net), .O(n27232));   // verilog/coms.v(152[5:27])
    defparam i1_2_lut_adj_1357.LUT_INIT = 16'heeee;
    SB_LUT4 i20866_4_lut (.I0(n8_adj_4729), .I1(\FRAME_MATCHER.i [31]), 
            .I2(n27025), .I3(\FRAME_MATCHER.i [3]), .O(n3303));   // verilog/coms.v(228[9:54])
    defparam i20866_4_lut.LUT_INIT = 16'h3230;
    SB_LUT4 i2_3_lut_4_lut_adj_1358 (.I0(\data_out_frame[13] [0]), .I1(n26718), 
            .I2(\data_out_frame[17] [4]), .I3(\data_out_frame[15] [2]), 
            .O(n44435));
    defparam i2_3_lut_4_lut_adj_1358.LUT_INIT = 16'h6996;
    SB_LUT4 n51552_bdd_4_lut (.I0(n51552), .I1(n51267), .I2(n7_adj_4730), 
            .I3(byte_transmit_counter[4]), .O(tx_data[7]));
    defparam n51552_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_3_lut_adj_1359 (.I0(n55), .I1(n43859), .I2(n3303), .I3(GND_net), 
            .O(n4_adj_4731));
    defparam i1_3_lut_adj_1359.LUT_INIT = 16'hcdcd;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_35903 (.I0(byte_transmit_counter[3]), 
            .I1(n51213), .I2(n49354), .I3(byte_transmit_counter[4]), .O(n51546));
    defparam byte_transmit_counter_3__bdd_4_lut_35903.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_4_lut_adj_1360 (.I0(\FRAME_MATCHER.state [0]), .I1(n44726), 
            .I2(n27061), .I3(n4_adj_4731), .O(n17_adj_4732));   // verilog/coms.v(202[5:24])
    defparam i1_4_lut_adj_1360.LUT_INIT = 16'haf23;
    SB_DFF current_limit_i0_i9 (.Q(current_limit[9]), .C(CLK_c), .D(n29584));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i1_4_lut_adj_1361 (.I0(\FRAME_MATCHER.state [3]), .I1(n17_adj_4732), 
            .I2(n44728), .I3(\FRAME_MATCHER.state [2]), .O(n43142));   // verilog/coms.v(202[5:24])
    defparam i1_4_lut_adj_1361.LUT_INIT = 16'hccce;
    SB_DFF current_limit_i0_i10 (.Q(current_limit[10]), .C(CLK_c), .D(n29583));   // verilog/coms.v(128[12] 303[6])
    SB_DFF current_limit_i0_i11 (.Q(current_limit[11]), .C(CLK_c), .D(n29582));   // verilog/coms.v(128[12] 303[6])
    SB_DFF current_limit_i0_i12 (.Q(current_limit[12]), .C(CLK_c), .D(n29581));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i1_2_lut_adj_1362 (.I0(\data_in_frame[13] [1]), .I1(n45300), 
            .I2(GND_net), .I3(GND_net), .O(n44161));
    defparam i1_2_lut_adj_1362.LUT_INIT = 16'h9999;
    SB_DFF current_limit_i0_i13 (.Q(current_limit[13]), .C(CLK_c), .D(n29580));   // verilog/coms.v(128[12] 303[6])
    SB_DFF current_limit_i0_i14 (.Q(current_limit[14]), .C(CLK_c), .D(n29579));   // verilog/coms.v(128[12] 303[6])
    SB_DFF current_limit_i0_i15 (.Q(current_limit[15]), .C(CLK_c), .D(n29578));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i1_2_lut_3_lut_adj_1363 (.I0(\data_out_frame[20] [4]), .I1(n41801), 
            .I2(n40636), .I3(GND_net), .O(n44257));
    defparam i1_2_lut_3_lut_adj_1363.LUT_INIT = 16'h6969;
    SB_LUT4 i15457_3_lut_4_lut (.I0(n8_adj_4681), .I1(n43832), .I2(rx_data[7]), 
            .I3(\data_in_frame[4] [7]), .O(n29405));
    defparam i15457_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF PWMLimit_i0_i1 (.Q(PWMLimit[1]), .C(CLK_c), .D(n29577));   // verilog/coms.v(128[12] 303[6])
    SB_DFF PWMLimit_i0_i2 (.Q(PWMLimit[2]), .C(CLK_c), .D(n29576));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i15458_3_lut_4_lut (.I0(n8_adj_4681), .I1(n43832), .I2(rx_data[6]), 
            .I3(\data_in_frame[4] [6]), .O(n29406));
    defparam i15458_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_4_lut_adj_1364 (.I0(\data_out_frame[20] [6]), .I1(\data_out_frame[20] [7]), 
            .I2(\data_out_frame[20] [5]), .I3(\data_out_frame[20] [1]), 
            .O(n43905));
    defparam i1_2_lut_4_lut_adj_1364.LUT_INIT = 16'h6996;
    SB_DFFE setpoint__i23 (.Q(setpoint[23]), .C(CLK_c), .E(n28531), .D(n7593));   // verilog/coms.v(128[12] 303[6])
    SB_DFFE setpoint__i22 (.Q(setpoint[22]), .C(CLK_c), .E(n28531), .D(n7592));   // verilog/coms.v(128[12] 303[6])
    SB_DFFE setpoint__i21 (.Q(setpoint[21]), .C(CLK_c), .E(n28531), .D(n7591));   // verilog/coms.v(128[12] 303[6])
    SB_DFFE setpoint__i20 (.Q(setpoint[20]), .C(CLK_c), .E(n28531), .D(n7590));   // verilog/coms.v(128[12] 303[6])
    SB_DFFE setpoint__i19 (.Q(setpoint[19]), .C(CLK_c), .E(n28531), .D(n7589));   // verilog/coms.v(128[12] 303[6])
    SB_DFFE setpoint__i18 (.Q(setpoint[18]), .C(CLK_c), .E(n28531), .D(n7588));   // verilog/coms.v(128[12] 303[6])
    SB_DFFE setpoint__i17 (.Q(setpoint[17]), .C(CLK_c), .E(n28531), .D(n7587));   // verilog/coms.v(128[12] 303[6])
    SB_DFFE setpoint__i16 (.Q(setpoint[16]), .C(CLK_c), .E(n28531), .D(n7586));   // verilog/coms.v(128[12] 303[6])
    SB_DFFE setpoint__i15 (.Q(setpoint[15]), .C(CLK_c), .E(n28531), .D(n7585));   // verilog/coms.v(128[12] 303[6])
    SB_DFFE setpoint__i14 (.Q(setpoint[14]), .C(CLK_c), .E(n28531), .D(n7584));   // verilog/coms.v(128[12] 303[6])
    SB_DFFE setpoint__i13 (.Q(setpoint[13]), .C(CLK_c), .E(n28531), .D(n7583));   // verilog/coms.v(128[12] 303[6])
    SB_DFFE setpoint__i12 (.Q(setpoint[12]), .C(CLK_c), .E(n28531), .D(n7582));   // verilog/coms.v(128[12] 303[6])
    SB_DFFE setpoint__i11 (.Q(setpoint[11]), .C(CLK_c), .E(n28531), .D(n7581));   // verilog/coms.v(128[12] 303[6])
    SB_DFFE setpoint__i10 (.Q(setpoint[10]), .C(CLK_c), .E(n28531), .D(n7580));   // verilog/coms.v(128[12] 303[6])
    SB_DFFE setpoint__i9 (.Q(setpoint[9]), .C(CLK_c), .E(n28531), .D(n7579));   // verilog/coms.v(128[12] 303[6])
    SB_DFFE setpoint__i8 (.Q(setpoint[8]), .C(CLK_c), .E(n28531), .D(n7578));   // verilog/coms.v(128[12] 303[6])
    SB_DFFE setpoint__i7 (.Q(setpoint[7]), .C(CLK_c), .E(n28531), .D(n7577));   // verilog/coms.v(128[12] 303[6])
    SB_DFFE setpoint__i6 (.Q(setpoint[6]), .C(CLK_c), .E(n28531), .D(n7576));   // verilog/coms.v(128[12] 303[6])
    SB_DFFE setpoint__i5 (.Q(setpoint[5]), .C(CLK_c), .E(n28531), .D(n7575));   // verilog/coms.v(128[12] 303[6])
    SB_DFFE setpoint__i4 (.Q(setpoint[4]), .C(CLK_c), .E(n28531), .D(n7574));   // verilog/coms.v(128[12] 303[6])
    SB_DFFE setpoint__i3 (.Q(setpoint[3]), .C(CLK_c), .E(n28531), .D(n7573));   // verilog/coms.v(128[12] 303[6])
    SB_DFFE setpoint__i2 (.Q(setpoint[2]), .C(CLK_c), .E(n28531), .D(n7572));   // verilog/coms.v(128[12] 303[6])
    SB_DFFE setpoint__i1 (.Q(setpoint[1]), .C(CLK_c), .E(n28531), .D(n7571));   // verilog/coms.v(128[12] 303[6])
    SB_DFFSS \FRAME_MATCHER.state_i31  (.Q(\FRAME_MATCHER.state [31]), .C(CLK_c), 
            .D(n43210), .S(n43086));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i15459_3_lut_4_lut (.I0(n8_adj_4681), .I1(n43832), .I2(rx_data[5]), 
            .I3(\data_in_frame[4] [5]), .O(n29407));
    defparam i15459_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15460_3_lut_4_lut (.I0(n8_adj_4681), .I1(n43832), .I2(rx_data[4]), 
            .I3(\data_in_frame[4] [4]), .O(n29408));
    defparam i15460_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_35686 (.I0(byte_transmit_counter[1]), 
            .I1(n48191), .I2(n48192), .I3(byte_transmit_counter[2]), .O(n51276));
    defparam byte_transmit_counter_1__bdd_4_lut_35686.LUT_INIT = 16'he4aa;
    SB_LUT4 i15461_3_lut_4_lut (.I0(n8_adj_4681), .I1(n43832), .I2(rx_data[3]), 
            .I3(\data_in_frame[4] [3]), .O(n29409));
    defparam i15461_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 n51474_bdd_4_lut (.I0(n51474), .I1(\data_out_frame[25] [3]), 
            .I2(\data_out_frame[24] [3]), .I3(byte_transmit_counter[1]), 
            .O(n51477));
    defparam n51474_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i15462_3_lut_4_lut (.I0(n8_adj_4681), .I1(n43832), .I2(rx_data[2]), 
            .I3(\data_in_frame[4] [2]), .O(n29410));
    defparam i15462_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_4_lut_adj_1365 (.I0(n27901), .I1(\data_out_frame[20] [5]), 
            .I2(n41801), .I3(n44257), .O(n41615));
    defparam i2_3_lut_4_lut_adj_1365.LUT_INIT = 16'h6996;
    SB_LUT4 i15463_3_lut_4_lut (.I0(n8_adj_4681), .I1(n43832), .I2(rx_data[1]), 
            .I3(\data_in_frame[4] [1]), .O(n29411));
    defparam i15463_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i32517_3_lut (.I0(\data_out_frame[8] [3]), .I1(\data_out_frame[9] [3]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n48104));
    defparam i32517_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15464_3_lut_4_lut (.I0(n8_adj_4681), .I1(n43832), .I2(rx_data[0]), 
            .I3(\data_in_frame[4] [0]), .O(n29412));
    defparam i15464_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i32518_3_lut (.I0(\data_out_frame[10] [3]), .I1(\data_out_frame[11] [3]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n48105));
    defparam i32518_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i32524_3_lut (.I0(\data_out_frame[14] [3]), .I1(\data_out_frame[15] [3]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n48111));
    defparam i32524_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF PWMLimit_i0_i3 (.Q(PWMLimit[3]), .C(CLK_c), .D(n29575));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i32523_3_lut (.I0(\data_out_frame[12] [3]), .I1(\data_out_frame[13] [3]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n48110));
    defparam i32523_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1366 (.I0(\data_in_frame[9] [7]), .I1(\data_in_frame[9] [6]), 
            .I2(n27544), .I3(n27554), .O(n28009));   // verilog/coms.v(86[17:28])
    defparam i1_2_lut_3_lut_4_lut_adj_1366.LUT_INIT = 16'h6996;
    SB_LUT4 i32535_3_lut (.I0(\data_out_frame[8] [4]), .I1(\data_out_frame[9] [4]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n48122));
    defparam i32535_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 equal_312_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8_adj_4681));   // verilog/coms.v(155[7:23])
    defparam equal_312_i8_2_lut_3_lut.LUT_INIT = 16'hfbfb;
    SB_LUT4 i32536_3_lut (.I0(\data_out_frame[10] [4]), .I1(\data_out_frame[11] [4]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n48123));
    defparam i32536_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14_2_lut (.I0(rx_data_ready), .I1(\FRAME_MATCHER.rx_data_ready_prev ), 
            .I2(GND_net), .I3(GND_net), .O(n161));   // verilog/coms.v(154[9:50])
    defparam i14_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i2_2_lut_3_lut (.I0(\data_out_frame[16] [0]), .I1(\data_out_frame[18] [1]), 
            .I2(n27885), .I3(GND_net), .O(n10_adj_4733));
    defparam i2_2_lut_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1367 (.I0(n27820), .I1(n27850), .I2(\data_in_frame[8] [7]), 
            .I3(n27933), .O(n44528));   // verilog/coms.v(74[16:42])
    defparam i1_2_lut_3_lut_4_lut_adj_1367.LUT_INIT = 16'h6996;
    SB_DFF PWMLimit_i0_i4 (.Q(PWMLimit[4]), .C(CLK_c), .D(n29574));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i3_4_lut_adj_1368 (.I0(n35014), .I1(\FRAME_MATCHER.i [5]), .I2(\FRAME_MATCHER.i [4]), 
            .I3(\FRAME_MATCHER.i [3]), .O(n43820));   // verilog/coms.v(155[7:23])
    defparam i3_4_lut_adj_1368.LUT_INIT = 16'hffdf;
    SB_LUT4 i2_2_lut_3_lut_4_lut (.I0(\data_in_frame[6] [7]), .I1(\data_in_frame[6] [6]), 
            .I2(n44394), .I3(n27948), .O(n10_adj_4734));   // verilog/coms.v(86[17:28])
    defparam i2_2_lut_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 n51546_bdd_4_lut (.I0(n51546), .I1(n51309), .I2(n7_adj_4735), 
            .I3(byte_transmit_counter[4]), .O(tx_data[6]));
    defparam n51546_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF PWMLimit_i0_i5 (.Q(PWMLimit[5]), .C(CLK_c), .D(n29573));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1369 (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(n43832), .I3(\FRAME_MATCHER.i [0]), .O(n43838));   // verilog/coms.v(155[7:23])
    defparam i1_2_lut_3_lut_4_lut_adj_1369.LUT_INIT = 16'hfbff;
    SB_LUT4 i1_2_lut_4_lut_adj_1370 (.I0(\data_out_frame[23] [4]), .I1(\data_out_frame[23] [6]), 
            .I2(n27406), .I3(\data_out_frame[24] [3]), .O(n30));
    defparam i1_2_lut_4_lut_adj_1370.LUT_INIT = 16'h6996;
    SB_DFF PWMLimit_i0_i6 (.Q(PWMLimit[6]), .C(CLK_c), .D(n29572));   // verilog/coms.v(128[12] 303[6])
    SB_DFF PWMLimit_i0_i7 (.Q(PWMLimit[7]), .C(CLK_c), .D(n29571));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1371 (.I0(\FRAME_MATCHER.state [1]), 
            .I1(\FRAME_MATCHER.state [2]), .I2(\FRAME_MATCHER.state [0]), 
            .I3(n27004), .O(n27235));
    defparam i1_2_lut_3_lut_4_lut_adj_1371.LUT_INIT = 16'hff7f;
    SB_DFF PWMLimit_i0_i8 (.Q(PWMLimit[8]), .C(CLK_c), .D(n29570));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i32545_3_lut (.I0(\data_out_frame[14] [4]), .I1(\data_out_frame[15] [4]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n48132));
    defparam i32545_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n51276_bdd_4_lut (.I0(n51276), .I1(n48084), .I2(n48083), .I3(byte_transmit_counter[2]), 
            .O(n51279));
    defparam n51276_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i32544_3_lut (.I0(\data_out_frame[12] [4]), .I1(\data_out_frame[13] [4]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n48131));
    defparam i32544_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF PWMLimit_i0_i9 (.Q(PWMLimit[9]), .C(CLK_c), .D(n29569));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i32541_3_lut (.I0(\data_out_frame[8] [5]), .I1(\data_out_frame[9] [5]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n48128));
    defparam i32541_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i32542_3_lut (.I0(\data_out_frame[10] [5]), .I1(\data_out_frame[11] [5]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n48129));
    defparam i32542_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF PWMLimit_i0_i10 (.Q(PWMLimit[10]), .C(CLK_c), .D(n29568));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i32515_3_lut (.I0(\data_out_frame[14] [5]), .I1(\data_out_frame[15] [5]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n48102));
    defparam i32515_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1372 (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(n43841), .I3(\FRAME_MATCHER.i [0]), .O(n43847));   // verilog/coms.v(155[7:23])
    defparam i1_2_lut_3_lut_4_lut_adj_1372.LUT_INIT = 16'hfbff;
    SB_LUT4 i32514_3_lut (.I0(\data_out_frame[12] [5]), .I1(\data_out_frame[13] [5]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n48101));
    defparam i32514_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_43_4 (.CI(n38555), .I0(\FRAME_MATCHER.i [2]), .I1(GND_net), 
            .CO(n38556));
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1373 (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(n43820), .I3(\FRAME_MATCHER.i [0]), .O(n43822));   // verilog/coms.v(155[7:23])
    defparam i1_2_lut_3_lut_4_lut_adj_1373.LUT_INIT = 16'hfbff;
    SB_LUT4 i32550_3_lut (.I0(\data_out_frame[8] [6]), .I1(\data_out_frame[9] [6]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n48137));
    defparam i32550_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i32551_3_lut (.I0(\data_out_frame[10] [6]), .I1(\data_out_frame[11] [6]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n48138));
    defparam i32551_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i32476_3_lut (.I0(\data_out_frame[14] [6]), .I1(\data_out_frame[15] [6]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n48063));
    defparam i32476_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i32475_3_lut (.I0(\data_out_frame[12] [6]), .I1(\data_out_frame[13] [6]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n48062));
    defparam i32475_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i32640_3_lut (.I0(\data_out_frame[8] [1]), .I1(\data_out_frame[9] [1]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n48227));
    defparam i32640_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i32641_3_lut (.I0(\data_out_frame[10] [1]), .I1(\data_out_frame[11] [1]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n48228));
    defparam i32641_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i32635_3_lut (.I0(\data_out_frame[14] [1]), .I1(\data_out_frame[15] [1]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n48222));
    defparam i32635_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_adj_1374 (.I0(\data_in_frame[7] [7]), .I1(n44052), 
            .I2(\data_in_frame[8] [0]), .I3(GND_net), .O(n44006));
    defparam i1_2_lut_3_lut_adj_1374.LUT_INIT = 16'h9696;
    SB_LUT4 i1_3_lut_4_lut_adj_1375 (.I0(n3303), .I1(n22132), .I2(n55), 
            .I3(n48_adj_4649), .O(n43829));   // verilog/coms.v(228[6] 230[9])
    defparam i1_3_lut_4_lut_adj_1375.LUT_INIT = 16'hff04;
    SB_LUT4 i32634_3_lut (.I0(\data_out_frame[12] [1]), .I1(\data_out_frame[13] [1]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n48221));
    defparam i32634_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2_2_lut_4_lut (.I0(n27809), .I1(n40665), .I2(\data_out_frame[17] [4]), 
            .I3(\data_out_frame[15] [2]), .O(n10_adj_4736));
    defparam i2_2_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1376 (.I0(\data_in_frame[4] [6]), .I1(\data_in_frame[5] [0]), 
            .I2(\data_in_frame[0] [7]), .I3(\data_in_frame[3] [3]), .O(n47357));   // verilog/coms.v(74[16:42])
    defparam i1_2_lut_3_lut_4_lut_adj_1376.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1377 (.I0(n40836), .I1(n45489), .I2(n44029), 
            .I3(\data_out_frame[20] [1]), .O(n41633));
    defparam i1_2_lut_4_lut_adj_1377.LUT_INIT = 16'h6996;
    SB_LUT4 i2_2_lut_3_lut_4_lut_adj_1378 (.I0(\data_out_frame[4] [6]), .I1(\data_out_frame[5] [0]), 
            .I2(\data_out_frame[7] [2]), .I3(\data_out_frame[5] [1]), .O(n27612));   // verilog/coms.v(86[17:28])
    defparam i2_2_lut_3_lut_4_lut_adj_1378.LUT_INIT = 16'h6996;
    SB_LUT4 i1_3_lut_adj_1379 (.I0(n44813), .I1(\FRAME_MATCHER.state [3]), 
            .I2(n35382), .I3(GND_net), .O(n27157));
    defparam i1_3_lut_adj_1379.LUT_INIT = 16'haeae;
    SB_DFF PWMLimit_i0_i11 (.Q(PWMLimit[11]), .C(CLK_c), .D(n29567));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1380 (.I0(\data_out_frame[22] [5]), .I1(\data_out_frame[20] [4]), 
            .I2(n41801), .I3(n40636), .O(n43960));
    defparam i1_2_lut_3_lut_4_lut_adj_1380.LUT_INIT = 16'h6996;
    SB_LUT4 i35539_3_lut (.I0(n44724), .I1(n44829), .I2(n27157), .I3(GND_net), 
            .O(n45257));
    defparam i35539_3_lut.LUT_INIT = 16'h0101;
    SB_LUT4 i1_2_lut_4_lut_adj_1381 (.I0(\data_out_frame[22] [3]), .I1(\data_out_frame[20] [2]), 
            .I2(n41171), .I3(n41829), .O(n41809));
    defparam i1_2_lut_4_lut_adj_1381.LUT_INIT = 16'h9669;
    SB_LUT4 add_43_3_lut (.I0(n3345), .I1(\FRAME_MATCHER.i [1]), .I2(GND_net), 
            .I3(n38554), .O(n2_adj_4594)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_3_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_4_lut_adj_1382 (.I0(\FRAME_MATCHER.state [0]), .I1(n24450), 
            .I2(\FRAME_MATCHER.state [2]), .I3(n23931), .O(n46039));
    defparam i1_4_lut_adj_1382.LUT_INIT = 16'h5040;
    SB_CARRY add_43_3 (.CI(n38554), .I0(\FRAME_MATCHER.i [1]), .I1(GND_net), 
            .CO(n38555));
    SB_LUT4 add_43_2_lut (.I0(n3345), .I1(\FRAME_MATCHER.i [0]), .I2(n161), 
            .I3(GND_net), .O(n2_adj_4596)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_43_2 (.CI(GND_net), .I0(\FRAME_MATCHER.i [0]), .I1(n161), 
            .CO(n38554));
    SB_LUT4 i35559_4_lut (.I0(n27157), .I1(n35382), .I2(n47279), .I3(n46039), 
            .O(n43762));
    defparam i35559_4_lut.LUT_INIT = 16'h1115;
    SB_LUT4 i1_2_lut_3_lut_adj_1383 (.I0(\data_in_frame[12] [5]), .I1(n27873), 
            .I2(n27574), .I3(GND_net), .O(n44290));
    defparam i1_2_lut_3_lut_adj_1383.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1384 (.I0(\data_in_frame[12] [5]), .I1(n27873), 
            .I2(\data_in_frame[12] [4]), .I3(GND_net), .O(n4_adj_4657));
    defparam i1_2_lut_3_lut_adj_1384.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1385 (.I0(\data_in_frame[7] [7]), .I1(n44052), 
            .I2(\data_in_frame[5] [7]), .I3(\data_in_frame[10] [3]), .O(n44589));
    defparam i2_3_lut_4_lut_adj_1385.LUT_INIT = 16'h6996;
    SB_LUT4 i15392_3_lut_4_lut (.I0(n8_adj_4681), .I1(n43841), .I2(rx_data[7]), 
            .I3(\data_in_frame[12] [7]), .O(n29340));
    defparam i15392_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF PWMLimit_i0_i12 (.Q(PWMLimit[12]), .C(CLK_c), .D(n29566));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_35676 (.I0(byte_transmit_counter[1]), 
            .I1(n48197), .I2(n48198), .I3(byte_transmit_counter[2]), .O(n51270));
    defparam byte_transmit_counter_1__bdd_4_lut_35676.LUT_INIT = 16'he4aa;
    SB_LUT4 n51270_bdd_4_lut (.I0(n51270), .I1(n48087), .I2(n48086), .I3(byte_transmit_counter[2]), 
            .O(n51273));
    defparam n51270_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_35671 (.I0(byte_transmit_counter[1]), 
            .I1(n48068), .I2(n48069), .I3(byte_transmit_counter[2]), .O(n51264));
    defparam byte_transmit_counter_1__bdd_4_lut_35671.LUT_INIT = 16'he4aa;
    SB_LUT4 n51264_bdd_4_lut (.I0(n51264), .I1(n48231), .I2(n48230), .I3(byte_transmit_counter[2]), 
            .O(n51267));
    defparam n51264_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_35711 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[22] [1]), .I2(\data_out_frame[23] [1]), 
            .I3(byte_transmit_counter[1]), .O(n51258));
    defparam byte_transmit_counter_0__bdd_4_lut_35711.LUT_INIT = 16'he4aa;
    SB_LUT4 n51258_bdd_4_lut (.I0(n51258), .I1(\data_out_frame[21] [1]), 
            .I2(\data_out_frame[20] [1]), .I3(byte_transmit_counter[1]), 
            .O(n51261));
    defparam n51258_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF data_out_frame_0___i103 (.Q(\data_out_frame[12] [6]), .C(CLK_c), 
           .D(n29021));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i1_2_lut_3_lut_adj_1386 (.I0(\data_out_frame[20] [2]), .I1(n41171), 
            .I2(n41829), .I3(GND_net), .O(n41805));
    defparam i1_2_lut_3_lut_adj_1386.LUT_INIT = 16'h6969;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_35666 (.I0(byte_transmit_counter[1]), 
            .I1(n48095), .I2(n48096), .I3(byte_transmit_counter[2]), .O(n51252));
    defparam byte_transmit_counter_1__bdd_4_lut_35666.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_2_lut_3_lut_adj_1387 (.I0(\data_out_frame[24] [1]), .I1(\data_out_frame[24] [2]), 
            .I2(n44140), .I3(GND_net), .O(n44142));   // verilog/coms.v(75[16:43])
    defparam i1_2_lut_3_lut_adj_1387.LUT_INIT = 16'h6969;
    SB_LUT4 n51252_bdd_4_lut (.I0(n51252), .I1(n48090), .I2(n48089), .I3(byte_transmit_counter[2]), 
            .O(n51255));
    defparam n51252_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_35657 (.I0(byte_transmit_counter[1]), 
            .I1(n48182), .I2(n48183), .I3(byte_transmit_counter[2]), .O(n51246));
    defparam byte_transmit_counter_1__bdd_4_lut_35657.LUT_INIT = 16'he4aa;
    SB_DFF PWMLimit_i0_i13 (.Q(PWMLimit[13]), .C(CLK_c), .D(n29565));   // verilog/coms.v(128[12] 303[6])
    SB_DFF PWMLimit_i0_i14 (.Q(PWMLimit[14]), .C(CLK_c), .D(n29564));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_35898 (.I0(byte_transmit_counter[3]), 
            .I1(n51231), .I2(n49352), .I3(byte_transmit_counter[4]), .O(n51540));
    defparam byte_transmit_counter_3__bdd_4_lut_35898.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_2_lut_3_lut_adj_1388 (.I0(\FRAME_MATCHER.state [2]), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.state [0]), .I3(GND_net), .O(n47567));
    defparam i1_2_lut_3_lut_adj_1388.LUT_INIT = 16'hfdfd;
    SB_LUT4 n51246_bdd_4_lut (.I0(n51246), .I1(n48093), .I2(n48092), .I3(byte_transmit_counter[2]), 
            .O(n51249));
    defparam n51246_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF PWMLimit_i0_i15 (.Q(PWMLimit[15]), .C(CLK_c), .D(n29563));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_35652 (.I0(byte_transmit_counter[1]), 
            .I1(n48146), .I2(n48147), .I3(byte_transmit_counter[2]), .O(n51240));
    defparam byte_transmit_counter_1__bdd_4_lut_35652.LUT_INIT = 16'he4aa;
    SB_DFF PWMLimit_i0_i16 (.Q(PWMLimit[16]), .C(CLK_c), .D(n29562));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 n51240_bdd_4_lut (.I0(n51240), .I1(n48120), .I2(n48119), .I3(byte_transmit_counter[2]), 
            .O(n51243));
    defparam n51240_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF PWMLimit_i0_i17 (.Q(PWMLimit[17]), .C(CLK_c), .D(n29561));   // verilog/coms.v(128[12] 303[6])
    SB_DFF PWMLimit_i0_i18 (.Q(PWMLimit[18]), .C(CLK_c), .D(n29560));   // verilog/coms.v(128[12] 303[6])
    SB_DFF PWMLimit_i0_i19 (.Q(PWMLimit[19]), .C(CLK_c), .D(n29559));   // verilog/coms.v(128[12] 303[6])
    SB_DFF PWMLimit_i0_i20 (.Q(PWMLimit[20]), .C(CLK_c), .D(n29558));   // verilog/coms.v(128[12] 303[6])
    SB_DFF PWMLimit_i0_i21 (.Q(PWMLimit[21]), .C(CLK_c), .D(n29557));   // verilog/coms.v(128[12] 303[6])
    SB_DFF PWMLimit_i0_i22 (.Q(PWMLimit[22]), .C(CLK_c), .D(n29556));   // verilog/coms.v(128[12] 303[6])
    SB_DFF PWMLimit_i0_i23 (.Q(PWMLimit[23]), .C(CLK_c), .D(n29555));   // verilog/coms.v(128[12] 303[6])
    SB_DFF \FRAME_MATCHER.state_i2  (.Q(\FRAME_MATCHER.state [2]), .C(CLK_c), 
           .D(n51605));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_35647 (.I0(byte_transmit_counter[1]), 
            .I1(n48113), .I2(n48114), .I3(byte_transmit_counter[2]), .O(n51234));
    defparam byte_transmit_counter_1__bdd_4_lut_35647.LUT_INIT = 16'he4aa;
    SB_DFFSS \FRAME_MATCHER.state_i30  (.Q(\FRAME_MATCHER.state [30]), .C(CLK_c), 
            .D(n43208), .S(n43088));   // verilog/coms.v(128[12] 303[6])
    SB_DFFSS \FRAME_MATCHER.state_i29  (.Q(\FRAME_MATCHER.state [29]), .C(CLK_c), 
            .D(n43206), .S(n35236));   // verilog/coms.v(128[12] 303[6])
    SB_DFFSS \FRAME_MATCHER.state_i28  (.Q(\FRAME_MATCHER.state [28]), .C(CLK_c), 
            .D(n43202), .S(n43092));   // verilog/coms.v(128[12] 303[6])
    SB_DFFSS \FRAME_MATCHER.state_i27  (.Q(\FRAME_MATCHER.state [27]), .C(CLK_c), 
            .D(n34596), .S(n35234));   // verilog/coms.v(128[12] 303[6])
    SB_DFFSS \FRAME_MATCHER.state_i26  (.Q(\FRAME_MATCHER.state [26]), .C(CLK_c), 
            .D(n43200), .S(n43094));   // verilog/coms.v(128[12] 303[6])
    SB_DFFSS \FRAME_MATCHER.state_i25  (.Q(\FRAME_MATCHER.state [25]), .C(CLK_c), 
            .D(n43198), .S(n43096));   // verilog/coms.v(128[12] 303[6])
    SB_DFFSS \FRAME_MATCHER.state_i24  (.Q(\FRAME_MATCHER.state [24]), .C(CLK_c), 
            .D(n43196), .S(n43098));   // verilog/coms.v(128[12] 303[6])
    SB_DFFSS \FRAME_MATCHER.state_i23  (.Q(\FRAME_MATCHER.state [23]), .C(CLK_c), 
            .D(n34594), .S(n35232));   // verilog/coms.v(128[12] 303[6])
    SB_DFFSS \FRAME_MATCHER.state_i22  (.Q(\FRAME_MATCHER.state [22]), .C(CLK_c), 
            .D(n43194), .S(n43102));   // verilog/coms.v(128[12] 303[6])
    SB_DFFSS \FRAME_MATCHER.state_i21  (.Q(\FRAME_MATCHER.state [21]), .C(CLK_c), 
            .D(n43192), .S(n43104));   // verilog/coms.v(128[12] 303[6])
    SB_DFFSS \FRAME_MATCHER.state_i20  (.Q(\FRAME_MATCHER.state [20]), .C(CLK_c), 
            .D(n43190), .S(n43106));   // verilog/coms.v(128[12] 303[6])
    SB_DFFSS \FRAME_MATCHER.state_i19  (.Q(\FRAME_MATCHER.state [19]), .C(CLK_c), 
            .D(n43188), .S(n43108));   // verilog/coms.v(128[12] 303[6])
    SB_DFFSS \FRAME_MATCHER.state_i18  (.Q(\FRAME_MATCHER.state [18]), .C(CLK_c), 
            .D(n43186), .S(n43110));   // verilog/coms.v(128[12] 303[6])
    SB_DFFSS \FRAME_MATCHER.state_i17  (.Q(\FRAME_MATCHER.state [17]), .C(CLK_c), 
            .D(n43184), .S(n43112));   // verilog/coms.v(128[12] 303[6])
    SB_DFFSS \FRAME_MATCHER.state_i16  (.Q(\FRAME_MATCHER.state [16]), .C(CLK_c), 
            .D(n43182), .S(n43114));   // verilog/coms.v(128[12] 303[6])
    SB_DFFSS \FRAME_MATCHER.state_i15  (.Q(\FRAME_MATCHER.state [15]), .C(CLK_c), 
            .D(n43180), .S(n43116));   // verilog/coms.v(128[12] 303[6])
    SB_DFFSS \FRAME_MATCHER.state_i14  (.Q(\FRAME_MATCHER.state [14]), .C(CLK_c), 
            .D(n43178), .S(n43118));   // verilog/coms.v(128[12] 303[6])
    SB_DFFSS \FRAME_MATCHER.state_i13  (.Q(\FRAME_MATCHER.state [13]), .C(CLK_c), 
            .D(n43172), .S(n43120));   // verilog/coms.v(128[12] 303[6])
    SB_DFFSS \FRAME_MATCHER.state_i12  (.Q(\FRAME_MATCHER.state [12]), .C(CLK_c), 
            .D(n43166), .S(n43122));   // verilog/coms.v(128[12] 303[6])
    SB_DFFSS \FRAME_MATCHER.state_i11  (.Q(\FRAME_MATCHER.state [11]), .C(CLK_c), 
            .D(n43164), .S(n43124));   // verilog/coms.v(128[12] 303[6])
    SB_DFFSS \FRAME_MATCHER.state_i10  (.Q(\FRAME_MATCHER.state [10]), .C(CLK_c), 
            .D(n43162), .S(n43126));   // verilog/coms.v(128[12] 303[6])
    SB_DFFSS \FRAME_MATCHER.state_i9  (.Q(\FRAME_MATCHER.state [9]), .C(CLK_c), 
            .D(n43160), .S(n43128));   // verilog/coms.v(128[12] 303[6])
    SB_DFFSS \FRAME_MATCHER.state_i8  (.Q(\FRAME_MATCHER.state [8]), .C(CLK_c), 
            .D(n43158), .S(n43130));   // verilog/coms.v(128[12] 303[6])
    SB_DFFSS \FRAME_MATCHER.state_i7  (.Q(\FRAME_MATCHER.state [7]), .C(CLK_c), 
            .D(n43156), .S(n43132));   // verilog/coms.v(128[12] 303[6])
    SB_DFFSS \FRAME_MATCHER.state_i6  (.Q(\FRAME_MATCHER.state [6]), .C(CLK_c), 
            .D(n43154), .S(n43134));   // verilog/coms.v(128[12] 303[6])
    SB_DFFSS \FRAME_MATCHER.state_i5  (.Q(\FRAME_MATCHER.state [5]), .C(CLK_c), 
            .D(n43150), .S(n35228));   // verilog/coms.v(128[12] 303[6])
    SB_DFFSS \FRAME_MATCHER.state_i4  (.Q(\FRAME_MATCHER.state [4]), .C(CLK_c), 
            .D(n43146), .S(n43026));   // verilog/coms.v(128[12] 303[6])
    SB_DFFSS \FRAME_MATCHER.state_i3  (.Q(\FRAME_MATCHER.state [3]), .C(CLK_c), 
            .D(n43036), .S(n10_adj_4627));   // verilog/coms.v(128[12] 303[6])
    SB_DFFSS \FRAME_MATCHER.state_i1  (.Q(\FRAME_MATCHER.state [1]), .C(CLK_c), 
            .D(n43032), .S(n51606));   // verilog/coms.v(128[12] 303[6])
    SB_DFFSS \FRAME_MATCHER.i_i9  (.Q(\FRAME_MATCHER.i [9]), .C(CLK_c), 
            .D(n2_adj_4701), .S(n3_adj_4624));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 n51540_bdd_4_lut (.I0(n51540), .I1(n51303), .I2(n7_adj_4737), 
            .I3(byte_transmit_counter[4]), .O(tx_data[5]));
    defparam n51540_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 select_686_Select_2_i3_2_lut (.I0(\FRAME_MATCHER.i [2]), .I1(n4141), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4593));
    defparam select_686_Select_2_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i15393_3_lut_4_lut (.I0(n8_adj_4681), .I1(n43841), .I2(rx_data[6]), 
            .I3(\data_in_frame[12] [6]), .O(n29341));
    defparam i15393_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFFSS \FRAME_MATCHER.i_i8  (.Q(\FRAME_MATCHER.i [8]), .C(CLK_c), 
            .D(n2_adj_4702), .S(n3_adj_4623));   // verilog/coms.v(128[12] 303[6])
    SB_DFFSS \FRAME_MATCHER.i_i7  (.Q(\FRAME_MATCHER.i [7]), .C(CLK_c), 
            .D(n2_adj_4704), .S(n3_adj_4622));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 select_686_Select_4_i3_2_lut (.I0(\FRAME_MATCHER.i [4]), .I1(n4141), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4591));
    defparam select_686_Select_4_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1389 (.I0(\data_in_frame[2] [4]), .I1(\data_in_frame[0] [3]), 
            .I2(\data_in_frame[0] [2]), .I3(n27948), .O(Kp_23__N_1059));   // verilog/coms.v(76[16:43])
    defparam i1_2_lut_3_lut_4_lut_adj_1389.LUT_INIT = 16'h6996;
    SB_DFFSS \FRAME_MATCHER.i_i6  (.Q(\FRAME_MATCHER.i [6]), .C(CLK_c), 
            .D(n2_adj_4706), .S(n3_adj_4621));   // verilog/coms.v(128[12] 303[6])
    SB_DFFSS \FRAME_MATCHER.i_i5  (.Q(\FRAME_MATCHER.i [5]), .C(CLK_c), 
            .D(n2_adj_4707), .S(n3_adj_4620));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1390 (.I0(n26875), .I1(\data_out_frame[14] [1]), 
            .I2(n44544), .I3(\data_out_frame[18] [4]), .O(n43964));
    defparam i1_2_lut_3_lut_4_lut_adj_1390.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1391 (.I0(\data_in_frame[0] [5]), .I1(\data_in_frame[0] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n44230));   // verilog/coms.v(78[16:27])
    defparam i1_2_lut_adj_1391.LUT_INIT = 16'h6666;
    SB_LUT4 i15432_3_lut_4_lut (.I0(n35263), .I1(n43832), .I2(rx_data[7]), 
            .I3(\data_in_frame[7] [7]), .O(n29380));
    defparam i15432_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4_4_lut_adj_1392 (.I0(\data_in_frame[0] [4]), .I1(\data_in_frame[0] [7]), 
            .I2(n43914), .I3(n6_adj_4738), .O(Kp_23__N_1008));   // verilog/coms.v(71[16:27])
    defparam i4_4_lut_adj_1392.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1393 (.I0(\data_in_frame[2] [0]), .I1(\data_in_frame[0] [0]), 
            .I2(Kp_23__N_1008), .I3(GND_net), .O(n45873));   // verilog/coms.v(71[16:69])
    defparam i2_3_lut_adj_1393.LUT_INIT = 16'h9696;
    SB_LUT4 i35536_3_lut (.I0(\FRAME_MATCHER.state [3]), .I1(n44813), .I2(n35382), 
            .I3(GND_net), .O(n45285));
    defparam i35536_3_lut.LUT_INIT = 16'h0101;
    SB_LUT4 i9_4_lut_adj_1394 (.I0(n45873), .I1(\data_in_frame[0] [7]), 
            .I2(\data_in_frame[1] [5]), .I3(\data_in_frame[1] [1]), .O(n26));
    defparam i9_4_lut_adj_1394.LUT_INIT = 16'h4010;
    SB_LUT4 i35611_4_lut (.I0(n44813), .I1(\FRAME_MATCHER.state [3]), .I2(n7477), 
            .I3(n35382), .O(n44841));
    defparam i35611_4_lut.LUT_INIT = 16'h5011;
    SB_LUT4 i13_4_lut (.I0(n27948), .I1(n26), .I2(\data_in_frame[2] [7]), 
            .I3(n44230), .O(n30_adj_4739));
    defparam i13_4_lut.LUT_INIT = 16'h4004;
    SB_LUT4 i6_4_lut_adj_1395 (.I0(\data_in_frame[0] [7]), .I1(Kp_23__N_1008), 
            .I2(n43944), .I3(n43989), .O(n23));
    defparam i6_4_lut_adj_1395.LUT_INIT = 16'h1248;
    SB_LUT4 i5_3_lut_adj_1396 (.I0(Kp_23__N_1008), .I1(n7), .I2(\data_in_frame[2] [1]), 
            .I3(GND_net), .O(n22));
    defparam i5_3_lut_adj_1396.LUT_INIT = 16'h1212;
    SB_LUT4 i32378_2_lut (.I0(n27952), .I1(n27461), .I2(GND_net), .I3(GND_net), 
            .O(n47901));
    defparam i32378_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i15_4_lut_adj_1397 (.I0(n23), .I1(n30_adj_4739), .I2(\data_in_frame[1] [6]), 
            .I3(n6_adj_4685), .O(n32));
    defparam i15_4_lut_adj_1397.LUT_INIT = 16'h0080;
    SB_LUT4 i15433_3_lut_4_lut (.I0(n35263), .I1(n43832), .I2(rx_data[6]), 
            .I3(\data_in_frame[7] [6]), .O(n29381));
    defparam i15433_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i34974_2_lut (.I0(\FRAME_MATCHER.state [1]), .I1(\FRAME_MATCHER.state [2]), 
            .I2(GND_net), .I3(GND_net), .O(n7477));   // verilog/coms.v(146[4] 302[11])
    defparam i34974_2_lut.LUT_INIT = 16'h1111;
    SB_LUT4 i10_4_lut_adj_1398 (.I0(\data_in_frame[1] [3]), .I1(n24450), 
            .I2(\data_in_frame[1] [4]), .I3(\data_in_frame[1] [2]), .O(n27));
    defparam i10_4_lut_adj_1398.LUT_INIT = 16'h2000;
    SB_LUT4 i16_4_lut_adj_1399 (.I0(n27), .I1(n32), .I2(n47901), .I3(n22), 
            .O(\FRAME_MATCHER.state_31__N_2872 [3]));
    defparam i16_4_lut_adj_1399.LUT_INIT = 16'h0800;
    SB_LUT4 i1_2_lut_adj_1400 (.I0(\FRAME_MATCHER.state [3]), .I1(n44724), 
            .I2(GND_net), .I3(GND_net), .O(n43727));
    defparam i1_2_lut_adj_1400.LUT_INIT = 16'h2222;
    SB_LUT4 i15434_3_lut_4_lut (.I0(n35263), .I1(n43832), .I2(rx_data[5]), 
            .I3(\data_in_frame[7] [5]), .O(n29382));
    defparam i15434_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_35893 (.I0(byte_transmit_counter[3]), 
            .I1(n51237), .I2(n49350), .I3(byte_transmit_counter[4]), .O(n51534));
    defparam byte_transmit_counter_3__bdd_4_lut_35893.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_4_lut_adj_1401 (.I0(n47565), .I1(n43727), .I2(\FRAME_MATCHER.state [1]), 
            .I3(\FRAME_MATCHER.state [2]), .O(n23975));
    defparam i1_4_lut_adj_1401.LUT_INIT = 16'hccdc;
    SB_LUT4 i2_4_lut_adj_1402 (.I0(\FRAME_MATCHER.state [1]), .I1(n43719), 
            .I2(n23975), .I3(\FRAME_MATCHER.state_31__N_2872 [3]), .O(n24278));
    defparam i2_4_lut_adj_1402.LUT_INIT = 16'h2000;
    SB_LUT4 i15435_3_lut_4_lut (.I0(n35263), .I1(n43832), .I2(rx_data[4]), 
            .I3(\data_in_frame[7] [4]), .O(n29383));
    defparam i15435_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i15436_3_lut_4_lut (.I0(n35263), .I1(n43832), .I2(rx_data[3]), 
            .I3(\data_in_frame[7] [3]), .O(n29384));
    defparam i15436_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF data_out_frame_0___i104 (.Q(\data_out_frame[12] [7]), .C(CLK_c), 
           .D(n29020));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 n51534_bdd_4_lut (.I0(n51534), .I1(n51297), .I2(n7_adj_4740), 
            .I3(byte_transmit_counter[4]), .O(tx_data[4]));
    defparam n51534_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i15437_3_lut_4_lut (.I0(n35263), .I1(n43832), .I2(rx_data[2]), 
            .I3(\data_in_frame[7] [2]), .O(n29385));
    defparam i15437_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_3_lut_adj_1403 (.I0(\data_out_frame[14] [1]), .I1(n26875), 
            .I2(\data_out_frame[11] [4]), .I3(GND_net), .O(n44409));
    defparam i1_2_lut_3_lut_adj_1403.LUT_INIT = 16'h9696;
    SB_DFF data_out_frame_0___i184 (.Q(\data_out_frame[22] [7]), .C(CLK_c), 
           .D(n29542));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i15438_3_lut_4_lut (.I0(n35263), .I1(n43832), .I2(rx_data[1]), 
            .I3(\data_in_frame[7] [1]), .O(n29386));
    defparam i15438_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2_3_lut_4_lut_adj_1404 (.I0(\data_out_frame[14] [1]), .I1(n26875), 
            .I2(n41611), .I3(\data_out_frame[16] [4]), .O(n46020));
    defparam i2_3_lut_4_lut_adj_1404.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1405 (.I0(n26888), .I1(\data_out_frame[11] [5]), 
            .I2(\data_out_frame[15] [7]), .I3(GND_net), .O(n41637));
    defparam i1_2_lut_3_lut_adj_1405.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1406 (.I0(n43714), .I1(n55_adj_4741), .I2(n63_adj_4742), 
            .I3(n45_adj_4743), .O(n43719));
    defparam i2_3_lut_4_lut_adj_1406.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_3_lut_4_lut_adj_1407 (.I0(n43714), .I1(n55_adj_4741), .I2(n45_adj_4743), 
            .I3(n63_adj_4742), .O(n44829));
    defparam i2_3_lut_4_lut_adj_1407.LUT_INIT = 16'hfffe;
    SB_DFF data_out_frame_0___i185 (.Q(\data_out_frame[23] [0]), .C(CLK_c), 
           .D(n29541));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i15394_3_lut_4_lut (.I0(n8_adj_4681), .I1(n43841), .I2(rx_data[5]), 
            .I3(\data_in_frame[12] [5]), .O(n29342));
    defparam i15394_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i5_3_lut_4_lut (.I0(\data_out_frame[8] [6]), .I1(n43974), .I2(n10_adj_4744), 
            .I3(n44325), .O(n27809));   // verilog/coms.v(76[16:43])
    defparam i5_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1408 (.I0(\data_out_frame[8] [6]), .I1(n43974), 
            .I2(n1247), .I3(\data_out_frame[10] [7]), .O(n44388));   // verilog/coms.v(76[16:43])
    defparam i2_3_lut_4_lut_adj_1408.LUT_INIT = 16'h6996;
    SB_LUT4 n51234_bdd_4_lut (.I0(n51234), .I1(n48126), .I2(n48125), .I3(byte_transmit_counter[2]), 
            .O(n51237));
    defparam n51234_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i2_2_lut_3_lut_adj_1409 (.I0(\data_out_frame[15] [5]), .I1(\data_out_frame[17] [7]), 
            .I2(\data_out_frame[13] [6]), .I3(GND_net), .O(n10_adj_4745));
    defparam i2_2_lut_3_lut_adj_1409.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1410 (.I0(\data_out_frame[15] [5]), .I1(\data_out_frame[17] [7]), 
            .I2(n40821), .I3(GND_net), .O(n44202));
    defparam i1_2_lut_3_lut_adj_1410.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1411 (.I0(n44172), .I1(n44456), .I2(n27406), 
            .I3(\data_out_frame[19] [5]), .O(n46018));
    defparam i2_3_lut_4_lut_adj_1411.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1412 (.I0(n44172), .I1(n44456), .I2(\data_out_frame[20] [0]), 
            .I3(GND_net), .O(n41816));
    defparam i1_2_lut_3_lut_adj_1412.LUT_INIT = 16'h9696;
    SB_LUT4 add_4114_9_lut (.I0(GND_net), .I1(byte_transmit_counter[7]), 
            .I2(GND_net), .I3(n38591), .O(n9046[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4114_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4114_8_lut (.I0(GND_net), .I1(byte_transmit_counter[6]), 
            .I2(GND_net), .I3(n38590), .O(n9046[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4114_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_4_lut_adj_1413 (.I0(n43905), .I1(n44319), .I2(\data_out_frame[20] [4]), 
            .I3(n27901), .O(n44482));
    defparam i1_2_lut_4_lut_adj_1413.LUT_INIT = 16'h6996;
    SB_LUT4 i5_2_lut_4_lut (.I0(n43905), .I1(n44319), .I2(\data_out_frame[20] [4]), 
            .I3(n40764), .O(n19_adj_4746));
    defparam i5_2_lut_4_lut.LUT_INIT = 16'h6996;
    SB_CARRY add_4114_8 (.CI(n38590), .I0(byte_transmit_counter[6]), .I1(GND_net), 
            .CO(n38591));
    SB_DFF data_out_frame_0___i186 (.Q(\data_out_frame[23] [1]), .C(CLK_c), 
           .D(n29540));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i5_3_lut_4_lut_adj_1414 (.I0(\data_out_frame[20] [3]), .I1(n41723), 
            .I2(n10_adj_4747), .I3(n44134), .O(n41718));
    defparam i5_3_lut_4_lut_adj_1414.LUT_INIT = 16'h9669;
    SB_LUT4 add_4114_7_lut (.I0(GND_net), .I1(byte_transmit_counter[5]), 
            .I2(GND_net), .I3(n38589), .O(n9046[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4114_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15439_3_lut_4_lut (.I0(n35263), .I1(n43832), .I2(rx_data[0]), 
            .I3(\data_in_frame[7] [0]), .O(n29387));
    defparam i15439_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF data_out_frame_0___i187 (.Q(\data_out_frame[23] [2]), .C(CLK_c), 
           .D(n29539));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i188 (.Q(\data_out_frame[23] [3]), .C(CLK_c), 
           .D(n29538));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i189 (.Q(\data_out_frame[23] [4]), .C(CLK_c), 
           .D(n29537));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i2_3_lut_4_lut_adj_1415 (.I0(\data_out_frame[20] [3]), .I1(n41723), 
            .I2(\data_out_frame[22] [4]), .I3(\data_out_frame[22] [3]), 
            .O(n44029));
    defparam i2_3_lut_4_lut_adj_1415.LUT_INIT = 16'h9669;
    SB_LUT4 i15395_3_lut_4_lut (.I0(n8_adj_4681), .I1(n43841), .I2(rx_data[4]), 
            .I3(\data_in_frame[12] [4]), .O(n29343));
    defparam i15395_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_CARRY add_4114_7 (.CI(n38589), .I0(byte_transmit_counter[5]), .I1(GND_net), 
            .CO(n38590));
    SB_DFF data_out_frame_0___i190 (.Q(\data_out_frame[23] [5]), .C(CLK_c), 
           .D(n29529));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i191 (.Q(\data_out_frame[23] [6]), .C(CLK_c), 
           .D(n29528));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i2_3_lut_4_lut_adj_1416 (.I0(n44482), .I1(n44571), .I2(n44187), 
            .I3(n45489), .O(n46161));
    defparam i2_3_lut_4_lut_adj_1416.LUT_INIT = 16'h9669;
    SB_LUT4 i15396_3_lut_4_lut (.I0(n8_adj_4681), .I1(n43841), .I2(rx_data[3]), 
            .I3(\data_in_frame[12] [3]), .O(n29344));
    defparam i15396_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_out_frame_0___i192 (.Q(\data_out_frame[23] [7]), .C(CLK_c), 
           .D(n29527));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 add_4114_6_lut (.I0(GND_net), .I1(byte_transmit_counter[4]), 
            .I2(GND_net), .I3(n38588), .O(n9046[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4114_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4114_6 (.CI(n38588), .I0(byte_transmit_counter[4]), .I1(GND_net), 
            .CO(n38589));
    SB_LUT4 i2_3_lut_4_lut_adj_1417 (.I0(\data_out_frame[24] [4]), .I1(n41809), 
            .I2(\data_out_frame[24] [5]), .I3(n45721), .O(n45385));
    defparam i2_3_lut_4_lut_adj_1417.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1418 (.I0(\data_out_frame[24] [4]), .I1(n41809), 
            .I2(n41718), .I3(\data_out_frame[24] [3]), .O(n44267));
    defparam i1_2_lut_3_lut_4_lut_adj_1418.LUT_INIT = 16'h6996;
    SB_LUT4 add_4114_5_lut (.I0(GND_net), .I1(byte_transmit_counter[3]), 
            .I2(GND_net), .I3(n38587), .O(n9046[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4114_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4114_5 (.CI(n38587), .I0(byte_transmit_counter[3]), .I1(GND_net), 
            .CO(n38588));
    SB_LUT4 add_4114_4_lut (.I0(GND_net), .I1(byte_transmit_counter[2]), 
            .I2(GND_net), .I3(n38586), .O(n9046[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4114_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i2_3_lut_4_lut_adj_1419 (.I0(\data_out_frame[24] [3]), .I1(n41718), 
            .I2(\data_out_frame[24] [2]), .I3(n2326), .O(n45560));
    defparam i2_3_lut_4_lut_adj_1419.LUT_INIT = 16'h9669;
    SB_DFF data_out_frame_0___i193 (.Q(\data_out_frame[24] [0]), .C(CLK_c), 
           .D(n29526));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i194 (.Q(\data_out_frame[24] [1]), .C(CLK_c), 
           .D(n29525));   // verilog/coms.v(128[12] 303[6])
    SB_CARRY add_4114_4 (.CI(n38586), .I0(byte_transmit_counter[2]), .I1(GND_net), 
            .CO(n38587));
    SB_DFF data_out_frame_0___i195 (.Q(\data_out_frame[24] [2]), .C(CLK_c), 
           .D(n29523));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i196 (.Q(\data_out_frame[24] [3]), .C(CLK_c), 
           .D(n29522));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i197 (.Q(\data_out_frame[24] [4]), .C(CLK_c), 
           .D(n29521));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i198 (.Q(\data_out_frame[24] [5]), .C(CLK_c), 
           .D(n29520));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i199 (.Q(\data_out_frame[24] [6]), .C(CLK_c), 
           .D(n29519));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i200 (.Q(\data_out_frame[24] [7]), .C(CLK_c), 
           .D(n29518));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i201 (.Q(\data_out_frame[25] [0]), .C(CLK_c), 
           .D(n29517));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 add_4114_3_lut (.I0(GND_net), .I1(byte_transmit_counter[1]), 
            .I2(GND_net), .I3(n38585), .O(n9046[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4114_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4114_3 (.CI(n38585), .I0(byte_transmit_counter[1]), .I1(GND_net), 
            .CO(n38586));
    SB_LUT4 add_4114_2_lut (.I0(GND_net), .I1(byte_transmit_counter[0]), 
            .I2(tx_transmit_N_3677), .I3(GND_net), .O(n9046[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4114_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4114_2 (.CI(GND_net), .I0(byte_transmit_counter[0]), .I1(tx_transmit_N_3677), 
            .CO(n38585));
    SB_DFF data_out_frame_0___i202 (.Q(\data_out_frame[25] [1]), .C(CLK_c), 
           .D(n29506));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i203 (.Q(\data_out_frame[25] [2]), .C(CLK_c), 
           .D(n29505));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i204 (.Q(\data_out_frame[25] [3]), .C(CLK_c), 
           .D(n29504));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i205 (.Q(\data_out_frame[25] [4]), .C(CLK_c), 
           .D(n29503));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i206 (.Q(\data_out_frame[25] [5]), .C(CLK_c), 
           .D(n29501));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i207 (.Q(\data_out_frame[25] [6]), .C(CLK_c), 
           .D(n29500));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i208 (.Q(\data_out_frame[25] [7]), .C(CLK_c), 
           .D(n29499));   // verilog/coms.v(128[12] 303[6])
    SB_DFF neopxl_color_i0_i1 (.Q(neopxl_color[1]), .C(CLK_c), .D(n29466));   // verilog/coms.v(128[12] 303[6])
    SB_DFF neopxl_color_i0_i2 (.Q(neopxl_color[2]), .C(CLK_c), .D(n29465));   // verilog/coms.v(128[12] 303[6])
    SB_DFF neopxl_color_i0_i3 (.Q(neopxl_color[3]), .C(CLK_c), .D(n29464));   // verilog/coms.v(128[12] 303[6])
    SB_DFF neopxl_color_i0_i4 (.Q(neopxl_color[4]), .C(CLK_c), .D(n29463));   // verilog/coms.v(128[12] 303[6])
    SB_DFF neopxl_color_i0_i5 (.Q(neopxl_color[5]), .C(CLK_c), .D(n29462));   // verilog/coms.v(128[12] 303[6])
    SB_DFF neopxl_color_i0_i6 (.Q(neopxl_color[6]), .C(CLK_c), .D(n29461));   // verilog/coms.v(128[12] 303[6])
    SB_DFF neopxl_color_i0_i7 (.Q(neopxl_color[7]), .C(CLK_c), .D(n29460));   // verilog/coms.v(128[12] 303[6])
    SB_DFF neopxl_color_i0_i8 (.Q(neopxl_color[8]), .C(CLK_c), .D(n29459));   // verilog/coms.v(128[12] 303[6])
    SB_DFF neopxl_color_i0_i9 (.Q(neopxl_color[9]), .C(CLK_c), .D(n29458));   // verilog/coms.v(128[12] 303[6])
    SB_DFF neopxl_color_i0_i10 (.Q(neopxl_color[10]), .C(CLK_c), .D(n29457));   // verilog/coms.v(128[12] 303[6])
    SB_DFF neopxl_color_i0_i11 (.Q(neopxl_color[11]), .C(CLK_c), .D(n29456));   // verilog/coms.v(128[12] 303[6])
    SB_DFF neopxl_color_i0_i12 (.Q(neopxl_color[12]), .C(CLK_c), .D(n29455));   // verilog/coms.v(128[12] 303[6])
    SB_DFF neopxl_color_i0_i13 (.Q(neopxl_color[13]), .C(CLK_c), .D(n29454));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_35888 (.I0(byte_transmit_counter[3]), 
            .I1(n51243), .I2(n49349), .I3(byte_transmit_counter[4]), .O(n51528));
    defparam byte_transmit_counter_3__bdd_4_lut_35888.LUT_INIT = 16'he4aa;
    SB_DFF neopxl_color_i0_i14 (.Q(neopxl_color[14]), .C(CLK_c), .D(n29453));   // verilog/coms.v(128[12] 303[6])
    SB_DFF neopxl_color_i0_i15 (.Q(neopxl_color[15]), .C(CLK_c), .D(n29452));   // verilog/coms.v(128[12] 303[6])
    SB_DFF neopxl_color_i0_i16 (.Q(neopxl_color[16]), .C(CLK_c), .D(n29451));   // verilog/coms.v(128[12] 303[6])
    SB_DFF neopxl_color_i0_i17 (.Q(neopxl_color[17]), .C(CLK_c), .D(n29450));   // verilog/coms.v(128[12] 303[6])
    SB_DFF neopxl_color_i0_i18 (.Q(neopxl_color[18]), .C(CLK_c), .D(n29449));   // verilog/coms.v(128[12] 303[6])
    SB_DFF neopxl_color_i0_i19 (.Q(neopxl_color[19]), .C(CLK_c), .D(n29448));   // verilog/coms.v(128[12] 303[6])
    SB_DFF neopxl_color_i0_i20 (.Q(neopxl_color[20]), .C(CLK_c), .D(n29447));   // verilog/coms.v(128[12] 303[6])
    SB_DFF neopxl_color_i0_i21 (.Q(neopxl_color[21]), .C(CLK_c), .D(n29446));   // verilog/coms.v(128[12] 303[6])
    SB_DFF neopxl_color_i0_i22 (.Q(neopxl_color[22]), .C(CLK_c), .D(n29445));   // verilog/coms.v(128[12] 303[6])
    SB_DFF neopxl_color_i0_i23 (.Q(neopxl_color[23]), .C(CLK_c), .D(n29444));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i2 (.Q(\data_in_frame[0] [1]), .C(CLK_c), .D(n29443));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i3 (.Q(\data_in_frame[0] [2]), .C(CLK_c), .D(n29442));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i4 (.Q(\data_in_frame[0] [3]), .C(CLK_c), .D(n29441));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i5 (.Q(\data_in_frame[0] [4]), .C(CLK_c), .D(n29440));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i6 (.Q(\data_in_frame[0] [5]), .C(CLK_c), .D(n29439));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i7 (.Q(\data_in_frame[0] [6]), .C(CLK_c), .D(n29438));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i8 (.Q(\data_in_frame[0] [7]), .C(CLK_c), .D(n29437));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i9 (.Q(\data_in_frame[1] [0]), .C(CLK_c), .D(n29436));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i2_3_lut_4_lut_adj_1420 (.I0(n31_adj_4748), .I1(n24450), .I2(\FRAME_MATCHER.state [2]), 
            .I3(n27227), .O(n28522));
    defparam i2_3_lut_4_lut_adj_1420.LUT_INIT = 16'h0010;
    SB_DFF data_in_frame_0__i10 (.Q(\data_in_frame[1] [1]), .C(CLK_c), .D(n29435));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i11 (.Q(\data_in_frame[1] [2]), .C(CLK_c), .D(n29434));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i12 (.Q(\data_in_frame[1] [3]), .C(CLK_c), .D(n29433));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i13 (.Q(\data_in_frame[1] [4]), .C(CLK_c), .D(n29432));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i14 (.Q(\data_in_frame[1] [5]), .C(CLK_c), .D(n29431));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i2094_2_lut_3_lut (.I0(n31_adj_4748), .I1(n24450), .I2(\FRAME_MATCHER.state [1]), 
            .I3(GND_net), .O(n7569));
    defparam i2094_2_lut_3_lut.LUT_INIT = 16'h1010;
    SB_DFF data_in_frame_0__i15 (.Q(\data_in_frame[1] [6]), .C(CLK_c), .D(n29430));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i16 (.Q(\data_in_frame[1] [7]), .C(CLK_c), .D(n29429));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i17 (.Q(\data_in_frame[2] [0]), .C(CLK_c), .D(n29428));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i18 (.Q(\data_in_frame[2] [1]), .C(CLK_c), .D(n29427));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i19 (.Q(\data_in_frame[2] [2]), .C(CLK_c), .D(n29426));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i20 (.Q(\data_in_frame[2] [3]), .C(CLK_c), .D(n29425));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i21 (.Q(\data_in_frame[2] [4]), .C(CLK_c), .D(n29424));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i22 (.Q(\data_in_frame[2] [5]), .C(CLK_c), .D(n29423));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i23 (.Q(\data_in_frame[2] [6]), .C(CLK_c), .D(n29422));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i24 (.Q(\data_in_frame[2] [7]), .C(CLK_c), .D(n29421));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i25 (.Q(\data_in_frame[3] [0]), .C(CLK_c), .D(n29420));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i26 (.Q(\data_in_frame[3] [1]), .C(CLK_c), .D(n29419));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i27 (.Q(\data_in_frame[3] [2]), .C(CLK_c), .D(n29418));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i28 (.Q(\data_in_frame[3] [3]), .C(CLK_c), .D(n29417));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i29 (.Q(\data_in_frame[3] [4]), .C(CLK_c), .D(n29416));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i30 (.Q(\data_in_frame[3] [5]), .C(CLK_c), .D(n29415));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i31 (.Q(\data_in_frame[3] [6]), .C(CLK_c), .D(n29414));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i32 (.Q(\data_in_frame[3] [7]), .C(CLK_c), .D(n29413));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i33 (.Q(\data_in_frame[4] [0]), .C(CLK_c), .D(n29412));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i34 (.Q(\data_in_frame[4] [1]), .C(CLK_c), .D(n29411));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i35 (.Q(\data_in_frame[4] [2]), .C(CLK_c), .D(n29410));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i36 (.Q(\data_in_frame[4] [3]), .C(CLK_c), .D(n29409));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i37 (.Q(\data_in_frame[4] [4]), .C(CLK_c), .D(n29408));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i38 (.Q(\data_in_frame[4] [5]), .C(CLK_c), .D(n29407));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i39 (.Q(\data_in_frame[4] [6]), .C(CLK_c), .D(n29406));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i40 (.Q(\data_in_frame[4] [7]), .C(CLK_c), .D(n29405));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i41 (.Q(\data_in_frame[5] [0]), .C(CLK_c), .D(n29403));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i42 (.Q(\data_in_frame[5] [1]), .C(CLK_c), .D(n29402));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i43 (.Q(\data_in_frame[5] [2]), .C(CLK_c), .D(n29401));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i44 (.Q(\data_in_frame[5] [3]), .C(CLK_c), .D(n29400));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i45 (.Q(\data_in_frame[5] [4]), .C(CLK_c), .D(n29399));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i46 (.Q(\data_in_frame[5] [5]), .C(CLK_c), .D(n29398));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i47 (.Q(\data_in_frame[5] [6]), .C(CLK_c), .D(n29397));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i48 (.Q(\data_in_frame[5] [7]), .C(CLK_c), .D(n29396));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i49 (.Q(\data_in_frame[6] [0]), .C(CLK_c), .D(n29395));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i50 (.Q(\data_in_frame[6] [1]), .C(CLK_c), .D(n29394));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i51 (.Q(\data_in_frame[6] [2]), .C(CLK_c), .D(n29393));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i52 (.Q(\data_in_frame[6] [3]), .C(CLK_c), .D(n29392));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i53 (.Q(\data_in_frame[6] [4]), .C(CLK_c), .D(n29391));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i54 (.Q(\data_in_frame[6] [5]), .C(CLK_c), .D(n29390));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 n51528_bdd_4_lut (.I0(n51528), .I1(n51291), .I2(n7_adj_4749), 
            .I3(byte_transmit_counter[4]), .O(tx_data[3]));
    defparam n51528_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF data_in_frame_0__i55 (.Q(\data_in_frame[6] [6]), .C(CLK_c), .D(n29389));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i56 (.Q(\data_in_frame[6] [7]), .C(CLK_c), .D(n29388));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i57 (.Q(\data_in_frame[7] [0]), .C(CLK_c), .D(n29387));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i58 (.Q(\data_in_frame[7] [1]), .C(CLK_c), .D(n29386));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i59 (.Q(\data_in_frame[7] [2]), .C(CLK_c), .D(n29385));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i60 (.Q(\data_in_frame[7] [3]), .C(CLK_c), .D(n29384));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i61 (.Q(\data_in_frame[7] [4]), .C(CLK_c), .D(n29383));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i62 (.Q(\data_in_frame[7] [5]), .C(CLK_c), .D(n29382));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i63 (.Q(\data_in_frame[7] [6]), .C(CLK_c), .D(n29381));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i64 (.Q(\data_in_frame[7] [7]), .C(CLK_c), .D(n29380));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i65 (.Q(\data_in_frame[8] [0]), .C(CLK_c), .D(n29379));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i66 (.Q(\data_in_frame[8] [1]), .C(CLK_c), .D(n29378));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i67 (.Q(\data_in_frame[8] [2]), .C(CLK_c), .D(n29377));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i68 (.Q(\data_in_frame[8] [3]), .C(CLK_c), .D(n29376));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i69 (.Q(\data_in_frame[8] [4]), .C(CLK_c), .D(n29375));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i70 (.Q(\data_in_frame[8] [5]), .C(CLK_c), .D(n29374));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i71 (.Q(\data_in_frame[8] [6]), .C(CLK_c), .D(n29373));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i72 (.Q(\data_in_frame[8] [7]), .C(CLK_c), .D(n29372));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i73 (.Q(\data_in_frame[9] [0]), .C(CLK_c), .D(n29371));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i74 (.Q(\data_in_frame[9] [1]), .C(CLK_c), .D(n29370));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i75 (.Q(\data_in_frame[9] [2]), .C(CLK_c), .D(n29369));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i76 (.Q(\data_in_frame[9] [3]), .C(CLK_c), .D(n29368));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i77 (.Q(\data_in_frame[9] [4]), .C(CLK_c), .D(n29367));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i78 (.Q(\data_in_frame[9] [5]), .C(CLK_c), .D(n29366));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i79 (.Q(\data_in_frame[9] [6]), .C(CLK_c), .D(n29365));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i80 (.Q(\data_in_frame[9] [7]), .C(CLK_c), .D(n29364));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i81 (.Q(\data_in_frame[10] [0]), .C(CLK_c), 
           .D(n29363));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i82 (.Q(\data_in_frame[10] [1]), .C(CLK_c), 
           .D(n29362));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i83 (.Q(\data_in_frame[10] [2]), .C(CLK_c), 
           .D(n29361));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i84 (.Q(\data_in_frame[10] [3]), .C(CLK_c), 
           .D(n29360));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i85 (.Q(\data_in_frame[10] [4]), .C(CLK_c), 
           .D(n29359));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i86 (.Q(\data_in_frame[10] [5]), .C(CLK_c), 
           .D(n29358));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i87 (.Q(\data_in_frame[10] [6]), .C(CLK_c), 
           .D(n29357));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i88 (.Q(\data_in_frame[10] [7]), .C(CLK_c), 
           .D(n29356));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i89 (.Q(\data_in_frame[11] [0]), .C(CLK_c), 
           .D(n29355));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i90 (.Q(\data_in_frame[11] [1]), .C(CLK_c), 
           .D(n29354));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i91 (.Q(\data_in_frame[11] [2]), .C(CLK_c), 
           .D(n29353));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i92 (.Q(\data_in_frame[11] [3]), .C(CLK_c), 
           .D(n29352));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i93 (.Q(\data_in_frame[11] [4]), .C(CLK_c), 
           .D(n29351));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i94 (.Q(\data_in_frame[11] [5]), .C(CLK_c), 
           .D(n29350));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i95 (.Q(\data_in_frame[11] [6]), .C(CLK_c), 
           .D(n29349));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 add_43_33_lut (.I0(n3345), .I1(\FRAME_MATCHER.i [31]), .I2(GND_net), 
            .I3(n38584), .O(n2_adj_4682)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_33_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1421 (.I0(\FRAME_MATCHER.state [1]), 
            .I1(\FRAME_MATCHER.state [0]), .I2(n27123), .I3(\FRAME_MATCHER.state [3]), 
            .O(n57));   // verilog/coms.v(264[5:27])
    defparam i1_2_lut_3_lut_4_lut_adj_1421.LUT_INIT = 16'hfffe;
    SB_DFF data_in_frame_0__i96 (.Q(\data_in_frame[11] [7]), .C(CLK_c), 
           .D(n29348));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i97 (.Q(\data_in_frame[12] [0]), .C(CLK_c), 
           .D(n29347));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i98 (.Q(\data_in_frame[12] [1]), .C(CLK_c), 
           .D(n29346));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i99 (.Q(\data_in_frame[12] [2]), .C(CLK_c), 
           .D(n29345));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i100 (.Q(\data_in_frame[12] [3]), .C(CLK_c), 
           .D(n29344));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i101 (.Q(\data_in_frame[12] [4]), .C(CLK_c), 
           .D(n29343));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 add_43_32_lut (.I0(n3345), .I1(\FRAME_MATCHER.i [30]), .I2(GND_net), 
            .I3(n38583), .O(n2_adj_4683)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_32_lut.LUT_INIT = 16'h8228;
    SB_DFF data_in_frame_0__i102 (.Q(\data_in_frame[12] [5]), .C(CLK_c), 
           .D(n29342));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i103 (.Q(\data_in_frame[12] [6]), .C(CLK_c), 
           .D(n29341));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i104 (.Q(\data_in_frame[12] [7]), .C(CLK_c), 
           .D(n29340));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i105 (.Q(\data_in_frame[13] [0]), .C(CLK_c), 
           .D(n29339));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i106 (.Q(\data_in_frame[13] [1]), .C(CLK_c), 
           .D(n29338));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i107 (.Q(\data_in_frame[13] [2]), .C(CLK_c), 
           .D(n29336));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i108 (.Q(\data_in_frame[13] [3]), .C(CLK_c), 
           .D(n29335));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i109 (.Q(\data_in_frame[13] [4]), .C(CLK_c), 
           .D(n29334));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i110 (.Q(\data_in_frame[13] [5]), .C(CLK_c), 
           .D(n29333));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i111 (.Q(\data_in_frame[13] [6]), .C(CLK_c), 
           .D(n29332));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i112 (.Q(\data_in_frame[13] [7]), .C(CLK_c), 
           .D(n29331));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i113 (.Q(\data_in_frame[14] [0]), .C(CLK_c), 
           .D(n29330));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i114 (.Q(\data_in_frame[14] [1]), .C(CLK_c), 
           .D(n29329));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i115 (.Q(\data_in_frame[14] [2]), .C(CLK_c), 
           .D(n29328));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i116 (.Q(\data_in_frame[14] [3]), .C(CLK_c), 
           .D(n29327));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i117 (.Q(\data_in_frame[14] [4]), .C(CLK_c), 
           .D(n29326));   // verilog/coms.v(128[12] 303[6])
    SB_CARRY add_43_32 (.CI(n38583), .I0(\FRAME_MATCHER.i [30]), .I1(GND_net), 
            .CO(n38584));
    SB_DFF data_in_frame_0__i118 (.Q(\data_in_frame[14] [5]), .C(CLK_c), 
           .D(n29325));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i119 (.Q(\data_in_frame[14] [6]), .C(CLK_c), 
           .D(n29322));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i120 (.Q(\data_in_frame[14] [7]), .C(CLK_c), 
           .D(n29321));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i121 (.Q(\data_in_frame[15] [0]), .C(CLK_c), 
           .D(n29320));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i122 (.Q(\data_in_frame[15] [1]), .C(CLK_c), 
           .D(n29319));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i123 (.Q(\data_in_frame[15] [2]), .C(CLK_c), 
           .D(n29318));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i124 (.Q(\data_in_frame[15] [3]), .C(CLK_c), 
           .D(n29317));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i125 (.Q(\data_in_frame[15] [4]), .C(CLK_c), 
           .D(n29316));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 add_43_31_lut (.I0(n3345), .I1(\FRAME_MATCHER.i [29]), .I2(GND_net), 
            .I3(n38582), .O(n2_adj_4688)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_31_lut.LUT_INIT = 16'h8228;
    SB_DFF data_in_frame_0__i126 (.Q(\data_in_frame[15] [5]), .C(CLK_c), 
           .D(n29315));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i127 (.Q(\data_in_frame[15] [6]), .C(CLK_c), 
           .D(n29314));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i128 (.Q(\data_in_frame[15] [7]), .C(CLK_c), 
           .D(n29313));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i129 (.Q(\data_in_frame[16] [0]), .C(CLK_c), 
           .D(n29312));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i130 (.Q(\data_in_frame[16] [1]), .C(CLK_c), 
           .D(n29311));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i131 (.Q(\data_in_frame[16] [2]), .C(CLK_c), 
           .D(n29310));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i132 (.Q(\data_in_frame[16] [3]), .C(CLK_c), 
           .D(n29309));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i133 (.Q(\data_in_frame[16] [4]), .C(CLK_c), 
           .D(n29308));   // verilog/coms.v(128[12] 303[6])
    SB_CARRY add_43_31 (.CI(n38582), .I0(\FRAME_MATCHER.i [29]), .I1(GND_net), 
            .CO(n38583));
    SB_DFF data_in_frame_0__i134 (.Q(\data_in_frame[16] [5]), .C(CLK_c), 
           .D(n29307));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i135 (.Q(\data_in_frame[16] [6]), .C(CLK_c), 
           .D(n29306));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i136 (.Q(\data_in_frame[16] [7]), .C(CLK_c), 
           .D(n29305));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 add_43_30_lut (.I0(n3345), .I1(\FRAME_MATCHER.i [28]), .I2(GND_net), 
            .I3(n38581), .O(n2_adj_4689)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_30_lut.LUT_INIT = 16'h8228;
    SB_DFF data_in_frame_0__i137 (.Q(\data_in_frame[17] [0]), .C(CLK_c), 
           .D(n29304));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i138 (.Q(\data_in_frame[17] [1]), .C(CLK_c), 
           .D(n29303));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i139 (.Q(\data_in_frame[17] [2]), .C(CLK_c), 
           .D(n29302));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i140 (.Q(\data_in_frame[17] [3]), .C(CLK_c), 
           .D(n29301));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i141 (.Q(\data_in_frame[17] [4]), .C(CLK_c), 
           .D(n29300));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i142 (.Q(\data_in_frame[17] [5]), .C(CLK_c), 
           .D(n29299));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i143 (.Q(\data_in_frame[17] [6]), .C(CLK_c), 
           .D(n29298));   // verilog/coms.v(128[12] 303[6])
    SB_CARRY add_43_30 (.CI(n38581), .I0(\FRAME_MATCHER.i [28]), .I1(GND_net), 
            .CO(n38582));
    SB_DFF data_in_frame_0__i144 (.Q(\data_in_frame[17] [7]), .C(CLK_c), 
           .D(n29297));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i145 (.Q(\data_in_frame[18] [0]), .C(CLK_c), 
           .D(n29296));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i146 (.Q(\data_in_frame[18] [1]), .C(CLK_c), 
           .D(n29295));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i147 (.Q(\data_in_frame[18] [2]), .C(CLK_c), 
           .D(n29294));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i148 (.Q(\data_in_frame[18] [3]), .C(CLK_c), 
           .D(n29293));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i149 (.Q(\data_in_frame[18] [4]), .C(CLK_c), 
           .D(n29292));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i150 (.Q(\data_in_frame[18] [5]), .C(CLK_c), 
           .D(n29291));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i151 (.Q(\data_in_frame[18] [6]), .C(CLK_c), 
           .D(n29289));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i152 (.Q(\data_in_frame[18] [7]), .C(CLK_c), 
           .D(n29287));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 add_43_29_lut (.I0(n3345), .I1(\FRAME_MATCHER.i [27]), .I2(GND_net), 
            .I3(n38580), .O(n2_adj_4690)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_29_lut.LUT_INIT = 16'h8228;
    SB_DFF data_in_frame_0__i153 (.Q(\data_in_frame[19] [0]), .C(CLK_c), 
           .D(n29286));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i154 (.Q(\data_in_frame[19] [1]), .C(CLK_c), 
           .D(n29285));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i155 (.Q(\data_in_frame[19] [2]), .C(CLK_c), 
           .D(n29284));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i156 (.Q(\data_in_frame[19] [3]), .C(CLK_c), 
           .D(n29283));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i157 (.Q(\data_in_frame[19] [4]), .C(CLK_c), 
           .D(n29282));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i158 (.Q(\data_in_frame[19] [5]), .C(CLK_c), 
           .D(n29281));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i159 (.Q(\data_in_frame[19] [6]), .C(CLK_c), 
           .D(n29280));   // verilog/coms.v(128[12] 303[6])
    SB_CARRY add_43_29 (.CI(n38580), .I0(\FRAME_MATCHER.i [27]), .I1(GND_net), 
            .CO(n38581));
    SB_DFF data_in_frame_0__i160 (.Q(\data_in_frame[19] [7]), .C(CLK_c), 
           .D(n29279));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i161 (.Q(\data_in_frame[20] [0]), .C(CLK_c), 
           .D(n29278));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i162 (.Q(\data_in_frame[20] [1]), .C(CLK_c), 
           .D(n29277));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i163 (.Q(\data_in_frame[20] [2]), .C(CLK_c), 
           .D(n29276));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i164 (.Q(\data_in_frame[20] [3]), .C(CLK_c), 
           .D(n29275));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i165 (.Q(\data_in_frame[20] [4]), .C(CLK_c), 
           .D(n29274));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i166 (.Q(\data_in_frame[20] [5]), .C(CLK_c), 
           .D(n29273));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i167 (.Q(\data_in_frame[20] [6]), .C(CLK_c), 
           .D(n29272));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i168 (.Q(\data_in_frame[20] [7]), .C(CLK_c), 
           .D(n29271));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i169 (.Q(\data_in_frame[21] [0]), .C(CLK_c), 
           .D(n29270));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i170 (.Q(\data_in_frame[21] [1]), .C(CLK_c), 
           .D(n29269));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i171 (.Q(\data_in_frame[21] [2]), .C(CLK_c), 
           .D(n29268));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i172 (.Q(\data_in_frame[21] [3]), .C(CLK_c), 
           .D(n29267));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i173 (.Q(\data_in_frame[21] [4]), .C(CLK_c), 
           .D(n29266));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i174 (.Q(\data_in_frame[21] [5]), .C(CLK_c), 
           .D(n29265));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i175 (.Q(\data_in_frame[21] [6]), .C(CLK_c), 
           .D(n29264));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i176 (.Q(\data_in_frame[21] [7]), .C(CLK_c), 
           .D(n29263));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i177 (.Q(\data_in_frame[22] [0]), .C(CLK_c), 
           .D(n29262));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i178 (.Q(\data_in_frame[22] [1]), .C(CLK_c), 
           .D(n29261));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i179 (.Q(\data_in_frame[22] [2]), .C(CLK_c), 
           .D(n29260));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i180 (.Q(\data_in_frame[22] [3]), .C(CLK_c), 
           .D(n29259));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i181 (.Q(\data_in_frame[22] [4]), .C(CLK_c), 
           .D(n29258));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i182 (.Q(\data_in_frame[22] [5]), .C(CLK_c), 
           .D(n29257));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i183 (.Q(\data_in_frame[22] [6]), .C(CLK_c), 
           .D(n29256));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i184 (.Q(\data_in_frame[22] [7]), .C(CLK_c), 
           .D(n29255));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i185 (.Q(\data_in_frame[23] [0]), .C(CLK_c), 
           .D(n29254));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i186 (.Q(\data_in_frame[23] [1]), .C(CLK_c), 
           .D(n29253));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 add_43_28_lut (.I0(n3345), .I1(\FRAME_MATCHER.i [26]), .I2(GND_net), 
            .I3(n38579), .O(n2_adj_4691)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_28_lut.LUT_INIT = 16'h8228;
    SB_DFF data_in_frame_0__i187 (.Q(\data_in_frame[23] [2]), .C(CLK_c), 
           .D(n29252));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i188 (.Q(\data_in_frame[23] [3]), .C(CLK_c), 
           .D(n29251));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i189 (.Q(\data_in_frame[23] [4]), .C(CLK_c), 
           .D(n29250));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_0___i2 (.Q(\data_in[0] [1]), .C(CLK_c), .D(n29244));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_0___i3 (.Q(\data_in[0] [2]), .C(CLK_c), .D(n29243));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_0___i4 (.Q(\data_in[0] [3]), .C(CLK_c), .D(n29242));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_0___i5 (.Q(\data_in[0] [4]), .C(CLK_c), .D(n29241));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_0___i6 (.Q(\data_in[0] [5]), .C(CLK_c), .D(n29240));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_0___i7 (.Q(\data_in[0] [6]), .C(CLK_c), .D(n29239));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_0___i8 (.Q(\data_in[0] [7]), .C(CLK_c), .D(n29225));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_0___i9 (.Q(\data_in[1] [0]), .C(CLK_c), .D(n29224));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_0___i10 (.Q(\data_in[1] [1]), .C(CLK_c), .D(n29223));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_0___i11 (.Q(\data_in[1] [2]), .C(CLK_c), .D(n29221));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_0___i12 (.Q(\data_in[1] [3]), .C(CLK_c), .D(n29220));   // verilog/coms.v(128[12] 303[6])
    SB_CARRY add_43_28 (.CI(n38579), .I0(\FRAME_MATCHER.i [26]), .I1(GND_net), 
            .CO(n38580));
    SB_DFF data_in_0___i13 (.Q(\data_in[1] [4]), .C(CLK_c), .D(n29219));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_0___i14 (.Q(\data_in[1] [5]), .C(CLK_c), .D(n29218));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_0___i15 (.Q(\data_in[1] [6]), .C(CLK_c), .D(n29217));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_0___i16 (.Q(\data_in[1] [7]), .C(CLK_c), .D(n29216));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_0___i17 (.Q(\data_in[2] [0]), .C(CLK_c), .D(n29215));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_0___i18 (.Q(\data_in[2] [1]), .C(CLK_c), .D(n29214));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_0___i19 (.Q(\data_in[2] [2]), .C(CLK_c), .D(n29213));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_0___i20 (.Q(\data_in[2] [3]), .C(CLK_c), .D(n29212));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_0___i21 (.Q(\data_in[2] [4]), .C(CLK_c), .D(n29211));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_0___i22 (.Q(\data_in[2] [5]), .C(CLK_c), .D(n29210));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_0___i23 (.Q(\data_in[2] [6]), .C(CLK_c), .D(n29209));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_0___i24 (.Q(\data_in[2] [7]), .C(CLK_c), .D(n29208));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_0___i25 (.Q(\data_in[3] [0]), .C(CLK_c), .D(n29207));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_0___i26 (.Q(\data_in[3] [1]), .C(CLK_c), .D(n29206));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_0___i27 (.Q(\data_in[3] [2]), .C(CLK_c), .D(n29205));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_0___i28 (.Q(\data_in[3] [3]), .C(CLK_c), .D(n29204));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_0___i29 (.Q(\data_in[3] [4]), .C(CLK_c), .D(n29203));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_0___i30 (.Q(\data_in[3] [5]), .C(CLK_c), .D(n29202));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_0___i31 (.Q(\data_in[3] [6]), .C(CLK_c), .D(n29201));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_0___i32 (.Q(\data_in[3] [7]), .C(CLK_c), .D(n29200));   // verilog/coms.v(128[12] 303[6])
    SB_DFF Kp_i1 (.Q(\Kp[1] ), .C(CLK_c), .D(n29199));   // verilog/coms.v(128[12] 303[6])
    SB_DFF Kp_i2 (.Q(\Kp[2] ), .C(CLK_c), .D(n29198));   // verilog/coms.v(128[12] 303[6])
    SB_DFF Kp_i3 (.Q(\Kp[3] ), .C(CLK_c), .D(n29197));   // verilog/coms.v(128[12] 303[6])
    SB_DFF Kp_i4 (.Q(\Kp[4] ), .C(CLK_c), .D(n29196));   // verilog/coms.v(128[12] 303[6])
    SB_DFF Kp_i5 (.Q(\Kp[5] ), .C(CLK_c), .D(n29195));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 add_43_27_lut (.I0(n3345), .I1(\FRAME_MATCHER.i [25]), .I2(GND_net), 
            .I3(n38578), .O(n2_adj_4692)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_27_lut.LUT_INIT = 16'h8228;
    SB_DFF Kp_i6 (.Q(\Kp[6] ), .C(CLK_c), .D(n29194));   // verilog/coms.v(128[12] 303[6])
    SB_DFF Kp_i7 (.Q(\Kp[7] ), .C(CLK_c), .D(n29193));   // verilog/coms.v(128[12] 303[6])
    SB_DFF Kp_i8 (.Q(\Kp[8] ), .C(CLK_c), .D(n29192));   // verilog/coms.v(128[12] 303[6])
    SB_DFF Kp_i9 (.Q(\Kp[9] ), .C(CLK_c), .D(n29191));   // verilog/coms.v(128[12] 303[6])
    SB_DFF Kp_i10 (.Q(\Kp[10] ), .C(CLK_c), .D(n29190));   // verilog/coms.v(128[12] 303[6])
    SB_DFF Kp_i11 (.Q(\Kp[11] ), .C(CLK_c), .D(n29189));   // verilog/coms.v(128[12] 303[6])
    SB_DFF Kp_i12 (.Q(\Kp[12] ), .C(CLK_c), .D(n29188));   // verilog/coms.v(128[12] 303[6])
    SB_DFF Kp_i13 (.Q(\Kp[13] ), .C(CLK_c), .D(n29187));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_35883 (.I0(byte_transmit_counter[3]), 
            .I1(n51249), .I2(n49347), .I3(byte_transmit_counter[4]), .O(n51522));
    defparam byte_transmit_counter_3__bdd_4_lut_35883.LUT_INIT = 16'he4aa;
    SB_DFF Kp_i14 (.Q(\Kp[14] ), .C(CLK_c), .D(n29183));   // verilog/coms.v(128[12] 303[6])
    SB_DFF Kp_i15 (.Q(\Kp[15] ), .C(CLK_c), .D(n29182));   // verilog/coms.v(128[12] 303[6])
    SB_DFF Ki_i1 (.Q(\Ki[1] ), .C(CLK_c), .D(n29181));   // verilog/coms.v(128[12] 303[6])
    SB_DFF Ki_i2 (.Q(\Ki[2] ), .C(CLK_c), .D(n29180));   // verilog/coms.v(128[12] 303[6])
    SB_DFF Ki_i3 (.Q(\Ki[3] ), .C(CLK_c), .D(n29179));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 n51522_bdd_4_lut (.I0(n51522), .I1(n51279), .I2(n7_adj_4750), 
            .I3(byte_transmit_counter[4]), .O(tx_data[2]));
    defparam n51522_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF Ki_i4 (.Q(\Ki[4] ), .C(CLK_c), .D(n29178));   // verilog/coms.v(128[12] 303[6])
    SB_DFF Ki_i5 (.Q(\Ki[5] ), .C(CLK_c), .D(n29177));   // verilog/coms.v(128[12] 303[6])
    SB_DFF Ki_i6 (.Q(\Ki[6] ), .C(CLK_c), .D(n29176));   // verilog/coms.v(128[12] 303[6])
    SB_DFF Ki_i7 (.Q(\Ki[7] ), .C(CLK_c), .D(n29175));   // verilog/coms.v(128[12] 303[6])
    SB_DFF Ki_i8 (.Q(\Ki[8] ), .C(CLK_c), .D(n29174));   // verilog/coms.v(128[12] 303[6])
    SB_DFF Ki_i9 (.Q(\Ki[9] ), .C(CLK_c), .D(n29173));   // verilog/coms.v(128[12] 303[6])
    SB_CARRY add_43_27 (.CI(n38578), .I0(\FRAME_MATCHER.i [25]), .I1(GND_net), 
            .CO(n38579));
    SB_DFF Ki_i10 (.Q(\Ki[10] ), .C(CLK_c), .D(n29172));   // verilog/coms.v(128[12] 303[6])
    SB_DFF Ki_i11 (.Q(\Ki[11] ), .C(CLK_c), .D(n29171));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_35878 (.I0(byte_transmit_counter[3]), 
            .I1(n50124), .I2(n49353), .I3(byte_transmit_counter[4]), .O(n51516));
    defparam byte_transmit_counter_3__bdd_4_lut_35878.LUT_INIT = 16'he4aa;
    SB_DFF data_out_frame_0___i105 (.Q(\data_out_frame[13] [0]), .C(CLK_c), 
           .D(n29019));   // verilog/coms.v(128[12] 303[6])
    SB_DFF Ki_i12 (.Q(\Ki[12] ), .C(CLK_c), .D(n29170));   // verilog/coms.v(128[12] 303[6])
    SB_DFF Ki_i13 (.Q(\Ki[13] ), .C(CLK_c), .D(n29169));   // verilog/coms.v(128[12] 303[6])
    SB_DFF Ki_i14 (.Q(\Ki[14] ), .C(CLK_c), .D(n29168));   // verilog/coms.v(128[12] 303[6])
    SB_DFF Ki_i15 (.Q(\Ki[15] ), .C(CLK_c), .D(n29167));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 add_43_26_lut (.I0(n3345), .I1(\FRAME_MATCHER.i [24]), .I2(GND_net), 
            .I3(n38577), .O(n2_adj_4693)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_26_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_43_26 (.CI(n38577), .I0(\FRAME_MATCHER.i [24]), .I1(GND_net), 
            .CO(n38578));
    SB_LUT4 i2_2_lut_adj_1422 (.I0(\FRAME_MATCHER.state [2]), .I1(\FRAME_MATCHER.state [0]), 
            .I2(GND_net), .I3(GND_net), .O(n34607));   // verilog/coms.v(146[4] 302[11])
    defparam i2_2_lut_adj_1422.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1423 (.I0(\FRAME_MATCHER.state [27]), .I1(\FRAME_MATCHER.state [23]), 
            .I2(GND_net), .I3(GND_net), .O(n55_adj_4741));   // verilog/coms.v(128[12] 303[6])
    defparam i1_2_lut_adj_1423.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_3_lut_adj_1424 (.I0(\data_in_frame[1] [7]), .I1(\data_in_frame[1] [6]), 
            .I2(\data_in_frame[4] [2]), .I3(GND_net), .O(n44305));   // verilog/coms.v(79[16:27])
    defparam i1_2_lut_3_lut_adj_1424.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_1425 (.I0(\FRAME_MATCHER.state [4]), .I1(\FRAME_MATCHER.state [5]), 
            .I2(\FRAME_MATCHER.state [7]), .I3(\FRAME_MATCHER.state [6]), 
            .O(n45_adj_4743));
    defparam i3_4_lut_adj_1425.LUT_INIT = 16'hfffe;
    SB_LUT4 i3_4_lut_adj_1426 (.I0(\FRAME_MATCHER.state [10]), .I1(\FRAME_MATCHER.state [9]), 
            .I2(\FRAME_MATCHER.state [14]), .I3(\FRAME_MATCHER.state [13]), 
            .O(n43817));   // verilog/coms.v(128[12] 303[6])
    defparam i3_4_lut_adj_1426.LUT_INIT = 16'hfffe;
    SB_LUT4 i4_2_lut_adj_1427 (.I0(\FRAME_MATCHER.state [25]), .I1(\FRAME_MATCHER.state [19]), 
            .I2(GND_net), .I3(GND_net), .O(n18_adj_4751));   // verilog/coms.v(213[5:16])
    defparam i4_2_lut_adj_1427.LUT_INIT = 16'heeee;
    SB_LUT4 i10_4_lut_adj_1428 (.I0(\FRAME_MATCHER.state [21]), .I1(\FRAME_MATCHER.state [22]), 
            .I2(\FRAME_MATCHER.state [20]), .I3(\FRAME_MATCHER.state [29]), 
            .O(n24));   // verilog/coms.v(213[5:16])
    defparam i10_4_lut_adj_1428.LUT_INIT = 16'hfffe;
    SB_LUT4 i8_4_lut_adj_1429 (.I0(\FRAME_MATCHER.state [18]), .I1(\FRAME_MATCHER.state [17]), 
            .I2(\FRAME_MATCHER.state [26]), .I3(\FRAME_MATCHER.state [16]), 
            .O(n22_adj_4752));   // verilog/coms.v(213[5:16])
    defparam i8_4_lut_adj_1429.LUT_INIT = 16'hfffe;
    SB_LUT4 i12_4_lut (.I0(\FRAME_MATCHER.state [30]), .I1(n24), .I2(n18_adj_4751), 
            .I3(\FRAME_MATCHER.state [28]), .O(n26_adj_4753));   // verilog/coms.v(213[5:16])
    defparam i12_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i21080_2_lut_2_lut_3_lut_4_lut (.I0(n55), .I1(n27230), .I2(rx_data_ready), 
            .I3(\FRAME_MATCHER.rx_data_ready_prev ), .O(n35014));
    defparam i21080_2_lut_2_lut_3_lut_4_lut.LUT_INIT = 16'h0070;
    SB_LUT4 i2_3_lut_4_lut_adj_1430 (.I0(\FRAME_MATCHER.state [1]), .I1(\FRAME_MATCHER.state [2]), 
            .I2(\FRAME_MATCHER.state [0]), .I3(n27004), .O(n55));
    defparam i2_3_lut_4_lut_adj_1430.LUT_INIT = 16'hffbf;
    SB_LUT4 i1_3_lut_4_lut_adj_1431 (.I0(\data_in_frame[1] [7]), .I1(\data_in_frame[1] [6]), 
            .I2(\data_in_frame[1] [4]), .I3(n27420), .O(n43938));   // verilog/coms.v(79[16:27])
    defparam i1_3_lut_4_lut_adj_1431.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1432 (.I0(\FRAME_MATCHER.state [2]), .I1(\FRAME_MATCHER.state [0]), 
            .I2(n27123), .I3(\FRAME_MATCHER.state [3]), .O(n27230));   // verilog/coms.v(255[5:25])
    defparam i2_3_lut_4_lut_adj_1432.LUT_INIT = 16'hfffb;
    SB_LUT4 i13_4_lut_adj_1433 (.I0(\FRAME_MATCHER.state [24]), .I1(n26_adj_4753), 
            .I2(n22_adj_4752), .I3(\FRAME_MATCHER.state [31]), .O(n43714));   // verilog/coms.v(213[5:16])
    defparam i13_4_lut_adj_1433.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1434 (.I0(n44482), .I1(\data_out_frame[19] [5]), 
            .I2(n41807), .I3(\data_out_frame[21] [7]), .O(n44134));
    defparam i1_2_lut_3_lut_4_lut_adj_1434.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1435 (.I0(\FRAME_MATCHER.state [11]), .I1(\FRAME_MATCHER.state [8]), 
            .I2(\FRAME_MATCHER.state [12]), .I3(\FRAME_MATCHER.state [15]), 
            .O(n43716));
    defparam i3_4_lut_adj_1435.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_adj_1436 (.I0(n43716), .I1(n43714), .I2(GND_net), 
            .I3(GND_net), .O(n4_adj_4754));   // verilog/coms.v(213[5:16])
    defparam i1_2_lut_adj_1436.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1437 (.I0(\data_out_frame[20] [3]), .I1(n41723), 
            .I2(\data_out_frame[22] [5]), .I3(n44257), .O(n27279));
    defparam i1_2_lut_3_lut_4_lut_adj_1437.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_3_lut_4_lut (.I0(n25208), .I1(\data_out_frame[11] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n45977));
    defparam i3_4_lut_3_lut_4_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i2_4_lut_adj_1438 (.I0(n43817), .I1(n45_adj_4743), .I2(n55_adj_4741), 
            .I3(n4_adj_4754), .O(n27123));   // verilog/coms.v(213[5:16])
    defparam i2_4_lut_adj_1438.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_adj_1439 (.I0(n27123), .I1(\FRAME_MATCHER.state [3]), 
            .I2(GND_net), .I3(GND_net), .O(n27004));
    defparam i1_2_lut_adj_1439.LUT_INIT = 16'heeee;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_35642 (.I0(byte_transmit_counter[1]), 
            .I1(n48080), .I2(n48081), .I3(byte_transmit_counter[2]), .O(n51228));
    defparam byte_transmit_counter_1__bdd_4_lut_35642.LUT_INIT = 16'he4aa;
    SB_LUT4 n51228_bdd_4_lut (.I0(n51228), .I1(n48135), .I2(n48134), .I3(byte_transmit_counter[2]), 
            .O(n51231));
    defparam n51228_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_3_lut_adj_1440 (.I0(\data_in_frame[0] [1]), .I1(\data_in_frame[0] [5]), 
            .I2(\data_in_frame[0] [6]), .I3(GND_net), .O(n6_adj_4738));   // verilog/coms.v(71[16:27])
    defparam i1_2_lut_3_lut_adj_1440.LUT_INIT = 16'h9696;
    SB_LUT4 i34966_2_lut_3_lut (.I0(\FRAME_MATCHER.state [1]), .I1(\FRAME_MATCHER.state [2]), 
            .I2(\FRAME_MATCHER.state [0]), .I3(GND_net), .O(n28824));
    defparam i34966_2_lut_3_lut.LUT_INIT = 16'h0e0e;
    SB_LUT4 i1_4_lut_4_lut (.I0(\FRAME_MATCHER.state [0]), .I1(\FRAME_MATCHER.state [1]), 
            .I2(\FRAME_MATCHER.state [2]), .I3(\FRAME_MATCHER.state_31__N_2872 [3]), 
            .O(n47279));
    defparam i1_4_lut_4_lut.LUT_INIT = 16'habaf;
    SB_LUT4 i21293_2_lut_3_lut_4_lut (.I0(n22132), .I1(n4120), .I2(n43829), 
            .I3(\FRAME_MATCHER.state [23]), .O(n35232));
    defparam i21293_2_lut_3_lut_4_lut.LUT_INIT = 16'hf800;
    SB_LUT4 i1_2_lut_3_lut_adj_1441 (.I0(\data_in_frame[2] [5]), .I1(\data_in_frame[0] [3]), 
            .I2(\data_in_frame[0] [4]), .I3(GND_net), .O(n6_adj_4685));   // verilog/coms.v(167[9:87])
    defparam i1_2_lut_3_lut_adj_1441.LUT_INIT = 16'h9696;
    SB_LUT4 i21290_2_lut_3_lut_4_lut (.I0(n22132), .I1(n4120), .I2(n43829), 
            .I3(\FRAME_MATCHER.state [5]), .O(n35228));
    defparam i21290_2_lut_3_lut_4_lut.LUT_INIT = 16'hf800;
    SB_LUT4 i3_3_lut_4_lut (.I0(n55), .I1(n27230), .I2(n63), .I3(n27235), 
            .O(n8_adj_4726));
    defparam i3_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i21289_1_lut_2_lut (.I0(n55), .I1(n27230), .I2(GND_net), .I3(GND_net), 
            .O(n3345));
    defparam i21289_1_lut_2_lut.LUT_INIT = 16'h7777;
    SB_LUT4 i1_3_lut_4_lut_adj_1442 (.I0(\FRAME_MATCHER.state [1]), .I1(n27230), 
            .I2(n43850), .I3(n771), .O(n43859));   // verilog/coms.v(202[5:24])
    defparam i1_3_lut_4_lut_adj_1442.LUT_INIT = 16'hf0f1;
    SB_LUT4 i1_3_lut_4_lut_adj_1443 (.I0(n55), .I1(n27230), .I2(n57), 
            .I3(\FRAME_MATCHER.state [2]), .O(n4141));
    defparam i1_3_lut_4_lut_adj_1443.LUT_INIT = 16'h8880;
    SB_LUT4 select_686_Select_0_i3_2_lut (.I0(\FRAME_MATCHER.i [0]), .I1(n4141), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4597));
    defparam select_686_Select_0_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_3_lut_4_lut_adj_1444 (.I0(\FRAME_MATCHER.i [0]), .I1(\FRAME_MATCHER.i [4]), 
            .I2(n27189), .I3(\FRAME_MATCHER.i [1]), .O(n5_adj_4727));
    defparam i1_3_lut_4_lut_adj_1444.LUT_INIT = 16'hfefc;
    SB_LUT4 i1_2_lut_3_lut_adj_1445 (.I0(\state[0] ), .I1(\state[2] ), .I2(\state[3] ), 
            .I3(GND_net), .O(n7754));
    defparam i1_2_lut_3_lut_adj_1445.LUT_INIT = 16'h0202;
    SB_LUT4 i1_3_lut_4_lut_adj_1446 (.I0(\data_in_frame[2] [5]), .I1(\data_in_frame[0] [3]), 
            .I2(\data_in_frame[2] [6]), .I3(\data_in_frame[0] [5]), .O(n44376));   // verilog/coms.v(167[9:87])
    defparam i1_3_lut_4_lut_adj_1446.LUT_INIT = 16'h6996;
    SB_LUT4 i15424_3_lut_4_lut (.I0(n8_adj_4729), .I1(n43841), .I2(rx_data[7]), 
            .I3(\data_in_frame[8] [7]), .O(n29372));
    defparam i15424_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_2_lut_4_lut_adj_1447 (.I0(n27123), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.state [0]), .I3(\FRAME_MATCHER.state [1]), 
            .O(n27227));   // verilog/coms.v(232[5:23])
    defparam i2_2_lut_4_lut_adj_1447.LUT_INIT = 16'hfeff;
    SB_LUT4 i29210_2_lut_3_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n27230), 
            .I2(n4452), .I3(GND_net), .O(n44726));
    defparam i29210_2_lut_3_lut.LUT_INIT = 16'hfdfd;
    SB_LUT4 i1_3_lut_4_lut_adj_1448 (.I0(\data_in_frame[0] [6]), .I1(\data_in_frame[1] [0]), 
            .I2(Kp_23__N_1027), .I3(\data_in_frame[3] [0]), .O(n28228));   // verilog/coms.v(78[16:27])
    defparam i1_3_lut_4_lut_adj_1448.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1449 (.I0(\data_in_frame[2] [4]), .I1(\data_in_frame[0] [3]), 
            .I2(\data_in_frame[0] [2]), .I3(GND_net), .O(n27461));   // verilog/coms.v(167[9:87])
    defparam i1_2_lut_3_lut_adj_1449.LUT_INIT = 16'h9696;
    SB_LUT4 i15425_3_lut_4_lut (.I0(n8_adj_4729), .I1(n43841), .I2(rx_data[6]), 
            .I3(\data_in_frame[8] [6]), .O(n29373));
    defparam i15425_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1450 (.I0(\data_in_frame[9] [4]), .I1(\data_in_frame[9] [5]), 
            .I2(\data_in_frame[11] [6]), .I3(GND_net), .O(n43971));
    defparam i1_2_lut_3_lut_adj_1450.LUT_INIT = 16'h9696;
    SB_LUT4 i15426_3_lut_4_lut (.I0(n8_adj_4729), .I1(n43841), .I2(rx_data[5]), 
            .I3(\data_in_frame[8] [5]), .O(n29374));
    defparam i15426_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 select_686_Select_3_i3_2_lut (.I0(\FRAME_MATCHER.i [3]), .I1(n4141), 
            .I2(GND_net), .I3(GND_net), .O(n3));
    defparam select_686_Select_3_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_3_lut_4_lut_adj_1451 (.I0(\data_in_frame[1] [1]), .I1(\data_in_frame[0] [6]), 
            .I2(\data_in_frame[1] [0]), .I3(\data_in_frame[3] [2]), .O(n28357));
    defparam i1_3_lut_4_lut_adj_1451.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1452 (.I0(\data_in_frame[5] [3]), .I1(n26199), 
            .I2(\data_in_frame[2] [7]), .I3(GND_net), .O(n44335));   // verilog/coms.v(86[17:63])
    defparam i1_2_lut_3_lut_adj_1452.LUT_INIT = 16'h9696;
    SB_LUT4 i1_3_lut_4_lut_adj_1453 (.I0(\data_in_frame[3] [1]), .I1(\data_in_frame[5] [1]), 
            .I2(n43899), .I3(n47351), .O(n47361));   // verilog/coms.v(74[16:42])
    defparam i1_3_lut_4_lut_adj_1453.LUT_INIT = 16'h6996;
    SB_LUT4 i1_3_lut_4_lut_adj_1454 (.I0(n40688), .I1(\data_in_frame[9] [1]), 
            .I2(n44574), .I3(\data_in_frame[9] [0]), .O(n47339));   // verilog/coms.v(86[17:63])
    defparam i1_3_lut_4_lut_adj_1454.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1455 (.I0(\FRAME_MATCHER.state [1]), .I1(\FRAME_MATCHER.state [0]), 
            .I2(n43719), .I3(\FRAME_MATCHER.state [2]), .O(n35382));   // verilog/coms.v(264[5:27])
    defparam i2_3_lut_4_lut_adj_1455.LUT_INIT = 16'hfffe;
    SB_LUT4 i29208_2_lut_3_lut (.I0(\FRAME_MATCHER.state [1]), .I1(\FRAME_MATCHER.state [0]), 
            .I2(\FRAME_MATCHER.state [2]), .I3(GND_net), .O(n44724));   // verilog/coms.v(264[5:27])
    defparam i29208_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i29212_2_lut_3_lut (.I0(\FRAME_MATCHER.state [1]), .I1(\FRAME_MATCHER.state [0]), 
            .I2(n27123), .I3(GND_net), .O(n44728));   // verilog/coms.v(264[5:27])
    defparam i29212_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_2_lut_3_lut_adj_1456 (.I0(\data_in_frame[9] [1]), .I1(\data_in_frame[9] [2]), 
            .I2(Kp_23__N_1253), .I3(GND_net), .O(n44419));   // verilog/coms.v(73[16:41])
    defparam i1_2_lut_3_lut_adj_1456.LUT_INIT = 16'h9696;
    SB_LUT4 i15427_3_lut_4_lut (.I0(n8_adj_4729), .I1(n43841), .I2(rx_data[4]), 
            .I3(\data_in_frame[8] [4]), .O(n29375));
    defparam i15427_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15428_3_lut_4_lut (.I0(n8_adj_4729), .I1(n43841), .I2(rx_data[3]), 
            .I3(\data_in_frame[8] [3]), .O(n29376));
    defparam i15428_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15429_3_lut_4_lut (.I0(n8_adj_4729), .I1(n43841), .I2(rx_data[2]), 
            .I3(\data_in_frame[8] [2]), .O(n29377));
    defparam i15429_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 n51516_bdd_4_lut (.I0(n51516), .I1(n51315), .I2(n7_adj_4755), 
            .I3(byte_transmit_counter[4]), .O(tx_data[1]));
    defparam n51516_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i15430_3_lut_4_lut (.I0(n8_adj_4729), .I1(n43841), .I2(rx_data[1]), 
            .I3(\data_in_frame[8] [1]), .O(n29378));
    defparam i15430_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15431_3_lut_4_lut (.I0(n8_adj_4729), .I1(n43841), .I2(rx_data[0]), 
            .I3(\data_in_frame[8] [0]), .O(n29379));
    defparam i15431_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_4_lut_adj_1457 (.I0(\data_out_frame[20] [7]), .I1(n41653), 
            .I2(n27901), .I3(n41677), .O(n44586));
    defparam i2_3_lut_4_lut_adj_1457.LUT_INIT = 16'h9669;
    SB_LUT4 i15302_3_lut_4_lut (.I0(n35263), .I1(n43820), .I2(rx_data[4]), 
            .I3(\data_in_frame[23] [4]), .O(n29250));
    defparam i15302_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_3_lut_4_lut_adj_1458 (.I0(\data_in_frame[3] [5]), .I1(\data_in_frame[5] [7]), 
            .I2(n44513), .I3(Kp_23__N_1103), .O(n27488));   // verilog/coms.v(79[16:27])
    defparam i1_3_lut_4_lut_adj_1458.LUT_INIT = 16'h6996;
    SB_LUT4 i15303_3_lut_4_lut (.I0(n35263), .I1(n43820), .I2(rx_data[3]), 
            .I3(\data_in_frame[23] [3]), .O(n29251));
    defparam i15303_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i15304_3_lut_4_lut (.I0(n35263), .I1(n43820), .I2(rx_data[2]), 
            .I3(\data_in_frame[23] [2]), .O(n29252));
    defparam i15304_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i15305_3_lut_4_lut (.I0(n35263), .I1(n43820), .I2(rx_data[1]), 
            .I3(\data_in_frame[23] [1]), .O(n29253));
    defparam i15305_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i15306_3_lut_4_lut (.I0(n35263), .I1(n43820), .I2(rx_data[0]), 
            .I3(\data_in_frame[23] [0]), .O(n29254));
    defparam i15306_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i15652_3_lut_4_lut (.I0(n35263), .I1(n43820), .I2(rx_data[6]), 
            .I3(\data_in_frame[23] [6]), .O(n29600));
    defparam i15652_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i15653_3_lut_4_lut (.I0(n35263), .I1(n43820), .I2(rx_data[7]), 
            .I3(\data_in_frame[23] [7]), .O(n29601));
    defparam i15653_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i15655_3_lut_4_lut (.I0(n35263), .I1(n43820), .I2(rx_data[5]), 
            .I3(\data_in_frame[23] [5]), .O(n29603));
    defparam i15655_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2_3_lut_4_lut_adj_1459 (.I0(\data_out_frame[20] [7]), .I1(n41653), 
            .I2(\data_out_frame[19] [0]), .I3(n44580), .O(n44175));
    defparam i2_3_lut_4_lut_adj_1459.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1460 (.I0(\data_in_frame[8] [3]), .I1(n27475), 
            .I2(n44513), .I3(Kp_23__N_1103), .O(n4_adj_4619));   // verilog/coms.v(74[16:42])
    defparam i1_2_lut_4_lut_adj_1460.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1461 (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(n43820), .I3(\FRAME_MATCHER.i [0]), .O(n43824));
    defparam i1_2_lut_3_lut_4_lut_adj_1461.LUT_INIT = 16'hfff7;
    SB_LUT4 i21321_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n35263));
    defparam i21321_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1462 (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(n43841), .I3(\FRAME_MATCHER.i [0]), .O(n43848));
    defparam i1_2_lut_3_lut_4_lut_adj_1462.LUT_INIT = 16'hfff7;
    SB_LUT4 i2_3_lut_4_lut_adj_1463 (.I0(n26875), .I1(n44026), .I2(\data_out_frame[18] [6]), 
            .I3(\data_out_frame[21] [1]), .O(n44580));
    defparam i2_3_lut_4_lut_adj_1463.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1464 (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(n43832), .I3(\FRAME_MATCHER.i [0]), .O(n43839));
    defparam i1_2_lut_3_lut_4_lut_adj_1464.LUT_INIT = 16'hfff7;
    SB_LUT4 i5_3_lut_4_lut_adj_1465 (.I0(\data_out_frame[6] [3]), .I1(n43874), 
            .I2(\data_out_frame[12] [5]), .I3(\data_out_frame[14] [7]), 
            .O(n14));   // verilog/coms.v(73[16:27])
    defparam i5_3_lut_4_lut_adj_1465.LUT_INIT = 16'h6996;
    SB_LUT4 i15416_3_lut_4_lut (.I0(n8_adj_4645), .I1(n43841), .I2(rx_data[7]), 
            .I3(\data_in_frame[9] [7]), .O(n29364));
    defparam i15416_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_3_lut_4_lut_adj_1466 (.I0(n43938), .I1(\data_in_frame[5] [3]), 
            .I2(n27730), .I3(n47759), .O(n40688));   // verilog/coms.v(86[17:63])
    defparam i1_3_lut_4_lut_adj_1466.LUT_INIT = 16'h6996;
    SB_LUT4 i3_3_lut_4_lut_adj_1467 (.I0(\data_in_frame[20] [4]), .I1(\data_in_frame[22] [6]), 
            .I2(n40631), .I3(n40620), .O(n8_adj_4696));
    defparam i3_3_lut_4_lut_adj_1467.LUT_INIT = 16'h6996;
    SB_LUT4 i1_3_lut_4_lut_adj_1468 (.I0(n22132), .I1(\FRAME_MATCHER.state [1]), 
            .I2(n27230), .I3(n4452), .O(n37));   // verilog/coms.v(255[5:25])
    defparam i1_3_lut_4_lut_adj_1468.LUT_INIT = 16'h0008;
    SB_LUT4 i15417_3_lut_4_lut (.I0(n8_adj_4645), .I1(n43841), .I2(rx_data[6]), 
            .I3(\data_in_frame[9] [6]), .O(n29365));
    defparam i15417_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_4_lut_adj_1469 (.I0(\data_in_frame[12] [4]), .I1(n27574), 
            .I2(\data_in_frame[14] [5]), .I3(n41760), .O(n44350));
    defparam i2_3_lut_4_lut_adj_1469.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_3_lut_adj_1470 (.I0(\data_in_frame[9] [1]), .I1(\data_in_frame[9] [0]), 
            .I2(\data_in_frame[10] [7]), .I3(GND_net), .O(n44538));
    defparam i1_2_lut_3_lut_adj_1470.LUT_INIT = 16'h9696;
    SB_LUT4 i4_4_lut_adj_1471 (.I0(n45244), .I1(n44049), .I2(n44400), 
            .I3(n6_adj_4756), .O(n45477));
    defparam i4_4_lut_adj_1471.LUT_INIT = 16'h9669;
    SB_LUT4 i5_4_lut_adj_1472 (.I0(n41718), .I1(n41809), .I2(n40779), 
            .I3(n41701), .O(n12_adj_4757));
    defparam i5_4_lut_adj_1472.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1473 (.I0(n47339), .I1(n26693), .I2(n27979), 
            .I3(n40688), .O(n40676));
    defparam i1_2_lut_4_lut_adj_1473.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1474 (.I0(n62), .I1(n65), .I2(\data_in[0] [3]), 
            .I3(GND_net), .O(n33811));
    defparam i1_2_lut_3_lut_adj_1474.LUT_INIT = 16'h1010;
    SB_LUT4 i1_2_lut_3_lut_adj_1475 (.I0(n46024), .I1(\data_in_frame[17] [5]), 
            .I2(n44284), .I3(GND_net), .O(Kp_23__N_1811));
    defparam i1_2_lut_3_lut_adj_1475.LUT_INIT = 16'h6969;
    SB_LUT4 i6_4_lut_adj_1476 (.I0(n44355), .I1(n27475), .I2(n43932), 
            .I3(\data_in_frame[8] [1]), .O(n14_adj_4758));   // verilog/coms.v(76[16:43])
    defparam i6_4_lut_adj_1476.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1477 (.I0(n27461), .I1(n14_adj_4758), .I2(n10_adj_4734), 
            .I3(\data_in_frame[1] [3]), .O(n45753));   // verilog/coms.v(76[16:43])
    defparam i7_4_lut_adj_1477.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1478 (.I0(n40972), .I1(\data_in_frame[8] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n41711));
    defparam i1_2_lut_adj_1478.LUT_INIT = 16'h6666;
    SB_LUT4 i12_4_lut_adj_1479 (.I0(n40728), .I1(n27544), .I2(n45753), 
            .I3(n27554), .O(n28));
    defparam i12_4_lut_adj_1479.LUT_INIT = 16'hf7ff;
    SB_LUT4 i6_4_lut_adj_1480 (.I0(\data_out_frame[25] [7]), .I1(n12_adj_4757), 
            .I2(n44140), .I3(n41633), .O(n46198));
    defparam i6_4_lut_adj_1480.LUT_INIT = 16'h9669;
    SB_LUT4 i10_4_lut_adj_1481 (.I0(n27976), .I1(n27817), .I2(n27933), 
            .I3(n4_adj_4659), .O(n26_adj_4759));
    defparam i10_4_lut_adj_1481.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_3_lut_4_lut_adj_1482 (.I0(n62), .I1(n65), .I2(n19692), 
            .I3(n53), .O(n27061));
    defparam i1_3_lut_4_lut_adj_1482.LUT_INIT = 16'hf0e0;
    SB_LUT4 i5_4_lut_adj_1483 (.I0(\data_out_frame[23] [6]), .I1(n44193), 
            .I2(\data_out_frame[24] [1]), .I3(n44263), .O(n12_adj_4760));
    defparam i5_4_lut_adj_1483.LUT_INIT = 16'h9669;
    SB_LUT4 i6_4_lut_adj_1484 (.I0(\data_out_frame[24] [0]), .I1(n12_adj_4760), 
            .I2(n44472), .I3(\data_out_frame[21] [6]), .O(n45472));
    defparam i6_4_lut_adj_1484.LUT_INIT = 16'h9669;
    SB_LUT4 i11_4_lut (.I0(n27979), .I1(n27506), .I2(n40688), .I3(n41711), 
            .O(n27_adj_4761));
    defparam i11_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i9_4_lut_adj_1485 (.I0(n27850), .I1(n27820), .I2(n44243), 
            .I3(n8_adj_4672), .O(n25));
    defparam i9_4_lut_adj_1485.LUT_INIT = 16'hffef;
    SB_LUT4 i15_4_lut_adj_1486 (.I0(n25), .I1(n27_adj_4761), .I2(n26_adj_4759), 
            .I3(n28), .O(n31_adj_4748));
    defparam i15_4_lut_adj_1486.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_3_lut_adj_1487 (.I0(n27457), .I1(n28288), .I2(\data_in_frame[12] [3]), 
            .I3(GND_net), .O(n6_adj_4674));
    defparam i1_2_lut_3_lut_adj_1487.LUT_INIT = 16'h9696;
    SB_LUT4 i1_3_lut_4_lut_adj_1488 (.I0(n27979), .I1(\data_in_frame[10] [6]), 
            .I2(\data_in_frame[12] [7]), .I3(n47519), .O(n47523));   // verilog/coms.v(72[16:27])
    defparam i1_3_lut_4_lut_adj_1488.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1489 (.I0(\FRAME_MATCHER.state [3]), .I1(\FRAME_MATCHER.state [0]), 
            .I2(GND_net), .I3(GND_net), .O(n47565));
    defparam i1_2_lut_adj_1489.LUT_INIT = 16'heeee;
    SB_LUT4 i4630_3_lut (.I0(n31), .I1(n31_adj_4748), .I2(\FRAME_MATCHER.state [1]), 
            .I3(GND_net), .O(n23931));
    defparam i4630_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34915_4_lut (.I0(n43719), .I1(n23931), .I2(n24450), .I3(n47567), 
            .O(n28531));
    defparam i34915_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 mux_2094_i1_3_lut (.I0(\data_in_frame[19] [0]), .I1(\data_in_frame[3] [0]), 
            .I2(n7569), .I3(GND_net), .O(n7570));
    defparam mux_2094_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut_4_lut_adj_1490 (.I0(Kp_23__N_1253), .I1(\data_in_frame[8] [7]), 
            .I2(n26693), .I3(n40676), .O(n44620));
    defparam i1_3_lut_4_lut_adj_1490.LUT_INIT = 16'h9669;
    SB_LUT4 i2_3_lut_4_lut_adj_1491 (.I0(\data_in_frame[18] [3]), .I1(\data_in_frame[18] [1]), 
            .I2(n44559), .I3(\data_in_frame[18] [5]), .O(n43992));   // verilog/coms.v(79[16:27])
    defparam i2_3_lut_4_lut_adj_1491.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1492 (.I0(\data_out_frame[21] [7]), .I1(n45503), 
            .I2(GND_net), .I3(GND_net), .O(n44193));
    defparam i1_2_lut_adj_1492.LUT_INIT = 16'h9999;
    SB_LUT4 i3_4_lut_adj_1493 (.I0(n2326), .I1(n46018), .I2(n44193), .I3(n43929), 
            .O(n44140));
    defparam i3_4_lut_adj_1493.LUT_INIT = 16'h9669;
    SB_LUT4 select_686_Select_10_i3_2_lut (.I0(\FRAME_MATCHER.i [10]), .I1(n4141), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4709));
    defparam select_686_Select_10_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_3_lut_adj_1494 (.I0(n27590), .I1(\data_in_frame[5] [6]), 
            .I2(n44589), .I3(GND_net), .O(n6_adj_4673));   // verilog/coms.v(97[12:25])
    defparam i1_2_lut_3_lut_adj_1494.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_4_lut_adj_1495 (.I0(\data_in_frame[20] [6]), .I1(\data_in_frame[20] [7]), 
            .I2(n40734), .I3(\data_in_frame[18] [7]), .O(n44459));
    defparam i1_2_lut_4_lut_adj_1495.LUT_INIT = 16'h6996;
    SB_LUT4 select_686_Select_11_i3_2_lut (.I0(\FRAME_MATCHER.i [11]), .I1(n4141), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4708));
    defparam select_686_Select_11_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i5_3_lut_4_lut_adj_1496 (.I0(\data_in_frame[13] [7]), .I1(n41598), 
            .I2(n10_adj_4665), .I3(n41644), .O(n44453));
    defparam i5_3_lut_4_lut_adj_1496.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1497 (.I0(\data_in[3] [4]), .I1(n10_adj_4717), 
            .I2(\data_in[2] [7]), .I3(\data_in[2] [4]), .O(n6_adj_4718));
    defparam i1_2_lut_4_lut_adj_1497.LUT_INIT = 16'hffdf;
    SB_LUT4 i1_2_lut_4_lut_adj_1498 (.I0(\data_in[3] [4]), .I1(n10_adj_4717), 
            .I2(\data_in[2] [7]), .I3(\data_in[1] [5]), .O(n12_adj_4712));
    defparam i1_2_lut_4_lut_adj_1498.LUT_INIT = 16'hffdf;
    SB_LUT4 i1_2_lut_4_lut_adj_1499 (.I0(\data_in[1] [0]), .I1(\data_in[0] [6]), 
            .I2(\data_in[3] [0]), .I3(n33811), .O(n33827));
    defparam i1_2_lut_4_lut_adj_1499.LUT_INIT = 16'hdfff;
    SB_LUT4 i1_2_lut_4_lut_adj_1500 (.I0(\data_in[1] [0]), .I1(\data_in[0] [6]), 
            .I2(\data_in[3] [0]), .I3(\data_in[0] [3]), .O(n53));
    defparam i1_2_lut_4_lut_adj_1500.LUT_INIT = 16'hdfff;
    SB_LUT4 select_686_Select_12_i3_2_lut (.I0(\FRAME_MATCHER.i [12]), .I1(n4141), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4705));
    defparam select_686_Select_12_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 equal_299_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8_adj_4645));   // verilog/coms.v(155[7:23])
    defparam equal_299_i8_2_lut_3_lut.LUT_INIT = 16'hefef;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_35873 (.I0(byte_transmit_counter[3]), 
            .I1(n51255), .I2(n49351), .I3(byte_transmit_counter[4]), .O(n51510));
    defparam byte_transmit_counter_3__bdd_4_lut_35873.LUT_INIT = 16'he4aa;
    SB_LUT4 equal_300_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8_adj_4729));   // verilog/coms.v(155[7:23])
    defparam equal_300_i8_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 n51510_bdd_4_lut (.I0(n51510), .I1(n51273), .I2(n7_adj_4762), 
            .I3(byte_transmit_counter[4]), .O(tx_data[0]));
    defparam n51510_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i15418_3_lut_4_lut (.I0(n8_adj_4645), .I1(n43841), .I2(rx_data[5]), 
            .I3(\data_in_frame[9] [5]), .O(n29366));
    defparam i15418_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15419_3_lut_4_lut (.I0(n8_adj_4645), .I1(n43841), .I2(rx_data[4]), 
            .I3(\data_in_frame[9] [4]), .O(n29367));
    defparam i15419_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15420_3_lut_4_lut (.I0(n8_adj_4645), .I1(n43841), .I2(rx_data[3]), 
            .I3(\data_in_frame[9] [3]), .O(n29368));
    defparam i15420_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15421_3_lut_4_lut (.I0(n8_adj_4645), .I1(n43841), .I2(rx_data[2]), 
            .I3(\data_in_frame[9] [2]), .O(n29369));
    defparam i15421_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15489_3_lut_4_lut (.I0(n8_adj_4729), .I1(n43832), .I2(rx_data[7]), 
            .I3(\data_in_frame[0] [7]), .O(n29437));
    defparam i15489_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15490_3_lut_4_lut (.I0(n8_adj_4729), .I1(n43832), .I2(rx_data[6]), 
            .I3(\data_in_frame[0] [6]), .O(n29438));
    defparam i15490_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15491_3_lut_4_lut (.I0(n8_adj_4729), .I1(n43832), .I2(rx_data[5]), 
            .I3(\data_in_frame[0] [5]), .O(n29439));
    defparam i15491_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 select_686_Select_13_i3_2_lut (.I0(\FRAME_MATCHER.i [13]), .I1(n4141), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4703));
    defparam select_686_Select_13_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i15422_3_lut_4_lut (.I0(n8_adj_4645), .I1(n43841), .I2(rx_data[1]), 
            .I3(\data_in_frame[9] [1]), .O(n29370));
    defparam i15422_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15492_3_lut_4_lut (.I0(n8_adj_4729), .I1(n43832), .I2(rx_data[4]), 
            .I3(\data_in_frame[0] [4]), .O(n29440));
    defparam i15492_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i4_4_lut_adj_1501 (.I0(n44211), .I1(n40764), .I2(n41801), 
            .I3(n44482), .O(n10_adj_4763));
    defparam i4_4_lut_adj_1501.LUT_INIT = 16'h9669;
    SB_LUT4 i5_3_lut_adj_1502 (.I0(n41171), .I1(n10_adj_4763), .I2(n41723), 
            .I3(GND_net), .O(n2326));
    defparam i5_3_lut_adj_1502.LUT_INIT = 16'h6969;
    SB_LUT4 i4_4_lut_adj_1503 (.I0(n44187), .I1(n41615), .I2(n41805), 
            .I3(n44468), .O(n10_adj_4747));
    defparam i4_4_lut_adj_1503.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_3_lut_adj_1504 (.I0(\data_in_frame[13] [4]), .I1(\data_in_frame[18] [0]), 
            .I2(n27536), .I3(GND_net), .O(n6_adj_4658));   // verilog/coms.v(71[16:27])
    defparam i1_2_lut_3_lut_adj_1504.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1505 (.I0(\data_in_frame[15] [6]), .I1(\data_in_frame[17] [7]), 
            .I2(\data_in_frame[17] [6]), .I3(GND_net), .O(n43954));   // verilog/coms.v(71[16:27])
    defparam i1_2_lut_3_lut_adj_1505.LUT_INIT = 16'h9696;
    SB_LUT4 select_686_Select_14_i3_2_lut (.I0(\FRAME_MATCHER.i [14]), .I1(n4141), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4700));
    defparam select_686_Select_14_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i15493_3_lut_4_lut (.I0(n8_adj_4729), .I1(n43832), .I2(rx_data[3]), 
            .I3(\data_in_frame[0] [3]), .O(n29441));
    defparam i15493_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15423_3_lut_4_lut (.I0(n8_adj_4645), .I1(n43841), .I2(rx_data[0]), 
            .I3(\data_in_frame[9] [0]), .O(n29371));
    defparam i15423_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15494_3_lut_4_lut (.I0(n8_adj_4729), .I1(n43832), .I2(rx_data[2]), 
            .I3(\data_in_frame[0] [2]), .O(n29442));
    defparam i15494_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1506 (.I0(\data_in_frame[13] [7]), .I1(\data_in_frame[13] [6]), 
            .I2(\data_in_frame[15] [1]), .I3(GND_net), .O(n47851));
    defparam i1_2_lut_3_lut_adj_1506.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_4_lut_adj_1507 (.I0(\data_in_frame[19] [2]), .I1(n27668), 
            .I2(n46393), .I3(\data_in_frame[19] [4]), .O(n44196));
    defparam i1_2_lut_4_lut_adj_1507.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1508 (.I0(\data_out_frame[4] [6]), .I1(\data_out_frame[5] [0]), 
            .I2(\data_out_frame[11] [2]), .I3(n4_adj_4764), .O(n44522));   // verilog/coms.v(86[17:28])
    defparam i2_3_lut_4_lut_adj_1508.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1509 (.I0(n45489), .I1(n44029), .I2(\data_out_frame[20] [1]), 
            .I3(GND_net), .O(n45721));
    defparam i2_3_lut_adj_1509.LUT_INIT = 16'h6969;
    SB_LUT4 i15495_3_lut_4_lut (.I0(n8_adj_4729), .I1(n43832), .I2(rx_data[1]), 
            .I3(\data_in_frame[0] [1]), .O(n29443));
    defparam i15495_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i3_4_lut_adj_1510 (.I0(n41633), .I1(n44281), .I2(\data_out_frame[25] [0]), 
            .I3(\data_out_frame[24] [5]), .O(n45796));
    defparam i3_4_lut_adj_1510.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1511 (.I0(n27599), .I1(n2520), .I2(GND_net), 
            .I3(GND_net), .O(n44281));
    defparam i1_2_lut_adj_1511.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1512 (.I0(n40836), .I1(n44281), .I2(n44149), 
            .I3(n41701), .O(n45804));
    defparam i3_4_lut_adj_1512.LUT_INIT = 16'h6996;
    SB_LUT4 i15096_3_lut_4_lut (.I0(n8_adj_4729), .I1(n43832), .I2(rx_data[0]), 
            .I3(\data_in_frame[0] [0]), .O(n29044));
    defparam i15096_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_4_lut_adj_1513 (.I0(\FRAME_MATCHER.i [4]), .I1(\FRAME_MATCHER.i [5]), 
            .I2(\FRAME_MATCHER.i [3]), .I3(n35014), .O(n43841));   // verilog/coms.v(155[7:23])
    defparam i2_3_lut_4_lut_adj_1513.LUT_INIT = 16'hefff;
    SB_LUT4 i2_3_lut_4_lut_adj_1514 (.I0(\FRAME_MATCHER.i [4]), .I1(\FRAME_MATCHER.i [5]), 
            .I2(\FRAME_MATCHER.i [3]), .I3(n35014), .O(n43832));   // verilog/coms.v(155[7:23])
    defparam i2_3_lut_4_lut_adj_1514.LUT_INIT = 16'hfeff;
    SB_LUT4 i1_2_lut_3_lut_adj_1515 (.I0(\data_in_frame[4] [6]), .I1(\data_in_frame[5] [0]), 
            .I2(n28228), .I3(GND_net), .O(n44000));   // verilog/coms.v(74[16:42])
    defparam i1_2_lut_3_lut_adj_1515.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1516 (.I0(\data_out_frame[25] [7]), .I1(\data_out_frame[25] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n44049));   // verilog/coms.v(72[16:27])
    defparam i1_2_lut_adj_1516.LUT_INIT = 16'h6666;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_35913 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [0]), .I2(\data_out_frame[27] [0]), 
            .I3(byte_transmit_counter[1]), .O(n51504));
    defparam byte_transmit_counter_0__bdd_4_lut_35913.LUT_INIT = 16'he4aa;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_0_i7_3_lut_4_lut (.I0(byte_transmit_counter[2]), 
            .I1(byte_transmit_counter[1]), .I2(n48187), .I3(n48185), .O(n7_adj_4762));   // verilog/coms.v(107[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_0_i7_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_1_i7_3_lut_4_lut (.I0(byte_transmit_counter[2]), 
            .I1(byte_transmit_counter[1]), .I2(n48055), .I3(n48053), .O(n7_adj_4755));   // verilog/coms.v(107[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_1_i7_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_2_i7_3_lut_4_lut (.I0(byte_transmit_counter[2]), 
            .I1(byte_transmit_counter[1]), .I2(n48049), .I3(n48047), .O(n7_adj_4750));   // verilog/coms.v(107[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_2_i7_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 i1_2_lut_adj_1517 (.I0(\data_out_frame[22] [1]), .I1(n41472), 
            .I2(GND_net), .I3(GND_net), .O(n44187));
    defparam i1_2_lut_adj_1517.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_3_lut_adj_1518 (.I0(n27756), .I1(\data_out_frame[18] [7]), 
            .I2(n40704), .I3(GND_net), .O(n41677));
    defparam i1_2_lut_3_lut_adj_1518.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_1519 (.I0(n43861), .I1(n44476), .I2(n44202), 
            .I3(n44084), .O(n45489));
    defparam i3_4_lut_adj_1519.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1520 (.I0(\data_out_frame[21] [5]), .I1(n44226), 
            .I2(n44406), .I3(\data_out_frame[19] [3]), .O(n44472));
    defparam i1_4_lut_adj_1520.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1521 (.I0(\data_out_frame[23] [7]), .I1(n44472), 
            .I2(GND_net), .I3(GND_net), .O(n43929));   // verilog/coms.v(79[16:27])
    defparam i1_2_lut_adj_1521.LUT_INIT = 16'h6666;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_3_i7_3_lut_4_lut (.I0(byte_transmit_counter[2]), 
            .I1(byte_transmit_counter[1]), .I2(n48307), .I3(n48305), .O(n7_adj_4749));   // verilog/coms.v(107[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_3_i7_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 n51504_bdd_4_lut (.I0(n51504), .I1(\data_out_frame[25] [0]), 
            .I2(\data_out_frame[24] [0]), .I3(byte_transmit_counter[1]), 
            .O(n51507));
    defparam n51504_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_adj_1522 (.I0(\data_out_frame[24] [1]), .I1(\data_out_frame[24] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n44032));   // verilog/coms.v(75[16:43])
    defparam i1_2_lut_adj_1522.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1523 (.I0(\data_out_frame[23] [4]), .I1(\data_out_frame[23] [6]), 
            .I2(n27406), .I3(GND_net), .O(n44400));   // verilog/coms.v(79[16:27])
    defparam i2_3_lut_adj_1523.LUT_INIT = 16'h9696;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_4_i7_3_lut_4_lut (.I0(byte_transmit_counter[2]), 
            .I1(byte_transmit_counter[1]), .I2(n48220), .I3(n48218), .O(n7_adj_4740));   // verilog/coms.v(107[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_4_i7_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 i1_2_lut_3_lut_adj_1524 (.I0(\data_in_frame[1] [2]), .I1(\data_in_frame[1] [1]), 
            .I2(n43938), .I3(GND_net), .O(Kp_23__N_1027));   // verilog/coms.v(86[17:63])
    defparam i1_2_lut_3_lut_adj_1524.LUT_INIT = 16'h9696;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_7_i7_3_lut_4_lut (.I0(byte_transmit_counter[2]), 
            .I1(byte_transmit_counter[1]), .I2(n48196), .I3(n48194), .O(n7_adj_4730));   // verilog/coms.v(107[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_7_i7_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 i5_3_lut_4_lut_adj_1525 (.I0(n27756), .I1(\data_out_frame[18] [7]), 
            .I2(\data_out_frame[16] [3]), .I3(n10_adj_4765), .O(n41472));
    defparam i5_3_lut_4_lut_adj_1525.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1526 (.I0(n27326), .I1(\data_out_frame[19] [6]), 
            .I2(\data_out_frame[19] [7]), .I3(\data_out_frame[20] [0]), 
            .O(n14_adj_4766));
    defparam i6_4_lut_adj_1526.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1527 (.I0(n44119), .I1(n14_adj_4766), .I2(n10_adj_4736), 
            .I3(\data_out_frame[22] [2]), .O(n41829));
    defparam i7_4_lut_adj_1527.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1528 (.I0(n40638), .I1(n28009), .I2(\data_in_frame[10] [0]), 
            .I3(GND_net), .O(n41814));
    defparam i1_2_lut_3_lut_adj_1528.LUT_INIT = 16'h9696;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_6_i7_3_lut_4_lut (.I0(byte_transmit_counter[2]), 
            .I1(byte_transmit_counter[1]), .I2(n48205), .I3(n48203), .O(n7_adj_4735));   // verilog/coms.v(107[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_6_i7_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 i1_2_lut_4_lut_adj_1529 (.I0(n43980), .I1(\data_out_frame[14] [4]), 
            .I2(n27265), .I3(\data_out_frame[16] [6]), .O(n44302));   // verilog/coms.v(76[16:43])
    defparam i1_2_lut_4_lut_adj_1529.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1530 (.I0(n44290), .I1(n44507), .I2(n44161), 
            .I3(GND_net), .O(n41598));
    defparam i2_3_lut_adj_1530.LUT_INIT = 16'h9696;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_5_i7_3_lut_4_lut (.I0(byte_transmit_counter[2]), 
            .I1(byte_transmit_counter[1]), .I2(n48214), .I3(n48212), .O(n7_adj_4737));   // verilog/coms.v(107[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_5_i7_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 i1_2_lut_4_lut_adj_1531 (.I0(n43980), .I1(\data_out_frame[14] [4]), 
            .I2(n27265), .I3(\data_out_frame[16] [5]), .O(n27834));   // verilog/coms.v(76[16:43])
    defparam i1_2_lut_4_lut_adj_1531.LUT_INIT = 16'h6996;
    SB_LUT4 i2_2_lut_4_lut_adj_1532 (.I0(n43932), .I1(n44516), .I2(\data_in_frame[6] [2]), 
            .I3(n4_adj_4619), .O(n27976));   // verilog/coms.v(79[16:27])
    defparam i2_2_lut_4_lut_adj_1532.LUT_INIT = 16'h6996;
    SB_LUT4 i15397_3_lut_4_lut (.I0(n8_adj_4681), .I1(n43841), .I2(rx_data[2]), 
            .I3(\data_in_frame[12] [2]), .O(n29345));
    defparam i15397_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_4_lut_adj_1533 (.I0(n43932), .I1(n44516), .I2(\data_in_frame[6] [2]), 
            .I3(n44358), .O(n27506));   // verilog/coms.v(79[16:27])
    defparam i1_2_lut_4_lut_adj_1533.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_35864 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [7]), .I2(\data_out_frame[27] [7]), 
            .I3(byte_transmit_counter[1]), .O(n51498));
    defparam byte_transmit_counter_0__bdd_4_lut_35864.LUT_INIT = 16'he4aa;
    SB_LUT4 i2_3_lut_4_lut_adj_1534 (.I0(\data_out_frame[6] [3]), .I1(\data_out_frame[4] [1]), 
            .I2(\data_out_frame[4] [2]), .I3(\data_out_frame[8] [4]), .O(n43920));   // verilog/coms.v(76[16:43])
    defparam i2_3_lut_4_lut_adj_1534.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1535 (.I0(\data_out_frame[17] [2]), .I1(n28070), 
            .I2(n26718), .I3(n28314), .O(n44406));
    defparam i3_4_lut_adj_1535.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1536 (.I0(n44287), .I1(n27326), .I2(\data_out_frame[17] [5]), 
            .I3(GND_net), .O(n45596));
    defparam i2_3_lut_adj_1536.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1537 (.I0(\data_out_frame[6] [3]), .I1(\data_out_frame[4] [1]), 
            .I2(\data_out_frame[6] [4]), .I3(\data_out_frame[4] [3]), .O(n1247));   // verilog/coms.v(76[16:43])
    defparam i1_2_lut_3_lut_4_lut_adj_1537.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1538 (.I0(n45596), .I1(n44172), .I2(\data_out_frame[22] [0]), 
            .I3(\data_out_frame[19] [6]), .O(n45503));
    defparam i3_4_lut_adj_1538.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1539 (.I0(n44406), .I1(n44456), .I2(\data_out_frame[19] [4]), 
            .I3(GND_net), .O(n27406));
    defparam i2_3_lut_adj_1539.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1540 (.I0(\data_in_frame[10] [4]), .I1(n27976), 
            .I2(n4_adj_4659), .I3(GND_net), .O(n27873));   // verilog/coms.v(75[16:43])
    defparam i1_2_lut_3_lut_adj_1540.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_1541 (.I0(n27406), .I1(n45503), .I2(n46161), 
            .I3(\data_out_frame[21] [6]), .O(n44211));
    defparam i3_4_lut_adj_1541.LUT_INIT = 16'h9669;
    SB_LUT4 i2_2_lut_3_lut_4_lut_adj_1542 (.I0(\FRAME_MATCHER.state [1]), 
            .I1(n34607), .I2(r_SM_Main_2__N_3780[0]), .I3(tx_active), 
            .O(n6_adj_4767));
    defparam i2_2_lut_3_lut_4_lut_adj_1542.LUT_INIT = 16'hfff7;
    SB_LUT4 i21_4_lut_adj_1543 (.I0(n44262), .I1(n44125), .I2(n44208), 
            .I3(n43960), .O(n50_adj_4768));
    defparam i21_4_lut_adj_1543.LUT_INIT = 16'h6996;
    SB_LUT4 i19_4_lut_adj_1544 (.I0(n44485), .I1(n44580), .I2(n43905), 
            .I3(n44211), .O(n48_adj_4769));
    defparam i19_4_lut_adj_1544.LUT_INIT = 16'h6996;
    SB_LUT4 i20_4_lut_adj_1545 (.I0(n44029), .I1(n41829), .I2(n41661), 
            .I3(n44498), .O(n49));
    defparam i20_4_lut_adj_1545.LUT_INIT = 16'h6996;
    SB_LUT4 i35567_3_lut_4_lut (.I0(tx_active), .I1(r_SM_Main_2__N_3780[0]), 
            .I2(n63), .I3(n27235), .O(n28546));
    defparam i35567_3_lut_4_lut.LUT_INIT = 16'h0f1f;
    SB_LUT4 i18_4_lut_adj_1546 (.I0(\data_out_frame[24] [5]), .I1(n41801), 
            .I2(\data_out_frame[23] [2]), .I3(n44134), .O(n47_adj_4770));
    defparam i18_4_lut_adj_1546.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1547 (.I0(\data_out_frame[4] [3]), .I1(\data_out_frame[6] [4]), 
            .I2(\data_out_frame[4] [2]), .I3(GND_net), .O(n43974));   // verilog/coms.v(76[16:43])
    defparam i1_2_lut_3_lut_adj_1547.LUT_INIT = 16'h9696;
    SB_LUT4 i17_4_lut_adj_1548 (.I0(\data_out_frame[24] [6]), .I1(n44032), 
            .I2(n44541), .I3(\data_out_frame[24] [4]), .O(n46_adj_4771));
    defparam i17_4_lut_adj_1548.LUT_INIT = 16'h6996;
    SB_LUT4 i2_2_lut_4_lut_adj_1549 (.I0(n44183), .I1(n44465), .I2(n41751), 
            .I3(\data_in_frame[18] [7]), .O(n6_adj_4637));
    defparam i2_2_lut_4_lut_adj_1549.LUT_INIT = 16'h6996;
    SB_LUT4 i16_4_lut_adj_1550 (.I0(\data_out_frame[23] [3]), .I1(n43929), 
            .I2(n44605), .I3(\data_out_frame[23] [5]), .O(n45_adj_4772));
    defparam i16_4_lut_adj_1550.LUT_INIT = 16'h6996;
    SB_LUT4 i27_4_lut (.I0(n47_adj_4770), .I1(n49), .I2(n48_adj_4769), 
            .I3(n50_adj_4768), .O(n56));
    defparam i27_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i22_4_lut (.I0(\data_out_frame[22] [6]), .I1(\data_out_frame[22] [7]), 
            .I2(n45244), .I3(n30), .O(n51));
    defparam i22_4_lut.LUT_INIT = 16'h9669;
    SB_LUT4 i15408_3_lut_4_lut (.I0(n8), .I1(n43841), .I2(rx_data[7]), 
            .I3(\data_in_frame[10] [7]), .O(n29356));
    defparam i15408_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1551 (.I0(tx_active), .I1(r_SM_Main_2__N_3780[0]), 
            .I2(tx_transmit_N_3677), .I3(GND_net), .O(n2263));
    defparam i1_2_lut_3_lut_adj_1551.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_3_lut_4_lut_adj_1552 (.I0(n44020), .I1(n44394), .I2(\data_in_frame[6] [0]), 
            .I3(n44355), .O(n44094));   // verilog/coms.v(86[17:28])
    defparam i1_3_lut_4_lut_adj_1552.LUT_INIT = 16'h6996;
    SB_LUT4 i28_4_lut (.I0(n51), .I1(n56), .I2(n45_adj_4772), .I3(n46_adj_4771), 
            .O(n40779));
    defparam i28_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i15409_3_lut_4_lut (.I0(n8), .I1(n43841), .I2(rx_data[6]), 
            .I3(\data_in_frame[10] [6]), .O(n29357));
    defparam i15409_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i3_4_lut_adj_1553 (.I0(\data_out_frame[24] [0]), .I1(n40779), 
            .I2(n27279), .I3(n27599), .O(n40836));
    defparam i3_4_lut_adj_1553.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1554 (.I0(\data_out_frame[25] [5]), .I1(n44447), 
            .I2(n44152), .I3(n44049), .O(n2520));   // verilog/coms.v(72[16:27])
    defparam i3_4_lut_adj_1554.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1555 (.I0(n44143), .I1(n2520), .I2(n40836), .I3(n44444), 
            .O(n10_adj_4773));
    defparam i4_4_lut_adj_1555.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_1556 (.I0(n41693), .I1(n10_adj_4773), .I2(n45499), 
            .I3(GND_net), .O(n45371));
    defparam i5_3_lut_adj_1556.LUT_INIT = 16'h6969;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1557 (.I0(n27820), .I1(n27850), .I2(\data_in_frame[9] [3]), 
            .I3(\data_in_frame[9] [2]), .O(Kp_23__N_1468));   // verilog/coms.v(74[16:42])
    defparam i1_2_lut_3_lut_4_lut_adj_1557.LUT_INIT = 16'h6996;
    SB_LUT4 i15410_3_lut_4_lut (.I0(n8), .I1(n43841), .I2(rx_data[5]), 
            .I3(\data_in_frame[10] [5]), .O(n29358));
    defparam i15410_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1558 (.I0(\data_out_frame[15] [5]), .I1(\data_out_frame[17] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n44119));
    defparam i1_2_lut_adj_1558.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_4_lut_adj_1559 (.I0(\data_in_frame[9] [2]), .I1(\data_in_frame[9] [3]), 
            .I2(n44491), .I3(\data_in_frame[9] [4]), .O(n44574));   // verilog/coms.v(74[16:42])
    defparam i2_3_lut_4_lut_adj_1559.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1560 (.I0(\data_in_frame[9] [7]), .I1(\data_in_frame[9] [6]), 
            .I2(\data_in_frame[9] [5]), .I3(GND_net), .O(n44491));   // verilog/coms.v(86[17:28])
    defparam i1_2_lut_3_lut_adj_1560.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1561 (.I0(n52_adj_4626), .I1(n37), .I2(\FRAME_MATCHER.state [4]), 
            .I3(GND_net), .O(n43146));
    defparam i1_2_lut_3_lut_adj_1561.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1562 (.I0(n52_adj_4626), .I1(n37), .I2(\FRAME_MATCHER.state [5]), 
            .I3(GND_net), .O(n43150));
    defparam i1_2_lut_3_lut_adj_1562.LUT_INIT = 16'he0e0;
    SB_LUT4 i6_4_lut_adj_1563 (.I0(n44583), .I1(\data_out_frame[15] [6]), 
            .I2(n44254), .I3(\data_out_frame[15] [4]), .O(n14_adj_4774));
    defparam i6_4_lut_adj_1563.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1564 (.I0(\data_out_frame[18] [0]), .I1(n14_adj_4774), 
            .I2(n10_adj_4733), .I3(n44119), .O(n41171));
    defparam i7_4_lut_adj_1564.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1565 (.I0(\data_out_frame[20] [2]), .I1(n41171), 
            .I2(GND_net), .I3(GND_net), .O(n41661));
    defparam i1_2_lut_adj_1565.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_3_lut_adj_1566 (.I0(n52_adj_4626), .I1(n37), .I2(\FRAME_MATCHER.state [6]), 
            .I3(GND_net), .O(n43154));
    defparam i1_2_lut_3_lut_adj_1566.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1567 (.I0(n52_adj_4626), .I1(n37), .I2(\FRAME_MATCHER.state [7]), 
            .I3(GND_net), .O(n43156));
    defparam i1_2_lut_3_lut_adj_1567.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_adj_1568 (.I0(\data_out_frame[24] [6]), .I1(\data_out_frame[25] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n44149));
    defparam i1_2_lut_adj_1568.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_3_lut_adj_1569 (.I0(n52_adj_4626), .I1(n37), .I2(\FRAME_MATCHER.state [8]), 
            .I3(GND_net), .O(n43158));
    defparam i1_2_lut_3_lut_adj_1569.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1570 (.I0(n52_adj_4626), .I1(n37), .I2(\FRAME_MATCHER.state [9]), 
            .I3(GND_net), .O(n43160));
    defparam i1_2_lut_3_lut_adj_1570.LUT_INIT = 16'he0e0;
    SB_LUT4 i3_4_lut_adj_1571 (.I0(\data_out_frame[25] [1]), .I1(n44149), 
            .I2(n41701), .I3(n41693), .O(n45888));
    defparam i3_4_lut_adj_1571.LUT_INIT = 16'h6996;
    SB_LUT4 i15411_3_lut_4_lut (.I0(n8), .I1(n43841), .I2(rx_data[4]), 
            .I3(\data_in_frame[10] [4]), .O(n29359));
    defparam i15411_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15412_3_lut_4_lut (.I0(n8), .I1(n43841), .I2(rx_data[3]), 
            .I3(\data_in_frame[10] [3]), .O(n29360));
    defparam i15412_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1572 (.I0(n52_adj_4626), .I1(n37), .I2(\FRAME_MATCHER.state [10]), 
            .I3(GND_net), .O(n43162));
    defparam i1_2_lut_3_lut_adj_1572.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_3_lut_4_lut_adj_1573 (.I0(\FRAME_MATCHER.state [3]), .I1(n22132), 
            .I2(n4120), .I3(n37), .O(n43036));
    defparam i1_3_lut_4_lut_adj_1573.LUT_INIT = 16'haa80;
    SB_LUT4 i15413_3_lut_4_lut (.I0(n8), .I1(n43841), .I2(rx_data[2]), 
            .I3(\data_in_frame[10] [2]), .O(n29361));
    defparam i15413_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1574 (.I0(n52_adj_4626), .I1(n37), .I2(\FRAME_MATCHER.state [11]), 
            .I3(GND_net), .O(n43164));
    defparam i1_2_lut_3_lut_adj_1574.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1575 (.I0(n52_adj_4626), .I1(n37), .I2(\FRAME_MATCHER.state [12]), 
            .I3(GND_net), .O(n43166));
    defparam i1_2_lut_3_lut_adj_1575.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1576 (.I0(n52_adj_4626), .I1(n37), .I2(\FRAME_MATCHER.state [17]), 
            .I3(GND_net), .O(n43184));
    defparam i1_2_lut_3_lut_adj_1576.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1577 (.I0(n52_adj_4626), .I1(n37), .I2(\FRAME_MATCHER.state [18]), 
            .I3(GND_net), .O(n43186));
    defparam i1_2_lut_3_lut_adj_1577.LUT_INIT = 16'he0e0;
    SB_LUT4 i15414_3_lut_4_lut (.I0(n8), .I1(n43841), .I2(rx_data[1]), 
            .I3(\data_in_frame[10] [1]), .O(n29362));
    defparam i15414_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1578 (.I0(n52_adj_4626), .I1(n37), .I2(\FRAME_MATCHER.state [19]), 
            .I3(GND_net), .O(n43188));
    defparam i1_2_lut_3_lut_adj_1578.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1579 (.I0(n52_adj_4626), .I1(n37), .I2(\FRAME_MATCHER.state [20]), 
            .I3(GND_net), .O(n43190));
    defparam i1_2_lut_3_lut_adj_1579.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1580 (.I0(n52_adj_4626), .I1(n37), .I2(\FRAME_MATCHER.state [21]), 
            .I3(GND_net), .O(n43192));
    defparam i1_2_lut_3_lut_adj_1580.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1581 (.I0(n52_adj_4626), .I1(n37), .I2(\FRAME_MATCHER.state [22]), 
            .I3(GND_net), .O(n43194));
    defparam i1_2_lut_3_lut_adj_1581.LUT_INIT = 16'he0e0;
    SB_LUT4 i15415_3_lut_4_lut (.I0(n8), .I1(n43841), .I2(rx_data[0]), 
            .I3(\data_in_frame[10] [0]), .O(n29363));
    defparam i15415_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i6_4_lut_adj_1582 (.I0(n41637), .I1(n44416), .I2(n44583), 
            .I3(n28221), .O(n14_adj_4775));
    defparam i6_4_lut_adj_1582.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1583 (.I0(\data_out_frame[18] [1]), .I1(n14_adj_4775), 
            .I2(n10_adj_4745), .I3(n40636), .O(n41723));
    defparam i7_4_lut_adj_1583.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_4_lut_adj_1584 (.I0(\data_out_frame[12] [7]), .I1(\data_out_frame[12] [6]), 
            .I2(n10), .I3(n1191), .O(n26718));   // verilog/coms.v(86[17:28])
    defparam i5_3_lut_4_lut_adj_1584.LUT_INIT = 16'h6996;
    SB_LUT4 i20665_2_lut_3_lut (.I0(n52_adj_4626), .I1(n37), .I2(\FRAME_MATCHER.state [23]), 
            .I3(GND_net), .O(n34594));
    defparam i20665_2_lut_3_lut.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1585 (.I0(n52_adj_4626), .I1(n37), .I2(\FRAME_MATCHER.state [24]), 
            .I3(GND_net), .O(n43196));
    defparam i1_2_lut_3_lut_adj_1585.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1586 (.I0(n52_adj_4626), .I1(n37), .I2(\FRAME_MATCHER.state [25]), 
            .I3(GND_net), .O(n43198));
    defparam i1_2_lut_3_lut_adj_1586.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1587 (.I0(n52_adj_4626), .I1(n37), .I2(\FRAME_MATCHER.state [26]), 
            .I3(GND_net), .O(n43200));
    defparam i1_2_lut_3_lut_adj_1587.LUT_INIT = 16'he0e0;
    SB_LUT4 i2_3_lut_4_lut_adj_1588 (.I0(\data_out_frame[12] [7]), .I1(\data_out_frame[12] [6]), 
            .I2(\data_out_frame[12] [3]), .I3(n27261), .O(n44495));   // verilog/coms.v(86[17:28])
    defparam i2_3_lut_4_lut_adj_1588.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1589 (.I0(\FRAME_MATCHER.state_31__N_2808 [1]), 
            .I1(n4120), .I2(n27235), .I3(n2263), .O(n43032));
    defparam i1_2_lut_4_lut_adj_1589.LUT_INIT = 16'h8a88;
    SB_LUT4 select_719_Select_1_i1_3_lut_4_lut (.I0(n771), .I1(\FRAME_MATCHER.state [1]), 
            .I2(n27230), .I3(\FRAME_MATCHER.state_31__N_2808 [1]), .O(n1));
    defparam select_719_Select_1_i1_3_lut_4_lut.LUT_INIT = 16'h0302;
    SB_LUT4 n51498_bdd_4_lut (.I0(n51498), .I1(\data_out_frame[25] [7]), 
            .I2(\data_out_frame[24] [7]), .I3(byte_transmit_counter[1]), 
            .O(n51501));
    defparam n51498_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1590 (.I0(\data_in_frame[13] [0]), .I1(n44290), 
            .I2(n41059), .I3(\data_in_frame[9] [4]), .O(n6_adj_4663));
    defparam i1_2_lut_3_lut_4_lut_adj_1590.LUT_INIT = 16'h6996;
    SB_LUT4 i20666_2_lut_3_lut (.I0(n52_adj_4626), .I1(n37), .I2(\FRAME_MATCHER.state [27]), 
            .I3(GND_net), .O(n34596));
    defparam i20666_2_lut_3_lut.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_adj_1591 (.I0(\data_out_frame[24] [7]), .I1(n27279), 
            .I2(GND_net), .I3(GND_net), .O(n44605));   // verilog/coms.v(79[16:27])
    defparam i1_2_lut_adj_1591.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_3_lut_adj_1592 (.I0(n44183), .I1(n44465), .I2(n41751), 
            .I3(GND_net), .O(n44450));
    defparam i1_2_lut_3_lut_adj_1592.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1593 (.I0(\data_out_frame[20] [5]), .I1(\data_out_frame[20] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n44568));
    defparam i1_2_lut_adj_1593.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1594 (.I0(\data_out_frame[20] [2]), .I1(\data_out_frame[20] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n44319));
    defparam i1_2_lut_adj_1594.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_4_lut_adj_1595 (.I0(\data_out_frame[4] [7]), .I1(\data_out_frame[7] [1]), 
            .I2(n1168), .I3(\data_out_frame[8] [7]), .O(n43917));   // verilog/coms.v(72[16:69])
    defparam i1_2_lut_4_lut_adj_1595.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1596 (.I0(n41302), .I1(\data_in_frame[17] [0]), 
            .I2(n44217), .I3(GND_net), .O(n41751));
    defparam i1_2_lut_3_lut_adj_1596.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1597 (.I0(n52_adj_4626), .I1(n37), .I2(\FRAME_MATCHER.state [28]), 
            .I3(GND_net), .O(n43202));
    defparam i1_2_lut_3_lut_adj_1597.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1598 (.I0(n52_adj_4626), .I1(n37), .I2(\FRAME_MATCHER.state [29]), 
            .I3(GND_net), .O(n43206));
    defparam i1_2_lut_3_lut_adj_1598.LUT_INIT = 16'he0e0;
    SB_LUT4 i9_4_lut_adj_1599 (.I0(n44319), .I1(n44519), .I2(n44586), 
            .I3(n44190), .O(n23_adj_4776));
    defparam i9_4_lut_adj_1599.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut_adj_1600 (.I0(\data_out_frame[23] [0]), .I1(n44568), 
            .I2(n28400), .I3(\data_out_frame[22] [7]), .O(n22_adj_4777));
    defparam i8_4_lut_adj_1600.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1601 (.I0(n52_adj_4626), .I1(n37), .I2(\FRAME_MATCHER.state [30]), 
            .I3(GND_net), .O(n43208));
    defparam i1_2_lut_3_lut_adj_1601.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1602 (.I0(n52_adj_4626), .I1(n37), .I2(\FRAME_MATCHER.state [31]), 
            .I3(GND_net), .O(n43210));
    defparam i1_2_lut_3_lut_adj_1602.LUT_INIT = 16'he0e0;
    SB_LUT4 i12_4_lut_adj_1603 (.I0(n23_adj_4776), .I1(n19_adj_4746), .I2(n41807), 
            .I3(n44278), .O(n26_adj_4778));
    defparam i12_4_lut_adj_1603.LUT_INIT = 16'h9669;
    SB_LUT4 i13_4_lut_adj_1604 (.I0(n46020), .I1(n26_adj_4778), .I2(n22_adj_4777), 
            .I3(n41642), .O(n41693));
    defparam i13_4_lut_adj_1604.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1605 (.I0(\data_out_frame[25] [1]), .I1(\data_out_frame[25] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n44447));
    defparam i1_2_lut_adj_1605.LUT_INIT = 16'h6666;
    SB_LUT4 i15398_3_lut_4_lut (.I0(n8_adj_4681), .I1(n43841), .I2(rx_data[1]), 
            .I3(\data_in_frame[12] [1]), .O(n29346));
    defparam i15398_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_4_lut_adj_1606 (.I0(\data_out_frame[4] [7]), .I1(\data_out_frame[7] [1]), 
            .I2(n1168), .I3(\data_out_frame[9] [4]), .O(n6_adj_4603));   // verilog/coms.v(72[16:69])
    defparam i1_2_lut_4_lut_adj_1606.LUT_INIT = 16'h6996;
    SB_LUT4 i1_3_lut_4_lut_adj_1607 (.I0(n33827), .I1(n19692), .I2(n27235), 
            .I3(n2263), .O(n52_adj_4626));
    defparam i1_3_lut_4_lut_adj_1607.LUT_INIT = 16'h0800;
    SB_LUT4 i3_4_lut_adj_1608 (.I0(\data_out_frame[22] [6]), .I1(n44605), 
            .I2(n41615), .I3(n41596), .O(n44143));
    defparam i3_4_lut_adj_1608.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1609 (.I0(n33827), .I1(n19692), .I2(n27232), 
            .I3(n771), .O(n48_adj_4649));
    defparam i1_2_lut_3_lut_4_lut_adj_1609.LUT_INIT = 16'h0008;
    SB_LUT4 i2_3_lut_adj_1610 (.I0(n44143), .I1(n44447), .I2(n41693), 
            .I3(GND_net), .O(n45375));
    defparam i2_3_lut_adj_1610.LUT_INIT = 16'h6969;
    SB_LUT4 i1_2_lut_adj_1611 (.I0(n27809), .I1(\data_out_frame[16] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n44416));
    defparam i1_2_lut_adj_1611.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_4_lut_adj_1612 (.I0(\FRAME_MATCHER.state [1]), .I1(n44829), 
            .I2(\FRAME_MATCHER.state [3]), .I3(n44724), .O(n28621));   // verilog/coms.v(128[12] 303[6])
    defparam i2_3_lut_4_lut_adj_1612.LUT_INIT = 16'h0010;
    SB_LUT4 i5_4_lut_adj_1613 (.I0(n44416), .I1(n44553), .I2(n45977), 
            .I3(n44275), .O(n12_adj_4779));
    defparam i5_4_lut_adj_1613.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1614 (.I0(n33827), .I1(n19692), .I2(n27230), 
            .I3(n771), .O(n4_adj_4647));
    defparam i1_2_lut_3_lut_4_lut_adj_1614.LUT_INIT = 16'h0008;
    SB_LUT4 i1_2_lut_3_lut_adj_1615 (.I0(n27004), .I1(n34607), .I2(n24234), 
            .I3(GND_net), .O(n43729));
    defparam i1_2_lut_3_lut_adj_1615.LUT_INIT = 16'h4040;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1616 (.I0(n27004), .I1(n34607), .I2(n22132), 
            .I3(n3303), .O(n43795));
    defparam i1_2_lut_3_lut_4_lut_adj_1616.LUT_INIT = 16'h0040;
    SB_LUT4 i1_2_lut_3_lut_adj_1617 (.I0(n44263), .I1(n27998), .I2(n44472), 
            .I3(GND_net), .O(n6_adj_4756));
    defparam i1_2_lut_3_lut_adj_1617.LUT_INIT = 16'h6969;
    SB_LUT4 i1_3_lut_4_lut_adj_1618 (.I0(\data_in_frame[13] [2]), .I1(\data_in_frame[13] [0]), 
            .I2(\data_in_frame[15] [2]), .I3(\data_in_frame[12] [6]), .O(n47743));
    defparam i1_3_lut_4_lut_adj_1618.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1619 (.I0(\data_out_frame[16] [1]), .I1(n12_adj_4779), 
            .I2(\data_out_frame[18] [2]), .I3(\data_out_frame[15] [6]), 
            .O(n40636));
    defparam i6_4_lut_adj_1619.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1620 (.I0(n41801), .I1(n40636), .I2(GND_net), 
            .I3(GND_net), .O(n40764));
    defparam i1_2_lut_adj_1620.LUT_INIT = 16'h9999;
    SB_LUT4 i1_2_lut_adj_1621 (.I0(\data_out_frame[20] [6]), .I1(\data_out_frame[20] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n44468));
    defparam i1_2_lut_adj_1621.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1622 (.I0(\data_out_frame[23] [1]), .I1(\data_out_frame[23] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n44541));   // verilog/coms.v(79[16:27])
    defparam i1_2_lut_adj_1622.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1623 (.I0(n43861), .I1(n44042), .I2(n27771), 
            .I3(\data_out_frame[17] [3]), .O(n44456));
    defparam i3_4_lut_adj_1623.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1624 (.I0(\data_out_frame[15] [3]), .I1(n44435), 
            .I2(n27885), .I3(GND_net), .O(n44172));
    defparam i2_3_lut_adj_1624.LUT_INIT = 16'h9696;
    SB_LUT4 i1_3_lut_4_lut_adj_1625 (.I0(\data_in_frame[0] [5]), .I1(n27454), 
            .I2(n43938), .I3(\data_in_frame[1] [0]), .O(n26199));   // verilog/coms.v(78[16:27])
    defparam i1_3_lut_4_lut_adj_1625.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1626 (.I0(\data_out_frame[16] [0]), .I1(\data_out_frame[18] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n44501));
    defparam i1_2_lut_adj_1626.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1627 (.I0(\data_out_frame[19] [7]), .I1(\data_out_frame[17] [5]), 
            .I2(\data_out_frame[18] [0]), .I3(GND_net), .O(n44476));
    defparam i2_3_lut_adj_1627.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_4_lut_adj_1628 (.I0(n27834), .I1(\data_out_frame[18] [5]), 
            .I2(\data_out_frame[16] [3]), .I3(n40704), .O(n41642));
    defparam i1_2_lut_4_lut_adj_1628.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1629 (.I0(\data_out_frame[15] [4]), .I1(\data_out_frame[15] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n27326));
    defparam i1_2_lut_adj_1629.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1630 (.I0(\data_out_frame[15] [1]), .I1(\data_out_frame[15] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n27771));
    defparam i1_2_lut_adj_1630.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1631 (.I0(\data_out_frame[13] [4]), .I1(n44522), 
            .I2(n43917), .I3(\data_out_frame[11] [3]), .O(n10_adj_4744));
    defparam i4_4_lut_adj_1631.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1632 (.I0(\data_in_frame[13] [2]), .I1(\data_in_frame[13] [0]), 
            .I2(\data_in_frame[15] [7]), .I3(GND_net), .O(n44507));
    defparam i1_2_lut_3_lut_adj_1632.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1633 (.I0(\data_out_frame[18] [5]), .I1(\data_out_frame[16] [3]), 
            .I2(n40704), .I3(GND_net), .O(n44208));
    defparam i1_2_lut_3_lut_adj_1633.LUT_INIT = 16'h9696;
    SB_LUT4 i5_3_lut_adj_1634 (.I0(\data_out_frame[10] [6]), .I1(\data_out_frame[9] [0]), 
            .I2(\data_out_frame[8] [6]), .I3(GND_net), .O(n14_adj_4780));   // verilog/coms.v(75[16:43])
    defparam i5_3_lut_adj_1634.LUT_INIT = 16'h9696;
    SB_LUT4 i6_4_lut_adj_1635 (.I0(n44322), .I1(\data_out_frame[13] [2]), 
            .I2(\data_out_frame[11] [0]), .I3(n43911), .O(n15_adj_4781));   // verilog/coms.v(75[16:43])
    defparam i6_4_lut_adj_1635.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut_adj_1636 (.I0(n15_adj_4781), .I1(\data_out_frame[8] [4]), 
            .I2(n14_adj_4780), .I3(n1130), .O(n27885));   // verilog/coms.v(75[16:43])
    defparam i8_4_lut_adj_1636.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1637 (.I0(n44263), .I1(n27998), .I2(\data_out_frame[23] [5]), 
            .I3(GND_net), .O(n27599));
    defparam i1_2_lut_3_lut_adj_1637.LUT_INIT = 16'h6969;
    SB_LUT4 i15365_3_lut_4_lut (.I0(n35263), .I1(n43841), .I2(rx_data[7]), 
            .I3(\data_in_frame[15] [7]), .O(n29313));
    defparam i15365_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5_3_lut_4_lut_adj_1638 (.I0(\data_out_frame[7] [5]), .I1(n28046), 
            .I2(n10_adj_4618), .I3(n44003), .O(n40704));
    defparam i5_3_lut_4_lut_adj_1638.LUT_INIT = 16'h6996;
    SB_LUT4 i15366_3_lut_4_lut (.I0(n35263), .I1(n43841), .I2(rx_data[6]), 
            .I3(\data_in_frame[15] [6]), .O(n29314));
    defparam i15366_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2_3_lut_4_lut_adj_1639 (.I0(\data_out_frame[4] [7]), .I1(\data_out_frame[5] [2]), 
            .I2(\data_out_frame[5] [1]), .I3(\data_out_frame[7] [3]), .O(n28046));
    defparam i2_3_lut_4_lut_adj_1639.LUT_INIT = 16'h6996;
    SB_LUT4 i15400_3_lut_4_lut (.I0(n8_adj_4655), .I1(n43841), .I2(rx_data[7]), 
            .I3(\data_in_frame[11] [7]), .O(n29348));
    defparam i15400_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_adj_1640 (.I0(\data_out_frame[11] [1]), .I1(\data_out_frame[8] [7]), 
            .I2(\data_out_frame[8] [5]), .I3(GND_net), .O(n43911));
    defparam i2_3_lut_adj_1640.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1641 (.I0(\data_out_frame[8] [0]), .I1(\data_out_frame[7] [7]), 
            .I2(\data_out_frame[7] [6]), .I3(GND_net), .O(n28177));   // verilog/coms.v(76[16:27])
    defparam i1_2_lut_3_lut_adj_1641.LUT_INIT = 16'h9696;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_35637 (.I0(byte_transmit_counter[1]), 
            .I1(n48041), .I2(n48042), .I3(byte_transmit_counter[2]), .O(n51210));
    defparam byte_transmit_counter_1__bdd_4_lut_35637.LUT_INIT = 16'he4aa;
    SB_LUT4 i15367_3_lut_4_lut (.I0(n35263), .I1(n43841), .I2(rx_data[5]), 
            .I3(\data_in_frame[15] [5]), .O(n29315));
    defparam i15367_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4_4_lut_adj_1642 (.I0(n44388), .I1(n43911), .I2(\data_out_frame[13] [3]), 
            .I3(n44522), .O(n10_adj_4728));
    defparam i4_4_lut_adj_1642.LUT_INIT = 16'h6996;
    SB_LUT4 i15368_3_lut_4_lut (.I0(n35263), .I1(n43841), .I2(rx_data[4]), 
            .I3(\data_in_frame[15] [4]), .O(n29316));
    defparam i15368_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i15401_3_lut_4_lut (.I0(n8_adj_4655), .I1(n43841), .I2(rx_data[6]), 
            .I3(\data_in_frame[11] [6]), .O(n29349));
    defparam i15401_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i5_3_lut_adj_1643 (.I0(n44015), .I1(n10_adj_4728), .I2(\data_out_frame[9] [1]), 
            .I3(GND_net), .O(n28221));
    defparam i5_3_lut_adj_1643.LUT_INIT = 16'h9696;
    SB_LUT4 i15369_3_lut_4_lut (.I0(n35263), .I1(n43841), .I2(rx_data[3]), 
            .I3(\data_in_frame[15] [3]), .O(n29317));
    defparam i15369_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i15370_3_lut_4_lut (.I0(n35263), .I1(n43841), .I2(rx_data[2]), 
            .I3(\data_in_frame[15] [2]), .O(n29318));
    defparam i15370_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i6_4_lut_adj_1644 (.I0(\data_out_frame[13] [1]), .I1(n43920), 
            .I2(n27745), .I3(n44388), .O(n16_adj_4782));   // verilog/coms.v(77[16:43])
    defparam i6_4_lut_adj_1644.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1645 (.I0(\data_out_frame[6] [1]), .I1(n44328), 
            .I2(\data_out_frame[8] [3]), .I3(\data_out_frame[4] [0]), .O(n17_adj_4783));   // verilog/coms.v(77[16:43])
    defparam i7_4_lut_adj_1645.LUT_INIT = 16'h6996;
    SB_LUT4 i9_4_lut_adj_1646 (.I0(n17_adj_4783), .I1(\data_out_frame[11] [0]), 
            .I2(n16_adj_4782), .I3(\data_out_frame[8] [5]), .O(n43861));   // verilog/coms.v(77[16:43])
    defparam i9_4_lut_adj_1646.LUT_INIT = 16'h6996;
    SB_LUT4 i15371_3_lut_4_lut (.I0(n35263), .I1(n43841), .I2(rx_data[1]), 
            .I3(\data_in_frame[15] [1]), .O(n29319));
    defparam i15371_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2_3_lut_adj_1647 (.I0(\data_out_frame[12] [7]), .I1(\data_out_frame[5] [7]), 
            .I2(\data_out_frame[10] [5]), .I3(GND_net), .O(n44328));   // verilog/coms.v(77[16:43])
    defparam i2_3_lut_adj_1647.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1648 (.I0(\data_out_frame[13] [0]), .I1(n26718), 
            .I2(GND_net), .I3(GND_net), .O(n40665));
    defparam i1_2_lut_adj_1648.LUT_INIT = 16'h6666;
    SB_LUT4 i15372_3_lut_4_lut (.I0(n35263), .I1(n43841), .I2(rx_data[0]), 
            .I3(\data_in_frame[15] [0]), .O(n29320));
    defparam i15372_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i10_4_lut_adj_1649 (.I0(n40665), .I1(n44328), .I2(n44055), 
            .I3(\data_out_frame[10] [3]), .O(n28_adj_4784));
    defparam i10_4_lut_adj_1649.LUT_INIT = 16'h6996;
    SB_LUT4 i15402_3_lut_4_lut (.I0(n8_adj_4655), .I1(n43841), .I2(rx_data[5]), 
            .I3(\data_in_frame[11] [5]), .O(n29350));
    defparam i15402_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13_4_lut_adj_1650 (.I0(n44026), .I1(n27756), .I2(n43896), 
            .I3(n27248), .O(n31_adj_4785));
    defparam i13_4_lut_adj_1650.LUT_INIT = 16'h6996;
    SB_LUT4 i12_4_lut_adj_1651 (.I0(\data_out_frame[14] [6]), .I1(n44287), 
            .I2(n44525), .I3(n44240), .O(n30_adj_4786));
    defparam i12_4_lut_adj_1651.LUT_INIT = 16'h6996;
    SB_LUT4 i16_4_lut_adj_1652 (.I0(n31_adj_4785), .I1(n27885), .I2(n28_adj_4784), 
            .I3(\data_out_frame[14] [4]), .O(n34));
    defparam i16_4_lut_adj_1652.LUT_INIT = 16'h6996;
    SB_LUT4 i1_3_lut_4_lut_adj_1653 (.I0(n44105), .I1(n44620), .I2(n44611), 
            .I3(n27933), .O(n44562));
    defparam i1_3_lut_4_lut_adj_1653.LUT_INIT = 16'h6996;
    SB_LUT4 i11_4_lut_adj_1654 (.I0(n27809), .I1(n43968), .I2(n44248), 
            .I3(\data_out_frame[11] [5]), .O(n29));
    defparam i11_4_lut_adj_1654.LUT_INIT = 16'h6996;
    SB_LUT4 i2_4_lut_adj_1655 (.I0(n29), .I1(\data_out_frame[15] [7]), .I2(n34), 
            .I3(n30_adj_4786), .O(n7_adj_4787));
    defparam i2_4_lut_adj_1655.LUT_INIT = 16'h9669;
    SB_LUT4 i5_4_lut_adj_1656 (.I0(\data_out_frame[16] [4]), .I1(\data_out_frame[16] [1]), 
            .I2(\data_out_frame[16] [7]), .I3(n27481), .O(n12_adj_4788));
    defparam i5_4_lut_adj_1656.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1657 (.I0(n7_adj_4787), .I1(n27771), .I2(\data_out_frame[15] [0]), 
            .I3(n44084), .O(n45747));
    defparam i4_4_lut_adj_1657.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1658 (.I0(n45747), .I1(n12_adj_4788), .I2(n44202), 
            .I3(n28400), .O(n45357));
    defparam i6_4_lut_adj_1658.LUT_INIT = 16'h9669;
    SB_LUT4 i12_4_lut_adj_1659 (.I0(\data_out_frame[17] [1]), .I1(\data_out_frame[18] [3]), 
            .I2(n45357), .I3(\data_out_frame[19] [4]), .O(n28_adj_4789));
    defparam i12_4_lut_adj_1659.LUT_INIT = 16'h9669;
    SB_LUT4 i10_4_lut_adj_1660 (.I0(n44476), .I1(\data_out_frame[17] [6]), 
            .I2(\data_out_frame[17] [3]), .I3(\data_out_frame[18] [7]), 
            .O(n26_adj_4790));
    defparam i10_4_lut_adj_1660.LUT_INIT = 16'h6996;
    SB_LUT4 i11_4_lut_adj_1661 (.I0(n44501), .I1(n43964), .I2(n44438), 
            .I3(\data_out_frame[19] [6]), .O(n27_adj_4791));
    defparam i11_4_lut_adj_1661.LUT_INIT = 16'h6996;
    SB_LUT4 i9_4_lut_adj_1662 (.I0(\data_out_frame[17] [4]), .I1(n44125), 
            .I2(\data_out_frame[18] [5]), .I3(\data_out_frame[18] [2]), 
            .O(n25_adj_4792));
    defparam i9_4_lut_adj_1662.LUT_INIT = 16'h6996;
    SB_LUT4 i1_3_lut_4_lut_adj_1663 (.I0(n44105), .I1(n44620), .I2(\data_in_frame[10] [7]), 
            .I3(\data_in_frame[11] [1]), .O(n43877));
    defparam i1_3_lut_4_lut_adj_1663.LUT_INIT = 16'h9669;
    SB_LUT4 i2_2_lut_4_lut_adj_1664 (.I0(\data_out_frame[4] [6]), .I1(\data_out_frame[5] [0]), 
            .I2(n4_c), .I3(\data_out_frame[5] [4]), .O(n10_adj_4613));   // verilog/coms.v(72[16:27])
    defparam i2_2_lut_4_lut_adj_1664.LUT_INIT = 16'h6996;
    SB_LUT4 i1_3_lut_4_lut_adj_1665 (.I0(n43877), .I1(n44012), .I2(n27520), 
            .I3(Kp_23__N_1561), .O(n40653));   // verilog/coms.v(72[16:27])
    defparam i1_3_lut_4_lut_adj_1665.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1666 (.I0(byte_transmit_counter[6]), .I1(byte_transmit_counter[7]), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_4793));   // verilog/coms.v(215[11:56])
    defparam i1_2_lut_adj_1666.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_1667 (.I0(byte_transmit_counter[4]), .I1(byte_transmit_counter[0]), 
            .I2(byte_transmit_counter[2]), .I3(byte_transmit_counter[1]), 
            .O(n4_adj_4794));
    defparam i1_4_lut_adj_1667.LUT_INIT = 16'ha8a0;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_35859 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [6]), .I2(\data_out_frame[27] [6]), 
            .I3(byte_transmit_counter[1]), .O(n51492));
    defparam byte_transmit_counter_0__bdd_4_lut_35859.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_4_lut_adj_1668 (.I0(n40676), .I1(n44556), .I2(n41814), 
            .I3(n47503), .O(n45300));
    defparam i1_4_lut_adj_1668.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1669 (.I0(n43877), .I1(n44012), .I2(n41606), 
            .I3(GND_net), .O(n41793));   // verilog/coms.v(72[16:27])
    defparam i1_2_lut_3_lut_adj_1669.LUT_INIT = 16'h9696;
    SB_LUT4 i15357_3_lut_4_lut (.I0(n8_adj_4729), .I1(n43820), .I2(rx_data[7]), 
            .I3(\data_in_frame[16] [7]), .O(n29305));
    defparam i15357_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15_4_lut_adj_1670 (.I0(n25_adj_4792), .I1(n27_adj_4791), .I2(n26_adj_4790), 
            .I3(n28_adj_4789), .O(n41609));
    defparam i15_4_lut_adj_1670.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1671 (.I0(\data_out_frame[18] [5]), .I1(\data_out_frame[19] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n44278));
    defparam i1_2_lut_adj_1671.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1672 (.I0(\data_out_frame[19] [3]), .I1(n41609), 
            .I2(GND_net), .I3(GND_net), .O(n44190));
    defparam i1_2_lut_adj_1672.LUT_INIT = 16'h6666;
    SB_LUT4 i35564_4_lut (.I0(byte_transmit_counter[3]), .I1(byte_transmit_counter[5]), 
            .I2(n4_adj_4794), .I3(n4_adj_4793), .O(tx_transmit_N_3677));
    defparam i35564_4_lut.LUT_INIT = 16'h0013;
    SB_LUT4 i1_2_lut_adj_1673 (.I0(n43716), .I1(n43817), .I2(GND_net), 
            .I3(GND_net), .O(n63_adj_4742));
    defparam i1_2_lut_adj_1673.LUT_INIT = 16'heeee;
    SB_LUT4 i4_4_lut_adj_1674 (.I0(n44190), .I1(n28186), .I2(n41653), 
            .I3(n44278), .O(n10_adj_4765));
    defparam i4_4_lut_adj_1674.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1675 (.I0(n41472), .I1(n41816), .I2(GND_net), 
            .I3(GND_net), .O(n41807));
    defparam i1_2_lut_adj_1675.LUT_INIT = 16'h9999;
    SB_LUT4 i15358_3_lut_4_lut (.I0(n8_adj_4729), .I1(n43820), .I2(rx_data[6]), 
            .I3(\data_in_frame[16] [6]), .O(n29306));
    defparam i15358_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15359_3_lut_4_lut (.I0(n8_adj_4729), .I1(n43820), .I2(rx_data[5]), 
            .I3(\data_in_frame[16] [5]), .O(n29307));
    defparam i15359_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15403_3_lut_4_lut (.I0(n8_adj_4655), .I1(n43841), .I2(rx_data[4]), 
            .I3(\data_in_frame[11] [4]), .O(n29351));
    defparam i15403_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15360_3_lut_4_lut (.I0(n8_adj_4729), .I1(n43820), .I2(rx_data[4]), 
            .I3(\data_in_frame[16] [4]), .O(n29308));
    defparam i15360_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_4_lut_adj_1676 (.I0(n26774), .I1(n44038), .I2(\data_in_frame[16] [2]), 
            .I3(\data_in_frame[14] [2]), .O(n40631));
    defparam i2_3_lut_4_lut_adj_1676.LUT_INIT = 16'h6996;
    SB_LUT4 i29293_3_lut (.I0(n44724), .I1(n43719), .I2(\FRAME_MATCHER.state [3]), 
            .I3(GND_net), .O(n44813));
    defparam i29293_3_lut.LUT_INIT = 16'hecec;
    SB_LUT4 i1_2_lut_4_lut_adj_1677 (.I0(\data_out_frame[8] [3]), .I1(\data_out_frame[8] [1]), 
            .I2(\data_out_frame[7] [7]), .I3(\data_out_frame[5] [5]), .O(n43908));   // verilog/coms.v(72[16:62])
    defparam i1_2_lut_4_lut_adj_1677.LUT_INIT = 16'h6996;
    SB_LUT4 mux_1428_i1_4_lut (.I0(tx_transmit_N_3677), .I1(\FRAME_MATCHER.state [3]), 
            .I2(n35382), .I3(n6_adj_4767), .O(n5403[0]));   // verilog/coms.v(146[4] 302[11])
    defparam mux_1428_i1_4_lut.LUT_INIT = 16'h0cac;
    SB_LUT4 i15361_3_lut_4_lut (.I0(n8_adj_4729), .I1(n43820), .I2(rx_data[3]), 
            .I3(\data_in_frame[16] [3]), .O(n29309));
    defparam i15361_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15362_3_lut_4_lut (.I0(n8_adj_4729), .I1(n43820), .I2(rx_data[2]), 
            .I3(\data_in_frame[16] [2]), .O(n29310));
    defparam i15362_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15363_3_lut_4_lut (.I0(n8_adj_4729), .I1(n43820), .I2(rx_data[1]), 
            .I3(\data_in_frame[16] [1]), .O(n29311));
    defparam i15363_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_adj_1678 (.I0(\data_out_frame[19] [2]), .I1(n41816), 
            .I2(\data_out_frame[22] [6]), .I3(GND_net), .O(n44519));
    defparam i2_3_lut_adj_1678.LUT_INIT = 16'h6969;
    SB_LUT4 n51492_bdd_4_lut (.I0(n51492), .I1(\data_out_frame[25] [6]), 
            .I2(\data_out_frame[24] [6]), .I3(byte_transmit_counter[1]), 
            .O(n51495));
    defparam n51492_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i15404_3_lut_4_lut (.I0(n8_adj_4655), .I1(n43841), .I2(rx_data[3]), 
            .I3(\data_in_frame[11] [3]), .O(n29352));
    defparam i15404_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15364_3_lut_4_lut (.I0(n8_adj_4729), .I1(n43820), .I2(rx_data[0]), 
            .I3(\data_in_frame[16] [0]), .O(n29312));
    defparam i15364_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i3_3_lut_4_lut_adj_1679 (.I0(\data_in_frame[18] [7]), .I1(\data_in_frame[18] [6]), 
            .I2(n44459), .I3(\data_in_frame[18] [4]), .O(n8_adj_4669));   // verilog/coms.v(79[16:27])
    defparam i3_3_lut_4_lut_adj_1679.LUT_INIT = 16'h6996;
    SB_LUT4 i15349_3_lut_4_lut (.I0(n8_adj_4645), .I1(n43820), .I2(rx_data[7]), 
            .I3(\data_in_frame[17] [7]), .O(n29297));
    defparam i15349_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i6_4_lut_adj_1680 (.I0(n44257), .I1(n41609), .I2(n44541), 
            .I3(n44468), .O(n16_adj_4795));
    defparam i6_4_lut_adj_1680.LUT_INIT = 16'h9669;
    SB_LUT4 i15350_3_lut_4_lut (.I0(n8_adj_4645), .I1(n43820), .I2(rx_data[6]), 
            .I3(\data_in_frame[17] [6]), .O(n29298));
    defparam i15350_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i7_4_lut_adj_1681 (.I0(n41642), .I1(n44519), .I2(n44571), 
            .I3(n44268), .O(n17_adj_4796));
    defparam i7_4_lut_adj_1681.LUT_INIT = 16'h9669;
    SB_LUT4 i9_4_lut_adj_1682 (.I0(n17_adj_4796), .I1(\data_out_frame[21] [0]), 
            .I2(n16_adj_4795), .I3(\data_out_frame[19] [3]), .O(n41596));
    defparam i9_4_lut_adj_1682.LUT_INIT = 16'h6996;
    SB_LUT4 n51210_bdd_4_lut (.I0(n51210), .I1(n48144), .I2(n48143), .I3(byte_transmit_counter[2]), 
            .O(n51213));
    defparam n51210_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3_4_lut_adj_1683 (.I0(\data_out_frame[25] [3]), .I1(n41682), 
            .I2(\data_out_frame[25] [2]), .I3(n41596), .O(n46011));
    defparam i3_4_lut_adj_1683.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1684 (.I0(\data_out_frame[4] [1]), .I1(\data_out_frame[4] [0]), 
            .I2(\data_out_frame[6] [2]), .I3(\data_out_frame[6] [6]), .O(n44322));   // verilog/coms.v(75[16:43])
    defparam i1_2_lut_4_lut_adj_1684.LUT_INIT = 16'h6996;
    SB_LUT4 i2_2_lut_3_lut_adj_1685 (.I0(n46118), .I1(\data_in_frame[16] [1]), 
            .I2(\data_in_frame[13] [5]), .I3(GND_net), .O(n10_adj_4604));
    defparam i2_2_lut_3_lut_adj_1685.LUT_INIT = 16'h6969;
    SB_LUT4 i15399_3_lut_4_lut (.I0(n8_adj_4681), .I1(n43841), .I2(rx_data[0]), 
            .I3(\data_in_frame[12] [0]), .O(n29347));
    defparam i15399_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15351_3_lut_4_lut (.I0(n8_adj_4645), .I1(n43820), .I2(rx_data[5]), 
            .I3(\data_in_frame[17] [5]), .O(n29299));
    defparam i15351_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15352_3_lut_4_lut (.I0(n8_adj_4645), .I1(n43820), .I2(rx_data[4]), 
            .I3(\data_in_frame[17] [4]), .O(n29300));
    defparam i15352_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i3_3_lut_adj_1686 (.I0(n28049), .I1(\data_out_frame[11] [3]), 
            .I2(\data_out_frame[9] [1]), .I3(GND_net), .O(n8_adj_4797));
    defparam i3_3_lut_adj_1686.LUT_INIT = 16'h9696;
    SB_LUT4 i15353_3_lut_4_lut (.I0(n8_adj_4645), .I1(n43820), .I2(rx_data[3]), 
            .I3(\data_in_frame[17] [3]), .O(n29301));
    defparam i15353_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_4_lut_adj_1687 (.I0(\data_out_frame[13] [5]), .I1(n27745), 
            .I2(n8_adj_4797), .I3(n43917), .O(n44583));
    defparam i1_4_lut_adj_1687.LUT_INIT = 16'h6996;
    SB_LUT4 i3_3_lut_adj_1688 (.I0(n44583), .I1(\data_out_frame[11] [4]), 
            .I2(n25208), .I3(GND_net), .O(n40821));
    defparam i3_3_lut_adj_1688.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1689 (.I0(\data_out_frame[10] [4]), .I1(\data_out_frame[6] [0]), 
            .I2(\data_out_frame[6] [1]), .I3(\data_out_frame[6] [2]), .O(n43874));   // verilog/coms.v(73[16:27])
    defparam i2_3_lut_4_lut_adj_1689.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1690 (.I0(\data_out_frame[19] [2]), .I1(n44302), 
            .I2(n44262), .I3(GND_net), .O(n44263));
    defparam i1_2_lut_3_lut_adj_1690.LUT_INIT = 16'h9696;
    SB_LUT4 i15354_3_lut_4_lut (.I0(n8_adj_4645), .I1(n43820), .I2(rx_data[2]), 
            .I3(\data_in_frame[17] [2]), .O(n29302));
    defparam i15354_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i4_4_lut_adj_1691 (.I0(n44254), .I1(\data_out_frame[16] [2]), 
            .I2(\data_out_frame[18] [3]), .I3(n44409), .O(n10_adj_4798));
    defparam i4_4_lut_adj_1691.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_1692 (.I0(n25208), .I1(n10_adj_4798), .I2(\data_out_frame[16] [1]), 
            .I3(GND_net), .O(n41801));
    defparam i5_3_lut_adj_1692.LUT_INIT = 16'h9696;
    SB_LUT4 i15355_3_lut_4_lut (.I0(n8_adj_4645), .I1(n43820), .I2(rx_data[1]), 
            .I3(\data_in_frame[17] [1]), .O(n29303));
    defparam i15355_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15356_3_lut_4_lut (.I0(n8_adj_4645), .I1(n43820), .I2(rx_data[0]), 
            .I3(\data_in_frame[17] [0]), .O(n29304));
    defparam i15356_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1693 (.I0(\data_out_frame[20] [5]), .I1(n41801), 
            .I2(GND_net), .I3(GND_net), .O(n44268));
    defparam i1_2_lut_adj_1693.LUT_INIT = 16'h9999;
    SB_LUT4 i5_4_lut_adj_1694 (.I0(\data_out_frame[23] [1]), .I1(n44268), 
            .I2(n41611), .I3(\data_out_frame[22] [7]), .O(n13_adj_4799));
    defparam i5_4_lut_adj_1694.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1695 (.I0(n13_adj_4799), .I1(n11_adj_4725), .I2(n46020), 
            .I3(n27834), .O(n41682));
    defparam i7_4_lut_adj_1695.LUT_INIT = 16'h9669;
    SB_LUT4 i15405_3_lut_4_lut (.I0(n8_adj_4655), .I1(n43841), .I2(rx_data[2]), 
            .I3(\data_in_frame[11] [2]), .O(n29353));
    defparam i15405_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15339_3_lut_4_lut (.I0(n8), .I1(n43820), .I2(rx_data[7]), 
            .I3(\data_in_frame[18] [7]), .O(n29287));
    defparam i15339_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1696 (.I0(n41682), .I1(n25338), .I2(GND_net), 
            .I3(GND_net), .O(n44444));
    defparam i1_2_lut_adj_1696.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1697 (.I0(\data_out_frame[25] [3]), .I1(\data_out_frame[25] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n44152));
    defparam i1_2_lut_adj_1697.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1698 (.I0(\data_out_frame[16] [5]), .I1(\data_out_frame[16] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n28400));
    defparam i1_2_lut_adj_1698.LUT_INIT = 16'h6666;
    SB_LUT4 i15341_3_lut_4_lut (.I0(n8), .I1(n43820), .I2(rx_data[6]), 
            .I3(\data_in_frame[18] [6]), .O(n29289));
    defparam i15341_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i342_2_lut (.I0(\data_out_frame[4] [5]), .I1(\data_out_frame[4] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n1130));   // verilog/coms.v(77[16:27])
    defparam i342_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1699 (.I0(n1130), .I1(n44015), .I2(\data_out_frame[9] [2]), 
            .I3(\data_out_frame[6] [6]), .O(n28049));
    defparam i3_4_lut_adj_1699.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1700 (.I0(\data_out_frame[7] [0]), .I1(n1168), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_4764));   // verilog/coms.v(86[17:70])
    defparam i1_2_lut_adj_1700.LUT_INIT = 16'h6666;
    SB_LUT4 i5_4_lut_adj_1701 (.I0(n44096), .I1(\data_out_frame[11] [6]), 
            .I2(\data_out_frame[14] [0]), .I3(\data_out_frame[5] [3]), .O(n12_adj_4800));
    defparam i5_4_lut_adj_1701.LUT_INIT = 16'h6996;
    SB_LUT4 i32538_3_lut (.I0(\data_out_frame[16] [4]), .I1(\data_out_frame[17] [4]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n48125));
    defparam i32538_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i32539_3_lut (.I0(\data_out_frame[18] [4]), .I1(\data_out_frame[19] [4]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n48126));
    defparam i32539_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_35854 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [5]), .I2(\data_out_frame[27] [5]), 
            .I3(byte_transmit_counter[1]), .O(n51486));
    defparam byte_transmit_counter_0__bdd_4_lut_35854.LUT_INIT = 16'he4aa;
    SB_LUT4 n51486_bdd_4_lut (.I0(n51486), .I1(\data_out_frame[25] [5]), 
            .I2(\data_out_frame[24] [5]), .I3(byte_transmit_counter[1]), 
            .O(n51489));
    defparam n51486_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i15406_3_lut_4_lut (.I0(n8_adj_4655), .I1(n43841), .I2(rx_data[1]), 
            .I3(\data_in_frame[11] [1]), .O(n29354));
    defparam i15406_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i6_4_lut_adj_1702 (.I0(n44137), .I1(n12_adj_4800), .I2(\data_out_frame[13] [7]), 
            .I3(n27612), .O(n44553));
    defparam i6_4_lut_adj_1702.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1703 (.I0(\data_out_frame[9] [3]), .I1(n4_adj_4764), 
            .I2(n4_c), .I3(n28049), .O(n25208));
    defparam i3_4_lut_adj_1703.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1704 (.I0(\data_out_frame[19] [1]), .I1(\data_out_frame[21] [3]), 
            .I2(n44226), .I3(GND_net), .O(n6_adj_4601));
    defparam i1_2_lut_3_lut_adj_1704.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1705 (.I0(\data_out_frame[16] [3]), .I1(\data_out_frame[16] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n27481));   // verilog/coms.v(86[17:28])
    defparam i1_2_lut_adj_1705.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_4_lut_adj_1706 (.I0(\data_in_frame[8] [7]), .I1(\data_in_frame[9] [1]), 
            .I2(n44072), .I3(n27817), .O(Kp_23__N_1465));   // verilog/coms.v(73[16:41])
    defparam i2_3_lut_4_lut_adj_1706.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1707 (.I0(\data_out_frame[21] [0]), .I1(\data_out_frame[16] [5]), 
            .I2(\data_out_frame[16] [6]), .I3(GND_net), .O(n44498));
    defparam i1_2_lut_3_lut_adj_1707.LUT_INIT = 16'h9696;
    uart_tx tx (.\r_Bit_Index[0] (\r_Bit_Index[0] ), .GND_net(GND_net), 
            .CLK_c(CLK_c), .tx_o(tx_o), .tx_data({tx_data}), .r_SM_Main({r_SM_Main}), 
            .VCC_net(VCC_net), .\r_SM_Main_2__N_3777[1] (\r_SM_Main_2__N_3777[1] ), 
            .n29230(n29230), .n51602(n51602), .n29066(n29066), .tx_active(tx_active), 
            .n28662(n28662), .n28970(n28970), .\r_SM_Main_2__N_3780[0] (r_SM_Main_2__N_3780[0]), 
            .n19541(n19541), .n4(n4), .tx_enable(tx_enable)) /* synthesis syn_module_defined=1 */ ;   // verilog/coms.v(108[10:70])
    uart_rx rx (.CLK_c(CLK_c), .\r_SM_Main_2__N_3706[2] (\r_SM_Main_2__N_3706[2] ), 
            .GND_net(GND_net), .n4(n4_adj_6), .r_SM_Main({r_SM_Main_adj_13}), 
            .r_Rx_Data(r_Rx_Data), .RX_N_10(RX_N_10), .VCC_net(VCC_net), 
            .\r_Bit_Index[0] (\r_Bit_Index[0]_adj_10 ), .n4_adj_4(n4_adj_11), 
            .n4_adj_5(n4_adj_12), .n34695(n34695), .n29233(n29233), .n43326(n43326), 
            .rx_data_ready(rx_data_ready), .n28666(n28666), .n28972(n28972), 
            .n28562(n28562), .n29524(n29524), .rx_data({rx_data}), .n29516(n29516), 
            .n29510(n29510), .n29508(n29508), .n29502(n29502), .n29467(n29467), 
            .n29404(n29404), .n43724(n43724), .n29237(n29237), .n27131(n27131), 
            .n27126(n27126)) /* synthesis syn_module_defined=1 */ ;   // verilog/coms.v(94[10:44])
    
endmodule
//
// Verilog Description of module uart_tx
//

module uart_tx (\r_Bit_Index[0] , GND_net, CLK_c, tx_o, tx_data, r_SM_Main, 
            VCC_net, \r_SM_Main_2__N_3777[1] , n29230, n51602, n29066, 
            tx_active, n28662, n28970, \r_SM_Main_2__N_3780[0] , n19541, 
            n4, tx_enable) /* synthesis syn_module_defined=1 */ ;
    output \r_Bit_Index[0] ;
    input GND_net;
    input CLK_c;
    output tx_o;
    input [7:0]tx_data;
    output [2:0]r_SM_Main;
    input VCC_net;
    output \r_SM_Main_2__N_3777[1] ;
    input n29230;
    input n51602;
    input n29066;
    output tx_active;
    output n28662;
    output n28970;
    input \r_SM_Main_2__N_3780[0] ;
    output n19541;
    output n4;
    output tx_enable;
    
    wire CLK_c /* synthesis SET_AS_NETWORK=CLK_c, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(3[9:12])
    wire [2:0]r_Bit_Index;   // verilog/uart_tx.v(33[16:27])
    wire [2:0]n307;
    wire [7:0]r_Tx_Data;   // verilog/uart_tx.v(34[16:25])
    
    wire n48059, n48060, n48066, n48065;
    wire [8:0]n41;
    
    wire n1;
    wire [8:0]r_Clock_Count;   // verilog/uart_tx.v(32[16:29])
    
    wire n28870, n3, n26628, n21834, n39439, n39438, n39437, n39436, 
        n39435, n39434, n39433, n39432, n45936, n10, n3_adj_4589, 
        n35159, n21833, o_Tx_Serial_N_3808, n51222;
    
    SB_LUT4 i2438_3_lut (.I0(r_Bit_Index[2]), .I1(r_Bit_Index[1]), .I2(\r_Bit_Index[0] ), 
            .I3(GND_net), .O(n307[2]));   // verilog/uart_tx.v(98[36:51])
    defparam i2438_3_lut.LUT_INIT = 16'h6a6a;
    SB_LUT4 i32472_3_lut (.I0(r_Tx_Data[0]), .I1(r_Tx_Data[1]), .I2(\r_Bit_Index[0] ), 
            .I3(GND_net), .O(n48059));
    defparam i32472_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i32473_3_lut (.I0(r_Tx_Data[2]), .I1(r_Tx_Data[3]), .I2(\r_Bit_Index[0] ), 
            .I3(GND_net), .O(n48060));
    defparam i32473_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i32479_3_lut (.I0(r_Tx_Data[6]), .I1(r_Tx_Data[7]), .I2(\r_Bit_Index[0] ), 
            .I3(GND_net), .O(n48066));
    defparam i32479_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i32478_3_lut (.I0(r_Tx_Data[4]), .I1(r_Tx_Data[5]), .I2(\r_Bit_Index[0] ), 
            .I3(GND_net), .O(n48065));
    defparam i32478_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFESR r_Clock_Count_2256__i1 (.Q(r_Clock_Count[1]), .C(CLK_c), .E(n1), 
            .D(n41[1]), .R(n28870));   // verilog/uart_tx.v(118[34:51])
    SB_DFFESR r_Clock_Count_2256__i2 (.Q(r_Clock_Count[2]), .C(CLK_c), .E(n1), 
            .D(n41[2]), .R(n28870));   // verilog/uart_tx.v(118[34:51])
    SB_DFFESR r_Clock_Count_2256__i3 (.Q(r_Clock_Count[3]), .C(CLK_c), .E(n1), 
            .D(n41[3]), .R(n28870));   // verilog/uart_tx.v(118[34:51])
    SB_DFFESR r_Clock_Count_2256__i4 (.Q(r_Clock_Count[4]), .C(CLK_c), .E(n1), 
            .D(n41[4]), .R(n28870));   // verilog/uart_tx.v(118[34:51])
    SB_DFFESR r_Clock_Count_2256__i5 (.Q(r_Clock_Count[5]), .C(CLK_c), .E(n1), 
            .D(n41[5]), .R(n28870));   // verilog/uart_tx.v(118[34:51])
    SB_DFFESR r_Clock_Count_2256__i6 (.Q(r_Clock_Count[6]), .C(CLK_c), .E(n1), 
            .D(n41[6]), .R(n28870));   // verilog/uart_tx.v(118[34:51])
    SB_DFFESR r_Clock_Count_2256__i7 (.Q(r_Clock_Count[7]), .C(CLK_c), .E(n1), 
            .D(n41[7]), .R(n28870));   // verilog/uart_tx.v(118[34:51])
    SB_DFFESR r_Clock_Count_2256__i8 (.Q(r_Clock_Count[8]), .C(CLK_c), .E(n1), 
            .D(n41[8]), .R(n28870));   // verilog/uart_tx.v(118[34:51])
    SB_DFFE o_Tx_Serial_45 (.Q(tx_o), .C(CLK_c), .E(n1), .D(n3));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i0 (.Q(r_Tx_Data[0]), .C(CLK_c), .E(n26628), .D(tx_data[0]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFSR r_SM_Main_i0 (.Q(r_SM_Main[0]), .C(CLK_c), .D(n21834), .R(r_SM_Main[2]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_LUT4 r_Clock_Count_2256_add_4_10_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[8]), .I3(n39439), .O(n41[8])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2256_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 r_Clock_Count_2256_add_4_9_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[7]), .I3(n39438), .O(n41[7])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2256_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2256_add_4_9 (.CI(n39438), .I0(GND_net), .I1(r_Clock_Count[7]), 
            .CO(n39439));
    SB_LUT4 r_Clock_Count_2256_add_4_8_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[6]), .I3(n39437), .O(n41[6])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2256_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2256_add_4_8 (.CI(n39437), .I0(GND_net), .I1(r_Clock_Count[6]), 
            .CO(n39438));
    SB_LUT4 r_Clock_Count_2256_add_4_7_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[5]), .I3(n39436), .O(n41[5])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2256_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2256_add_4_7 (.CI(n39436), .I0(GND_net), .I1(r_Clock_Count[5]), 
            .CO(n39437));
    SB_LUT4 r_Clock_Count_2256_add_4_6_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[4]), .I3(n39435), .O(n41[4])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2256_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2256_add_4_6 (.CI(n39435), .I0(GND_net), .I1(r_Clock_Count[4]), 
            .CO(n39436));
    SB_LUT4 r_Clock_Count_2256_add_4_5_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[3]), .I3(n39434), .O(n41[3])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2256_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2256_add_4_5 (.CI(n39434), .I0(GND_net), .I1(r_Clock_Count[3]), 
            .CO(n39435));
    SB_LUT4 r_Clock_Count_2256_add_4_4_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[2]), .I3(n39433), .O(n41[2])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2256_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2256_add_4_4 (.CI(n39433), .I0(GND_net), .I1(r_Clock_Count[2]), 
            .CO(n39434));
    SB_LUT4 i2431_2_lut (.I0(r_Bit_Index[1]), .I1(\r_Bit_Index[0] ), .I2(GND_net), 
            .I3(GND_net), .O(n307[1]));   // verilog/uart_tx.v(98[36:51])
    defparam i2431_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 r_Clock_Count_2256_add_4_3_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[1]), .I3(n39432), .O(n41[1])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2256_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2256_add_4_3 (.CI(n39432), .I0(GND_net), .I1(r_Clock_Count[1]), 
            .CO(n39433));
    SB_LUT4 r_Clock_Count_2256_add_4_2_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[0]), .I3(VCC_net), .O(n41[0])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2256_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2256_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(r_Clock_Count[0]), 
            .CO(n39432));
    SB_DFFESR r_Clock_Count_2256__i0 (.Q(r_Clock_Count[0]), .C(CLK_c), .E(n1), 
            .D(n41[0]), .R(n28870));   // verilog/uart_tx.v(118[34:51])
    SB_LUT4 i3_4_lut (.I0(r_Clock_Count[0]), .I1(r_Clock_Count[3]), .I2(r_Clock_Count[1]), 
            .I3(r_Clock_Count[2]), .O(n45936));
    defparam i3_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i4_4_lut (.I0(r_Clock_Count[4]), .I1(r_Clock_Count[5]), .I2(n45936), 
            .I3(r_Clock_Count[8]), .O(n10));
    defparam i4_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i5_3_lut (.I0(r_Clock_Count[6]), .I1(n10), .I2(r_Clock_Count[7]), 
            .I3(GND_net), .O(\r_SM_Main_2__N_3777[1] ));
    defparam i5_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i34921_4_lut (.I0(r_SM_Main[2]), .I1(\r_SM_Main_2__N_3777[1] ), 
            .I2(r_SM_Main[1]), .I3(r_SM_Main[0]), .O(n28870));
    defparam i34921_4_lut.LUT_INIT = 16'h4445;
    SB_LUT4 i1_1_lut (.I0(r_SM_Main[2]), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n1));
    defparam i1_1_lut.LUT_INIT = 16'h5555;
    SB_DFF r_Bit_Index_i0 (.Q(\r_Bit_Index[0] ), .C(CLK_c), .D(n29230));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_SM_Main_i2 (.Q(r_SM_Main[2]), .C(CLK_c), .D(n51602));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Tx_Active_47 (.Q(tx_active), .C(CLK_c), .D(n29066));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFSR r_SM_Main_i1 (.Q(r_SM_Main[1]), .C(CLK_c), .D(n3_adj_4589), 
            .R(r_SM_Main[2]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i7 (.Q(r_Tx_Data[7]), .C(CLK_c), .E(n26628), .D(tx_data[7]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i6 (.Q(r_Tx_Data[6]), .C(CLK_c), .E(n26628), .D(tx_data[6]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i5 (.Q(r_Tx_Data[5]), .C(CLK_c), .E(n26628), .D(tx_data[5]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i4 (.Q(r_Tx_Data[4]), .C(CLK_c), .E(n26628), .D(tx_data[4]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i3 (.Q(r_Tx_Data[3]), .C(CLK_c), .E(n26628), .D(tx_data[3]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i2 (.Q(r_Tx_Data[2]), .C(CLK_c), .E(n26628), .D(tx_data[2]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i1 (.Q(r_Tx_Data[1]), .C(CLK_c), .E(n26628), .D(tx_data[1]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFESR r_Bit_Index_i1 (.Q(r_Bit_Index[1]), .C(CLK_c), .E(n28662), 
            .D(n307[1]), .R(n28970));   // verilog/uart_tx.v(40[10] 143[8])
    SB_LUT4 i5717_2_lut (.I0(\r_SM_Main_2__N_3780[0] ), .I1(r_SM_Main[0]), 
            .I2(GND_net), .I3(GND_net), .O(n19541));   // verilog/uart_tx.v(43[7] 142[14])
    defparam i5717_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i2_3_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), .I2(\r_Bit_Index[0] ), 
            .I3(GND_net), .O(n35159));
    defparam i2_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i8002_4_lut (.I0(\r_SM_Main_2__N_3780[0] ), .I1(n35159), .I2(r_SM_Main[1]), 
            .I3(\r_SM_Main_2__N_3777[1] ), .O(n21833));   // verilog/uart_tx.v(43[7] 142[14])
    defparam i8002_4_lut.LUT_INIT = 16'hca0a;
    SB_LUT4 i8003_3_lut (.I0(n21833), .I1(\r_SM_Main_2__N_3777[1] ), .I2(r_SM_Main[0]), 
            .I3(GND_net), .O(n21834));   // verilog/uart_tx.v(43[7] 142[14])
    defparam i8003_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 r_SM_Main_2__I_0_56_i3_3_lut (.I0(r_SM_Main[0]), .I1(o_Tx_Serial_N_3808), 
            .I2(r_SM_Main[1]), .I3(GND_net), .O(n3));   // verilog/uart_tx.v(43[7] 142[14])
    defparam r_SM_Main_2__I_0_56_i3_3_lut.LUT_INIT = 16'he5e5;
    SB_LUT4 i1_3_lut_4_lut_4_lut (.I0(\r_SM_Main_2__N_3777[1] ), .I1(r_SM_Main[0]), 
            .I2(r_SM_Main[1]), .I3(r_SM_Main[2]), .O(n4));
    defparam i1_3_lut_4_lut_4_lut.LUT_INIT = 16'h008f;
    SB_DFFESR r_Bit_Index_i2 (.Q(r_Bit_Index[2]), .C(CLK_c), .E(n28662), 
            .D(n307[2]), .R(n28970));   // verilog/uart_tx.v(40[10] 143[8])
    SB_LUT4 i1_3_lut_4_lut (.I0(r_SM_Main[2]), .I1(r_SM_Main[0]), .I2(r_SM_Main[1]), 
            .I3(\r_SM_Main_2__N_3777[1] ), .O(n28662));
    defparam i1_3_lut_4_lut.LUT_INIT = 16'h1101;
    SB_LUT4 i2_3_lut_4_lut (.I0(r_SM_Main[2]), .I1(r_SM_Main[0]), .I2(\r_SM_Main_2__N_3780[0] ), 
            .I3(r_SM_Main[1]), .O(n26628));
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h0010;
    SB_LUT4 i9984_2_lut_3_lut (.I0(\r_SM_Main_2__N_3777[1] ), .I1(r_SM_Main[0]), 
            .I2(r_SM_Main[1]), .I3(GND_net), .O(n3_adj_4589));
    defparam i9984_2_lut_3_lut.LUT_INIT = 16'h7878;
    SB_LUT4 i15022_3_lut (.I0(n28662), .I1(n35159), .I2(r_SM_Main[1]), 
            .I3(GND_net), .O(n28970));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i15022_3_lut.LUT_INIT = 16'h8a8a;
    SB_LUT4 r_Bit_Index_1__bdd_4_lut (.I0(r_Bit_Index[1]), .I1(n48065), 
            .I2(n48066), .I3(r_Bit_Index[2]), .O(n51222));
    defparam r_Bit_Index_1__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n51222_bdd_4_lut (.I0(n51222), .I1(n48060), .I2(n48059), .I3(r_Bit_Index[2]), 
            .O(o_Tx_Serial_N_3808));
    defparam n51222_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 o_Tx_Serial_I_0_1_lut (.I0(tx_o), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(tx_enable));   // verilog/uart_tx.v(38[24:36])
    defparam o_Tx_Serial_I_0_1_lut.LUT_INIT = 16'h5555;
    
endmodule
//
// Verilog Description of module uart_rx
//

module uart_rx (CLK_c, \r_SM_Main_2__N_3706[2] , GND_net, n4, r_SM_Main, 
            r_Rx_Data, RX_N_10, VCC_net, \r_Bit_Index[0] , n4_adj_4, 
            n4_adj_5, n34695, n29233, n43326, rx_data_ready, n28666, 
            n28972, n28562, n29524, rx_data, n29516, n29510, n29508, 
            n29502, n29467, n29404, n43724, n29237, n27131, n27126) /* synthesis syn_module_defined=1 */ ;
    input CLK_c;
    output \r_SM_Main_2__N_3706[2] ;
    input GND_net;
    output n4;
    output [2:0]r_SM_Main;
    output r_Rx_Data;
    input RX_N_10;
    input VCC_net;
    output \r_Bit_Index[0] ;
    output n4_adj_4;
    output n4_adj_5;
    output n34695;
    input n29233;
    input n43326;
    output rx_data_ready;
    output n28666;
    output n28972;
    output n28562;
    input n29524;
    output [7:0]rx_data;
    input n29516;
    input n29510;
    input n29508;
    input n29502;
    input n29467;
    input n29404;
    input n43724;
    input n29237;
    output n27131;
    output n27126;
    
    wire CLK_c /* synthesis SET_AS_NETWORK=CLK_c, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(3[9:12])
    wire [7:0]r_Clock_Count;   // verilog/uart_rx.v(32[17:30])
    
    wire n27023;
    wire [7:0]n37;
    
    wire n28612, n28879, n43790, n43725;
    wire [2:0]r_Bit_Index;   // verilog/uart_rx.v(33[17:28])
    
    wire n33, r_Rx_Data_R, n49361, n39431, n39430, n39429, n39428, 
        n39427, n31604, n39426, n39425;
    wire [2:0]n326;
    
    wire n35340, n43478, n35155, n31, n29, n6;
    
    SB_LUT4 i3_4_lut (.I0(r_Clock_Count[4]), .I1(r_Clock_Count[7]), .I2(r_Clock_Count[6]), 
            .I3(r_Clock_Count[5]), .O(n27023));   // verilog/uart_rx.v(68[17:52])
    defparam i3_4_lut.LUT_INIT = 16'hfffe;
    SB_DFFESR r_Clock_Count_2254__i1 (.Q(r_Clock_Count[1]), .C(CLK_c), .E(n28612), 
            .D(n37[1]), .R(n28879));   // verilog/uart_rx.v(120[34:51])
    SB_DFFESR r_Clock_Count_2254__i2 (.Q(r_Clock_Count[2]), .C(CLK_c), .E(n28612), 
            .D(n37[2]), .R(n28879));   // verilog/uart_rx.v(120[34:51])
    SB_DFFESR r_Clock_Count_2254__i3 (.Q(r_Clock_Count[3]), .C(CLK_c), .E(n28612), 
            .D(n37[3]), .R(n28879));   // verilog/uart_rx.v(120[34:51])
    SB_DFFESR r_Clock_Count_2254__i4 (.Q(r_Clock_Count[4]), .C(CLK_c), .E(n28612), 
            .D(n37[4]), .R(n28879));   // verilog/uart_rx.v(120[34:51])
    SB_DFFESR r_Clock_Count_2254__i5 (.Q(r_Clock_Count[5]), .C(CLK_c), .E(n28612), 
            .D(n37[5]), .R(n28879));   // verilog/uart_rx.v(120[34:51])
    SB_DFFESR r_Clock_Count_2254__i6 (.Q(r_Clock_Count[6]), .C(CLK_c), .E(n28612), 
            .D(n37[6]), .R(n28879));   // verilog/uart_rx.v(120[34:51])
    SB_DFFESR r_Clock_Count_2254__i7 (.Q(r_Clock_Count[7]), .C(CLK_c), .E(n28612), 
            .D(n37[7]), .R(n28879));   // verilog/uart_rx.v(120[34:51])
    SB_LUT4 i21223_3_lut (.I0(r_Clock_Count[3]), .I1(n27023), .I2(n43790), 
            .I3(GND_net), .O(\r_SM_Main_2__N_3706[2] ));
    defparam i21223_3_lut.LUT_INIT = 16'hecec;
    SB_LUT4 i2_3_lut (.I0(n27023), .I1(r_Clock_Count[3]), .I2(n43790), 
            .I3(GND_net), .O(n43725));
    defparam i2_3_lut.LUT_INIT = 16'h1010;
    SB_LUT4 equal_347_i4_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(GND_net), .I3(GND_net), .O(n4));   // verilog/uart_rx.v(97[17:39])
    defparam equal_347_i4_2_lut.LUT_INIT = 16'heeee;
    SB_DFFSR r_SM_Main_i0 (.Q(r_SM_Main[0]), .C(CLK_c), .D(n33), .R(r_SM_Main[2]));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Data_50 (.Q(r_Rx_Data), .C(CLK_c), .D(r_Rx_Data_R));   // verilog/uart_rx.v(41[10] 45[8])
    SB_DFF r_Rx_Data_R_49 (.Q(r_Rx_Data_R), .C(CLK_c), .D(RX_N_10));   // verilog/uart_rx.v(41[10] 45[8])
    SB_LUT4 i34399_3_lut (.I0(r_Rx_Data), .I1(r_SM_Main[0]), .I2(n43725), 
            .I3(GND_net), .O(n49361));
    defparam i34399_3_lut.LUT_INIT = 16'h7373;
    SB_LUT4 i1_4_lut (.I0(r_SM_Main[2]), .I1(n49361), .I2(\r_SM_Main_2__N_3706[2] ), 
            .I3(r_SM_Main[1]), .O(n28879));
    defparam i1_4_lut.LUT_INIT = 16'h5044;
    SB_LUT4 r_Clock_Count_2254_add_4_9_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[7]), .I3(n39431), .O(n37[7])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2254_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 r_Clock_Count_2254_add_4_8_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[6]), .I3(n39430), .O(n37[6])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2254_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2254_add_4_8 (.CI(n39430), .I0(GND_net), .I1(r_Clock_Count[6]), 
            .CO(n39431));
    SB_LUT4 r_Clock_Count_2254_add_4_7_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[5]), .I3(n39429), .O(n37[5])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2254_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2254_add_4_7 (.CI(n39429), .I0(GND_net), .I1(r_Clock_Count[5]), 
            .CO(n39430));
    SB_LUT4 r_Clock_Count_2254_add_4_6_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[4]), .I3(n39428), .O(n37[4])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2254_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2254_add_4_6 (.CI(n39428), .I0(GND_net), .I1(r_Clock_Count[4]), 
            .CO(n39429));
    SB_LUT4 r_Clock_Count_2254_add_4_5_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[3]), .I3(n39427), .O(n37[3])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2254_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2254_add_4_5 (.CI(n39427), .I0(GND_net), .I1(r_Clock_Count[3]), 
            .CO(n39428));
    SB_LUT4 i35570_4_lut (.I0(r_Rx_Data), .I1(r_SM_Main[2]), .I2(r_SM_Main[1]), 
            .I3(n31604), .O(n28612));
    defparam i35570_4_lut.LUT_INIT = 16'h3133;
    SB_LUT4 r_Clock_Count_2254_add_4_4_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[2]), .I3(n39426), .O(n37[2])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2254_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2254_add_4_4 (.CI(n39426), .I0(GND_net), .I1(r_Clock_Count[2]), 
            .CO(n39427));
    SB_LUT4 r_Clock_Count_2254_add_4_3_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[1]), .I3(n39425), .O(n37[1])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2254_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2254_add_4_3 (.CI(n39425), .I0(GND_net), .I1(r_Clock_Count[1]), 
            .CO(n39426));
    SB_LUT4 r_Clock_Count_2254_add_4_2_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[0]), .I3(VCC_net), .O(n37[0])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2254_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2254_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(r_Clock_Count[0]), 
            .CO(n39425));
    SB_LUT4 i2416_3_lut (.I0(r_Bit_Index[2]), .I1(r_Bit_Index[1]), .I2(\r_Bit_Index[0] ), 
            .I3(GND_net), .O(n326[2]));   // verilog/uart_rx.v(102[36:51])
    defparam i2416_3_lut.LUT_INIT = 16'h6a6a;
    SB_LUT4 i21395_2_lut (.I0(\r_SM_Main_2__N_3706[2] ), .I1(r_SM_Main[0]), 
            .I2(GND_net), .I3(GND_net), .O(n35340));
    defparam i21395_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i13_4_lut (.I0(n31604), .I1(n35340), .I2(r_SM_Main[1]), .I3(r_Rx_Data), 
            .O(n43478));   // verilog/uart_rx.v(30[17:26])
    defparam i13_4_lut.LUT_INIT = 16'h303a;
    SB_LUT4 i2409_2_lut (.I0(r_Bit_Index[1]), .I1(\r_Bit_Index[0] ), .I2(GND_net), 
            .I3(GND_net), .O(n326[1]));   // verilog/uart_rx.v(102[36:51])
    defparam i2409_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 equal_345_i4_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_4));   // verilog/uart_rx.v(97[17:39])
    defparam equal_345_i4_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 i1_2_lut (.I0(r_SM_Main[0]), .I1(n43725), .I2(GND_net), .I3(GND_net), 
            .O(n31604));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i1_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 equal_344_i4_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_5));   // verilog/uart_rx.v(97[17:39])
    defparam equal_344_i4_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 i20765_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), .I2(GND_net), 
            .I3(GND_net), .O(n34695));
    defparam i20765_2_lut.LUT_INIT = 16'h8888;
    SB_DFF r_Bit_Index_i0 (.Q(\r_Bit_Index[0] ), .C(CLK_c), .D(n29233));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_DV_52 (.Q(rx_data_ready), .C(CLK_c), .D(n43326));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFFESR r_Clock_Count_2254__i0 (.Q(r_Clock_Count[0]), .C(CLK_c), .E(n28612), 
            .D(n37[0]), .R(n28879));   // verilog/uart_rx.v(120[34:51])
    SB_DFFESR r_Bit_Index_i1 (.Q(r_Bit_Index[1]), .C(CLK_c), .E(n28666), 
            .D(n326[1]), .R(n28972));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFFSR r_SM_Main_i1 (.Q(r_SM_Main[1]), .C(CLK_c), .D(n43478), .R(r_SM_Main[2]));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFFESR r_Bit_Index_i2 (.Q(r_Bit_Index[2]), .C(CLK_c), .E(n28666), 
            .D(n326[2]), .R(n28972));   // verilog/uart_rx.v(49[10] 144[8])
    SB_LUT4 i1_3_lut_4_lut (.I0(\r_SM_Main_2__N_3706[2] ), .I1(r_SM_Main[0]), 
            .I2(r_SM_Main[2]), .I3(r_SM_Main[1]), .O(n28666));
    defparam i1_3_lut_4_lut.LUT_INIT = 16'h0203;
    SB_LUT4 i13_3_lut_4_lut (.I0(r_SM_Main[1]), .I1(r_SM_Main[2]), .I2(\r_SM_Main_2__N_3706[2] ), 
            .I3(r_SM_Main[0]), .O(n28562));
    defparam i13_3_lut_4_lut.LUT_INIT = 16'h2055;
    SB_DFF r_Rx_Byte_i7 (.Q(rx_data[7]), .C(CLK_c), .D(n29524));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i6 (.Q(rx_data[6]), .C(CLK_c), .D(n29516));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i5 (.Q(rx_data[5]), .C(CLK_c), .D(n29510));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i4 (.Q(rx_data[4]), .C(CLK_c), .D(n29508));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i3 (.Q(rx_data[3]), .C(CLK_c), .D(n29502));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i2 (.Q(rx_data[2]), .C(CLK_c), .D(n29467));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i1 (.Q(rx_data[1]), .C(CLK_c), .D(n29404));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_SM_Main_i2 (.Q(r_SM_Main[2]), .C(CLK_c), .D(n43724));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i0 (.Q(rx_data[0]), .C(CLK_c), .D(n29237));   // verilog/uart_rx.v(49[10] 144[8])
    SB_LUT4 i2_3_lut_adj_954 (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(\r_Bit_Index[0] ), .I3(GND_net), .O(n35155));
    defparam i2_3_lut_adj_954.LUT_INIT = 16'h8080;
    SB_LUT4 i33_3_lut (.I0(n35155), .I1(\r_SM_Main_2__N_3706[2] ), .I2(r_SM_Main[0]), 
            .I3(GND_net), .O(n31));   // verilog/uart_rx.v(30[17:26])
    defparam i33_3_lut.LUT_INIT = 16'hc7c7;
    SB_LUT4 i34_3_lut (.I0(r_Rx_Data), .I1(n43725), .I2(r_SM_Main[0]), 
            .I3(GND_net), .O(n29));   // verilog/uart_rx.v(30[17:26])
    defparam i34_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i32_3_lut (.I0(n29), .I1(n31), .I2(r_SM_Main[1]), .I3(GND_net), 
            .O(n33));   // verilog/uart_rx.v(30[17:26])
    defparam i32_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i2_3_lut_adj_955 (.I0(r_Clock_Count[0]), .I1(r_Clock_Count[1]), 
            .I2(r_Clock_Count[2]), .I3(GND_net), .O(n43790));
    defparam i2_3_lut_adj_955.LUT_INIT = 16'h8080;
    SB_LUT4 i2_2_lut (.I0(r_SM_Main[0]), .I1(r_SM_Main[2]), .I2(GND_net), 
            .I3(GND_net), .O(n6));
    defparam i2_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i15024_3_lut (.I0(n28666), .I1(n35155), .I2(r_SM_Main[1]), 
            .I3(GND_net), .O(n28972));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i15024_3_lut.LUT_INIT = 16'h8a8a;
    SB_LUT4 i1_2_lut_4_lut (.I0(n6), .I1(\r_SM_Main_2__N_3706[2] ), .I2(r_SM_Main[1]), 
            .I3(\r_Bit_Index[0] ), .O(n27131));
    defparam i1_2_lut_4_lut.LUT_INIT = 16'hffbf;
    SB_LUT4 i1_2_lut_4_lut_adj_956 (.I0(n6), .I1(\r_SM_Main_2__N_3706[2] ), 
            .I2(r_SM_Main[1]), .I3(\r_Bit_Index[0] ), .O(n27126));
    defparam i1_2_lut_4_lut_adj_956.LUT_INIT = 16'hbfff;
    
endmodule
//
// Verilog Description of module \quadrature_decoder(1,500000) 
//

module \quadrature_decoder(1,500000)  (n1891, b_prev, GND_net, a_new, 
            direction_N_4071, ENCODER1_B_N_keep, ENCODER1_A_N_keep, encoder1_position, 
            VCC_net, n29245, n1896) /* synthesis lattice_noprune=1 */ ;
    input n1891;
    output b_prev;
    input GND_net;
    output [1:0]a_new;
    output direction_N_4071;
    input ENCODER1_B_N_keep;
    input ENCODER1_A_N_keep;
    output [31:0]encoder1_position;
    input VCC_net;
    input n29245;
    output n1896;
    
    
    wire n29165, a_prev;
    wire [1:0]b_new;   // vhdl/quadrature_decoder.vhd(41[9:14])
    
    wire direction_N_4074, debounce_cnt;
    wire [1:0]a_new_c;   // vhdl/quadrature_decoder.vhd(40[9:14])
    
    wire a_prev_N_4077;
    wire [31:0]n133;
    
    wire direction_N_4070, n39407, n39406, n39405, n39404, n39403, 
        n39402, n39401, n39400, n39399, n39398, n39397, n39396, 
        n39395, n39394, n39393, n39392, n39391, n39390, n39389, 
        n39388, n39387, n39386, n39385, n39384, n39383, n39382, 
        n39381, n39380, n39379, n39378, n39377, n29222;
    
    SB_DFF a_prev_51 (.Q(a_prev), .C(n1891), .D(n29165));   // vhdl/quadrature_decoder.vhd(52[3] 89[10])
    SB_LUT4 b_prev_I_0_65_2_lut (.I0(b_prev), .I1(b_new[1]), .I2(GND_net), 
            .I3(GND_net), .O(direction_N_4074));   // vhdl/quadrature_decoder.vhd(80[37:56])
    defparam b_prev_I_0_65_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 debounce_cnt_I_0_4_lut (.I0(debounce_cnt), .I1(a_prev), .I2(direction_N_4074), 
            .I3(a_new[1]), .O(direction_N_4071));   // vhdl/quadrature_decoder.vhd(79[10] 80[64])
    defparam debounce_cnt_I_0_4_lut.LUT_INIT = 16'ha2a8;
    SB_DFF b_new_i0 (.Q(b_new[0]), .C(n1891), .D(ENCODER1_B_N_keep));   // vhdl/quadrature_decoder.vhd(52[3] 89[10])
    SB_DFF a_new_i0 (.Q(a_new_c[0]), .C(n1891), .D(ENCODER1_A_N_keep));   // vhdl/quadrature_decoder.vhd(52[3] 89[10])
    SB_DFF debounce_cnt_50 (.Q(debounce_cnt), .C(n1891), .D(a_prev_N_4077));   // vhdl/quadrature_decoder.vhd(52[3] 89[10])
    SB_DFFE position_2248__i31 (.Q(encoder1_position[31]), .C(n1891), .E(direction_N_4071), 
            .D(n133[31]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2248__i30 (.Q(encoder1_position[30]), .C(n1891), .E(direction_N_4071), 
            .D(n133[30]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2248__i29 (.Q(encoder1_position[29]), .C(n1891), .E(direction_N_4071), 
            .D(n133[29]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2248__i28 (.Q(encoder1_position[28]), .C(n1891), .E(direction_N_4071), 
            .D(n133[28]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2248__i27 (.Q(encoder1_position[27]), .C(n1891), .E(direction_N_4071), 
            .D(n133[27]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2248__i26 (.Q(encoder1_position[26]), .C(n1891), .E(direction_N_4071), 
            .D(n133[26]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2248__i25 (.Q(encoder1_position[25]), .C(n1891), .E(direction_N_4071), 
            .D(n133[25]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2248__i24 (.Q(encoder1_position[24]), .C(n1891), .E(direction_N_4071), 
            .D(n133[24]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2248__i23 (.Q(encoder1_position[23]), .C(n1891), .E(direction_N_4071), 
            .D(n133[23]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2248__i22 (.Q(encoder1_position[22]), .C(n1891), .E(direction_N_4071), 
            .D(n133[22]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2248__i21 (.Q(encoder1_position[21]), .C(n1891), .E(direction_N_4071), 
            .D(n133[21]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2248__i20 (.Q(encoder1_position[20]), .C(n1891), .E(direction_N_4071), 
            .D(n133[20]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2248__i19 (.Q(encoder1_position[19]), .C(n1891), .E(direction_N_4071), 
            .D(n133[19]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2248__i18 (.Q(encoder1_position[18]), .C(n1891), .E(direction_N_4071), 
            .D(n133[18]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2248__i17 (.Q(encoder1_position[17]), .C(n1891), .E(direction_N_4071), 
            .D(n133[17]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2248__i16 (.Q(encoder1_position[16]), .C(n1891), .E(direction_N_4071), 
            .D(n133[16]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2248__i15 (.Q(encoder1_position[15]), .C(n1891), .E(direction_N_4071), 
            .D(n133[15]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2248__i14 (.Q(encoder1_position[14]), .C(n1891), .E(direction_N_4071), 
            .D(n133[14]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2248__i13 (.Q(encoder1_position[13]), .C(n1891), .E(direction_N_4071), 
            .D(n133[13]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2248__i12 (.Q(encoder1_position[12]), .C(n1891), .E(direction_N_4071), 
            .D(n133[12]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2248__i11 (.Q(encoder1_position[11]), .C(n1891), .E(direction_N_4071), 
            .D(n133[11]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2248__i10 (.Q(encoder1_position[10]), .C(n1891), .E(direction_N_4071), 
            .D(n133[10]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2248__i9 (.Q(encoder1_position[9]), .C(n1891), .E(direction_N_4071), 
            .D(n133[9]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2248__i8 (.Q(encoder1_position[8]), .C(n1891), .E(direction_N_4071), 
            .D(n133[8]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2248__i7 (.Q(encoder1_position[7]), .C(n1891), .E(direction_N_4071), 
            .D(n133[7]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2248__i6 (.Q(encoder1_position[6]), .C(n1891), .E(direction_N_4071), 
            .D(n133[6]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2248__i5 (.Q(encoder1_position[5]), .C(n1891), .E(direction_N_4071), 
            .D(n133[5]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2248__i4 (.Q(encoder1_position[4]), .C(n1891), .E(direction_N_4071), 
            .D(n133[4]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2248__i3 (.Q(encoder1_position[3]), .C(n1891), .E(direction_N_4071), 
            .D(n133[3]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2248__i2 (.Q(encoder1_position[2]), .C(n1891), .E(direction_N_4071), 
            .D(n133[2]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2248__i1 (.Q(encoder1_position[1]), .C(n1891), .E(direction_N_4071), 
            .D(n133[1]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_LUT4 position_2248_add_4_33_lut (.I0(GND_net), .I1(direction_N_4070), 
            .I2(encoder1_position[31]), .I3(n39407), .O(n133[31])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2248_add_4_33_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 position_2248_add_4_32_lut (.I0(GND_net), .I1(direction_N_4070), 
            .I2(encoder1_position[30]), .I3(n39406), .O(n133[30])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2248_add_4_32_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2248_add_4_32 (.CI(n39406), .I0(direction_N_4070), 
            .I1(encoder1_position[30]), .CO(n39407));
    SB_LUT4 position_2248_add_4_31_lut (.I0(GND_net), .I1(direction_N_4070), 
            .I2(encoder1_position[29]), .I3(n39405), .O(n133[29])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2248_add_4_31_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2248_add_4_31 (.CI(n39405), .I0(direction_N_4070), 
            .I1(encoder1_position[29]), .CO(n39406));
    SB_LUT4 position_2248_add_4_30_lut (.I0(GND_net), .I1(direction_N_4070), 
            .I2(encoder1_position[28]), .I3(n39404), .O(n133[28])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2248_add_4_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2248_add_4_30 (.CI(n39404), .I0(direction_N_4070), 
            .I1(encoder1_position[28]), .CO(n39405));
    SB_LUT4 position_2248_add_4_29_lut (.I0(GND_net), .I1(direction_N_4070), 
            .I2(encoder1_position[27]), .I3(n39403), .O(n133[27])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2248_add_4_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2248_add_4_29 (.CI(n39403), .I0(direction_N_4070), 
            .I1(encoder1_position[27]), .CO(n39404));
    SB_LUT4 position_2248_add_4_28_lut (.I0(GND_net), .I1(direction_N_4070), 
            .I2(encoder1_position[26]), .I3(n39402), .O(n133[26])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2248_add_4_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2248_add_4_28 (.CI(n39402), .I0(direction_N_4070), 
            .I1(encoder1_position[26]), .CO(n39403));
    SB_LUT4 position_2248_add_4_27_lut (.I0(GND_net), .I1(direction_N_4070), 
            .I2(encoder1_position[25]), .I3(n39401), .O(n133[25])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2248_add_4_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2248_add_4_27 (.CI(n39401), .I0(direction_N_4070), 
            .I1(encoder1_position[25]), .CO(n39402));
    SB_LUT4 position_2248_add_4_26_lut (.I0(GND_net), .I1(direction_N_4070), 
            .I2(encoder1_position[24]), .I3(n39400), .O(n133[24])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2248_add_4_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2248_add_4_26 (.CI(n39400), .I0(direction_N_4070), 
            .I1(encoder1_position[24]), .CO(n39401));
    SB_LUT4 position_2248_add_4_25_lut (.I0(GND_net), .I1(direction_N_4070), 
            .I2(encoder1_position[23]), .I3(n39399), .O(n133[23])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2248_add_4_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2248_add_4_25 (.CI(n39399), .I0(direction_N_4070), 
            .I1(encoder1_position[23]), .CO(n39400));
    SB_LUT4 position_2248_add_4_24_lut (.I0(GND_net), .I1(direction_N_4070), 
            .I2(encoder1_position[22]), .I3(n39398), .O(n133[22])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2248_add_4_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2248_add_4_24 (.CI(n39398), .I0(direction_N_4070), 
            .I1(encoder1_position[22]), .CO(n39399));
    SB_LUT4 position_2248_add_4_23_lut (.I0(GND_net), .I1(direction_N_4070), 
            .I2(encoder1_position[21]), .I3(n39397), .O(n133[21])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2248_add_4_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2248_add_4_23 (.CI(n39397), .I0(direction_N_4070), 
            .I1(encoder1_position[21]), .CO(n39398));
    SB_LUT4 position_2248_add_4_22_lut (.I0(GND_net), .I1(direction_N_4070), 
            .I2(encoder1_position[20]), .I3(n39396), .O(n133[20])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2248_add_4_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2248_add_4_22 (.CI(n39396), .I0(direction_N_4070), 
            .I1(encoder1_position[20]), .CO(n39397));
    SB_LUT4 position_2248_add_4_21_lut (.I0(GND_net), .I1(direction_N_4070), 
            .I2(encoder1_position[19]), .I3(n39395), .O(n133[19])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2248_add_4_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2248_add_4_21 (.CI(n39395), .I0(direction_N_4070), 
            .I1(encoder1_position[19]), .CO(n39396));
    SB_LUT4 position_2248_add_4_20_lut (.I0(GND_net), .I1(direction_N_4070), 
            .I2(encoder1_position[18]), .I3(n39394), .O(n133[18])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2248_add_4_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2248_add_4_20 (.CI(n39394), .I0(direction_N_4070), 
            .I1(encoder1_position[18]), .CO(n39395));
    SB_LUT4 position_2248_add_4_19_lut (.I0(GND_net), .I1(direction_N_4070), 
            .I2(encoder1_position[17]), .I3(n39393), .O(n133[17])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2248_add_4_19_lut.LUT_INIT = 16'hC33C;
    SB_DFFE position_2248__i0 (.Q(encoder1_position[0]), .C(n1891), .E(direction_N_4071), 
            .D(n133[0]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFF a_new_i1 (.Q(a_new[1]), .C(n1891), .D(a_new_c[0]));   // vhdl/quadrature_decoder.vhd(52[3] 89[10])
    SB_DFF b_new_i1 (.Q(b_new[1]), .C(n1891), .D(b_new[0]));   // vhdl/quadrature_decoder.vhd(52[3] 89[10])
    SB_CARRY position_2248_add_4_19 (.CI(n39393), .I0(direction_N_4070), 
            .I1(encoder1_position[17]), .CO(n39394));
    SB_LUT4 position_2248_add_4_18_lut (.I0(GND_net), .I1(direction_N_4070), 
            .I2(encoder1_position[16]), .I3(n39392), .O(n133[16])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2248_add_4_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2248_add_4_18 (.CI(n39392), .I0(direction_N_4070), 
            .I1(encoder1_position[16]), .CO(n39393));
    SB_LUT4 position_2248_add_4_17_lut (.I0(GND_net), .I1(direction_N_4070), 
            .I2(encoder1_position[15]), .I3(n39391), .O(n133[15])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2248_add_4_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2248_add_4_17 (.CI(n39391), .I0(direction_N_4070), 
            .I1(encoder1_position[15]), .CO(n39392));
    SB_LUT4 position_2248_add_4_16_lut (.I0(GND_net), .I1(direction_N_4070), 
            .I2(encoder1_position[14]), .I3(n39390), .O(n133[14])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2248_add_4_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2248_add_4_16 (.CI(n39390), .I0(direction_N_4070), 
            .I1(encoder1_position[14]), .CO(n39391));
    SB_LUT4 position_2248_add_4_15_lut (.I0(GND_net), .I1(direction_N_4070), 
            .I2(encoder1_position[13]), .I3(n39389), .O(n133[13])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2248_add_4_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2248_add_4_15 (.CI(n39389), .I0(direction_N_4070), 
            .I1(encoder1_position[13]), .CO(n39390));
    SB_LUT4 position_2248_add_4_14_lut (.I0(GND_net), .I1(direction_N_4070), 
            .I2(encoder1_position[12]), .I3(n39388), .O(n133[12])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2248_add_4_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2248_add_4_14 (.CI(n39388), .I0(direction_N_4070), 
            .I1(encoder1_position[12]), .CO(n39389));
    SB_LUT4 position_2248_add_4_13_lut (.I0(GND_net), .I1(direction_N_4070), 
            .I2(encoder1_position[11]), .I3(n39387), .O(n133[11])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2248_add_4_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2248_add_4_13 (.CI(n39387), .I0(direction_N_4070), 
            .I1(encoder1_position[11]), .CO(n39388));
    SB_LUT4 position_2248_add_4_12_lut (.I0(GND_net), .I1(direction_N_4070), 
            .I2(encoder1_position[10]), .I3(n39386), .O(n133[10])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2248_add_4_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2248_add_4_12 (.CI(n39386), .I0(direction_N_4070), 
            .I1(encoder1_position[10]), .CO(n39387));
    SB_LUT4 position_2248_add_4_11_lut (.I0(GND_net), .I1(direction_N_4070), 
            .I2(encoder1_position[9]), .I3(n39385), .O(n133[9])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2248_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2248_add_4_11 (.CI(n39385), .I0(direction_N_4070), 
            .I1(encoder1_position[9]), .CO(n39386));
    SB_LUT4 position_2248_add_4_10_lut (.I0(GND_net), .I1(direction_N_4070), 
            .I2(encoder1_position[8]), .I3(n39384), .O(n133[8])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2248_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2248_add_4_10 (.CI(n39384), .I0(direction_N_4070), 
            .I1(encoder1_position[8]), .CO(n39385));
    SB_LUT4 position_2248_add_4_9_lut (.I0(GND_net), .I1(direction_N_4070), 
            .I2(encoder1_position[7]), .I3(n39383), .O(n133[7])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2248_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2248_add_4_9 (.CI(n39383), .I0(direction_N_4070), 
            .I1(encoder1_position[7]), .CO(n39384));
    SB_LUT4 position_2248_add_4_8_lut (.I0(GND_net), .I1(direction_N_4070), 
            .I2(encoder1_position[6]), .I3(n39382), .O(n133[6])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2248_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2248_add_4_8 (.CI(n39382), .I0(direction_N_4070), 
            .I1(encoder1_position[6]), .CO(n39383));
    SB_LUT4 position_2248_add_4_7_lut (.I0(GND_net), .I1(direction_N_4070), 
            .I2(encoder1_position[5]), .I3(n39381), .O(n133[5])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2248_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2248_add_4_7 (.CI(n39381), .I0(direction_N_4070), 
            .I1(encoder1_position[5]), .CO(n39382));
    SB_LUT4 position_2248_add_4_6_lut (.I0(GND_net), .I1(direction_N_4070), 
            .I2(encoder1_position[4]), .I3(n39380), .O(n133[4])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2248_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2248_add_4_6 (.CI(n39380), .I0(direction_N_4070), 
            .I1(encoder1_position[4]), .CO(n39381));
    SB_LUT4 position_2248_add_4_5_lut (.I0(GND_net), .I1(direction_N_4070), 
            .I2(encoder1_position[3]), .I3(n39379), .O(n133[3])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2248_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2248_add_4_5 (.CI(n39379), .I0(direction_N_4070), 
            .I1(encoder1_position[3]), .CO(n39380));
    SB_LUT4 position_2248_add_4_4_lut (.I0(GND_net), .I1(direction_N_4070), 
            .I2(encoder1_position[2]), .I3(n39378), .O(n133[2])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2248_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2248_add_4_4 (.CI(n39378), .I0(direction_N_4070), 
            .I1(encoder1_position[2]), .CO(n39379));
    SB_LUT4 position_2248_add_4_3_lut (.I0(GND_net), .I1(direction_N_4070), 
            .I2(encoder1_position[1]), .I3(n39377), .O(n133[1])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2248_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2248_add_4_3 (.CI(n39377), .I0(direction_N_4070), 
            .I1(encoder1_position[1]), .CO(n39378));
    SB_LUT4 position_2248_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(encoder1_position[0]), 
            .I3(VCC_net), .O(n133[0])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2248_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2248_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(encoder1_position[0]), 
            .CO(n39377));
    SB_DFF direction_57 (.Q(n1896), .C(n1891), .D(n29245));   // vhdl/quadrature_decoder.vhd(52[3] 89[10])
    SB_DFF b_prev_52 (.Q(b_prev), .C(n1891), .D(n29222));   // vhdl/quadrature_decoder.vhd(52[3] 89[10])
    SB_LUT4 i15217_3_lut_4_lut (.I0(debounce_cnt), .I1(a_prev_N_4077), .I2(a_new[1]), 
            .I3(a_prev), .O(n29165));   // vhdl/quadrature_decoder.vhd(52[3] 89[10])
    defparam i15217_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i15274_3_lut_4_lut (.I0(debounce_cnt), .I1(a_prev_N_4077), .I2(b_new[1]), 
            .I3(b_prev), .O(n29222));   // vhdl/quadrature_decoder.vhd(52[3] 89[10])
    defparam i15274_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i34962_4_lut (.I0(a_new_c[0]), .I1(b_new[0]), .I2(a_new[1]), 
            .I3(b_new[1]), .O(a_prev_N_4077));   // vhdl/quadrature_decoder.vhd(52[3] 89[10])
    defparam i34962_4_lut.LUT_INIT = 16'h8421;
    SB_LUT4 b_prev_I_0_63_2_lut (.I0(b_prev), .I1(a_new[1]), .I2(GND_net), 
            .I3(GND_net), .O(direction_N_4070));   // vhdl/quadrature_decoder.vhd(81[18:37])
    defparam b_prev_I_0_63_2_lut.LUT_INIT = 16'h9999;
    
endmodule
//
// Verilog Description of module EEPROM
//

module EEPROM (GND_net, CLK_c, n6129, \state[1] , \state[0] , n43386, 
            read, \state[2] , n7, n29054, rw, n43506, data_ready, 
            enable_slow_N_4354, n43380, n34717, n44748, n44835, \state[3] , 
            n6, n29159, data, \state_7__N_4251[0] , n7210, sda_enable, 
            n29146, \saved_addr[0] , scl_enable, \state_7__N_4267[3] , 
            \state[0]_adj_2 , n4, n4_adj_3, n27152, n34660, scl, 
            n10, n29033, n29032, n29031, n29030, n29029, n29028, 
            n29027, n7754, sda_out, VCC_net, n27147, n8, n49357, 
            n34664) /* synthesis syn_noprune=1, syn_module_defined=1 */ ;
    input GND_net;
    input CLK_c;
    output [0:0]n6129;
    output \state[1] ;
    output \state[0] ;
    input n43386;
    input read;
    output \state[2] ;
    output n7;
    input n29054;
    output rw;
    input n43506;
    output data_ready;
    output enable_slow_N_4354;
    input n43380;
    output n34717;
    input n44748;
    output n44835;
    output \state[3] ;
    output n6;
    input n29159;
    output [7:0]data;
    output \state_7__N_4251[0] ;
    output n7210;
    output sda_enable;
    input n29146;
    output \saved_addr[0] ;
    output scl_enable;
    input \state_7__N_4267[3] ;
    output \state[0]_adj_2 ;
    output n4;
    output n4_adj_3;
    output n27152;
    output n34660;
    output scl;
    output n10;
    input n29033;
    input n29032;
    input n29031;
    input n29030;
    input n29029;
    input n29028;
    input n29027;
    input n7754;
    output sda_out;
    input VCC_net;
    output n27147;
    input n8;
    output n49357;
    output n34664;
    
    wire CLK_c /* synthesis SET_AS_NETWORK=CLK_c, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(3[9:12])
    wire [15:0]delay_counter_15__N_4153;
    wire [15:0]delay_counter;   // verilog/eeprom.v(24[12:25])
    wire [15:0]n4787;
    
    wire n38649, n38650, n38648, n28725, n29004, n38647, n38646, 
        enable, n38645, n38644, n38643, n38642, n38641, n38640, 
        n38639, n38638;
    wire [7:0]state;   // verilog/i2c_controller.v(33[12:17])
    
    wire n28, n26, n27, n25, n27021, n38652, n38651;
    
    SB_LUT4 add_1012_14_lut (.I0(GND_net), .I1(delay_counter[12]), .I2(n4787[6]), 
            .I3(n38649), .O(delay_counter_15__N_4153[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1012_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1012_14 (.CI(n38649), .I0(delay_counter[12]), .I1(n4787[6]), 
            .CO(n38650));
    SB_LUT4 add_1012_13_lut (.I0(GND_net), .I1(delay_counter[11]), .I2(n4787[6]), 
            .I3(n38648), .O(delay_counter_15__N_4153[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1012_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1012_13 (.CI(n38648), .I0(delay_counter[11]), .I1(n4787[6]), 
            .CO(n38649));
    SB_DFFESR delay_counter_i0_i1 (.Q(delay_counter[1]), .C(CLK_c), .E(n28725), 
            .D(delay_counter_15__N_4153[1]), .R(n29004));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFFESR delay_counter_i0_i2 (.Q(delay_counter[2]), .C(CLK_c), .E(n28725), 
            .D(delay_counter_15__N_4153[2]), .R(n29004));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFFESR delay_counter_i0_i3 (.Q(delay_counter[3]), .C(CLK_c), .E(n28725), 
            .D(delay_counter_15__N_4153[3]), .R(n29004));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFFESS delay_counter_i0_i4 (.Q(delay_counter[4]), .C(CLK_c), .E(n28725), 
            .D(delay_counter_15__N_4153[4]), .S(n29004));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFFESR delay_counter_i0_i5 (.Q(delay_counter[5]), .C(CLK_c), .E(n28725), 
            .D(delay_counter_15__N_4153[5]), .R(n29004));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFFESS delay_counter_i0_i6 (.Q(delay_counter[6]), .C(CLK_c), .E(n28725), 
            .D(delay_counter_15__N_4153[6]), .S(n29004));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFFESS delay_counter_i0_i7 (.Q(delay_counter[7]), .C(CLK_c), .E(n28725), 
            .D(delay_counter_15__N_4153[7]), .S(n29004));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFFESS delay_counter_i0_i8 (.Q(delay_counter[8]), .C(CLK_c), .E(n28725), 
            .D(delay_counter_15__N_4153[8]), .S(n29004));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFFESS delay_counter_i0_i9 (.Q(delay_counter[9]), .C(CLK_c), .E(n28725), 
            .D(delay_counter_15__N_4153[9]), .S(n29004));   // verilog/eeprom.v(26[8] 58[4])
    SB_LUT4 add_1012_12_lut (.I0(GND_net), .I1(delay_counter[10]), .I2(n4787[6]), 
            .I3(n38647), .O(delay_counter_15__N_4153[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1012_12_lut.LUT_INIT = 16'hC33C;
    SB_DFFESS delay_counter_i0_i10 (.Q(delay_counter[10]), .C(CLK_c), .E(n28725), 
            .D(delay_counter_15__N_4153[10]), .S(n29004));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFFESR delay_counter_i0_i11 (.Q(delay_counter[11]), .C(CLK_c), .E(n28725), 
            .D(delay_counter_15__N_4153[11]), .R(n29004));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFFESR delay_counter_i0_i12 (.Q(delay_counter[12]), .C(CLK_c), .E(n28725), 
            .D(delay_counter_15__N_4153[12]), .R(n29004));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFFESR delay_counter_i0_i13 (.Q(delay_counter[13]), .C(CLK_c), .E(n28725), 
            .D(delay_counter_15__N_4153[13]), .R(n29004));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFFESR delay_counter_i0_i14 (.Q(delay_counter[14]), .C(CLK_c), .E(n28725), 
            .D(delay_counter_15__N_4153[14]), .R(n29004));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFFESR delay_counter_i0_i15 (.Q(delay_counter[15]), .C(CLK_c), .E(n28725), 
            .D(delay_counter_15__N_4153[15]), .R(n29004));   // verilog/eeprom.v(26[8] 58[4])
    SB_CARRY add_1012_12 (.CI(n38647), .I0(delay_counter[10]), .I1(n4787[6]), 
            .CO(n38648));
    SB_LUT4 add_1012_11_lut (.I0(GND_net), .I1(delay_counter[9]), .I2(n4787[6]), 
            .I3(n38646), .O(delay_counter_15__N_4153[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1012_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1012_11 (.CI(n38646), .I0(delay_counter[9]), .I1(n4787[6]), 
            .CO(n38647));
    SB_DFFSR enable_39 (.Q(enable), .C(CLK_c), .D(n6129[0]), .R(\state[1] ));   // verilog/eeprom.v(26[8] 58[4])
    SB_LUT4 add_1012_10_lut (.I0(GND_net), .I1(delay_counter[8]), .I2(n4787[6]), 
            .I3(n38645), .O(delay_counter_15__N_4153[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1012_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1012_10 (.CI(n38645), .I0(delay_counter[8]), .I1(n4787[6]), 
            .CO(n38646));
    SB_LUT4 add_1012_9_lut (.I0(GND_net), .I1(delay_counter[7]), .I2(n4787[6]), 
            .I3(n38644), .O(delay_counter_15__N_4153[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1012_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1012_9 (.CI(n38644), .I0(delay_counter[7]), .I1(n4787[6]), 
            .CO(n38645));
    SB_LUT4 add_1012_8_lut (.I0(GND_net), .I1(delay_counter[6]), .I2(n4787[6]), 
            .I3(n38643), .O(delay_counter_15__N_4153[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1012_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1012_8 (.CI(n38643), .I0(delay_counter[6]), .I1(n4787[6]), 
            .CO(n38644));
    SB_LUT4 add_1012_7_lut (.I0(GND_net), .I1(delay_counter[5]), .I2(n4787[6]), 
            .I3(n38642), .O(delay_counter_15__N_4153[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1012_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1012_7 (.CI(n38642), .I0(delay_counter[5]), .I1(n4787[6]), 
            .CO(n38643));
    SB_LUT4 add_1012_6_lut (.I0(GND_net), .I1(delay_counter[4]), .I2(n4787[6]), 
            .I3(n38641), .O(delay_counter_15__N_4153[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1012_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1012_6 (.CI(n38641), .I0(delay_counter[4]), .I1(n4787[6]), 
            .CO(n38642));
    SB_LUT4 add_1012_5_lut (.I0(GND_net), .I1(delay_counter[3]), .I2(n4787[6]), 
            .I3(n38640), .O(delay_counter_15__N_4153[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1012_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1012_5 (.CI(n38640), .I0(delay_counter[3]), .I1(n4787[6]), 
            .CO(n38641));
    SB_LUT4 add_1012_4_lut (.I0(GND_net), .I1(delay_counter[2]), .I2(n4787[6]), 
            .I3(n38639), .O(delay_counter_15__N_4153[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1012_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1012_4 (.CI(n38639), .I0(delay_counter[2]), .I1(n4787[6]), 
            .CO(n38640));
    SB_LUT4 add_1012_3_lut (.I0(GND_net), .I1(delay_counter[1]), .I2(n4787[6]), 
            .I3(n38638), .O(delay_counter_15__N_4153[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1012_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1012_3 (.CI(n38638), .I0(delay_counter[1]), .I1(n4787[6]), 
            .CO(n38639));
    SB_LUT4 add_1012_2_lut (.I0(GND_net), .I1(delay_counter[0]), .I2(n4787[6]), 
            .I3(GND_net), .O(delay_counter_15__N_4153[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1012_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1012_2 (.CI(GND_net), .I0(delay_counter[0]), .I1(n4787[6]), 
            .CO(n38638));
    SB_DFFESR delay_counter_i0_i0 (.Q(delay_counter[0]), .C(CLK_c), .E(n28725), 
            .D(delay_counter_15__N_4153[0]), .R(n29004));   // verilog/eeprom.v(26[8] 58[4])
    SB_LUT4 i15069_2_lut (.I0(n28725), .I1(\state[0] ), .I2(GND_net), 
            .I3(GND_net), .O(n29004));   // verilog/eeprom.v(26[8] 58[4])
    defparam i15069_2_lut.LUT_INIT = 16'h2222;
    SB_DFF state__i0 (.Q(\state[0] ), .C(CLK_c), .D(n43386));   // verilog/eeprom.v(26[8] 58[4])
    SB_LUT4 i1_3_lut (.I0(read), .I1(\state[1] ), .I2(\state[0] ), .I3(GND_net), 
            .O(n28725));
    defparam i1_3_lut.LUT_INIT = 16'h3232;
    SB_LUT4 i2_2_lut (.I0(state[1]), .I1(\state[2] ), .I2(GND_net), .I3(GND_net), 
            .O(n7));   // verilog/eeprom.v(42[12:28])
    defparam i2_2_lut.LUT_INIT = 16'heeee;
    SB_DFF rw_43 (.Q(rw), .C(CLK_c), .D(n29054));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFF data_ready_42 (.Q(data_ready), .C(CLK_c), .D(n43506));   // verilog/eeprom.v(26[8] 58[4])
    SB_LUT4 i12_4_lut (.I0(delay_counter[6]), .I1(delay_counter[10]), .I2(delay_counter[12]), 
            .I3(delay_counter[8]), .O(n28));   // verilog/eeprom.v(42[12:28])
    defparam i12_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i10_4_lut (.I0(delay_counter[11]), .I1(delay_counter[2]), .I2(delay_counter[7]), 
            .I3(delay_counter[5]), .O(n26));   // verilog/eeprom.v(42[12:28])
    defparam i10_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i11_4_lut (.I0(delay_counter[15]), .I1(delay_counter[3]), .I2(delay_counter[14]), 
            .I3(delay_counter[1]), .O(n27));   // verilog/eeprom.v(42[12:28])
    defparam i11_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i9_4_lut (.I0(delay_counter[4]), .I1(delay_counter[9]), .I2(delay_counter[13]), 
            .I3(delay_counter[0]), .O(n25));   // verilog/eeprom.v(42[12:28])
    defparam i9_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut (.I0(n25), .I1(n27), .I2(n26), .I3(n28), .O(n27021));   // verilog/eeprom.v(42[12:28])
    defparam i15_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i34969_2_lut (.I0(n27021), .I1(enable_slow_N_4354), .I2(GND_net), 
            .I3(GND_net), .O(n4787[6]));   // verilog/eeprom.v(46[18] 48[12])
    defparam i34969_2_lut.LUT_INIT = 16'h2222;
    SB_DFF state__i1 (.Q(\state[1] ), .C(CLK_c), .D(n43380));   // verilog/eeprom.v(26[8] 58[4])
    SB_LUT4 add_1012_17_lut (.I0(GND_net), .I1(delay_counter[15]), .I2(n4787[6]), 
            .I3(n38652), .O(delay_counter_15__N_4153[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1012_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_1012_16_lut (.I0(GND_net), .I1(delay_counter[14]), .I2(n4787[6]), 
            .I3(n38651), .O(delay_counter_15__N_4153[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1012_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1012_16 (.CI(n38651), .I0(delay_counter[14]), .I1(n4787[6]), 
            .CO(n38652));
    SB_LUT4 add_1012_15_lut (.I0(GND_net), .I1(delay_counter[13]), .I2(n4787[6]), 
            .I3(n38650), .O(delay_counter_15__N_4153[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1012_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1012_15 (.CI(n38650), .I0(delay_counter[13]), .I1(n4787[6]), 
            .CO(n38651));
    SB_LUT4 i21329_2_lut_3_lut (.I0(\state[0] ), .I1(\state[1] ), .I2(enable_slow_N_4354), 
            .I3(GND_net), .O(n34717));   // verilog/eeprom.v(51[5:9])
    defparam i21329_2_lut_3_lut.LUT_INIT = 16'hfbfb;
    SB_LUT4 i29315_4_lut_4_lut (.I0(\state[0] ), .I1(\state[1] ), .I2(n44748), 
            .I3(enable_slow_N_4354), .O(n44835));   // verilog/eeprom.v(51[5:9])
    defparam i29315_4_lut_4_lut.LUT_INIT = 16'hfcf8;
    SB_LUT4 i2_2_lut_adj_953 (.I0(\state[3] ), .I1(n27021), .I2(GND_net), 
            .I3(GND_net), .O(n6));   // verilog/eeprom.v(42[12:28])
    defparam i2_2_lut_adj_953.LUT_INIT = 16'heeee;
    SB_LUT4 mux_1460_Mux_0_i1_4_lut (.I0(read), .I1(n27021), .I2(\state[0] ), 
            .I3(enable_slow_N_4354), .O(n6129[0]));   // verilog/eeprom.v(29[3] 57[10])
    defparam mux_1460_Mux_0_i1_4_lut.LUT_INIT = 16'h0a3a;
    i2c_controller i2c (.n29159(n29159), .data({data}), .\state_7__N_4251[0] (\state_7__N_4251[0] ), 
            .enable_slow_N_4354(enable_slow_N_4354), .GND_net(GND_net), 
            .n7210(n7210), .\state[1] (state[1]), .\state[2] (\state[2] ), 
            .CLK_c(CLK_c), .sda_enable(sda_enable), .n29146(n29146), .\saved_addr[0] (\saved_addr[0] ), 
            .scl_enable(scl_enable), .\state[3] (\state[3] ), .\state_7__N_4267[3] (\state_7__N_4267[3] ), 
            .\state[0] (\state[0]_adj_2 ), .n4(n4), .n4_adj_1(n4_adj_3), 
            .n27152(n27152), .n34660(n34660), .scl(scl), .n10(n10), 
            .n29033(n29033), .n29032(n29032), .n29031(n29031), .n29030(n29030), 
            .n29029(n29029), .n29028(n29028), .n29027(n29027), .n7754(n7754), 
            .sda_out(sda_out), .VCC_net(VCC_net), .n27147(n27147), .n8(n8), 
            .n49357(n49357), .n34664(n34664), .enable(enable)) /* synthesis syn_noprune=1, syn_module_defined=1 */ ;   // verilog/eeprom.v(60[16] 74[4])
    
endmodule
//
// Verilog Description of module i2c_controller
//

module i2c_controller (n29159, data, \state_7__N_4251[0] , enable_slow_N_4354, 
            GND_net, n7210, \state[1] , \state[2] , CLK_c, sda_enable, 
            n29146, \saved_addr[0] , scl_enable, \state[3] , \state_7__N_4267[3] , 
            \state[0] , n4, n4_adj_1, n27152, n34660, scl, n10, 
            n29033, n29032, n29031, n29030, n29029, n29028, n29027, 
            n7754, sda_out, VCC_net, n27147, n8, n49357, n34664, 
            enable) /* synthesis syn_noprune=1, syn_module_defined=1 */ ;
    input n29159;
    output [7:0]data;
    output \state_7__N_4251[0] ;
    output enable_slow_N_4354;
    input GND_net;
    output n7210;
    output \state[1] ;
    output \state[2] ;
    input CLK_c;
    output sda_enable;
    input n29146;
    output \saved_addr[0] ;
    output scl_enable;
    output \state[3] ;
    input \state_7__N_4267[3] ;
    output \state[0] ;
    output n4;
    output n4_adj_1;
    output n27152;
    output n34660;
    output scl;
    output n10;
    input n29033;
    input n29032;
    input n29031;
    input n29030;
    input n29029;
    input n29028;
    input n29027;
    input n7754;
    output sda_out;
    input VCC_net;
    output n27147;
    input n8;
    output n49357;
    output n34664;
    input enable;
    
    wire i2c_clk /* synthesis is_clock=1, SET_AS_NETWORK=\eeprom/i2c/i2c_clk */ ;   // verilog/i2c_controller.v(41[6:13])
    wire CLK_c /* synthesis SET_AS_NETWORK=CLK_c, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(3[9:12])
    wire [7:0]n119;
    
    wire n28652;
    wire [7:0]counter;   // verilog/i2c_controller.v(36[12:19])
    
    wire n28919, enable_slow_N_4353, n5, n34873, n34863, n34871;
    wire [5:0]n29;
    wire [7:0]counter2;   // verilog/i2c_controller.v(37[12:20])
    
    wire n28864, n19508, n7616, n28861, i2c_clk_N_4340;
    wire [0:0]n7053;
    
    wire n43412, sda_out_adj_4574, scl_enable_N_4341, n43608, n45729, 
        n28594, n34673, n10_c, n13, n16, n9, n49300, n49288, 
        n7017, n15, n12, n7203, n15_adj_4577, n44752, n37, n33_adj_4578, 
        n34_adj_4579, n39, n10_adj_4580, n11, n11_adj_4581, n38827, 
        n38826, n38825, n38824, n38823, n38822, n38821, n39482, 
        n39481, n39480, n39479, n39478, state_7__N_4250, n11_adj_4582, 
        n11_adj_4583;
    
    SB_DFF data_out_i0_i0 (.Q(data[0]), .C(i2c_clk), .D(n29159));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESS counter_i1 (.Q(counter[1]), .C(i2c_clk), .E(n28652), .D(n119[1]), 
            .S(n28919));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESS counter_i2 (.Q(counter[2]), .C(i2c_clk), .E(n28652), .D(n119[2]), 
            .S(n28919));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESR counter_i3 (.Q(counter[3]), .C(i2c_clk), .E(n28652), .D(n119[3]), 
            .R(n28919));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESR counter_i4 (.Q(counter[4]), .C(i2c_clk), .E(n28652), .D(n119[4]), 
            .R(n28919));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESR counter_i5 (.Q(counter[5]), .C(i2c_clk), .E(n28652), .D(n119[5]), 
            .R(n28919));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESR counter_i6 (.Q(counter[6]), .C(i2c_clk), .E(n28652), .D(n119[6]), 
            .R(n28919));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESR counter_i7 (.Q(counter[7]), .C(i2c_clk), .E(n28652), .D(n119[7]), 
            .R(n28919));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_LUT4 i34902_2_lut (.I0(\state_7__N_4251[0] ), .I1(enable_slow_N_4354), 
            .I2(GND_net), .I3(GND_net), .O(enable_slow_N_4353));   // verilog/i2c_controller.v(62[6:32])
    defparam i34902_2_lut.LUT_INIT = 16'h7777;
    SB_DFFESS state_i0_i1 (.Q(\state[1] ), .C(i2c_clk), .E(n7210), .D(n5), 
            .S(n34873));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESS state_i0_i2 (.Q(\state[2] ), .C(i2c_clk), .E(n7210), .D(n34863), 
            .S(n34871));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFSR counter2_2259_2260__i6 (.Q(counter2[5]), .C(CLK_c), .D(n29[5]), 
            .R(n28864));   // verilog/i2c_controller.v(69[20:35])
    SB_DFFNESS write_enable_131 (.Q(sda_enable), .C(i2c_clk), .E(n7616), 
            .D(n19508), .S(n28861));   // verilog/i2c_controller.v(180[12] 215[6])
    SB_DFF saved_addr__i1 (.Q(\saved_addr[0] ), .C(i2c_clk), .D(n29146));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFF i2c_clk_121 (.Q(i2c_clk), .C(CLK_c), .D(i2c_clk_N_4340));   // verilog/i2c_controller.v(58[9] 71[5])
    SB_DFFNE sda_out_132 (.Q(sda_out_adj_4574), .C(i2c_clk), .E(n43412), 
            .D(n7053[0]));   // verilog/i2c_controller.v(180[12] 215[6])
    SB_DFFESS counter_i0 (.Q(counter[0]), .C(i2c_clk), .E(n28652), .D(n119[0]), 
            .S(n28919));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFN i2c_scl_enable_123 (.Q(scl_enable), .C(i2c_clk), .D(scl_enable_N_4341));   // verilog/i2c_controller.v(76[12] 82[6])
    SB_DFFESS state_i0_i3 (.Q(\state[3] ), .C(i2c_clk), .E(n7210), .D(n43608), 
            .S(n45729));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFE enable_slow_120 (.Q(\state_7__N_4251[0] ), .C(CLK_c), .E(n28594), 
            .D(enable_slow_N_4353));   // verilog/i2c_controller.v(58[9] 71[5])
    SB_LUT4 i1_4_lut (.I0(n34673), .I1(n10_c), .I2(n13), .I3(\state_7__N_4267[3] ), 
            .O(n16));   // verilog/i2c_controller.v(92[4] 172[11])
    defparam i1_4_lut.LUT_INIT = 16'ha2a0;
    SB_LUT4 i1_4_lut_adj_947 (.I0(\state[2] ), .I1(n16), .I2(\state[3] ), 
            .I3(n9), .O(n43608));   // verilog/i2c_controller.v(92[4] 172[11])
    defparam i1_4_lut_adj_947.LUT_INIT = 16'hccdc;
    SB_LUT4 i33783_2_lut (.I0(counter[1]), .I1(\saved_addr[0] ), .I2(GND_net), 
            .I3(GND_net), .O(n49300));   // verilog/i2c_controller.v(198[28:35])
    defparam i33783_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i33801_4_lut (.I0(n49300), .I1(\state[1] ), .I2(counter[0]), 
            .I3(counter[2]), .O(n49288));   // verilog/i2c_controller.v(181[4] 214[11])
    defparam i33801_4_lut.LUT_INIT = 16'hc008;
    SB_LUT4 mux_1671_i1_4_lut (.I0(n49288), .I1(\state[0] ), .I2(n7017), 
            .I3(\state[2] ), .O(n7053[0]));   // verilog/i2c_controller.v(181[4] 214[11])
    defparam mux_1671_i1_4_lut.LUT_INIT = 16'h303a;
    SB_DFFSR counter2_2259_2260__i5 (.Q(counter2[4]), .C(CLK_c), .D(n29[4]), 
            .R(n28864));   // verilog/i2c_controller.v(69[20:35])
    SB_LUT4 i1_2_lut (.I0(i2c_clk), .I1(n28864), .I2(GND_net), .I3(GND_net), 
            .O(i2c_clk_N_4340));
    defparam i1_2_lut.LUT_INIT = 16'h6666;
    SB_DFFSR counter2_2259_2260__i4 (.Q(counter2[3]), .C(CLK_c), .D(n29[3]), 
            .R(n28864));   // verilog/i2c_controller.v(69[20:35])
    SB_DFFSR counter2_2259_2260__i3 (.Q(counter2[2]), .C(CLK_c), .D(n29[2]), 
            .R(n28864));   // verilog/i2c_controller.v(69[20:35])
    SB_DFFSR counter2_2259_2260__i2 (.Q(counter2[1]), .C(CLK_c), .D(n29[1]), 
            .R(n28864));   // verilog/i2c_controller.v(69[20:35])
    SB_LUT4 equal_354_i4_2_lut (.I0(counter[1]), .I1(counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n4));   // verilog/i2c_controller.v(153[6:23])
    defparam equal_354_i4_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 equal_352_i4_2_lut (.I0(counter[1]), .I1(counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n4_adj_1));   // verilog/i2c_controller.v(153[6:23])
    defparam equal_352_i4_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 i1_2_lut_adj_948 (.I0(n15), .I1(counter[0]), .I2(GND_net), 
            .I3(GND_net), .O(n27152));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i1_2_lut_adj_948.LUT_INIT = 16'hbbbb;
    SB_LUT4 i20730_2_lut (.I0(counter[1]), .I1(counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n34660));
    defparam i20730_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i20714_2_lut (.I0(i2c_clk), .I1(scl_enable), .I2(GND_net), 
            .I3(GND_net), .O(scl));   // verilog/i2c_controller.v(45[19:61])
    defparam i20714_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 equal_277_i10_2_lut (.I0(\state[2] ), .I1(\state[3] ), .I2(GND_net), 
            .I3(GND_net), .O(n10_c));   // verilog/i2c_controller.v(77[27:43])
    defparam equal_277_i10_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i5_4_lut (.I0(counter[3]), .I1(counter[5]), .I2(counter[0]), 
            .I3(counter[4]), .O(n12));   // verilog/i2c_controller.v(110[10:22])
    defparam i5_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i6_4_lut (.I0(counter[6]), .I1(n12), .I2(counter[7]), .I3(n10), 
            .O(n7203));   // verilog/i2c_controller.v(110[10:22])
    defparam i6_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i29236_2_lut (.I0(\state_7__N_4267[3] ), .I1(n15_adj_4577), 
            .I2(GND_net), .I3(GND_net), .O(n44752));
    defparam i29236_2_lut.LUT_INIT = 16'h8888;
    SB_DFF data_out_i0_i7 (.Q(data[7]), .C(i2c_clk), .D(n29033));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFF data_out_i0_i6 (.Q(data[6]), .C(i2c_clk), .D(n29032));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFF data_out_i0_i5 (.Q(data[5]), .C(i2c_clk), .D(n29031));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFF data_out_i0_i4 (.Q(data[4]), .C(i2c_clk), .D(n29030));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFF data_out_i0_i3 (.Q(data[3]), .C(i2c_clk), .D(n29029));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFF data_out_i0_i2 (.Q(data[2]), .C(i2c_clk), .D(n29028));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFF data_out_i0_i1 (.Q(data[1]), .C(i2c_clk), .D(n29027));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFSR counter2_2259_2260__i1 (.Q(counter2[0]), .C(CLK_c), .D(n29[0]), 
            .R(n28864));   // verilog/i2c_controller.v(69[20:35])
    SB_LUT4 i17_4_lut (.I0(n7203), .I1(n44752), .I2(n7754), .I3(n37), 
            .O(n28652));
    defparam i17_4_lut.LUT_INIT = 16'h3a30;
    SB_LUT4 equal_277_i11_2_lut_3_lut_4_lut (.I0(\state[0] ), .I1(\state[1] ), 
            .I2(\state[2] ), .I3(\state[3] ), .O(n15_adj_4577));   // verilog/i2c_controller.v(77[27:43])
    defparam equal_277_i11_2_lut_3_lut_4_lut.LUT_INIT = 16'hfffd;
    SB_LUT4 i56_3_lut (.I0(\state[2] ), .I1(\state[0] ), .I2(\state[3] ), 
            .I3(GND_net), .O(n33_adj_4578));
    defparam i56_3_lut.LUT_INIT = 16'h1c1c;
    SB_LUT4 i1_3_lut (.I0(\state[1] ), .I1(n33_adj_4578), .I2(n37), .I3(GND_net), 
            .O(n28861));
    defparam i1_3_lut.LUT_INIT = 16'h5454;
    SB_LUT4 i2684_2_lut (.I0(sda_out_adj_4574), .I1(sda_enable), .I2(GND_net), 
            .I3(GND_net), .O(sda_out));   // verilog/i2c_controller.v(46[9:20])
    defparam i2684_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_949 (.I0(n34_adj_4579), .I1(n37), .I2(GND_net), 
            .I3(GND_net), .O(n39));
    defparam i1_2_lut_adj_949.LUT_INIT = 16'heeee;
    SB_LUT4 i35014_4_lut (.I0(n7017), .I1(n39), .I2(\state[2] ), .I3(\state[1] ), 
            .O(n7616));
    defparam i35014_4_lut.LUT_INIT = 16'hc8cc;
    SB_LUT4 i34976_2_lut (.I0(\state[0] ), .I1(n7017), .I2(GND_net), .I3(GND_net), 
            .O(n19508));   // verilog/i2c_controller.v(181[4] 214[11])
    defparam i34976_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i4_4_lut (.I0(counter2[3]), .I1(counter2[5]), .I2(counter2[2]), 
            .I3(counter2[4]), .O(n10_adj_4580));
    defparam i4_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i5_3_lut (.I0(counter2[1]), .I1(n10_adj_4580), .I2(counter2[0]), 
            .I3(GND_net), .O(n28864));
    defparam i5_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 equal_2238_i19_2_lut_3_lut_4_lut (.I0(\state[0] ), .I1(\state[1] ), 
            .I2(\state[2] ), .I3(\state[3] ), .O(enable_slow_N_4354));   // verilog/i2c_controller.v(77[47:62])
    defparam equal_2238_i19_2_lut_3_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i35550_3_lut (.I0(n7210), .I1(n15), .I2(n11), .I3(GND_net), 
            .O(n34871));
    defparam i35550_3_lut.LUT_INIT = 16'h2a2a;
    SB_LUT4 i35543_2_lut (.I0(\state_7__N_4267[3] ), .I1(n11_adj_4581), 
            .I2(GND_net), .I3(GND_net), .O(n34863));
    defparam i35543_2_lut.LUT_INIT = 16'h1111;
    SB_LUT4 state_7__I_0_143_i11_2_lut_3_lut_4_lut (.I0(\state[2] ), .I1(\state[3] ), 
            .I2(\state[0] ), .I3(\state[1] ), .O(n15));   // verilog/i2c_controller.v(151[5:14])
    defparam state_7__I_0_143_i11_2_lut_3_lut_4_lut.LUT_INIT = 16'hfdff;
    SB_LUT4 state_7__I_0_143_i9_2_lut (.I0(\state[0] ), .I1(\state[1] ), 
            .I2(GND_net), .I3(GND_net), .O(n9));   // verilog/i2c_controller.v(151[5:14])
    defparam state_7__I_0_143_i9_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 sub_39_add_2_9_lut (.I0(GND_net), .I1(counter[7]), .I2(VCC_net), 
            .I3(n38827), .O(n119[7])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_39_add_2_8_lut (.I0(GND_net), .I1(counter[6]), .I2(VCC_net), 
            .I3(n38826), .O(n119[6])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_39_add_2_8 (.CI(n38826), .I0(counter[6]), .I1(VCC_net), 
            .CO(n38827));
    SB_LUT4 sub_39_add_2_7_lut (.I0(GND_net), .I1(counter[5]), .I2(VCC_net), 
            .I3(n38825), .O(n119[5])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_39_add_2_7 (.CI(n38825), .I0(counter[5]), .I1(VCC_net), 
            .CO(n38826));
    SB_LUT4 sub_39_add_2_6_lut (.I0(GND_net), .I1(counter[4]), .I2(VCC_net), 
            .I3(n38824), .O(n119[4])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_39_add_2_6 (.CI(n38824), .I0(counter[4]), .I1(VCC_net), 
            .CO(n38825));
    SB_LUT4 sub_39_add_2_5_lut (.I0(GND_net), .I1(counter[3]), .I2(VCC_net), 
            .I3(n38823), .O(n119[3])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_39_add_2_5 (.CI(n38823), .I0(counter[3]), .I1(VCC_net), 
            .CO(n38824));
    SB_LUT4 sub_39_add_2_4_lut (.I0(GND_net), .I1(counter[2]), .I2(VCC_net), 
            .I3(n38822), .O(n119[2])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_39_add_2_4 (.CI(n38822), .I0(counter[2]), .I1(VCC_net), 
            .CO(n38823));
    SB_LUT4 sub_39_add_2_3_lut (.I0(GND_net), .I1(counter[1]), .I2(VCC_net), 
            .I3(n38821), .O(n119[1])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_39_add_2_3 (.CI(n38821), .I0(counter[1]), .I1(VCC_net), 
            .CO(n38822));
    SB_LUT4 sub_39_add_2_2_lut (.I0(GND_net), .I1(counter[0]), .I2(GND_net), 
            .I3(VCC_net), .O(n119[0])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_39_add_2_2 (.CI(VCC_net), .I0(counter[0]), .I1(GND_net), 
            .CO(n38821));
    SB_LUT4 counter2_2259_2260_add_4_7_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter2[5]), .I3(n39482), .O(n29[5])) /* synthesis syn_instantiated=1 */ ;
    defparam counter2_2259_2260_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 counter2_2259_2260_add_4_6_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter2[4]), .I3(n39481), .O(n29[4])) /* synthesis syn_instantiated=1 */ ;
    defparam counter2_2259_2260_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter2_2259_2260_add_4_6 (.CI(n39481), .I0(GND_net), .I1(counter2[4]), 
            .CO(n39482));
    SB_LUT4 counter2_2259_2260_add_4_5_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter2[3]), .I3(n39480), .O(n29[3])) /* synthesis syn_instantiated=1 */ ;
    defparam counter2_2259_2260_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter2_2259_2260_add_4_5 (.CI(n39480), .I0(GND_net), .I1(counter2[3]), 
            .CO(n39481));
    SB_LUT4 counter2_2259_2260_add_4_4_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter2[2]), .I3(n39479), .O(n29[2])) /* synthesis syn_instantiated=1 */ ;
    defparam counter2_2259_2260_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter2_2259_2260_add_4_4 (.CI(n39479), .I0(GND_net), .I1(counter2[2]), 
            .CO(n39480));
    SB_LUT4 counter2_2259_2260_add_4_3_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter2[1]), .I3(n39478), .O(n29[1])) /* synthesis syn_instantiated=1 */ ;
    defparam counter2_2259_2260_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter2_2259_2260_add_4_3 (.CI(n39478), .I0(GND_net), .I1(counter2[1]), 
            .CO(n39479));
    SB_LUT4 counter2_2259_2260_add_4_2_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter2[0]), .I3(VCC_net), .O(n29[0])) /* synthesis syn_instantiated=1 */ ;
    defparam counter2_2259_2260_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter2_2259_2260_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(counter2[0]), 
            .CO(n39478));
    SB_LUT4 i1_2_lut_adj_950 (.I0(counter[0]), .I1(n15), .I2(GND_net), 
            .I3(GND_net), .O(n27147));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i1_2_lut_adj_950.LUT_INIT = 16'heeee;
    SB_LUT4 i2_2_lut (.I0(counter[2]), .I1(counter[1]), .I2(GND_net), 
            .I3(GND_net), .O(n10));   // verilog/i2c_controller.v(110[10:22])
    defparam i2_2_lut.LUT_INIT = 16'heeee;
    SB_DFFE state_i0_i0 (.Q(\state[0] ), .C(i2c_clk), .E(VCC_net), .D(n8));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_LUT4 i21308_3_lut_4_lut (.I0(\state[3] ), .I1(\state[2] ), .I2(\state[0] ), 
            .I3(\state[1] ), .O(state_7__N_4250));
    defparam i21308_3_lut_4_lut.LUT_INIT = 16'ha888;
    SB_LUT4 state_7__I_0_138_i11_2_lut_4_lut (.I0(\state[0] ), .I1(\state[1] ), 
            .I2(\state[2] ), .I3(\state[3] ), .O(n11_adj_4582));   // verilog/i2c_controller.v(109[5:12])
    defparam state_7__I_0_138_i11_2_lut_4_lut.LUT_INIT = 16'hfffb;
    SB_LUT4 state_7__I_0_139_i11_2_lut_4_lut (.I0(\state[0] ), .I1(\state[1] ), 
            .I2(\state[2] ), .I3(\state[3] ), .O(n11_adj_4581));   // verilog/i2c_controller.v(117[5:13])
    defparam state_7__I_0_139_i11_2_lut_4_lut.LUT_INIT = 16'hfff7;
    SB_LUT4 i35012_4_lut_4_lut (.I0(\state[1] ), .I1(\state[2] ), .I2(\state[0] ), 
            .I3(\state[3] ), .O(n43412));
    defparam i35012_4_lut_4_lut.LUT_INIT = 16'h0156;
    SB_LUT4 i1_2_lut_4_lut (.I0(\state[1] ), .I1(\state[2] ), .I2(\state[0] ), 
            .I3(\state[3] ), .O(n34_adj_4579));
    defparam i1_2_lut_4_lut.LUT_INIT = 16'h0150;
    SB_LUT4 i29189_2_lut_4_lut (.I0(\state[0] ), .I1(\state[2] ), .I2(\state[3] ), 
            .I3(n44752), .O(n28919));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i29189_2_lut_4_lut.LUT_INIT = 16'h0002;
    SB_LUT4 i33867_3_lut_4_lut (.I0(n11_adj_4582), .I1(n11), .I2(enable_slow_N_4354), 
            .I3(\state_7__N_4251[0] ), .O(n49357));
    defparam i33867_3_lut_4_lut.LUT_INIT = 16'h8088;
    SB_LUT4 i35552_3_lut_4_lut (.I0(n11_adj_4582), .I1(n11), .I2(n15_adj_4577), 
            .I3(n7210), .O(n34873));
    defparam i35552_3_lut_4_lut.LUT_INIT = 16'h7f00;
    SB_LUT4 i1_2_lut_4_lut_adj_951 (.I0(\state[3] ), .I1(\state[1] ), .I2(\state[2] ), 
            .I3(\state[0] ), .O(n37));
    defparam i1_2_lut_4_lut_adj_951.LUT_INIT = 16'h0554;
    SB_LUT4 i20743_2_lut (.I0(\state[0] ), .I1(\state[1] ), .I2(GND_net), 
            .I3(GND_net), .O(n34673));
    defparam i20743_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i34910_4_lut (.I0(state_7__N_4250), .I1(n7203), .I2(n11_adj_4582), 
            .I3(n34664), .O(n7210));
    defparam i34910_4_lut.LUT_INIT = 16'h5111;
    SB_LUT4 i1_4_lut_adj_952 (.I0(n11_adj_4583), .I1(n11_adj_4581), .I2(\state_7__N_4267[3] ), 
            .I3(\saved_addr[0] ), .O(n5));   // verilog/i2c_controller.v(92[4] 172[11])
    defparam i1_4_lut_adj_952.LUT_INIT = 16'h5755;
    SB_LUT4 i35548_3_lut_4_lut (.I0(\state[2] ), .I1(\state[3] ), .I2(n7210), 
            .I3(\state[1] ), .O(n45729));   // verilog/i2c_controller.v(151[5:14])
    defparam i35548_3_lut_4_lut.LUT_INIT = 16'h0020;
    SB_LUT4 i1_3_lut_4_lut (.I0(\state[2] ), .I1(\state[3] ), .I2(enable), 
            .I3(\state_7__N_4267[3] ), .O(n13));   // verilog/i2c_controller.v(151[5:14])
    defparam i1_3_lut_4_lut.LUT_INIT = 16'h2202;
    SB_LUT4 i21320_2_lut_3_lut (.I0(\state[2] ), .I1(\state[3] ), .I2(\state[0] ), 
            .I3(GND_net), .O(n34664));   // verilog/i2c_controller.v(151[5:14])
    defparam i21320_2_lut_3_lut.LUT_INIT = 16'hfdfd;
    SB_LUT4 state_7__I_0_144_i11_2_lut_3_lut_4_lut (.I0(\state[2] ), .I1(\state[3] ), 
            .I2(\state[1] ), .I3(\state[0] ), .O(n11_adj_4583));   // verilog/i2c_controller.v(151[5:14])
    defparam state_7__I_0_144_i11_2_lut_3_lut_4_lut.LUT_INIT = 16'hfdff;
    SB_LUT4 i21426_3_lut_4_lut (.I0(\state[0] ), .I1(\state[1] ), .I2(\state[2] ), 
            .I3(n15_adj_4577), .O(scl_enable_N_4341));   // verilog/i2c_controller.v(77[47:62])
    defparam i21426_3_lut_4_lut.LUT_INIT = 16'hfe00;
    SB_LUT4 i3_4_lut_4_lut (.I0(\state[0] ), .I1(\state[1] ), .I2(\state[3] ), 
            .I3(\state[2] ), .O(n7017));   // verilog/i2c_controller.v(77[47:62])
    defparam i3_4_lut_4_lut.LUT_INIT = 16'h001a;
    SB_LUT4 i2_3_lut_4_lut (.I0(\state[0] ), .I1(\state[1] ), .I2(\state[2] ), 
            .I3(\state[3] ), .O(n11));   // verilog/i2c_controller.v(77[27:43])
    defparam i2_3_lut_4_lut.LUT_INIT = 16'hfdff;
    SB_LUT4 i1_2_lut_3_lut (.I0(enable), .I1(\state_7__N_4251[0] ), .I2(enable_slow_N_4354), 
            .I3(GND_net), .O(n28594));
    defparam i1_2_lut_3_lut.LUT_INIT = 16'heaea;
    
endmodule
//
// Verilog Description of module pwm
//

module pwm (pwm_out, clk32MHz, GND_net, pwm_setpoint, VCC_net) /* synthesis syn_module_defined=1 */ ;
    output pwm_out;
    input clk32MHz;
    input GND_net;
    input [23:0]pwm_setpoint;
    input VCC_net;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    
    wire pwm_out_N_821;
    wire [23:0]pwm_counter;   // verilog/pwm.v(11[19:30])
    
    wire n45276, n14, n13, n8, n10, pwm_counter_23__N_819, n17, 
        n19, n21, n9, n49679, n27, n15, n13_adj_4571, n11, n49673, 
        n12, n35, n30, n49690, n49996;
    wire [23:0]n101;
    
    wire n49992, n25, n23, n50370, n31, n29, n50188, n37, n33, 
        n50420, n6, n50292, n50293, n16, n45, n24, n43, n49658, 
        n8_adj_4572, n49655, n50232, n49752, n4, n50288, n50289, 
        n49669, n10_adj_4573, n49667, n50378, n49754, n50456, n50457, 
        n39, n50445, n41, n49660, n50388, n49760, n50390, n39367, 
        n39366, n39365, n39364, n39363, n39362, n39361, n39360, 
        n39359, n39358, n39357, n39356, n39355, n39354, n39353, 
        n39352, n39351, n39350, n39349, n39348, n39347, n39346, 
        n39345;
    
    SB_DFF pwm_out_12 (.Q(pwm_out), .C(clk32MHz), .D(pwm_out_N_821));   // verilog/pwm.v(16[12] 26[6])
    SB_LUT4 i2_3_lut (.I0(pwm_counter[6]), .I1(pwm_counter[8]), .I2(pwm_counter[7]), 
            .I3(GND_net), .O(n45276));
    defparam i2_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i6_4_lut (.I0(pwm_counter[17]), .I1(pwm_counter[19]), .I2(pwm_counter[16]), 
            .I3(pwm_counter[14]), .O(n14));
    defparam i6_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i5_4_lut (.I0(pwm_counter[11]), .I1(pwm_counter[18]), .I2(pwm_counter[22]), 
            .I3(pwm_counter[15]), .O(n13));
    defparam i5_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_4_lut (.I0(n45276), .I1(pwm_counter[13]), .I2(pwm_counter[10]), 
            .I3(pwm_counter[9]), .O(n8));
    defparam i2_4_lut.LUT_INIT = 16'heccc;
    SB_LUT4 i4_4_lut (.I0(pwm_counter[21]), .I1(n8), .I2(n13), .I3(n14), 
            .O(n10));
    defparam i4_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i35619_4_lut (.I0(pwm_counter[23]), .I1(pwm_counter[12]), .I2(n10), 
            .I3(pwm_counter[20]), .O(pwm_counter_23__N_819));   // verilog/pwm.v(18[8:40])
    defparam i35619_4_lut.LUT_INIT = 16'h5554;
    SB_LUT4 duty_23__I_0_i17_2_lut (.I0(pwm_counter[8]), .I1(pwm_setpoint[8]), 
            .I2(GND_net), .I3(GND_net), .O(n17));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i19_2_lut (.I0(pwm_counter[9]), .I1(pwm_setpoint[9]), 
            .I2(GND_net), .I3(GND_net), .O(n19));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i21_2_lut (.I0(pwm_counter[10]), .I1(pwm_setpoint[10]), 
            .I2(GND_net), .I3(GND_net), .O(n21));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i34092_4_lut (.I0(n21), .I1(n19), .I2(n17), .I3(n9), .O(n49679));
    defparam i34092_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i34086_4_lut (.I0(n27), .I1(n15), .I2(n13_adj_4571), .I3(n11), 
            .O(n49673));
    defparam i34086_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 duty_23__I_0_i30_3_lut (.I0(n12), .I1(pwm_setpoint[17]), .I2(n35), 
            .I3(GND_net), .O(n30));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34408_4_lut (.I0(n13_adj_4571), .I1(n11), .I2(n9), .I3(n49690), 
            .O(n49996));
    defparam i34408_4_lut.LUT_INIT = 16'heeef;
    SB_DFFSR pwm_counter_2246__i23 (.Q(pwm_counter[23]), .C(clk32MHz), .D(n101[23]), 
            .R(pwm_counter_23__N_819));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_2246__i22 (.Q(pwm_counter[22]), .C(clk32MHz), .D(n101[22]), 
            .R(pwm_counter_23__N_819));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_2246__i21 (.Q(pwm_counter[21]), .C(clk32MHz), .D(n101[21]), 
            .R(pwm_counter_23__N_819));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_2246__i20 (.Q(pwm_counter[20]), .C(clk32MHz), .D(n101[20]), 
            .R(pwm_counter_23__N_819));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_2246__i19 (.Q(pwm_counter[19]), .C(clk32MHz), .D(n101[19]), 
            .R(pwm_counter_23__N_819));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_2246__i18 (.Q(pwm_counter[18]), .C(clk32MHz), .D(n101[18]), 
            .R(pwm_counter_23__N_819));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_2246__i17 (.Q(pwm_counter[17]), .C(clk32MHz), .D(n101[17]), 
            .R(pwm_counter_23__N_819));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_2246__i16 (.Q(pwm_counter[16]), .C(clk32MHz), .D(n101[16]), 
            .R(pwm_counter_23__N_819));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_2246__i15 (.Q(pwm_counter[15]), .C(clk32MHz), .D(n101[15]), 
            .R(pwm_counter_23__N_819));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_2246__i14 (.Q(pwm_counter[14]), .C(clk32MHz), .D(n101[14]), 
            .R(pwm_counter_23__N_819));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_2246__i13 (.Q(pwm_counter[13]), .C(clk32MHz), .D(n101[13]), 
            .R(pwm_counter_23__N_819));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_2246__i12 (.Q(pwm_counter[12]), .C(clk32MHz), .D(n101[12]), 
            .R(pwm_counter_23__N_819));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_2246__i11 (.Q(pwm_counter[11]), .C(clk32MHz), .D(n101[11]), 
            .R(pwm_counter_23__N_819));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_2246__i10 (.Q(pwm_counter[10]), .C(clk32MHz), .D(n101[10]), 
            .R(pwm_counter_23__N_819));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_2246__i9 (.Q(pwm_counter[9]), .C(clk32MHz), .D(n101[9]), 
            .R(pwm_counter_23__N_819));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_2246__i8 (.Q(pwm_counter[8]), .C(clk32MHz), .D(n101[8]), 
            .R(pwm_counter_23__N_819));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_2246__i7 (.Q(pwm_counter[7]), .C(clk32MHz), .D(n101[7]), 
            .R(pwm_counter_23__N_819));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_2246__i6 (.Q(pwm_counter[6]), .C(clk32MHz), .D(n101[6]), 
            .R(pwm_counter_23__N_819));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_2246__i5 (.Q(pwm_counter[5]), .C(clk32MHz), .D(n101[5]), 
            .R(pwm_counter_23__N_819));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_2246__i4 (.Q(pwm_counter[4]), .C(clk32MHz), .D(n101[4]), 
            .R(pwm_counter_23__N_819));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_2246__i3 (.Q(pwm_counter[3]), .C(clk32MHz), .D(n101[3]), 
            .R(pwm_counter_23__N_819));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_2246__i2 (.Q(pwm_counter[2]), .C(clk32MHz), .D(n101[2]), 
            .R(pwm_counter_23__N_819));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_2246__i1 (.Q(pwm_counter[1]), .C(clk32MHz), .D(n101[1]), 
            .R(pwm_counter_23__N_819));   // verilog/pwm.v(17[20:33])
    SB_LUT4 i34404_4_lut (.I0(n19), .I1(n17), .I2(n15), .I3(n49996), 
            .O(n49992));
    defparam i34404_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i34782_4_lut (.I0(n25), .I1(n23), .I2(n21), .I3(n49992), 
            .O(n50370));
    defparam i34782_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i34600_4_lut (.I0(n31), .I1(n29), .I2(n27), .I3(n50370), 
            .O(n50188));
    defparam i34600_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i34832_4_lut (.I0(n37), .I1(n35), .I2(n33), .I3(n50188), 
            .O(n50420));
    defparam i34832_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i34704_3_lut (.I0(n6), .I1(pwm_setpoint[10]), .I2(n21), .I3(GND_net), 
            .O(n50292));   // verilog/pwm.v(21[8:24])
    defparam i34704_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34705_3_lut (.I0(n50292), .I1(pwm_setpoint[11]), .I2(n23), 
            .I3(GND_net), .O(n50293));   // verilog/pwm.v(21[8:24])
    defparam i34705_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i24_3_lut (.I0(n16), .I1(pwm_setpoint[22]), .I2(n45), 
            .I3(GND_net), .O(n24));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34071_4_lut (.I0(n43), .I1(n25), .I2(n23), .I3(n49679), 
            .O(n49658));
    defparam i34071_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i34644_4_lut (.I0(n24), .I1(n8_adj_4572), .I2(n45), .I3(n49655), 
            .O(n50232));   // verilog/pwm.v(21[8:24])
    defparam i34644_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i34164_3_lut (.I0(n50293), .I1(pwm_setpoint[12]), .I2(n25), 
            .I3(GND_net), .O(n49752));   // verilog/pwm.v(21[8:24])
    defparam i34164_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i4_4_lut (.I0(pwm_counter[0]), .I1(pwm_setpoint[1]), 
            .I2(pwm_counter[1]), .I3(pwm_setpoint[0]), .O(n4));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i4_4_lut.LUT_INIT = 16'h4d0c;
    SB_LUT4 i34700_3_lut (.I0(n4), .I1(pwm_setpoint[13]), .I2(n27), .I3(GND_net), 
            .O(n50288));   // verilog/pwm.v(21[8:24])
    defparam i34700_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34701_3_lut (.I0(n50288), .I1(pwm_setpoint[14]), .I2(n29), 
            .I3(GND_net), .O(n50289));   // verilog/pwm.v(21[8:24])
    defparam i34701_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34082_4_lut (.I0(n33), .I1(n31), .I2(n29), .I3(n49673), 
            .O(n49669));
    defparam i34082_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i34790_4_lut (.I0(n30), .I1(n10_adj_4573), .I2(n35), .I3(n49667), 
            .O(n50378));   // verilog/pwm.v(21[8:24])
    defparam i34790_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i34166_3_lut (.I0(n50289), .I1(pwm_setpoint[15]), .I2(n31), 
            .I3(GND_net), .O(n49754));   // verilog/pwm.v(21[8:24])
    defparam i34166_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34868_4_lut (.I0(n49754), .I1(n50378), .I2(n35), .I3(n49669), 
            .O(n50456));   // verilog/pwm.v(21[8:24])
    defparam i34868_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i34869_3_lut (.I0(n50456), .I1(pwm_setpoint[18]), .I2(n37), 
            .I3(GND_net), .O(n50457));   // verilog/pwm.v(21[8:24])
    defparam i34869_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34857_3_lut (.I0(n50457), .I1(pwm_setpoint[19]), .I2(n39), 
            .I3(GND_net), .O(n50445));   // verilog/pwm.v(21[8:24])
    defparam i34857_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34073_4_lut (.I0(n43), .I1(n41), .I2(n39), .I3(n50420), 
            .O(n49660));
    defparam i34073_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i34800_4_lut (.I0(n49752), .I1(n50232), .I2(n45), .I3(n49658), 
            .O(n50388));   // verilog/pwm.v(21[8:24])
    defparam i34800_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i34172_3_lut (.I0(n50445), .I1(pwm_setpoint[20]), .I2(n41), 
            .I3(GND_net), .O(n49760));   // verilog/pwm.v(21[8:24])
    defparam i34172_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34802_4_lut (.I0(n49760), .I1(n50388), .I2(n45), .I3(n49660), 
            .O(n50390));   // verilog/pwm.v(21[8:24])
    defparam i34802_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i34803_3_lut (.I0(n50390), .I1(pwm_counter[23]), .I2(pwm_setpoint[23]), 
            .I3(GND_net), .O(pwm_out_N_821));   // verilog/pwm.v(21[8:24])
    defparam i34803_3_lut.LUT_INIT = 16'h8e8e;
    SB_DFFSR pwm_counter_2246__i0 (.Q(pwm_counter[0]), .C(clk32MHz), .D(n101[0]), 
            .R(pwm_counter_23__N_819));   // verilog/pwm.v(17[20:33])
    SB_LUT4 pwm_counter_2246_add_4_25_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[23]), 
            .I3(n39367), .O(n101[23])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2246_add_4_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 pwm_counter_2246_add_4_24_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[22]), 
            .I3(n39366), .O(n101[22])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2246_add_4_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_2246_add_4_24 (.CI(n39366), .I0(GND_net), .I1(pwm_counter[22]), 
            .CO(n39367));
    SB_LUT4 pwm_counter_2246_add_4_23_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[21]), 
            .I3(n39365), .O(n101[21])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2246_add_4_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_2246_add_4_23 (.CI(n39365), .I0(GND_net), .I1(pwm_counter[21]), 
            .CO(n39366));
    SB_LUT4 pwm_counter_2246_add_4_22_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[20]), 
            .I3(n39364), .O(n101[20])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2246_add_4_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_2246_add_4_22 (.CI(n39364), .I0(GND_net), .I1(pwm_counter[20]), 
            .CO(n39365));
    SB_LUT4 pwm_counter_2246_add_4_21_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[19]), 
            .I3(n39363), .O(n101[19])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2246_add_4_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_2246_add_4_21 (.CI(n39363), .I0(GND_net), .I1(pwm_counter[19]), 
            .CO(n39364));
    SB_LUT4 pwm_counter_2246_add_4_20_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[18]), 
            .I3(n39362), .O(n101[18])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2246_add_4_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_2246_add_4_20 (.CI(n39362), .I0(GND_net), .I1(pwm_counter[18]), 
            .CO(n39363));
    SB_LUT4 pwm_counter_2246_add_4_19_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[17]), 
            .I3(n39361), .O(n101[17])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2246_add_4_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_2246_add_4_19 (.CI(n39361), .I0(GND_net), .I1(pwm_counter[17]), 
            .CO(n39362));
    SB_LUT4 pwm_counter_2246_add_4_18_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[16]), 
            .I3(n39360), .O(n101[16])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2246_add_4_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_2246_add_4_18 (.CI(n39360), .I0(GND_net), .I1(pwm_counter[16]), 
            .CO(n39361));
    SB_LUT4 pwm_counter_2246_add_4_17_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[15]), 
            .I3(n39359), .O(n101[15])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2246_add_4_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_2246_add_4_17 (.CI(n39359), .I0(GND_net), .I1(pwm_counter[15]), 
            .CO(n39360));
    SB_LUT4 pwm_counter_2246_add_4_16_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[14]), 
            .I3(n39358), .O(n101[14])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2246_add_4_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_2246_add_4_16 (.CI(n39358), .I0(GND_net), .I1(pwm_counter[14]), 
            .CO(n39359));
    SB_LUT4 pwm_counter_2246_add_4_15_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[13]), 
            .I3(n39357), .O(n101[13])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2246_add_4_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_2246_add_4_15 (.CI(n39357), .I0(GND_net), .I1(pwm_counter[13]), 
            .CO(n39358));
    SB_LUT4 pwm_counter_2246_add_4_14_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[12]), 
            .I3(n39356), .O(n101[12])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2246_add_4_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_2246_add_4_14 (.CI(n39356), .I0(GND_net), .I1(pwm_counter[12]), 
            .CO(n39357));
    SB_LUT4 pwm_counter_2246_add_4_13_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[11]), 
            .I3(n39355), .O(n101[11])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2246_add_4_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_2246_add_4_13 (.CI(n39355), .I0(GND_net), .I1(pwm_counter[11]), 
            .CO(n39356));
    SB_LUT4 pwm_counter_2246_add_4_12_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[10]), 
            .I3(n39354), .O(n101[10])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2246_add_4_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_2246_add_4_12 (.CI(n39354), .I0(GND_net), .I1(pwm_counter[10]), 
            .CO(n39355));
    SB_LUT4 pwm_counter_2246_add_4_11_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[9]), 
            .I3(n39353), .O(n101[9])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2246_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_2246_add_4_11 (.CI(n39353), .I0(GND_net), .I1(pwm_counter[9]), 
            .CO(n39354));
    SB_LUT4 pwm_counter_2246_add_4_10_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[8]), 
            .I3(n39352), .O(n101[8])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2246_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_2246_add_4_10 (.CI(n39352), .I0(GND_net), .I1(pwm_counter[8]), 
            .CO(n39353));
    SB_LUT4 pwm_counter_2246_add_4_9_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[7]), 
            .I3(n39351), .O(n101[7])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2246_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_2246_add_4_9 (.CI(n39351), .I0(GND_net), .I1(pwm_counter[7]), 
            .CO(n39352));
    SB_LUT4 pwm_counter_2246_add_4_8_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[6]), 
            .I3(n39350), .O(n101[6])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2246_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_2246_add_4_8 (.CI(n39350), .I0(GND_net), .I1(pwm_counter[6]), 
            .CO(n39351));
    SB_LUT4 pwm_counter_2246_add_4_7_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[5]), 
            .I3(n39349), .O(n101[5])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2246_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_2246_add_4_7 (.CI(n39349), .I0(GND_net), .I1(pwm_counter[5]), 
            .CO(n39350));
    SB_LUT4 pwm_counter_2246_add_4_6_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[4]), 
            .I3(n39348), .O(n101[4])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2246_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_2246_add_4_6 (.CI(n39348), .I0(GND_net), .I1(pwm_counter[4]), 
            .CO(n39349));
    SB_LUT4 pwm_counter_2246_add_4_5_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[3]), 
            .I3(n39347), .O(n101[3])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2246_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_2246_add_4_5 (.CI(n39347), .I0(GND_net), .I1(pwm_counter[3]), 
            .CO(n39348));
    SB_LUT4 pwm_counter_2246_add_4_4_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[2]), 
            .I3(n39346), .O(n101[2])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2246_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_2246_add_4_4 (.CI(n39346), .I0(GND_net), .I1(pwm_counter[2]), 
            .CO(n39347));
    SB_LUT4 pwm_counter_2246_add_4_3_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[1]), 
            .I3(n39345), .O(n101[1])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2246_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_2246_add_4_3 (.CI(n39345), .I0(GND_net), .I1(pwm_counter[1]), 
            .CO(n39346));
    SB_LUT4 pwm_counter_2246_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[0]), 
            .I3(VCC_net), .O(n101[0])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2246_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_2246_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(pwm_counter[0]), 
            .CO(n39345));
    SB_LUT4 i34103_3_lut_4_lut (.I0(pwm_counter[3]), .I1(pwm_setpoint[3]), 
            .I2(pwm_setpoint[2]), .I3(pwm_counter[2]), .O(n49690));   // verilog/pwm.v(21[8:24])
    defparam i34103_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 duty_23__I_0_i6_3_lut_3_lut (.I0(pwm_counter[3]), .I1(pwm_setpoint[3]), 
            .I2(pwm_setpoint[2]), .I3(GND_net), .O(n6));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 duty_23__I_0_i41_2_lut (.I0(pwm_counter[20]), .I1(pwm_setpoint[20]), 
            .I2(GND_net), .I3(GND_net), .O(n41));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i39_2_lut (.I0(pwm_counter[19]), .I1(pwm_setpoint[19]), 
            .I2(GND_net), .I3(GND_net), .O(n39));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i45_2_lut (.I0(pwm_counter[22]), .I1(pwm_setpoint[22]), 
            .I2(GND_net), .I3(GND_net), .O(n45));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i45_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i43_2_lut (.I0(pwm_counter[21]), .I1(pwm_setpoint[21]), 
            .I2(GND_net), .I3(GND_net), .O(n43));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i37_2_lut (.I0(pwm_counter[18]), .I1(pwm_setpoint[18]), 
            .I2(GND_net), .I3(GND_net), .O(n37));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i29_2_lut (.I0(pwm_counter[14]), .I1(pwm_setpoint[14]), 
            .I2(GND_net), .I3(GND_net), .O(n29));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i8_3_lut_3_lut (.I0(pwm_setpoint[4]), .I1(pwm_setpoint[8]), 
            .I2(pwm_counter[8]), .I3(GND_net), .O(n8_adj_4572));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i8_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 duty_23__I_0_i31_2_lut (.I0(pwm_counter[15]), .I1(pwm_setpoint[15]), 
            .I2(GND_net), .I3(GND_net), .O(n31));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i34068_2_lut_4_lut (.I0(pwm_counter[21]), .I1(pwm_setpoint[21]), 
            .I2(pwm_counter[9]), .I3(pwm_setpoint[9]), .O(n49655));
    defparam i34068_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 duty_23__I_0_i16_3_lut_3_lut (.I0(pwm_setpoint[9]), .I1(pwm_setpoint[21]), 
            .I2(pwm_counter[21]), .I3(GND_net), .O(n16));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i16_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 duty_23__I_0_i23_2_lut (.I0(pwm_counter[11]), .I1(pwm_setpoint[11]), 
            .I2(GND_net), .I3(GND_net), .O(n23));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i25_2_lut (.I0(pwm_counter[12]), .I1(pwm_setpoint[12]), 
            .I2(GND_net), .I3(GND_net), .O(n25));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i10_3_lut_3_lut (.I0(pwm_setpoint[5]), .I1(pwm_setpoint[6]), 
            .I2(pwm_counter[6]), .I3(GND_net), .O(n10_adj_4573));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i10_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i34080_2_lut_4_lut (.I0(pwm_counter[16]), .I1(pwm_setpoint[16]), 
            .I2(pwm_counter[7]), .I3(pwm_setpoint[7]), .O(n49667));
    defparam i34080_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 duty_23__I_0_i12_3_lut_3_lut (.I0(pwm_setpoint[7]), .I1(pwm_setpoint[16]), 
            .I2(pwm_counter[16]), .I3(GND_net), .O(n12));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i12_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 duty_23__I_0_i35_2_lut (.I0(pwm_counter[17]), .I1(pwm_setpoint[17]), 
            .I2(GND_net), .I3(GND_net), .O(n35));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i33_2_lut (.I0(pwm_counter[16]), .I1(pwm_setpoint[16]), 
            .I2(GND_net), .I3(GND_net), .O(n33));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i11_2_lut (.I0(pwm_counter[5]), .I1(pwm_setpoint[5]), 
            .I2(GND_net), .I3(GND_net), .O(n11));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i13_2_lut (.I0(pwm_counter[6]), .I1(pwm_setpoint[6]), 
            .I2(GND_net), .I3(GND_net), .O(n13_adj_4571));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i15_2_lut (.I0(pwm_counter[7]), .I1(pwm_setpoint[7]), 
            .I2(GND_net), .I3(GND_net), .O(n15));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i27_2_lut (.I0(pwm_counter[13]), .I1(pwm_setpoint[13]), 
            .I2(GND_net), .I3(GND_net), .O(n27));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i9_2_lut (.I0(pwm_counter[4]), .I1(pwm_setpoint[4]), 
            .I2(GND_net), .I3(GND_net), .O(n9));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i9_2_lut.LUT_INIT = 16'h6666;
    
endmodule
