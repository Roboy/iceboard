-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2017.08.27940

-- Build Date:         Sep 12 2017 08:26:01

-- File Generated:     Jan 29 2020 12:28:04

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "TinyFPGA_B" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of TinyFPGA_B
entity TinyFPGA_B is
port (
    USBPU : out std_logic;
    TX : out std_logic;
    SDA : inout std_logic;
    SCL : inout std_logic;
    RX : in std_logic;
    NEOPXL : out std_logic;
    LED : out std_logic;
    INLC : out std_logic;
    INLB : out std_logic;
    INLA : out std_logic;
    INHC : out std_logic;
    INHB : out std_logic;
    INHA : out std_logic;
    HALL3 : in std_logic;
    HALL2 : in std_logic;
    HALL1 : in std_logic;
    FAULT_N : in std_logic;
    ENCODER1_B : in std_logic;
    ENCODER1_A : in std_logic;
    ENCODER0_B : in std_logic;
    ENCODER0_A : in std_logic;
    DE : out std_logic;
    CS_MISO : in std_logic;
    CS_CLK : out std_logic;
    CS : out std_logic;
    CLK : in std_logic);
end TinyFPGA_B;

-- Architecture of TinyFPGA_B
-- View name is \INTERFACE\
architecture \INTERFACE\ of TinyFPGA_B is

signal \N__28245\ : std_logic;
signal \N__28244\ : std_logic;
signal \N__28243\ : std_logic;
signal \N__28236\ : std_logic;
signal \N__28235\ : std_logic;
signal \N__28234\ : std_logic;
signal \N__28227\ : std_logic;
signal \N__28226\ : std_logic;
signal \N__28225\ : std_logic;
signal \N__28218\ : std_logic;
signal \N__28217\ : std_logic;
signal \N__28216\ : std_logic;
signal \N__28209\ : std_logic;
signal \N__28208\ : std_logic;
signal \N__28207\ : std_logic;
signal \N__28200\ : std_logic;
signal \N__28199\ : std_logic;
signal \N__28198\ : std_logic;
signal \N__28191\ : std_logic;
signal \N__28190\ : std_logic;
signal \N__28189\ : std_logic;
signal \N__28182\ : std_logic;
signal \N__28181\ : std_logic;
signal \N__28180\ : std_logic;
signal \N__28173\ : std_logic;
signal \N__28172\ : std_logic;
signal \N__28171\ : std_logic;
signal \N__28164\ : std_logic;
signal \N__28163\ : std_logic;
signal \N__28162\ : std_logic;
signal \N__28155\ : std_logic;
signal \N__28154\ : std_logic;
signal \N__28153\ : std_logic;
signal \N__28146\ : std_logic;
signal \N__28145\ : std_logic;
signal \N__28144\ : std_logic;
signal \N__28137\ : std_logic;
signal \N__28136\ : std_logic;
signal \N__28135\ : std_logic;
signal \N__28128\ : std_logic;
signal \N__28127\ : std_logic;
signal \N__28126\ : std_logic;
signal \N__28119\ : std_logic;
signal \N__28118\ : std_logic;
signal \N__28117\ : std_logic;
signal \N__28110\ : std_logic;
signal \N__28109\ : std_logic;
signal \N__28108\ : std_logic;
signal \N__28091\ : std_logic;
signal \N__28088\ : std_logic;
signal \N__28085\ : std_logic;
signal \N__28082\ : std_logic;
signal \N__28079\ : std_logic;
signal \N__28076\ : std_logic;
signal \N__28073\ : std_logic;
signal \N__28072\ : std_logic;
signal \N__28069\ : std_logic;
signal \N__28066\ : std_logic;
signal \N__28063\ : std_logic;
signal \N__28062\ : std_logic;
signal \N__28057\ : std_logic;
signal \N__28054\ : std_logic;
signal \N__28049\ : std_logic;
signal \N__28046\ : std_logic;
signal \N__28043\ : std_logic;
signal \N__28040\ : std_logic;
signal \N__28037\ : std_logic;
signal \N__28034\ : std_logic;
signal \N__28031\ : std_logic;
signal \N__28030\ : std_logic;
signal \N__28027\ : std_logic;
signal \N__28026\ : std_logic;
signal \N__28023\ : std_logic;
signal \N__28020\ : std_logic;
signal \N__28015\ : std_logic;
signal \N__28010\ : std_logic;
signal \N__28007\ : std_logic;
signal \N__28004\ : std_logic;
signal \N__28001\ : std_logic;
signal \N__27998\ : std_logic;
signal \N__27995\ : std_logic;
signal \N__27994\ : std_logic;
signal \N__27991\ : std_logic;
signal \N__27988\ : std_logic;
signal \N__27987\ : std_logic;
signal \N__27984\ : std_logic;
signal \N__27981\ : std_logic;
signal \N__27978\ : std_logic;
signal \N__27975\ : std_logic;
signal \N__27970\ : std_logic;
signal \N__27965\ : std_logic;
signal \N__27962\ : std_logic;
signal \N__27959\ : std_logic;
signal \N__27956\ : std_logic;
signal \N__27953\ : std_logic;
signal \N__27950\ : std_logic;
signal \N__27947\ : std_logic;
signal \N__27944\ : std_logic;
signal \N__27943\ : std_logic;
signal \N__27940\ : std_logic;
signal \N__27937\ : std_logic;
signal \N__27934\ : std_logic;
signal \N__27931\ : std_logic;
signal \N__27928\ : std_logic;
signal \N__27925\ : std_logic;
signal \N__27920\ : std_logic;
signal \N__27919\ : std_logic;
signal \N__27916\ : std_logic;
signal \N__27915\ : std_logic;
signal \N__27912\ : std_logic;
signal \N__27911\ : std_logic;
signal \N__27910\ : std_logic;
signal \N__27909\ : std_logic;
signal \N__27908\ : std_logic;
signal \N__27907\ : std_logic;
signal \N__27904\ : std_logic;
signal \N__27903\ : std_logic;
signal \N__27902\ : std_logic;
signal \N__27899\ : std_logic;
signal \N__27894\ : std_logic;
signal \N__27891\ : std_logic;
signal \N__27890\ : std_logic;
signal \N__27889\ : std_logic;
signal \N__27888\ : std_logic;
signal \N__27887\ : std_logic;
signal \N__27886\ : std_logic;
signal \N__27883\ : std_logic;
signal \N__27882\ : std_logic;
signal \N__27881\ : std_logic;
signal \N__27878\ : std_logic;
signal \N__27875\ : std_logic;
signal \N__27874\ : std_logic;
signal \N__27871\ : std_logic;
signal \N__27864\ : std_logic;
signal \N__27861\ : std_logic;
signal \N__27856\ : std_logic;
signal \N__27851\ : std_logic;
signal \N__27848\ : std_logic;
signal \N__27839\ : std_logic;
signal \N__27832\ : std_logic;
signal \N__27829\ : std_logic;
signal \N__27824\ : std_logic;
signal \N__27809\ : std_logic;
signal \N__27806\ : std_logic;
signal \N__27805\ : std_logic;
signal \N__27802\ : std_logic;
signal \N__27799\ : std_logic;
signal \N__27794\ : std_logic;
signal \N__27791\ : std_logic;
signal \N__27788\ : std_logic;
signal \N__27787\ : std_logic;
signal \N__27786\ : std_logic;
signal \N__27785\ : std_logic;
signal \N__27784\ : std_logic;
signal \N__27783\ : std_logic;
signal \N__27782\ : std_logic;
signal \N__27781\ : std_logic;
signal \N__27780\ : std_logic;
signal \N__27779\ : std_logic;
signal \N__27778\ : std_logic;
signal \N__27777\ : std_logic;
signal \N__27776\ : std_logic;
signal \N__27775\ : std_logic;
signal \N__27774\ : std_logic;
signal \N__27773\ : std_logic;
signal \N__27770\ : std_logic;
signal \N__27769\ : std_logic;
signal \N__27768\ : std_logic;
signal \N__27767\ : std_logic;
signal \N__27766\ : std_logic;
signal \N__27765\ : std_logic;
signal \N__27762\ : std_logic;
signal \N__27761\ : std_logic;
signal \N__27760\ : std_logic;
signal \N__27757\ : std_logic;
signal \N__27756\ : std_logic;
signal \N__27755\ : std_logic;
signal \N__27754\ : std_logic;
signal \N__27753\ : std_logic;
signal \N__27752\ : std_logic;
signal \N__27751\ : std_logic;
signal \N__27750\ : std_logic;
signal \N__27749\ : std_logic;
signal \N__27748\ : std_logic;
signal \N__27747\ : std_logic;
signal \N__27746\ : std_logic;
signal \N__27745\ : std_logic;
signal \N__27744\ : std_logic;
signal \N__27743\ : std_logic;
signal \N__27742\ : std_logic;
signal \N__27739\ : std_logic;
signal \N__27736\ : std_logic;
signal \N__27733\ : std_logic;
signal \N__27732\ : std_logic;
signal \N__27731\ : std_logic;
signal \N__27730\ : std_logic;
signal \N__27729\ : std_logic;
signal \N__27728\ : std_logic;
signal \N__27727\ : std_logic;
signal \N__27726\ : std_logic;
signal \N__27725\ : std_logic;
signal \N__27724\ : std_logic;
signal \N__27723\ : std_logic;
signal \N__27722\ : std_logic;
signal \N__27721\ : std_logic;
signal \N__27716\ : std_logic;
signal \N__27715\ : std_logic;
signal \N__27714\ : std_logic;
signal \N__27713\ : std_logic;
signal \N__27712\ : std_logic;
signal \N__27711\ : std_logic;
signal \N__27710\ : std_logic;
signal \N__27709\ : std_logic;
signal \N__27708\ : std_logic;
signal \N__27707\ : std_logic;
signal \N__27706\ : std_logic;
signal \N__27701\ : std_logic;
signal \N__27694\ : std_logic;
signal \N__27683\ : std_logic;
signal \N__27680\ : std_logic;
signal \N__27677\ : std_logic;
signal \N__27674\ : std_logic;
signal \N__27671\ : std_logic;
signal \N__27670\ : std_logic;
signal \N__27659\ : std_logic;
signal \N__27654\ : std_logic;
signal \N__27653\ : std_logic;
signal \N__27650\ : std_logic;
signal \N__27649\ : std_logic;
signal \N__27648\ : std_logic;
signal \N__27647\ : std_logic;
signal \N__27644\ : std_logic;
signal \N__27643\ : std_logic;
signal \N__27642\ : std_logic;
signal \N__27641\ : std_logic;
signal \N__27638\ : std_logic;
signal \N__27635\ : std_logic;
signal \N__27630\ : std_logic;
signal \N__27629\ : std_logic;
signal \N__27628\ : std_logic;
signal \N__27627\ : std_logic;
signal \N__27624\ : std_logic;
signal \N__27621\ : std_logic;
signal \N__27620\ : std_logic;
signal \N__27617\ : std_logic;
signal \N__27614\ : std_logic;
signal \N__27613\ : std_logic;
signal \N__27612\ : std_logic;
signal \N__27611\ : std_logic;
signal \N__27608\ : std_logic;
signal \N__27607\ : std_logic;
signal \N__27606\ : std_logic;
signal \N__27605\ : std_logic;
signal \N__27604\ : std_logic;
signal \N__27599\ : std_logic;
signal \N__27596\ : std_logic;
signal \N__27591\ : std_logic;
signal \N__27590\ : std_logic;
signal \N__27589\ : std_logic;
signal \N__27588\ : std_logic;
signal \N__27587\ : std_logic;
signal \N__27586\ : std_logic;
signal \N__27583\ : std_logic;
signal \N__27582\ : std_logic;
signal \N__27581\ : std_logic;
signal \N__27578\ : std_logic;
signal \N__27575\ : std_logic;
signal \N__27570\ : std_logic;
signal \N__27569\ : std_logic;
signal \N__27566\ : std_logic;
signal \N__27565\ : std_logic;
signal \N__27564\ : std_logic;
signal \N__27561\ : std_logic;
signal \N__27560\ : std_logic;
signal \N__27557\ : std_logic;
signal \N__27556\ : std_logic;
signal \N__27553\ : std_logic;
signal \N__27550\ : std_logic;
signal \N__27547\ : std_logic;
signal \N__27546\ : std_logic;
signal \N__27545\ : std_logic;
signal \N__27544\ : std_logic;
signal \N__27543\ : std_logic;
signal \N__27542\ : std_logic;
signal \N__27541\ : std_logic;
signal \N__27538\ : std_logic;
signal \N__27529\ : std_logic;
signal \N__27520\ : std_logic;
signal \N__27519\ : std_logic;
signal \N__27518\ : std_logic;
signal \N__27515\ : std_logic;
signal \N__27514\ : std_logic;
signal \N__27513\ : std_logic;
signal \N__27510\ : std_logic;
signal \N__27509\ : std_logic;
signal \N__27504\ : std_logic;
signal \N__27501\ : std_logic;
signal \N__27490\ : std_logic;
signal \N__27485\ : std_logic;
signal \N__27476\ : std_logic;
signal \N__27467\ : std_logic;
signal \N__27460\ : std_logic;
signal \N__27459\ : std_logic;
signal \N__27456\ : std_logic;
signal \N__27453\ : std_logic;
signal \N__27448\ : std_logic;
signal \N__27443\ : std_logic;
signal \N__27436\ : std_logic;
signal \N__27431\ : std_logic;
signal \N__27428\ : std_logic;
signal \N__27423\ : std_logic;
signal \N__27422\ : std_logic;
signal \N__27421\ : std_logic;
signal \N__27418\ : std_logic;
signal \N__27415\ : std_logic;
signal \N__27412\ : std_logic;
signal \N__27411\ : std_logic;
signal \N__27410\ : std_logic;
signal \N__27407\ : std_logic;
signal \N__27402\ : std_logic;
signal \N__27397\ : std_logic;
signal \N__27394\ : std_logic;
signal \N__27393\ : std_logic;
signal \N__27390\ : std_logic;
signal \N__27387\ : std_logic;
signal \N__27386\ : std_logic;
signal \N__27385\ : std_logic;
signal \N__27384\ : std_logic;
signal \N__27383\ : std_logic;
signal \N__27382\ : std_logic;
signal \N__27381\ : std_logic;
signal \N__27378\ : std_logic;
signal \N__27375\ : std_logic;
signal \N__27372\ : std_logic;
signal \N__27371\ : std_logic;
signal \N__27368\ : std_logic;
signal \N__27365\ : std_logic;
signal \N__27362\ : std_logic;
signal \N__27357\ : std_logic;
signal \N__27348\ : std_logic;
signal \N__27345\ : std_logic;
signal \N__27342\ : std_logic;
signal \N__27335\ : std_logic;
signal \N__27334\ : std_logic;
signal \N__27333\ : std_logic;
signal \N__27332\ : std_logic;
signal \N__27331\ : std_logic;
signal \N__27330\ : std_logic;
signal \N__27327\ : std_logic;
signal \N__27326\ : std_logic;
signal \N__27325\ : std_logic;
signal \N__27322\ : std_logic;
signal \N__27319\ : std_logic;
signal \N__27318\ : std_logic;
signal \N__27315\ : std_logic;
signal \N__27312\ : std_logic;
signal \N__27311\ : std_logic;
signal \N__27310\ : std_logic;
signal \N__27307\ : std_logic;
signal \N__27306\ : std_logic;
signal \N__27305\ : std_logic;
signal \N__27304\ : std_logic;
signal \N__27303\ : std_logic;
signal \N__27302\ : std_logic;
signal \N__27295\ : std_logic;
signal \N__27290\ : std_logic;
signal \N__27279\ : std_logic;
signal \N__27272\ : std_logic;
signal \N__27263\ : std_logic;
signal \N__27260\ : std_logic;
signal \N__27255\ : std_logic;
signal \N__27252\ : std_logic;
signal \N__27247\ : std_logic;
signal \N__27240\ : std_logic;
signal \N__27235\ : std_logic;
signal \N__27226\ : std_logic;
signal \N__27223\ : std_logic;
signal \N__27218\ : std_logic;
signal \N__27215\ : std_logic;
signal \N__27206\ : std_logic;
signal \N__27205\ : std_logic;
signal \N__27202\ : std_logic;
signal \N__27199\ : std_logic;
signal \N__27196\ : std_logic;
signal \N__27195\ : std_logic;
signal \N__27194\ : std_logic;
signal \N__27193\ : std_logic;
signal \N__27192\ : std_logic;
signal \N__27191\ : std_logic;
signal \N__27190\ : std_logic;
signal \N__27189\ : std_logic;
signal \N__27188\ : std_logic;
signal \N__27187\ : std_logic;
signal \N__27186\ : std_logic;
signal \N__27185\ : std_logic;
signal \N__27182\ : std_logic;
signal \N__27181\ : std_logic;
signal \N__27180\ : std_logic;
signal \N__27179\ : std_logic;
signal \N__27176\ : std_logic;
signal \N__27175\ : std_logic;
signal \N__27174\ : std_logic;
signal \N__27171\ : std_logic;
signal \N__27166\ : std_logic;
signal \N__27163\ : std_logic;
signal \N__27160\ : std_logic;
signal \N__27155\ : std_logic;
signal \N__27142\ : std_logic;
signal \N__27139\ : std_logic;
signal \N__27136\ : std_logic;
signal \N__27133\ : std_logic;
signal \N__27130\ : std_logic;
signal \N__27127\ : std_logic;
signal \N__27126\ : std_logic;
signal \N__27123\ : std_logic;
signal \N__27118\ : std_logic;
signal \N__27109\ : std_logic;
signal \N__27106\ : std_logic;
signal \N__27103\ : std_logic;
signal \N__27098\ : std_logic;
signal \N__27095\ : std_logic;
signal \N__27092\ : std_logic;
signal \N__27091\ : std_logic;
signal \N__27088\ : std_logic;
signal \N__27085\ : std_logic;
signal \N__27084\ : std_logic;
signal \N__27081\ : std_logic;
signal \N__27080\ : std_logic;
signal \N__27079\ : std_logic;
signal \N__27078\ : std_logic;
signal \N__27077\ : std_logic;
signal \N__27076\ : std_logic;
signal \N__27075\ : std_logic;
signal \N__27074\ : std_logic;
signal \N__27073\ : std_logic;
signal \N__27066\ : std_logic;
signal \N__27059\ : std_logic;
signal \N__27048\ : std_logic;
signal \N__27043\ : std_logic;
signal \N__27036\ : std_logic;
signal \N__27031\ : std_logic;
signal \N__27026\ : std_logic;
signal \N__27025\ : std_logic;
signal \N__27024\ : std_logic;
signal \N__27021\ : std_logic;
signal \N__27018\ : std_logic;
signal \N__27017\ : std_logic;
signal \N__27016\ : std_logic;
signal \N__27013\ : std_logic;
signal \N__27010\ : std_logic;
signal \N__27009\ : std_logic;
signal \N__27008\ : std_logic;
signal \N__27005\ : std_logic;
signal \N__27002\ : std_logic;
signal \N__26999\ : std_logic;
signal \N__26998\ : std_logic;
signal \N__26995\ : std_logic;
signal \N__26992\ : std_logic;
signal \N__26989\ : std_logic;
signal \N__26988\ : std_logic;
signal \N__26987\ : std_logic;
signal \N__26984\ : std_logic;
signal \N__26981\ : std_logic;
signal \N__26978\ : std_logic;
signal \N__26973\ : std_logic;
signal \N__26964\ : std_logic;
signal \N__26957\ : std_logic;
signal \N__26952\ : std_logic;
signal \N__26947\ : std_logic;
signal \N__26938\ : std_logic;
signal \N__26937\ : std_logic;
signal \N__26936\ : std_logic;
signal \N__26933\ : std_logic;
signal \N__26922\ : std_logic;
signal \N__26919\ : std_logic;
signal \N__26904\ : std_logic;
signal \N__26901\ : std_logic;
signal \N__26898\ : std_logic;
signal \N__26895\ : std_logic;
signal \N__26892\ : std_logic;
signal \N__26889\ : std_logic;
signal \N__26886\ : std_logic;
signal \N__26885\ : std_logic;
signal \N__26882\ : std_logic;
signal \N__26881\ : std_logic;
signal \N__26880\ : std_logic;
signal \N__26877\ : std_logic;
signal \N__26870\ : std_logic;
signal \N__26863\ : std_logic;
signal \N__26858\ : std_logic;
signal \N__26849\ : std_logic;
signal \N__26840\ : std_logic;
signal \N__26833\ : std_logic;
signal \N__26822\ : std_logic;
signal \N__26817\ : std_logic;
signal \N__26800\ : std_logic;
signal \N__26795\ : std_logic;
signal \N__26786\ : std_logic;
signal \N__26779\ : std_logic;
signal \N__26768\ : std_logic;
signal \N__26765\ : std_logic;
signal \N__26764\ : std_logic;
signal \N__26761\ : std_logic;
signal \N__26756\ : std_logic;
signal \N__26753\ : std_logic;
signal \N__26740\ : std_logic;
signal \N__26735\ : std_logic;
signal \N__26728\ : std_logic;
signal \N__26725\ : std_logic;
signal \N__26720\ : std_logic;
signal \N__26705\ : std_logic;
signal \N__26704\ : std_logic;
signal \N__26703\ : std_logic;
signal \N__26700\ : std_logic;
signal \N__26697\ : std_logic;
signal \N__26694\ : std_logic;
signal \N__26691\ : std_logic;
signal \N__26684\ : std_logic;
signal \N__26681\ : std_logic;
signal \N__26678\ : std_logic;
signal \N__26675\ : std_logic;
signal \N__26672\ : std_logic;
signal \N__26671\ : std_logic;
signal \N__26668\ : std_logic;
signal \N__26667\ : std_logic;
signal \N__26664\ : std_logic;
signal \N__26661\ : std_logic;
signal \N__26658\ : std_logic;
signal \N__26651\ : std_logic;
signal \N__26648\ : std_logic;
signal \N__26645\ : std_logic;
signal \N__26642\ : std_logic;
signal \N__26639\ : std_logic;
signal \N__26636\ : std_logic;
signal \N__26635\ : std_logic;
signal \N__26634\ : std_logic;
signal \N__26631\ : std_logic;
signal \N__26628\ : std_logic;
signal \N__26625\ : std_logic;
signal \N__26620\ : std_logic;
signal \N__26617\ : std_logic;
signal \N__26614\ : std_logic;
signal \N__26611\ : std_logic;
signal \N__26606\ : std_logic;
signal \N__26603\ : std_logic;
signal \N__26600\ : std_logic;
signal \N__26597\ : std_logic;
signal \N__26594\ : std_logic;
signal \N__26593\ : std_logic;
signal \N__26590\ : std_logic;
signal \N__26587\ : std_logic;
signal \N__26586\ : std_logic;
signal \N__26583\ : std_logic;
signal \N__26580\ : std_logic;
signal \N__26577\ : std_logic;
signal \N__26574\ : std_logic;
signal \N__26571\ : std_logic;
signal \N__26568\ : std_logic;
signal \N__26561\ : std_logic;
signal \N__26558\ : std_logic;
signal \N__26555\ : std_logic;
signal \N__26552\ : std_logic;
signal \N__26549\ : std_logic;
signal \N__26546\ : std_logic;
signal \N__26543\ : std_logic;
signal \N__26540\ : std_logic;
signal \N__26539\ : std_logic;
signal \N__26538\ : std_logic;
signal \N__26535\ : std_logic;
signal \N__26532\ : std_logic;
signal \N__26529\ : std_logic;
signal \N__26522\ : std_logic;
signal \N__26519\ : std_logic;
signal \N__26516\ : std_logic;
signal \N__26513\ : std_logic;
signal \N__26512\ : std_logic;
signal \N__26511\ : std_logic;
signal \N__26508\ : std_logic;
signal \N__26505\ : std_logic;
signal \N__26502\ : std_logic;
signal \N__26499\ : std_logic;
signal \N__26496\ : std_logic;
signal \N__26493\ : std_logic;
signal \N__26490\ : std_logic;
signal \N__26483\ : std_logic;
signal \N__26480\ : std_logic;
signal \N__26477\ : std_logic;
signal \N__26474\ : std_logic;
signal \N__26471\ : std_logic;
signal \N__26468\ : std_logic;
signal \N__26467\ : std_logic;
signal \N__26464\ : std_logic;
signal \N__26461\ : std_logic;
signal \N__26460\ : std_logic;
signal \N__26457\ : std_logic;
signal \N__26454\ : std_logic;
signal \N__26451\ : std_logic;
signal \N__26444\ : std_logic;
signal \N__26441\ : std_logic;
signal \N__26438\ : std_logic;
signal \N__26435\ : std_logic;
signal \N__26432\ : std_logic;
signal \N__26429\ : std_logic;
signal \N__26426\ : std_logic;
signal \N__26423\ : std_logic;
signal \N__26420\ : std_logic;
signal \N__26419\ : std_logic;
signal \N__26418\ : std_logic;
signal \N__26415\ : std_logic;
signal \N__26410\ : std_logic;
signal \N__26407\ : std_logic;
signal \N__26404\ : std_logic;
signal \N__26399\ : std_logic;
signal \N__26396\ : std_logic;
signal \N__26393\ : std_logic;
signal \N__26390\ : std_logic;
signal \N__26387\ : std_logic;
signal \N__26386\ : std_logic;
signal \N__26385\ : std_logic;
signal \N__26382\ : std_logic;
signal \N__26379\ : std_logic;
signal \N__26376\ : std_logic;
signal \N__26369\ : std_logic;
signal \N__26366\ : std_logic;
signal \N__26363\ : std_logic;
signal \N__26360\ : std_logic;
signal \N__26357\ : std_logic;
signal \N__26354\ : std_logic;
signal \N__26351\ : std_logic;
signal \N__26348\ : std_logic;
signal \N__26345\ : std_logic;
signal \N__26342\ : std_logic;
signal \N__26339\ : std_logic;
signal \N__26336\ : std_logic;
signal \N__26335\ : std_logic;
signal \N__26332\ : std_logic;
signal \N__26331\ : std_logic;
signal \N__26328\ : std_logic;
signal \N__26325\ : std_logic;
signal \N__26322\ : std_logic;
signal \N__26319\ : std_logic;
signal \N__26312\ : std_logic;
signal \N__26309\ : std_logic;
signal \N__26306\ : std_logic;
signal \N__26303\ : std_logic;
signal \N__26300\ : std_logic;
signal \N__26297\ : std_logic;
signal \N__26294\ : std_logic;
signal \N__26293\ : std_logic;
signal \N__26290\ : std_logic;
signal \N__26287\ : std_logic;
signal \N__26284\ : std_logic;
signal \N__26283\ : std_logic;
signal \N__26278\ : std_logic;
signal \N__26275\ : std_logic;
signal \N__26272\ : std_logic;
signal \N__26267\ : std_logic;
signal \N__26264\ : std_logic;
signal \N__26261\ : std_logic;
signal \N__26258\ : std_logic;
signal \N__26255\ : std_logic;
signal \N__26252\ : std_logic;
signal \N__26249\ : std_logic;
signal \N__26246\ : std_logic;
signal \N__26245\ : std_logic;
signal \N__26244\ : std_logic;
signal \N__26241\ : std_logic;
signal \N__26238\ : std_logic;
signal \N__26235\ : std_logic;
signal \N__26232\ : std_logic;
signal \N__26229\ : std_logic;
signal \N__26224\ : std_logic;
signal \N__26221\ : std_logic;
signal \N__26218\ : std_logic;
signal \N__26213\ : std_logic;
signal \N__26210\ : std_logic;
signal \N__26207\ : std_logic;
signal \N__26204\ : std_logic;
signal \N__26201\ : std_logic;
signal \N__26198\ : std_logic;
signal \N__26195\ : std_logic;
signal \N__26192\ : std_logic;
signal \N__26191\ : std_logic;
signal \N__26188\ : std_logic;
signal \N__26185\ : std_logic;
signal \N__26184\ : std_logic;
signal \N__26181\ : std_logic;
signal \N__26178\ : std_logic;
signal \N__26175\ : std_logic;
signal \N__26172\ : std_logic;
signal \N__26165\ : std_logic;
signal \N__26162\ : std_logic;
signal \N__26159\ : std_logic;
signal \N__26156\ : std_logic;
signal \N__26153\ : std_logic;
signal \N__26150\ : std_logic;
signal \N__26147\ : std_logic;
signal \N__26146\ : std_logic;
signal \N__26145\ : std_logic;
signal \N__26142\ : std_logic;
signal \N__26139\ : std_logic;
signal \N__26136\ : std_logic;
signal \N__26133\ : std_logic;
signal \N__26130\ : std_logic;
signal \N__26125\ : std_logic;
signal \N__26120\ : std_logic;
signal \N__26117\ : std_logic;
signal \N__26114\ : std_logic;
signal \N__26111\ : std_logic;
signal \N__26108\ : std_logic;
signal \N__26105\ : std_logic;
signal \N__26102\ : std_logic;
signal \N__26099\ : std_logic;
signal \N__26096\ : std_logic;
signal \N__26093\ : std_logic;
signal \N__26092\ : std_logic;
signal \N__26089\ : std_logic;
signal \N__26088\ : std_logic;
signal \N__26085\ : std_logic;
signal \N__26082\ : std_logic;
signal \N__26077\ : std_logic;
signal \N__26074\ : std_logic;
signal \N__26069\ : std_logic;
signal \N__26066\ : std_logic;
signal \N__26063\ : std_logic;
signal \N__26060\ : std_logic;
signal \N__26057\ : std_logic;
signal \N__26056\ : std_logic;
signal \N__26055\ : std_logic;
signal \N__26052\ : std_logic;
signal \N__26049\ : std_logic;
signal \N__26046\ : std_logic;
signal \N__26043\ : std_logic;
signal \N__26040\ : std_logic;
signal \N__26033\ : std_logic;
signal \N__26030\ : std_logic;
signal \N__26027\ : std_logic;
signal \N__26024\ : std_logic;
signal \N__26021\ : std_logic;
signal \N__26018\ : std_logic;
signal \N__26015\ : std_logic;
signal \N__26014\ : std_logic;
signal \N__26011\ : std_logic;
signal \N__26008\ : std_logic;
signal \N__26003\ : std_logic;
signal \N__26000\ : std_logic;
signal \N__25997\ : std_logic;
signal \N__25994\ : std_logic;
signal \N__25993\ : std_logic;
signal \N__25990\ : std_logic;
signal \N__25987\ : std_logic;
signal \N__25984\ : std_logic;
signal \N__25981\ : std_logic;
signal \N__25980\ : std_logic;
signal \N__25975\ : std_logic;
signal \N__25972\ : std_logic;
signal \N__25967\ : std_logic;
signal \N__25964\ : std_logic;
signal \N__25961\ : std_logic;
signal \N__25958\ : std_logic;
signal \N__25955\ : std_logic;
signal \N__25952\ : std_logic;
signal \N__25949\ : std_logic;
signal \N__25948\ : std_logic;
signal \N__25945\ : std_logic;
signal \N__25942\ : std_logic;
signal \N__25939\ : std_logic;
signal \N__25934\ : std_logic;
signal \N__25931\ : std_logic;
signal \N__25928\ : std_logic;
signal \N__25925\ : std_logic;
signal \N__25922\ : std_logic;
signal \N__25919\ : std_logic;
signal \N__25916\ : std_logic;
signal \N__25913\ : std_logic;
signal \N__25912\ : std_logic;
signal \N__25909\ : std_logic;
signal \N__25906\ : std_logic;
signal \N__25901\ : std_logic;
signal \N__25898\ : std_logic;
signal \N__25895\ : std_logic;
signal \N__25892\ : std_logic;
signal \N__25889\ : std_logic;
signal \N__25886\ : std_logic;
signal \N__25883\ : std_logic;
signal \N__25880\ : std_logic;
signal \N__25877\ : std_logic;
signal \N__25876\ : std_logic;
signal \N__25875\ : std_logic;
signal \N__25872\ : std_logic;
signal \N__25869\ : std_logic;
signal \N__25866\ : std_logic;
signal \N__25863\ : std_logic;
signal \N__25860\ : std_logic;
signal \N__25857\ : std_logic;
signal \N__25852\ : std_logic;
signal \N__25849\ : std_logic;
signal \N__25846\ : std_logic;
signal \N__25843\ : std_logic;
signal \N__25840\ : std_logic;
signal \N__25835\ : std_logic;
signal \N__25834\ : std_logic;
signal \N__25833\ : std_logic;
signal \N__25832\ : std_logic;
signal \N__25829\ : std_logic;
signal \N__25826\ : std_logic;
signal \N__25825\ : std_logic;
signal \N__25824\ : std_logic;
signal \N__25821\ : std_logic;
signal \N__25818\ : std_logic;
signal \N__25817\ : std_logic;
signal \N__25816\ : std_logic;
signal \N__25807\ : std_logic;
signal \N__25804\ : std_logic;
signal \N__25799\ : std_logic;
signal \N__25796\ : std_logic;
signal \N__25793\ : std_logic;
signal \N__25784\ : std_logic;
signal \N__25781\ : std_logic;
signal \N__25778\ : std_logic;
signal \N__25775\ : std_logic;
signal \N__25772\ : std_logic;
signal \N__25769\ : std_logic;
signal \N__25766\ : std_logic;
signal \N__25763\ : std_logic;
signal \N__25762\ : std_logic;
signal \N__25759\ : std_logic;
signal \N__25756\ : std_logic;
signal \N__25753\ : std_logic;
signal \N__25750\ : std_logic;
signal \N__25747\ : std_logic;
signal \N__25744\ : std_logic;
signal \N__25739\ : std_logic;
signal \N__25736\ : std_logic;
signal \N__25733\ : std_logic;
signal \N__25730\ : std_logic;
signal \N__25727\ : std_logic;
signal \N__25724\ : std_logic;
signal \N__25723\ : std_logic;
signal \N__25720\ : std_logic;
signal \N__25717\ : std_logic;
signal \N__25714\ : std_logic;
signal \N__25711\ : std_logic;
signal \N__25706\ : std_logic;
signal \N__25705\ : std_logic;
signal \N__25704\ : std_logic;
signal \N__25703\ : std_logic;
signal \N__25700\ : std_logic;
signal \N__25697\ : std_logic;
signal \N__25696\ : std_logic;
signal \N__25693\ : std_logic;
signal \N__25690\ : std_logic;
signal \N__25689\ : std_logic;
signal \N__25686\ : std_logic;
signal \N__25685\ : std_logic;
signal \N__25684\ : std_logic;
signal \N__25683\ : std_logic;
signal \N__25682\ : std_logic;
signal \N__25681\ : std_logic;
signal \N__25680\ : std_logic;
signal \N__25679\ : std_logic;
signal \N__25678\ : std_logic;
signal \N__25673\ : std_logic;
signal \N__25672\ : std_logic;
signal \N__25665\ : std_logic;
signal \N__25664\ : std_logic;
signal \N__25663\ : std_logic;
signal \N__25662\ : std_logic;
signal \N__25661\ : std_logic;
signal \N__25660\ : std_logic;
signal \N__25659\ : std_logic;
signal \N__25656\ : std_logic;
signal \N__25649\ : std_logic;
signal \N__25642\ : std_logic;
signal \N__25637\ : std_logic;
signal \N__25634\ : std_logic;
signal \N__25633\ : std_logic;
signal \N__25632\ : std_logic;
signal \N__25629\ : std_logic;
signal \N__25628\ : std_logic;
signal \N__25625\ : std_logic;
signal \N__25616\ : std_logic;
signal \N__25613\ : std_logic;
signal \N__25610\ : std_logic;
signal \N__25599\ : std_logic;
signal \N__25590\ : std_logic;
signal \N__25587\ : std_logic;
signal \N__25574\ : std_logic;
signal \N__25571\ : std_logic;
signal \N__25568\ : std_logic;
signal \N__25565\ : std_logic;
signal \N__25562\ : std_logic;
signal \N__25559\ : std_logic;
signal \N__25558\ : std_logic;
signal \N__25555\ : std_logic;
signal \N__25552\ : std_logic;
signal \N__25549\ : std_logic;
signal \N__25544\ : std_logic;
signal \N__25541\ : std_logic;
signal \N__25538\ : std_logic;
signal \N__25535\ : std_logic;
signal \N__25532\ : std_logic;
signal \N__25529\ : std_logic;
signal \N__25526\ : std_logic;
signal \N__25525\ : std_logic;
signal \N__25522\ : std_logic;
signal \N__25519\ : std_logic;
signal \N__25514\ : std_logic;
signal \N__25511\ : std_logic;
signal \N__25508\ : std_logic;
signal \N__25505\ : std_logic;
signal \N__25502\ : std_logic;
signal \N__25501\ : std_logic;
signal \N__25498\ : std_logic;
signal \N__25495\ : std_logic;
signal \N__25494\ : std_logic;
signal \N__25491\ : std_logic;
signal \N__25488\ : std_logic;
signal \N__25485\ : std_logic;
signal \N__25478\ : std_logic;
signal \N__25475\ : std_logic;
signal \N__25472\ : std_logic;
signal \N__25469\ : std_logic;
signal \N__25466\ : std_logic;
signal \N__25463\ : std_logic;
signal \N__25462\ : std_logic;
signal \N__25459\ : std_logic;
signal \N__25456\ : std_logic;
signal \N__25453\ : std_logic;
signal \N__25450\ : std_logic;
signal \N__25445\ : std_logic;
signal \N__25442\ : std_logic;
signal \N__25439\ : std_logic;
signal \N__25436\ : std_logic;
signal \N__25433\ : std_logic;
signal \N__25430\ : std_logic;
signal \N__25429\ : std_logic;
signal \N__25426\ : std_logic;
signal \N__25425\ : std_logic;
signal \N__25422\ : std_logic;
signal \N__25419\ : std_logic;
signal \N__25416\ : std_logic;
signal \N__25409\ : std_logic;
signal \N__25406\ : std_logic;
signal \N__25403\ : std_logic;
signal \N__25400\ : std_logic;
signal \N__25397\ : std_logic;
signal \N__25394\ : std_logic;
signal \N__25393\ : std_logic;
signal \N__25390\ : std_logic;
signal \N__25389\ : std_logic;
signal \N__25386\ : std_logic;
signal \N__25383\ : std_logic;
signal \N__25380\ : std_logic;
signal \N__25377\ : std_logic;
signal \N__25374\ : std_logic;
signal \N__25371\ : std_logic;
signal \N__25368\ : std_logic;
signal \N__25361\ : std_logic;
signal \N__25358\ : std_logic;
signal \N__25355\ : std_logic;
signal \N__25352\ : std_logic;
signal \N__25349\ : std_logic;
signal \N__25348\ : std_logic;
signal \N__25345\ : std_logic;
signal \N__25342\ : std_logic;
signal \N__25341\ : std_logic;
signal \N__25336\ : std_logic;
signal \N__25333\ : std_logic;
signal \N__25328\ : std_logic;
signal \N__25325\ : std_logic;
signal \N__25322\ : std_logic;
signal \N__25319\ : std_logic;
signal \N__25316\ : std_logic;
signal \N__25313\ : std_logic;
signal \N__25312\ : std_logic;
signal \N__25309\ : std_logic;
signal \N__25308\ : std_logic;
signal \N__25305\ : std_logic;
signal \N__25302\ : std_logic;
signal \N__25299\ : std_logic;
signal \N__25292\ : std_logic;
signal \N__25289\ : std_logic;
signal \N__25286\ : std_logic;
signal \N__25283\ : std_logic;
signal \N__25280\ : std_logic;
signal \N__25277\ : std_logic;
signal \N__25276\ : std_logic;
signal \N__25273\ : std_logic;
signal \N__25270\ : std_logic;
signal \N__25267\ : std_logic;
signal \N__25264\ : std_logic;
signal \N__25261\ : std_logic;
signal \N__25256\ : std_logic;
signal \N__25253\ : std_logic;
signal \N__25250\ : std_logic;
signal \N__25247\ : std_logic;
signal \N__25244\ : std_logic;
signal \N__25241\ : std_logic;
signal \N__25240\ : std_logic;
signal \N__25239\ : std_logic;
signal \N__25236\ : std_logic;
signal \N__25233\ : std_logic;
signal \N__25230\ : std_logic;
signal \N__25227\ : std_logic;
signal \N__25224\ : std_logic;
signal \N__25217\ : std_logic;
signal \N__25214\ : std_logic;
signal \N__25211\ : std_logic;
signal \N__25208\ : std_logic;
signal \N__25205\ : std_logic;
signal \N__25202\ : std_logic;
signal \N__25199\ : std_logic;
signal \N__25198\ : std_logic;
signal \N__25195\ : std_logic;
signal \N__25192\ : std_logic;
signal \N__25187\ : std_logic;
signal \N__25186\ : std_logic;
signal \N__25183\ : std_logic;
signal \N__25180\ : std_logic;
signal \N__25175\ : std_logic;
signal \N__25174\ : std_logic;
signal \N__25171\ : std_logic;
signal \N__25168\ : std_logic;
signal \N__25165\ : std_logic;
signal \N__25162\ : std_logic;
signal \N__25161\ : std_logic;
signal \N__25158\ : std_logic;
signal \N__25155\ : std_logic;
signal \N__25152\ : std_logic;
signal \N__25149\ : std_logic;
signal \N__25144\ : std_logic;
signal \N__25139\ : std_logic;
signal \N__25136\ : std_logic;
signal \N__25133\ : std_logic;
signal \N__25130\ : std_logic;
signal \N__25127\ : std_logic;
signal \N__25124\ : std_logic;
signal \N__25123\ : std_logic;
signal \N__25120\ : std_logic;
signal \N__25117\ : std_logic;
signal \N__25114\ : std_logic;
signal \N__25113\ : std_logic;
signal \N__25110\ : std_logic;
signal \N__25107\ : std_logic;
signal \N__25104\ : std_logic;
signal \N__25097\ : std_logic;
signal \N__25094\ : std_logic;
signal \N__25091\ : std_logic;
signal \N__25088\ : std_logic;
signal \N__25085\ : std_logic;
signal \N__25082\ : std_logic;
signal \N__25079\ : std_logic;
signal \N__25076\ : std_logic;
signal \N__25073\ : std_logic;
signal \N__25072\ : std_logic;
signal \N__25071\ : std_logic;
signal \N__25068\ : std_logic;
signal \N__25065\ : std_logic;
signal \N__25062\ : std_logic;
signal \N__25059\ : std_logic;
signal \N__25052\ : std_logic;
signal \N__25049\ : std_logic;
signal \N__25046\ : std_logic;
signal \N__25043\ : std_logic;
signal \N__25040\ : std_logic;
signal \N__25037\ : std_logic;
signal \N__25034\ : std_logic;
signal \N__25033\ : std_logic;
signal \N__25030\ : std_logic;
signal \N__25027\ : std_logic;
signal \N__25026\ : std_logic;
signal \N__25023\ : std_logic;
signal \N__25018\ : std_logic;
signal \N__25013\ : std_logic;
signal \N__25010\ : std_logic;
signal \N__25007\ : std_logic;
signal \N__25004\ : std_logic;
signal \N__25001\ : std_logic;
signal \N__24998\ : std_logic;
signal \N__24995\ : std_logic;
signal \N__24994\ : std_logic;
signal \N__24991\ : std_logic;
signal \N__24988\ : std_logic;
signal \N__24985\ : std_logic;
signal \N__24984\ : std_logic;
signal \N__24981\ : std_logic;
signal \N__24978\ : std_logic;
signal \N__24975\ : std_logic;
signal \N__24968\ : std_logic;
signal \N__24965\ : std_logic;
signal \N__24962\ : std_logic;
signal \N__24959\ : std_logic;
signal \N__24956\ : std_logic;
signal \N__24953\ : std_logic;
signal \N__24950\ : std_logic;
signal \N__24947\ : std_logic;
signal \N__24946\ : std_logic;
signal \N__24943\ : std_logic;
signal \N__24940\ : std_logic;
signal \N__24935\ : std_logic;
signal \N__24932\ : std_logic;
signal \N__24929\ : std_logic;
signal \N__24926\ : std_logic;
signal \N__24923\ : std_logic;
signal \N__24922\ : std_logic;
signal \N__24919\ : std_logic;
signal \N__24918\ : std_logic;
signal \N__24915\ : std_logic;
signal \N__24912\ : std_logic;
signal \N__24907\ : std_logic;
signal \N__24902\ : std_logic;
signal \N__24899\ : std_logic;
signal \N__24896\ : std_logic;
signal \N__24893\ : std_logic;
signal \N__24890\ : std_logic;
signal \N__24887\ : std_logic;
signal \N__24884\ : std_logic;
signal \N__24883\ : std_logic;
signal \N__24880\ : std_logic;
signal \N__24877\ : std_logic;
signal \N__24874\ : std_logic;
signal \N__24871\ : std_logic;
signal \N__24870\ : std_logic;
signal \N__24865\ : std_logic;
signal \N__24862\ : std_logic;
signal \N__24857\ : std_logic;
signal \N__24854\ : std_logic;
signal \N__24851\ : std_logic;
signal \N__24848\ : std_logic;
signal \N__24845\ : std_logic;
signal \N__24842\ : std_logic;
signal \N__24839\ : std_logic;
signal \N__24836\ : std_logic;
signal \N__24833\ : std_logic;
signal \N__24832\ : std_logic;
signal \N__24829\ : std_logic;
signal \N__24826\ : std_logic;
signal \N__24825\ : std_logic;
signal \N__24822\ : std_logic;
signal \N__24819\ : std_logic;
signal \N__24816\ : std_logic;
signal \N__24811\ : std_logic;
signal \N__24808\ : std_logic;
signal \N__24803\ : std_logic;
signal \N__24800\ : std_logic;
signal \N__24797\ : std_logic;
signal \N__24796\ : std_logic;
signal \N__24793\ : std_logic;
signal \N__24790\ : std_logic;
signal \N__24787\ : std_logic;
signal \N__24784\ : std_logic;
signal \N__24781\ : std_logic;
signal \N__24776\ : std_logic;
signal \N__24773\ : std_logic;
signal \N__24770\ : std_logic;
signal \N__24767\ : std_logic;
signal \N__24764\ : std_logic;
signal \N__24763\ : std_logic;
signal \N__24762\ : std_logic;
signal \N__24761\ : std_logic;
signal \N__24760\ : std_logic;
signal \N__24759\ : std_logic;
signal \N__24758\ : std_logic;
signal \N__24757\ : std_logic;
signal \N__24754\ : std_logic;
signal \N__24753\ : std_logic;
signal \N__24750\ : std_logic;
signal \N__24747\ : std_logic;
signal \N__24742\ : std_logic;
signal \N__24741\ : std_logic;
signal \N__24738\ : std_logic;
signal \N__24737\ : std_logic;
signal \N__24736\ : std_logic;
signal \N__24735\ : std_logic;
signal \N__24732\ : std_logic;
signal \N__24729\ : std_logic;
signal \N__24728\ : std_logic;
signal \N__24727\ : std_logic;
signal \N__24722\ : std_logic;
signal \N__24719\ : std_logic;
signal \N__24714\ : std_logic;
signal \N__24707\ : std_logic;
signal \N__24706\ : std_logic;
signal \N__24705\ : std_logic;
signal \N__24702\ : std_logic;
signal \N__24701\ : std_logic;
signal \N__24698\ : std_logic;
signal \N__24689\ : std_logic;
signal \N__24680\ : std_logic;
signal \N__24671\ : std_logic;
signal \N__24668\ : std_logic;
signal \N__24659\ : std_logic;
signal \N__24658\ : std_logic;
signal \N__24655\ : std_logic;
signal \N__24654\ : std_logic;
signal \N__24651\ : std_logic;
signal \N__24648\ : std_logic;
signal \N__24645\ : std_logic;
signal \N__24642\ : std_logic;
signal \N__24639\ : std_logic;
signal \N__24636\ : std_logic;
signal \N__24633\ : std_logic;
signal \N__24630\ : std_logic;
signal \N__24625\ : std_logic;
signal \N__24620\ : std_logic;
signal \N__24617\ : std_logic;
signal \N__24614\ : std_logic;
signal \N__24611\ : std_logic;
signal \N__24608\ : std_logic;
signal \N__24605\ : std_logic;
signal \N__24604\ : std_logic;
signal \N__24601\ : std_logic;
signal \N__24600\ : std_logic;
signal \N__24597\ : std_logic;
signal \N__24594\ : std_logic;
signal \N__24591\ : std_logic;
signal \N__24584\ : std_logic;
signal \N__24581\ : std_logic;
signal \N__24578\ : std_logic;
signal \N__24575\ : std_logic;
signal \N__24574\ : std_logic;
signal \N__24571\ : std_logic;
signal \N__24568\ : std_logic;
signal \N__24565\ : std_logic;
signal \N__24560\ : std_logic;
signal \N__24557\ : std_logic;
signal \N__24554\ : std_logic;
signal \N__24551\ : std_logic;
signal \N__24550\ : std_logic;
signal \N__24547\ : std_logic;
signal \N__24544\ : std_logic;
signal \N__24543\ : std_logic;
signal \N__24540\ : std_logic;
signal \N__24537\ : std_logic;
signal \N__24534\ : std_logic;
signal \N__24527\ : std_logic;
signal \N__24524\ : std_logic;
signal \N__24521\ : std_logic;
signal \N__24518\ : std_logic;
signal \N__24517\ : std_logic;
signal \N__24514\ : std_logic;
signal \N__24511\ : std_logic;
signal \N__24508\ : std_logic;
signal \N__24503\ : std_logic;
signal \N__24500\ : std_logic;
signal \N__24497\ : std_logic;
signal \N__24494\ : std_logic;
signal \N__24491\ : std_logic;
signal \N__24488\ : std_logic;
signal \N__24487\ : std_logic;
signal \N__24484\ : std_logic;
signal \N__24483\ : std_logic;
signal \N__24480\ : std_logic;
signal \N__24477\ : std_logic;
signal \N__24474\ : std_logic;
signal \N__24471\ : std_logic;
signal \N__24466\ : std_logic;
signal \N__24461\ : std_logic;
signal \N__24458\ : std_logic;
signal \N__24455\ : std_logic;
signal \N__24452\ : std_logic;
signal \N__24449\ : std_logic;
signal \N__24446\ : std_logic;
signal \N__24443\ : std_logic;
signal \N__24440\ : std_logic;
signal \N__24437\ : std_logic;
signal \N__24434\ : std_logic;
signal \N__24431\ : std_logic;
signal \N__24428\ : std_logic;
signal \N__24425\ : std_logic;
signal \N__24422\ : std_logic;
signal \N__24419\ : std_logic;
signal \N__24416\ : std_logic;
signal \N__24413\ : std_logic;
signal \N__24410\ : std_logic;
signal \N__24407\ : std_logic;
signal \N__24404\ : std_logic;
signal \N__24401\ : std_logic;
signal \N__24398\ : std_logic;
signal \N__24395\ : std_logic;
signal \N__24392\ : std_logic;
signal \N__24389\ : std_logic;
signal \N__24386\ : std_logic;
signal \N__24383\ : std_logic;
signal \N__24380\ : std_logic;
signal \N__24377\ : std_logic;
signal \N__24374\ : std_logic;
signal \N__24371\ : std_logic;
signal \N__24368\ : std_logic;
signal \N__24365\ : std_logic;
signal \N__24362\ : std_logic;
signal \N__24359\ : std_logic;
signal \N__24356\ : std_logic;
signal \N__24353\ : std_logic;
signal \N__24350\ : std_logic;
signal \N__24349\ : std_logic;
signal \N__24348\ : std_logic;
signal \N__24347\ : std_logic;
signal \N__24346\ : std_logic;
signal \N__24345\ : std_logic;
signal \N__24344\ : std_logic;
signal \N__24343\ : std_logic;
signal \N__24342\ : std_logic;
signal \N__24323\ : std_logic;
signal \N__24320\ : std_logic;
signal \N__24317\ : std_logic;
signal \N__24314\ : std_logic;
signal \N__24311\ : std_logic;
signal \N__24308\ : std_logic;
signal \N__24305\ : std_logic;
signal \N__24302\ : std_logic;
signal \N__24299\ : std_logic;
signal \N__24296\ : std_logic;
signal \N__24293\ : std_logic;
signal \N__24290\ : std_logic;
signal \N__24287\ : std_logic;
signal \N__24284\ : std_logic;
signal \N__24283\ : std_logic;
signal \N__24280\ : std_logic;
signal \N__24277\ : std_logic;
signal \N__24274\ : std_logic;
signal \N__24273\ : std_logic;
signal \N__24270\ : std_logic;
signal \N__24267\ : std_logic;
signal \N__24264\ : std_logic;
signal \N__24261\ : std_logic;
signal \N__24258\ : std_logic;
signal \N__24255\ : std_logic;
signal \N__24248\ : std_logic;
signal \N__24245\ : std_logic;
signal \N__24244\ : std_logic;
signal \N__24241\ : std_logic;
signal \N__24238\ : std_logic;
signal \N__24235\ : std_logic;
signal \N__24232\ : std_logic;
signal \N__24231\ : std_logic;
signal \N__24228\ : std_logic;
signal \N__24225\ : std_logic;
signal \N__24222\ : std_logic;
signal \N__24215\ : std_logic;
signal \N__24212\ : std_logic;
signal \N__24209\ : std_logic;
signal \N__24208\ : std_logic;
signal \N__24205\ : std_logic;
signal \N__24202\ : std_logic;
signal \N__24201\ : std_logic;
signal \N__24198\ : std_logic;
signal \N__24195\ : std_logic;
signal \N__24192\ : std_logic;
signal \N__24185\ : std_logic;
signal \N__24182\ : std_logic;
signal \N__24179\ : std_logic;
signal \N__24178\ : std_logic;
signal \N__24175\ : std_logic;
signal \N__24172\ : std_logic;
signal \N__24171\ : std_logic;
signal \N__24168\ : std_logic;
signal \N__24165\ : std_logic;
signal \N__24162\ : std_logic;
signal \N__24155\ : std_logic;
signal \N__24152\ : std_logic;
signal \N__24149\ : std_logic;
signal \N__24146\ : std_logic;
signal \N__24143\ : std_logic;
signal \N__24140\ : std_logic;
signal \N__24137\ : std_logic;
signal \N__24134\ : std_logic;
signal \N__24131\ : std_logic;
signal \N__24128\ : std_logic;
signal \N__24125\ : std_logic;
signal \N__24122\ : std_logic;
signal \N__24119\ : std_logic;
signal \N__24116\ : std_logic;
signal \N__24113\ : std_logic;
signal \N__24110\ : std_logic;
signal \N__24107\ : std_logic;
signal \N__24104\ : std_logic;
signal \N__24101\ : std_logic;
signal \N__24098\ : std_logic;
signal \N__24095\ : std_logic;
signal \N__24092\ : std_logic;
signal \N__24091\ : std_logic;
signal \N__24088\ : std_logic;
signal \N__24085\ : std_logic;
signal \N__24080\ : std_logic;
signal \N__24077\ : std_logic;
signal \N__24076\ : std_logic;
signal \N__24075\ : std_logic;
signal \N__24074\ : std_logic;
signal \N__24071\ : std_logic;
signal \N__24070\ : std_logic;
signal \N__24067\ : std_logic;
signal \N__24066\ : std_logic;
signal \N__24063\ : std_logic;
signal \N__24062\ : std_logic;
signal \N__24061\ : std_logic;
signal \N__24060\ : std_logic;
signal \N__24059\ : std_logic;
signal \N__24044\ : std_logic;
signal \N__24043\ : std_logic;
signal \N__24042\ : std_logic;
signal \N__24041\ : std_logic;
signal \N__24038\ : std_logic;
signal \N__24037\ : std_logic;
signal \N__24034\ : std_logic;
signal \N__24033\ : std_logic;
signal \N__24030\ : std_logic;
signal \N__24027\ : std_logic;
signal \N__24024\ : std_logic;
signal \N__24011\ : std_logic;
signal \N__24008\ : std_logic;
signal \N__24005\ : std_logic;
signal \N__24004\ : std_logic;
signal \N__23999\ : std_logic;
signal \N__23996\ : std_logic;
signal \N__23993\ : std_logic;
signal \N__23990\ : std_logic;
signal \N__23987\ : std_logic;
signal \N__23984\ : std_logic;
signal \N__23981\ : std_logic;
signal \N__23978\ : std_logic;
signal \N__23969\ : std_logic;
signal \N__23966\ : std_logic;
signal \N__23963\ : std_logic;
signal \N__23960\ : std_logic;
signal \N__23959\ : std_logic;
signal \N__23956\ : std_logic;
signal \N__23951\ : std_logic;
signal \N__23948\ : std_logic;
signal \N__23945\ : std_logic;
signal \N__23942\ : std_logic;
signal \N__23939\ : std_logic;
signal \N__23936\ : std_logic;
signal \N__23933\ : std_logic;
signal \N__23930\ : std_logic;
signal \N__23927\ : std_logic;
signal \N__23924\ : std_logic;
signal \N__23921\ : std_logic;
signal \N__23918\ : std_logic;
signal \N__23915\ : std_logic;
signal \N__23912\ : std_logic;
signal \N__23909\ : std_logic;
signal \N__23908\ : std_logic;
signal \N__23905\ : std_logic;
signal \N__23902\ : std_logic;
signal \N__23901\ : std_logic;
signal \N__23898\ : std_logic;
signal \N__23895\ : std_logic;
signal \N__23892\ : std_logic;
signal \N__23891\ : std_logic;
signal \N__23886\ : std_logic;
signal \N__23883\ : std_logic;
signal \N__23880\ : std_logic;
signal \N__23877\ : std_logic;
signal \N__23874\ : std_logic;
signal \N__23867\ : std_logic;
signal \N__23864\ : std_logic;
signal \N__23861\ : std_logic;
signal \N__23858\ : std_logic;
signal \N__23855\ : std_logic;
signal \N__23852\ : std_logic;
signal \N__23849\ : std_logic;
signal \N__23846\ : std_logic;
signal \N__23845\ : std_logic;
signal \N__23842\ : std_logic;
signal \N__23839\ : std_logic;
signal \N__23838\ : std_logic;
signal \N__23835\ : std_logic;
signal \N__23832\ : std_logic;
signal \N__23829\ : std_logic;
signal \N__23828\ : std_logic;
signal \N__23823\ : std_logic;
signal \N__23820\ : std_logic;
signal \N__23817\ : std_logic;
signal \N__23814\ : std_logic;
signal \N__23811\ : std_logic;
signal \N__23804\ : std_logic;
signal \N__23801\ : std_logic;
signal \N__23798\ : std_logic;
signal \N__23795\ : std_logic;
signal \N__23792\ : std_logic;
signal \N__23789\ : std_logic;
signal \N__23788\ : std_logic;
signal \N__23785\ : std_logic;
signal \N__23782\ : std_logic;
signal \N__23779\ : std_logic;
signal \N__23776\ : std_logic;
signal \N__23773\ : std_logic;
signal \N__23772\ : std_logic;
signal \N__23769\ : std_logic;
signal \N__23768\ : std_logic;
signal \N__23765\ : std_logic;
signal \N__23762\ : std_logic;
signal \N__23759\ : std_logic;
signal \N__23756\ : std_logic;
signal \N__23747\ : std_logic;
signal \N__23744\ : std_logic;
signal \N__23741\ : std_logic;
signal \N__23738\ : std_logic;
signal \N__23735\ : std_logic;
signal \N__23732\ : std_logic;
signal \N__23729\ : std_logic;
signal \N__23726\ : std_logic;
signal \N__23723\ : std_logic;
signal \N__23722\ : std_logic;
signal \N__23719\ : std_logic;
signal \N__23716\ : std_logic;
signal \N__23711\ : std_logic;
signal \N__23710\ : std_logic;
signal \N__23707\ : std_logic;
signal \N__23704\ : std_logic;
signal \N__23703\ : std_logic;
signal \N__23698\ : std_logic;
signal \N__23695\ : std_logic;
signal \N__23692\ : std_logic;
signal \N__23687\ : std_logic;
signal \N__23684\ : std_logic;
signal \N__23681\ : std_logic;
signal \N__23678\ : std_logic;
signal \N__23675\ : std_logic;
signal \N__23672\ : std_logic;
signal \N__23669\ : std_logic;
signal \N__23666\ : std_logic;
signal \N__23665\ : std_logic;
signal \N__23662\ : std_logic;
signal \N__23659\ : std_logic;
signal \N__23658\ : std_logic;
signal \N__23653\ : std_logic;
signal \N__23650\ : std_logic;
signal \N__23649\ : std_logic;
signal \N__23646\ : std_logic;
signal \N__23643\ : std_logic;
signal \N__23640\ : std_logic;
signal \N__23635\ : std_logic;
signal \N__23630\ : std_logic;
signal \N__23627\ : std_logic;
signal \N__23624\ : std_logic;
signal \N__23621\ : std_logic;
signal \N__23618\ : std_logic;
signal \N__23615\ : std_logic;
signal \N__23612\ : std_logic;
signal \N__23611\ : std_logic;
signal \N__23608\ : std_logic;
signal \N__23605\ : std_logic;
signal \N__23600\ : std_logic;
signal \N__23599\ : std_logic;
signal \N__23596\ : std_logic;
signal \N__23595\ : std_logic;
signal \N__23592\ : std_logic;
signal \N__23589\ : std_logic;
signal \N__23586\ : std_logic;
signal \N__23579\ : std_logic;
signal \N__23576\ : std_logic;
signal \N__23573\ : std_logic;
signal \N__23570\ : std_logic;
signal \N__23567\ : std_logic;
signal \N__23564\ : std_logic;
signal \N__23561\ : std_logic;
signal \N__23558\ : std_logic;
signal \N__23555\ : std_logic;
signal \N__23552\ : std_logic;
signal \N__23549\ : std_logic;
signal \N__23546\ : std_logic;
signal \N__23543\ : std_logic;
signal \N__23540\ : std_logic;
signal \N__23537\ : std_logic;
signal \N__23534\ : std_logic;
signal \N__23531\ : std_logic;
signal \N__23528\ : std_logic;
signal \N__23525\ : std_logic;
signal \N__23522\ : std_logic;
signal \N__23519\ : std_logic;
signal \N__23516\ : std_logic;
signal \N__23513\ : std_logic;
signal \N__23510\ : std_logic;
signal \N__23507\ : std_logic;
signal \N__23504\ : std_logic;
signal \N__23501\ : std_logic;
signal \N__23498\ : std_logic;
signal \N__23495\ : std_logic;
signal \N__23492\ : std_logic;
signal \N__23489\ : std_logic;
signal \N__23488\ : std_logic;
signal \N__23485\ : std_logic;
signal \N__23482\ : std_logic;
signal \N__23481\ : std_logic;
signal \N__23476\ : std_logic;
signal \N__23475\ : std_logic;
signal \N__23472\ : std_logic;
signal \N__23469\ : std_logic;
signal \N__23466\ : std_logic;
signal \N__23459\ : std_logic;
signal \N__23456\ : std_logic;
signal \N__23453\ : std_logic;
signal \N__23450\ : std_logic;
signal \N__23447\ : std_logic;
signal \N__23444\ : std_logic;
signal \N__23441\ : std_logic;
signal \N__23438\ : std_logic;
signal \N__23435\ : std_logic;
signal \N__23432\ : std_logic;
signal \N__23429\ : std_logic;
signal \N__23426\ : std_logic;
signal \N__23425\ : std_logic;
signal \N__23422\ : std_logic;
signal \N__23421\ : std_logic;
signal \N__23418\ : std_logic;
signal \N__23415\ : std_logic;
signal \N__23412\ : std_logic;
signal \N__23409\ : std_logic;
signal \N__23406\ : std_logic;
signal \N__23403\ : std_logic;
signal \N__23400\ : std_logic;
signal \N__23397\ : std_logic;
signal \N__23392\ : std_logic;
signal \N__23387\ : std_logic;
signal \N__23384\ : std_logic;
signal \N__23381\ : std_logic;
signal \N__23378\ : std_logic;
signal \N__23375\ : std_logic;
signal \N__23374\ : std_logic;
signal \N__23373\ : std_logic;
signal \N__23372\ : std_logic;
signal \N__23371\ : std_logic;
signal \N__23370\ : std_logic;
signal \N__23369\ : std_logic;
signal \N__23366\ : std_logic;
signal \N__23365\ : std_logic;
signal \N__23364\ : std_logic;
signal \N__23363\ : std_logic;
signal \N__23362\ : std_logic;
signal \N__23361\ : std_logic;
signal \N__23354\ : std_logic;
signal \N__23353\ : std_logic;
signal \N__23352\ : std_logic;
signal \N__23349\ : std_logic;
signal \N__23348\ : std_logic;
signal \N__23347\ : std_logic;
signal \N__23346\ : std_logic;
signal \N__23345\ : std_logic;
signal \N__23342\ : std_logic;
signal \N__23341\ : std_logic;
signal \N__23338\ : std_logic;
signal \N__23333\ : std_logic;
signal \N__23332\ : std_logic;
signal \N__23331\ : std_logic;
signal \N__23328\ : std_logic;
signal \N__23325\ : std_logic;
signal \N__23324\ : std_logic;
signal \N__23319\ : std_logic;
signal \N__23316\ : std_logic;
signal \N__23313\ : std_logic;
signal \N__23306\ : std_logic;
signal \N__23299\ : std_logic;
signal \N__23294\ : std_logic;
signal \N__23291\ : std_logic;
signal \N__23288\ : std_logic;
signal \N__23277\ : std_logic;
signal \N__23272\ : std_logic;
signal \N__23255\ : std_logic;
signal \N__23254\ : std_logic;
signal \N__23251\ : std_logic;
signal \N__23248\ : std_logic;
signal \N__23245\ : std_logic;
signal \N__23244\ : std_logic;
signal \N__23239\ : std_logic;
signal \N__23236\ : std_logic;
signal \N__23231\ : std_logic;
signal \N__23228\ : std_logic;
signal \N__23225\ : std_logic;
signal \N__23222\ : std_logic;
signal \N__23221\ : std_logic;
signal \N__23220\ : std_logic;
signal \N__23217\ : std_logic;
signal \N__23214\ : std_logic;
signal \N__23211\ : std_logic;
signal \N__23208\ : std_logic;
signal \N__23205\ : std_logic;
signal \N__23202\ : std_logic;
signal \N__23199\ : std_logic;
signal \N__23194\ : std_logic;
signal \N__23189\ : std_logic;
signal \N__23188\ : std_logic;
signal \N__23185\ : std_logic;
signal \N__23182\ : std_logic;
signal \N__23179\ : std_logic;
signal \N__23178\ : std_logic;
signal \N__23175\ : std_logic;
signal \N__23172\ : std_logic;
signal \N__23169\ : std_logic;
signal \N__23166\ : std_logic;
signal \N__23159\ : std_logic;
signal \N__23156\ : std_logic;
signal \N__23153\ : std_logic;
signal \N__23150\ : std_logic;
signal \N__23147\ : std_logic;
signal \N__23144\ : std_logic;
signal \N__23141\ : std_logic;
signal \N__23140\ : std_logic;
signal \N__23139\ : std_logic;
signal \N__23136\ : std_logic;
signal \N__23131\ : std_logic;
signal \N__23126\ : std_logic;
signal \N__23123\ : std_logic;
signal \N__23120\ : std_logic;
signal \N__23117\ : std_logic;
signal \N__23114\ : std_logic;
signal \N__23113\ : std_logic;
signal \N__23110\ : std_logic;
signal \N__23107\ : std_logic;
signal \N__23106\ : std_logic;
signal \N__23103\ : std_logic;
signal \N__23100\ : std_logic;
signal \N__23097\ : std_logic;
signal \N__23092\ : std_logic;
signal \N__23087\ : std_logic;
signal \N__23084\ : std_logic;
signal \N__23081\ : std_logic;
signal \N__23078\ : std_logic;
signal \N__23077\ : std_logic;
signal \N__23074\ : std_logic;
signal \N__23073\ : std_logic;
signal \N__23070\ : std_logic;
signal \N__23067\ : std_logic;
signal \N__23064\ : std_logic;
signal \N__23059\ : std_logic;
signal \N__23054\ : std_logic;
signal \N__23051\ : std_logic;
signal \N__23048\ : std_logic;
signal \N__23045\ : std_logic;
signal \N__23042\ : std_logic;
signal \N__23039\ : std_logic;
signal \N__23036\ : std_logic;
signal \N__23035\ : std_logic;
signal \N__23032\ : std_logic;
signal \N__23031\ : std_logic;
signal \N__23028\ : std_logic;
signal \N__23025\ : std_logic;
signal \N__23022\ : std_logic;
signal \N__23017\ : std_logic;
signal \N__23012\ : std_logic;
signal \N__23009\ : std_logic;
signal \N__23006\ : std_logic;
signal \N__23003\ : std_logic;
signal \N__23000\ : std_logic;
signal \N__22997\ : std_logic;
signal \N__22994\ : std_logic;
signal \N__22991\ : std_logic;
signal \N__22990\ : std_logic;
signal \N__22987\ : std_logic;
signal \N__22984\ : std_logic;
signal \N__22983\ : std_logic;
signal \N__22980\ : std_logic;
signal \N__22979\ : std_logic;
signal \N__22978\ : std_logic;
signal \N__22977\ : std_logic;
signal \N__22974\ : std_logic;
signal \N__22971\ : std_logic;
signal \N__22970\ : std_logic;
signal \N__22969\ : std_logic;
signal \N__22966\ : std_logic;
signal \N__22963\ : std_logic;
signal \N__22960\ : std_logic;
signal \N__22959\ : std_logic;
signal \N__22958\ : std_logic;
signal \N__22957\ : std_logic;
signal \N__22956\ : std_logic;
signal \N__22955\ : std_logic;
signal \N__22954\ : std_logic;
signal \N__22951\ : std_logic;
signal \N__22950\ : std_logic;
signal \N__22949\ : std_logic;
signal \N__22944\ : std_logic;
signal \N__22943\ : std_logic;
signal \N__22942\ : std_logic;
signal \N__22939\ : std_logic;
signal \N__22938\ : std_logic;
signal \N__22935\ : std_logic;
signal \N__22930\ : std_logic;
signal \N__22927\ : std_logic;
signal \N__22924\ : std_logic;
signal \N__22923\ : std_logic;
signal \N__22922\ : std_logic;
signal \N__22921\ : std_logic;
signal \N__22920\ : std_logic;
signal \N__22917\ : std_logic;
signal \N__22912\ : std_logic;
signal \N__22907\ : std_logic;
signal \N__22906\ : std_logic;
signal \N__22903\ : std_logic;
signal \N__22898\ : std_logic;
signal \N__22895\ : std_logic;
signal \N__22892\ : std_logic;
signal \N__22889\ : std_logic;
signal \N__22888\ : std_logic;
signal \N__22885\ : std_logic;
signal \N__22882\ : std_logic;
signal \N__22879\ : std_logic;
signal \N__22874\ : std_logic;
signal \N__22871\ : std_logic;
signal \N__22862\ : std_logic;
signal \N__22855\ : std_logic;
signal \N__22854\ : std_logic;
signal \N__22853\ : std_logic;
signal \N__22852\ : std_logic;
signal \N__22851\ : std_logic;
signal \N__22850\ : std_logic;
signal \N__22849\ : std_logic;
signal \N__22848\ : std_logic;
signal \N__22847\ : std_logic;
signal \N__22846\ : std_logic;
signal \N__22845\ : std_logic;
signal \N__22842\ : std_logic;
signal \N__22831\ : std_logic;
signal \N__22828\ : std_logic;
signal \N__22819\ : std_logic;
signal \N__22812\ : std_logic;
signal \N__22803\ : std_logic;
signal \N__22794\ : std_logic;
signal \N__22789\ : std_logic;
signal \N__22772\ : std_logic;
signal \N__22769\ : std_logic;
signal \N__22766\ : std_logic;
signal \N__22763\ : std_logic;
signal \N__22760\ : std_logic;
signal \N__22757\ : std_logic;
signal \N__22754\ : std_logic;
signal \N__22751\ : std_logic;
signal \N__22748\ : std_logic;
signal \N__22745\ : std_logic;
signal \N__22742\ : std_logic;
signal \N__22739\ : std_logic;
signal \N__22736\ : std_logic;
signal \N__22733\ : std_logic;
signal \N__22732\ : std_logic;
signal \N__22729\ : std_logic;
signal \N__22726\ : std_logic;
signal \N__22723\ : std_logic;
signal \N__22720\ : std_logic;
signal \N__22715\ : std_logic;
signal \N__22712\ : std_logic;
signal \N__22709\ : std_logic;
signal \N__22706\ : std_logic;
signal \N__22703\ : std_logic;
signal \N__22700\ : std_logic;
signal \N__22697\ : std_logic;
signal \N__22694\ : std_logic;
signal \N__22691\ : std_logic;
signal \N__22688\ : std_logic;
signal \N__22685\ : std_logic;
signal \N__22684\ : std_logic;
signal \N__22681\ : std_logic;
signal \N__22678\ : std_logic;
signal \N__22675\ : std_logic;
signal \N__22674\ : std_logic;
signal \N__22669\ : std_logic;
signal \N__22666\ : std_logic;
signal \N__22661\ : std_logic;
signal \N__22658\ : std_logic;
signal \N__22655\ : std_logic;
signal \N__22652\ : std_logic;
signal \N__22649\ : std_logic;
signal \N__22646\ : std_logic;
signal \N__22645\ : std_logic;
signal \N__22642\ : std_logic;
signal \N__22639\ : std_logic;
signal \N__22636\ : std_logic;
signal \N__22635\ : std_logic;
signal \N__22630\ : std_logic;
signal \N__22627\ : std_logic;
signal \N__22622\ : std_logic;
signal \N__22619\ : std_logic;
signal \N__22616\ : std_logic;
signal \N__22613\ : std_logic;
signal \N__22610\ : std_logic;
signal \N__22607\ : std_logic;
signal \N__22606\ : std_logic;
signal \N__22605\ : std_logic;
signal \N__22602\ : std_logic;
signal \N__22597\ : std_logic;
signal \N__22592\ : std_logic;
signal \N__22589\ : std_logic;
signal \N__22586\ : std_logic;
signal \N__22583\ : std_logic;
signal \N__22580\ : std_logic;
signal \N__22577\ : std_logic;
signal \N__22574\ : std_logic;
signal \N__22571\ : std_logic;
signal \N__22570\ : std_logic;
signal \N__22567\ : std_logic;
signal \N__22564\ : std_logic;
signal \N__22563\ : std_logic;
signal \N__22560\ : std_logic;
signal \N__22555\ : std_logic;
signal \N__22552\ : std_logic;
signal \N__22549\ : std_logic;
signal \N__22544\ : std_logic;
signal \N__22541\ : std_logic;
signal \N__22538\ : std_logic;
signal \N__22535\ : std_logic;
signal \N__22532\ : std_logic;
signal \N__22529\ : std_logic;
signal \N__22528\ : std_logic;
signal \N__22525\ : std_logic;
signal \N__22524\ : std_logic;
signal \N__22521\ : std_logic;
signal \N__22518\ : std_logic;
signal \N__22515\ : std_logic;
signal \N__22510\ : std_logic;
signal \N__22507\ : std_logic;
signal \N__22502\ : std_logic;
signal \N__22499\ : std_logic;
signal \N__22496\ : std_logic;
signal \N__22493\ : std_logic;
signal \N__22490\ : std_logic;
signal \N__22489\ : std_logic;
signal \N__22486\ : std_logic;
signal \N__22483\ : std_logic;
signal \N__22480\ : std_logic;
signal \N__22479\ : std_logic;
signal \N__22476\ : std_logic;
signal \N__22473\ : std_logic;
signal \N__22470\ : std_logic;
signal \N__22463\ : std_logic;
signal \N__22460\ : std_logic;
signal \N__22457\ : std_logic;
signal \N__22454\ : std_logic;
signal \N__22451\ : std_logic;
signal \N__22448\ : std_logic;
signal \N__22445\ : std_logic;
signal \N__22444\ : std_logic;
signal \N__22443\ : std_logic;
signal \N__22440\ : std_logic;
signal \N__22437\ : std_logic;
signal \N__22434\ : std_logic;
signal \N__22431\ : std_logic;
signal \N__22428\ : std_logic;
signal \N__22425\ : std_logic;
signal \N__22418\ : std_logic;
signal \N__22415\ : std_logic;
signal \N__22412\ : std_logic;
signal \N__22409\ : std_logic;
signal \N__22406\ : std_logic;
signal \N__22405\ : std_logic;
signal \N__22402\ : std_logic;
signal \N__22399\ : std_logic;
signal \N__22396\ : std_logic;
signal \N__22393\ : std_logic;
signal \N__22388\ : std_logic;
signal \N__22385\ : std_logic;
signal \N__22382\ : std_logic;
signal \N__22379\ : std_logic;
signal \N__22376\ : std_logic;
signal \N__22373\ : std_logic;
signal \N__22370\ : std_logic;
signal \N__22369\ : std_logic;
signal \N__22366\ : std_logic;
signal \N__22363\ : std_logic;
signal \N__22360\ : std_logic;
signal \N__22355\ : std_logic;
signal \N__22352\ : std_logic;
signal \N__22349\ : std_logic;
signal \N__22346\ : std_logic;
signal \N__22343\ : std_logic;
signal \N__22340\ : std_logic;
signal \N__22339\ : std_logic;
signal \N__22338\ : std_logic;
signal \N__22335\ : std_logic;
signal \N__22332\ : std_logic;
signal \N__22329\ : std_logic;
signal \N__22326\ : std_logic;
signal \N__22319\ : std_logic;
signal \N__22316\ : std_logic;
signal \N__22313\ : std_logic;
signal \N__22310\ : std_logic;
signal \N__22307\ : std_logic;
signal \N__22304\ : std_logic;
signal \N__22301\ : std_logic;
signal \N__22298\ : std_logic;
signal \N__22297\ : std_logic;
signal \N__22294\ : std_logic;
signal \N__22291\ : std_logic;
signal \N__22286\ : std_logic;
signal \N__22283\ : std_logic;
signal \N__22280\ : std_logic;
signal \N__22277\ : std_logic;
signal \N__22274\ : std_logic;
signal \N__22271\ : std_logic;
signal \N__22270\ : std_logic;
signal \N__22269\ : std_logic;
signal \N__22266\ : std_logic;
signal \N__22261\ : std_logic;
signal \N__22258\ : std_logic;
signal \N__22253\ : std_logic;
signal \N__22250\ : std_logic;
signal \N__22247\ : std_logic;
signal \N__22244\ : std_logic;
signal \N__22241\ : std_logic;
signal \N__22240\ : std_logic;
signal \N__22237\ : std_logic;
signal \N__22234\ : std_logic;
signal \N__22231\ : std_logic;
signal \N__22230\ : std_logic;
signal \N__22227\ : std_logic;
signal \N__22224\ : std_logic;
signal \N__22221\ : std_logic;
signal \N__22214\ : std_logic;
signal \N__22211\ : std_logic;
signal \N__22208\ : std_logic;
signal \N__22205\ : std_logic;
signal \N__22202\ : std_logic;
signal \N__22199\ : std_logic;
signal \N__22198\ : std_logic;
signal \N__22195\ : std_logic;
signal \N__22192\ : std_logic;
signal \N__22189\ : std_logic;
signal \N__22186\ : std_logic;
signal \N__22183\ : std_logic;
signal \N__22178\ : std_logic;
signal \N__22175\ : std_logic;
signal \N__22172\ : std_logic;
signal \N__22169\ : std_logic;
signal \N__22166\ : std_logic;
signal \N__22165\ : std_logic;
signal \N__22162\ : std_logic;
signal \N__22159\ : std_logic;
signal \N__22156\ : std_logic;
signal \N__22155\ : std_logic;
signal \N__22150\ : std_logic;
signal \N__22147\ : std_logic;
signal \N__22142\ : std_logic;
signal \N__22139\ : std_logic;
signal \N__22136\ : std_logic;
signal \N__22133\ : std_logic;
signal \N__22130\ : std_logic;
signal \N__22127\ : std_logic;
signal \N__22126\ : std_logic;
signal \N__22125\ : std_logic;
signal \N__22122\ : std_logic;
signal \N__22119\ : std_logic;
signal \N__22116\ : std_logic;
signal \N__22113\ : std_logic;
signal \N__22110\ : std_logic;
signal \N__22107\ : std_logic;
signal \N__22100\ : std_logic;
signal \N__22097\ : std_logic;
signal \N__22094\ : std_logic;
signal \N__22091\ : std_logic;
signal \N__22088\ : std_logic;
signal \N__22085\ : std_logic;
signal \N__22082\ : std_logic;
signal \N__22081\ : std_logic;
signal \N__22080\ : std_logic;
signal \N__22077\ : std_logic;
signal \N__22074\ : std_logic;
signal \N__22071\ : std_logic;
signal \N__22068\ : std_logic;
signal \N__22065\ : std_logic;
signal \N__22062\ : std_logic;
signal \N__22055\ : std_logic;
signal \N__22052\ : std_logic;
signal \N__22049\ : std_logic;
signal \N__22046\ : std_logic;
signal \N__22043\ : std_logic;
signal \N__22042\ : std_logic;
signal \N__22039\ : std_logic;
signal \N__22038\ : std_logic;
signal \N__22035\ : std_logic;
signal \N__22030\ : std_logic;
signal \N__22025\ : std_logic;
signal \N__22022\ : std_logic;
signal \N__22019\ : std_logic;
signal \N__22016\ : std_logic;
signal \N__22013\ : std_logic;
signal \N__22012\ : std_logic;
signal \N__22009\ : std_logic;
signal \N__22006\ : std_logic;
signal \N__22003\ : std_logic;
signal \N__22002\ : std_logic;
signal \N__21999\ : std_logic;
signal \N__21996\ : std_logic;
signal \N__21993\ : std_logic;
signal \N__21986\ : std_logic;
signal \N__21983\ : std_logic;
signal \N__21980\ : std_logic;
signal \N__21977\ : std_logic;
signal \N__21976\ : std_logic;
signal \N__21973\ : std_logic;
signal \N__21970\ : std_logic;
signal \N__21967\ : std_logic;
signal \N__21962\ : std_logic;
signal \N__21959\ : std_logic;
signal \N__21956\ : std_logic;
signal \N__21953\ : std_logic;
signal \N__21952\ : std_logic;
signal \N__21951\ : std_logic;
signal \N__21948\ : std_logic;
signal \N__21945\ : std_logic;
signal \N__21942\ : std_logic;
signal \N__21937\ : std_logic;
signal \N__21932\ : std_logic;
signal \N__21929\ : std_logic;
signal \N__21926\ : std_logic;
signal \N__21925\ : std_logic;
signal \N__21922\ : std_logic;
signal \N__21919\ : std_logic;
signal \N__21916\ : std_logic;
signal \N__21913\ : std_logic;
signal \N__21912\ : std_logic;
signal \N__21909\ : std_logic;
signal \N__21906\ : std_logic;
signal \N__21903\ : std_logic;
signal \N__21896\ : std_logic;
signal \N__21893\ : std_logic;
signal \N__21890\ : std_logic;
signal \N__21889\ : std_logic;
signal \N__21886\ : std_logic;
signal \N__21883\ : std_logic;
signal \N__21880\ : std_logic;
signal \N__21877\ : std_logic;
signal \N__21876\ : std_logic;
signal \N__21873\ : std_logic;
signal \N__21870\ : std_logic;
signal \N__21867\ : std_logic;
signal \N__21860\ : std_logic;
signal \N__21857\ : std_logic;
signal \N__21854\ : std_logic;
signal \N__21851\ : std_logic;
signal \N__21848\ : std_logic;
signal \N__21845\ : std_logic;
signal \N__21844\ : std_logic;
signal \N__21841\ : std_logic;
signal \N__21838\ : std_logic;
signal \N__21835\ : std_logic;
signal \N__21832\ : std_logic;
signal \N__21831\ : std_logic;
signal \N__21826\ : std_logic;
signal \N__21823\ : std_logic;
signal \N__21818\ : std_logic;
signal \N__21817\ : std_logic;
signal \N__21814\ : std_logic;
signal \N__21811\ : std_logic;
signal \N__21808\ : std_logic;
signal \N__21803\ : std_logic;
signal \N__21800\ : std_logic;
signal \N__21797\ : std_logic;
signal \N__21794\ : std_logic;
signal \N__21793\ : std_logic;
signal \N__21792\ : std_logic;
signal \N__21791\ : std_logic;
signal \N__21790\ : std_logic;
signal \N__21789\ : std_logic;
signal \N__21788\ : std_logic;
signal \N__21785\ : std_logic;
signal \N__21784\ : std_logic;
signal \N__21781\ : std_logic;
signal \N__21778\ : std_logic;
signal \N__21777\ : std_logic;
signal \N__21776\ : std_logic;
signal \N__21773\ : std_logic;
signal \N__21772\ : std_logic;
signal \N__21771\ : std_logic;
signal \N__21766\ : std_logic;
signal \N__21765\ : std_logic;
signal \N__21764\ : std_logic;
signal \N__21763\ : std_logic;
signal \N__21762\ : std_logic;
signal \N__21761\ : std_logic;
signal \N__21758\ : std_logic;
signal \N__21753\ : std_logic;
signal \N__21750\ : std_logic;
signal \N__21747\ : std_logic;
signal \N__21746\ : std_logic;
signal \N__21743\ : std_logic;
signal \N__21742\ : std_logic;
signal \N__21741\ : std_logic;
signal \N__21738\ : std_logic;
signal \N__21731\ : std_logic;
signal \N__21728\ : std_logic;
signal \N__21721\ : std_logic;
signal \N__21716\ : std_logic;
signal \N__21711\ : std_logic;
signal \N__21706\ : std_logic;
signal \N__21697\ : std_logic;
signal \N__21680\ : std_logic;
signal \N__21677\ : std_logic;
signal \N__21676\ : std_logic;
signal \N__21673\ : std_logic;
signal \N__21670\ : std_logic;
signal \N__21667\ : std_logic;
signal \N__21664\ : std_logic;
signal \N__21661\ : std_logic;
signal \N__21658\ : std_logic;
signal \N__21653\ : std_logic;
signal \N__21650\ : std_logic;
signal \N__21647\ : std_logic;
signal \N__21644\ : std_logic;
signal \N__21643\ : std_logic;
signal \N__21640\ : std_logic;
signal \N__21637\ : std_logic;
signal \N__21632\ : std_logic;
signal \N__21629\ : std_logic;
signal \N__21626\ : std_logic;
signal \N__21623\ : std_logic;
signal \N__21620\ : std_logic;
signal \N__21617\ : std_logic;
signal \N__21616\ : std_logic;
signal \N__21615\ : std_logic;
signal \N__21612\ : std_logic;
signal \N__21609\ : std_logic;
signal \N__21606\ : std_logic;
signal \N__21603\ : std_logic;
signal \N__21598\ : std_logic;
signal \N__21593\ : std_logic;
signal \N__21590\ : std_logic;
signal \N__21587\ : std_logic;
signal \N__21584\ : std_logic;
signal \N__21581\ : std_logic;
signal \N__21580\ : std_logic;
signal \N__21577\ : std_logic;
signal \N__21574\ : std_logic;
signal \N__21571\ : std_logic;
signal \N__21568\ : std_logic;
signal \N__21563\ : std_logic;
signal \N__21560\ : std_logic;
signal \N__21559\ : std_logic;
signal \N__21556\ : std_logic;
signal \N__21553\ : std_logic;
signal \N__21552\ : std_logic;
signal \N__21549\ : std_logic;
signal \N__21546\ : std_logic;
signal \N__21543\ : std_logic;
signal \N__21536\ : std_logic;
signal \N__21533\ : std_logic;
signal \N__21530\ : std_logic;
signal \N__21527\ : std_logic;
signal \N__21524\ : std_logic;
signal \N__21521\ : std_logic;
signal \N__21518\ : std_logic;
signal \N__21517\ : std_logic;
signal \N__21514\ : std_logic;
signal \N__21511\ : std_logic;
signal \N__21510\ : std_logic;
signal \N__21507\ : std_logic;
signal \N__21504\ : std_logic;
signal \N__21501\ : std_logic;
signal \N__21494\ : std_logic;
signal \N__21493\ : std_logic;
signal \N__21490\ : std_logic;
signal \N__21487\ : std_logic;
signal \N__21482\ : std_logic;
signal \N__21481\ : std_logic;
signal \N__21478\ : std_logic;
signal \N__21475\ : std_logic;
signal \N__21470\ : std_logic;
signal \N__21467\ : std_logic;
signal \N__21464\ : std_logic;
signal \N__21461\ : std_logic;
signal \N__21458\ : std_logic;
signal \N__21455\ : std_logic;
signal \N__21454\ : std_logic;
signal \N__21453\ : std_logic;
signal \N__21450\ : std_logic;
signal \N__21447\ : std_logic;
signal \N__21444\ : std_logic;
signal \N__21441\ : std_logic;
signal \N__21438\ : std_logic;
signal \N__21435\ : std_logic;
signal \N__21428\ : std_logic;
signal \N__21427\ : std_logic;
signal \N__21424\ : std_logic;
signal \N__21421\ : std_logic;
signal \N__21416\ : std_logic;
signal \N__21413\ : std_logic;
signal \N__21410\ : std_logic;
signal \N__21407\ : std_logic;
signal \N__21404\ : std_logic;
signal \N__21401\ : std_logic;
signal \N__21398\ : std_logic;
signal \N__21395\ : std_logic;
signal \N__21392\ : std_logic;
signal \N__21391\ : std_logic;
signal \N__21390\ : std_logic;
signal \N__21387\ : std_logic;
signal \N__21384\ : std_logic;
signal \N__21381\ : std_logic;
signal \N__21378\ : std_logic;
signal \N__21371\ : std_logic;
signal \N__21370\ : std_logic;
signal \N__21367\ : std_logic;
signal \N__21364\ : std_logic;
signal \N__21361\ : std_logic;
signal \N__21356\ : std_logic;
signal \N__21353\ : std_logic;
signal \N__21350\ : std_logic;
signal \N__21347\ : std_logic;
signal \N__21344\ : std_logic;
signal \N__21341\ : std_logic;
signal \N__21340\ : std_logic;
signal \N__21337\ : std_logic;
signal \N__21334\ : std_logic;
signal \N__21331\ : std_logic;
signal \N__21326\ : std_logic;
signal \N__21323\ : std_logic;
signal \N__21320\ : std_logic;
signal \N__21317\ : std_logic;
signal \N__21314\ : std_logic;
signal \N__21311\ : std_logic;
signal \N__21310\ : std_logic;
signal \N__21307\ : std_logic;
signal \N__21306\ : std_logic;
signal \N__21303\ : std_logic;
signal \N__21300\ : std_logic;
signal \N__21297\ : std_logic;
signal \N__21294\ : std_logic;
signal \N__21291\ : std_logic;
signal \N__21288\ : std_logic;
signal \N__21285\ : std_logic;
signal \N__21278\ : std_logic;
signal \N__21275\ : std_logic;
signal \N__21272\ : std_logic;
signal \N__21269\ : std_logic;
signal \N__21266\ : std_logic;
signal \N__21265\ : std_logic;
signal \N__21264\ : std_logic;
signal \N__21261\ : std_logic;
signal \N__21258\ : std_logic;
signal \N__21255\ : std_logic;
signal \N__21252\ : std_logic;
signal \N__21249\ : std_logic;
signal \N__21246\ : std_logic;
signal \N__21241\ : std_logic;
signal \N__21238\ : std_logic;
signal \N__21233\ : std_logic;
signal \N__21230\ : std_logic;
signal \N__21227\ : std_logic;
signal \N__21224\ : std_logic;
signal \N__21221\ : std_logic;
signal \N__21218\ : std_logic;
signal \N__21215\ : std_logic;
signal \N__21212\ : std_logic;
signal \N__21209\ : std_logic;
signal \N__21206\ : std_logic;
signal \N__21203\ : std_logic;
signal \N__21200\ : std_logic;
signal \N__21197\ : std_logic;
signal \N__21194\ : std_logic;
signal \N__21191\ : std_logic;
signal \N__21188\ : std_logic;
signal \N__21185\ : std_logic;
signal \N__21182\ : std_logic;
signal \N__21179\ : std_logic;
signal \N__21176\ : std_logic;
signal \N__21173\ : std_logic;
signal \N__21170\ : std_logic;
signal \N__21167\ : std_logic;
signal \N__21164\ : std_logic;
signal \N__21161\ : std_logic;
signal \N__21158\ : std_logic;
signal \N__21155\ : std_logic;
signal \N__21152\ : std_logic;
signal \N__21149\ : std_logic;
signal \N__21146\ : std_logic;
signal \N__21143\ : std_logic;
signal \N__21140\ : std_logic;
signal \N__21137\ : std_logic;
signal \N__21134\ : std_logic;
signal \N__21131\ : std_logic;
signal \N__21128\ : std_logic;
signal \N__21125\ : std_logic;
signal \N__21122\ : std_logic;
signal \N__21119\ : std_logic;
signal \N__21116\ : std_logic;
signal \N__21113\ : std_logic;
signal \N__21110\ : std_logic;
signal \N__21107\ : std_logic;
signal \N__21106\ : std_logic;
signal \N__21103\ : std_logic;
signal \N__21100\ : std_logic;
signal \N__21095\ : std_logic;
signal \N__21092\ : std_logic;
signal \N__21089\ : std_logic;
signal \N__21086\ : std_logic;
signal \N__21083\ : std_logic;
signal \N__21080\ : std_logic;
signal \N__21077\ : std_logic;
signal \N__21076\ : std_logic;
signal \N__21073\ : std_logic;
signal \N__21072\ : std_logic;
signal \N__21069\ : std_logic;
signal \N__21066\ : std_logic;
signal \N__21063\ : std_logic;
signal \N__21056\ : std_logic;
signal \N__21053\ : std_logic;
signal \N__21050\ : std_logic;
signal \N__21047\ : std_logic;
signal \N__21044\ : std_logic;
signal \N__21041\ : std_logic;
signal \N__21038\ : std_logic;
signal \N__21035\ : std_logic;
signal \N__21032\ : std_logic;
signal \N__21029\ : std_logic;
signal \N__21026\ : std_logic;
signal \N__21023\ : std_logic;
signal \N__21020\ : std_logic;
signal \N__21017\ : std_logic;
signal \N__21014\ : std_logic;
signal \N__21011\ : std_logic;
signal \N__21008\ : std_logic;
signal \N__21005\ : std_logic;
signal \N__21002\ : std_logic;
signal \N__20999\ : std_logic;
signal \N__20996\ : std_logic;
signal \N__20993\ : std_logic;
signal \N__20990\ : std_logic;
signal \N__20987\ : std_logic;
signal \N__20984\ : std_logic;
signal \N__20981\ : std_logic;
signal \N__20978\ : std_logic;
signal \N__20975\ : std_logic;
signal \N__20974\ : std_logic;
signal \N__20971\ : std_logic;
signal \N__20968\ : std_logic;
signal \N__20965\ : std_logic;
signal \N__20960\ : std_logic;
signal \N__20957\ : std_logic;
signal \N__20954\ : std_logic;
signal \N__20951\ : std_logic;
signal \N__20948\ : std_logic;
signal \N__20945\ : std_logic;
signal \N__20942\ : std_logic;
signal \N__20939\ : std_logic;
signal \N__20936\ : std_logic;
signal \N__20933\ : std_logic;
signal \N__20930\ : std_logic;
signal \N__20927\ : std_logic;
signal \N__20924\ : std_logic;
signal \N__20921\ : std_logic;
signal \N__20918\ : std_logic;
signal \N__20917\ : std_logic;
signal \N__20914\ : std_logic;
signal \N__20911\ : std_logic;
signal \N__20906\ : std_logic;
signal \N__20903\ : std_logic;
signal \N__20900\ : std_logic;
signal \N__20897\ : std_logic;
signal \N__20894\ : std_logic;
signal \N__20891\ : std_logic;
signal \N__20888\ : std_logic;
signal \N__20885\ : std_logic;
signal \N__20882\ : std_logic;
signal \N__20879\ : std_logic;
signal \N__20876\ : std_logic;
signal \N__20873\ : std_logic;
signal \N__20870\ : std_logic;
signal \N__20867\ : std_logic;
signal \N__20864\ : std_logic;
signal \N__20861\ : std_logic;
signal \N__20858\ : std_logic;
signal \N__20855\ : std_logic;
signal \N__20852\ : std_logic;
signal \N__20849\ : std_logic;
signal \N__20846\ : std_logic;
signal \N__20843\ : std_logic;
signal \N__20840\ : std_logic;
signal \N__20837\ : std_logic;
signal \N__20834\ : std_logic;
signal \N__20831\ : std_logic;
signal \N__20830\ : std_logic;
signal \N__20829\ : std_logic;
signal \N__20826\ : std_logic;
signal \N__20823\ : std_logic;
signal \N__20820\ : std_logic;
signal \N__20817\ : std_logic;
signal \N__20814\ : std_logic;
signal \N__20811\ : std_logic;
signal \N__20804\ : std_logic;
signal \N__20803\ : std_logic;
signal \N__20800\ : std_logic;
signal \N__20797\ : std_logic;
signal \N__20796\ : std_logic;
signal \N__20793\ : std_logic;
signal \N__20790\ : std_logic;
signal \N__20787\ : std_logic;
signal \N__20782\ : std_logic;
signal \N__20779\ : std_logic;
signal \N__20776\ : std_logic;
signal \N__20773\ : std_logic;
signal \N__20768\ : std_logic;
signal \N__20767\ : std_logic;
signal \N__20764\ : std_logic;
signal \N__20763\ : std_logic;
signal \N__20760\ : std_logic;
signal \N__20757\ : std_logic;
signal \N__20754\ : std_logic;
signal \N__20751\ : std_logic;
signal \N__20748\ : std_logic;
signal \N__20745\ : std_logic;
signal \N__20742\ : std_logic;
signal \N__20737\ : std_logic;
signal \N__20734\ : std_logic;
signal \N__20731\ : std_logic;
signal \N__20726\ : std_logic;
signal \N__20723\ : std_logic;
signal \N__20720\ : std_logic;
signal \N__20717\ : std_logic;
signal \N__20714\ : std_logic;
signal \N__20711\ : std_logic;
signal \N__20708\ : std_logic;
signal \N__20705\ : std_logic;
signal \N__20702\ : std_logic;
signal \N__20699\ : std_logic;
signal \N__20696\ : std_logic;
signal \N__20693\ : std_logic;
signal \N__20692\ : std_logic;
signal \N__20689\ : std_logic;
signal \N__20688\ : std_logic;
signal \N__20685\ : std_logic;
signal \N__20682\ : std_logic;
signal \N__20679\ : std_logic;
signal \N__20674\ : std_logic;
signal \N__20671\ : std_logic;
signal \N__20666\ : std_logic;
signal \N__20663\ : std_logic;
signal \N__20660\ : std_logic;
signal \N__20657\ : std_logic;
signal \N__20654\ : std_logic;
signal \N__20651\ : std_logic;
signal \N__20648\ : std_logic;
signal \N__20647\ : std_logic;
signal \N__20644\ : std_logic;
signal \N__20643\ : std_logic;
signal \N__20640\ : std_logic;
signal \N__20637\ : std_logic;
signal \N__20634\ : std_logic;
signal \N__20631\ : std_logic;
signal \N__20626\ : std_logic;
signal \N__20623\ : std_logic;
signal \N__20620\ : std_logic;
signal \N__20615\ : std_logic;
signal \N__20612\ : std_logic;
signal \N__20611\ : std_logic;
signal \N__20610\ : std_logic;
signal \N__20609\ : std_logic;
signal \N__20608\ : std_logic;
signal \N__20607\ : std_logic;
signal \N__20606\ : std_logic;
signal \N__20603\ : std_logic;
signal \N__20600\ : std_logic;
signal \N__20599\ : std_logic;
signal \N__20598\ : std_logic;
signal \N__20597\ : std_logic;
signal \N__20596\ : std_logic;
signal \N__20595\ : std_logic;
signal \N__20592\ : std_logic;
signal \N__20589\ : std_logic;
signal \N__20588\ : std_logic;
signal \N__20587\ : std_logic;
signal \N__20586\ : std_logic;
signal \N__20585\ : std_logic;
signal \N__20582\ : std_logic;
signal \N__20581\ : std_logic;
signal \N__20580\ : std_logic;
signal \N__20579\ : std_logic;
signal \N__20578\ : std_logic;
signal \N__20573\ : std_logic;
signal \N__20570\ : std_logic;
signal \N__20567\ : std_logic;
signal \N__20564\ : std_logic;
signal \N__20561\ : std_logic;
signal \N__20558\ : std_logic;
signal \N__20557\ : std_logic;
signal \N__20554\ : std_logic;
signal \N__20551\ : std_logic;
signal \N__20544\ : std_logic;
signal \N__20539\ : std_logic;
signal \N__20532\ : std_logic;
signal \N__20527\ : std_logic;
signal \N__20524\ : std_logic;
signal \N__20519\ : std_logic;
signal \N__20516\ : std_logic;
signal \N__20507\ : std_logic;
signal \N__20486\ : std_logic;
signal \N__20483\ : std_logic;
signal \N__20482\ : std_logic;
signal \N__20479\ : std_logic;
signal \N__20476\ : std_logic;
signal \N__20473\ : std_logic;
signal \N__20470\ : std_logic;
signal \N__20469\ : std_logic;
signal \N__20466\ : std_logic;
signal \N__20463\ : std_logic;
signal \N__20460\ : std_logic;
signal \N__20453\ : std_logic;
signal \N__20450\ : std_logic;
signal \N__20449\ : std_logic;
signal \N__20446\ : std_logic;
signal \N__20443\ : std_logic;
signal \N__20438\ : std_logic;
signal \N__20437\ : std_logic;
signal \N__20434\ : std_logic;
signal \N__20431\ : std_logic;
signal \N__20426\ : std_logic;
signal \N__20425\ : std_logic;
signal \N__20422\ : std_logic;
signal \N__20419\ : std_logic;
signal \N__20416\ : std_logic;
signal \N__20415\ : std_logic;
signal \N__20412\ : std_logic;
signal \N__20409\ : std_logic;
signal \N__20406\ : std_logic;
signal \N__20399\ : std_logic;
signal \N__20396\ : std_logic;
signal \N__20393\ : std_logic;
signal \N__20390\ : std_logic;
signal \N__20387\ : std_logic;
signal \N__20386\ : std_logic;
signal \N__20385\ : std_logic;
signal \N__20382\ : std_logic;
signal \N__20379\ : std_logic;
signal \N__20376\ : std_logic;
signal \N__20369\ : std_logic;
signal \N__20366\ : std_logic;
signal \N__20363\ : std_logic;
signal \N__20360\ : std_logic;
signal \N__20357\ : std_logic;
signal \N__20354\ : std_logic;
signal \N__20353\ : std_logic;
signal \N__20352\ : std_logic;
signal \N__20349\ : std_logic;
signal \N__20346\ : std_logic;
signal \N__20343\ : std_logic;
signal \N__20340\ : std_logic;
signal \N__20337\ : std_logic;
signal \N__20334\ : std_logic;
signal \N__20331\ : std_logic;
signal \N__20328\ : std_logic;
signal \N__20321\ : std_logic;
signal \N__20318\ : std_logic;
signal \N__20315\ : std_logic;
signal \N__20312\ : std_logic;
signal \N__20309\ : std_logic;
signal \N__20306\ : std_logic;
signal \N__20303\ : std_logic;
signal \N__20300\ : std_logic;
signal \N__20297\ : std_logic;
signal \N__20294\ : std_logic;
signal \N__20291\ : std_logic;
signal \N__20288\ : std_logic;
signal \N__20285\ : std_logic;
signal \N__20282\ : std_logic;
signal \N__20281\ : std_logic;
signal \N__20278\ : std_logic;
signal \N__20275\ : std_logic;
signal \N__20274\ : std_logic;
signal \N__20269\ : std_logic;
signal \N__20266\ : std_logic;
signal \N__20263\ : std_logic;
signal \N__20260\ : std_logic;
signal \N__20257\ : std_logic;
signal \N__20254\ : std_logic;
signal \N__20249\ : std_logic;
signal \N__20248\ : std_logic;
signal \N__20245\ : std_logic;
signal \N__20244\ : std_logic;
signal \N__20241\ : std_logic;
signal \N__20238\ : std_logic;
signal \N__20235\ : std_logic;
signal \N__20230\ : std_logic;
signal \N__20227\ : std_logic;
signal \N__20224\ : std_logic;
signal \N__20219\ : std_logic;
signal \N__20216\ : std_logic;
signal \N__20213\ : std_logic;
signal \N__20210\ : std_logic;
signal \N__20207\ : std_logic;
signal \N__20206\ : std_logic;
signal \N__20203\ : std_logic;
signal \N__20200\ : std_logic;
signal \N__20197\ : std_logic;
signal \N__20194\ : std_logic;
signal \N__20189\ : std_logic;
signal \N__20186\ : std_logic;
signal \N__20183\ : std_logic;
signal \N__20180\ : std_logic;
signal \N__20177\ : std_logic;
signal \N__20174\ : std_logic;
signal \N__20171\ : std_logic;
signal \N__20168\ : std_logic;
signal \N__20165\ : std_logic;
signal \N__20162\ : std_logic;
signal \N__20159\ : std_logic;
signal \N__20156\ : std_logic;
signal \N__20155\ : std_logic;
signal \N__20152\ : std_logic;
signal \N__20151\ : std_logic;
signal \N__20148\ : std_logic;
signal \N__20145\ : std_logic;
signal \N__20142\ : std_logic;
signal \N__20139\ : std_logic;
signal \N__20132\ : std_logic;
signal \N__20131\ : std_logic;
signal \N__20130\ : std_logic;
signal \N__20127\ : std_logic;
signal \N__20124\ : std_logic;
signal \N__20121\ : std_logic;
signal \N__20118\ : std_logic;
signal \N__20115\ : std_logic;
signal \N__20112\ : std_logic;
signal \N__20107\ : std_logic;
signal \N__20104\ : std_logic;
signal \N__20101\ : std_logic;
signal \N__20096\ : std_logic;
signal \N__20093\ : std_logic;
signal \N__20090\ : std_logic;
signal \N__20087\ : std_logic;
signal \N__20084\ : std_logic;
signal \N__20081\ : std_logic;
signal \N__20078\ : std_logic;
signal \N__20075\ : std_logic;
signal \N__20072\ : std_logic;
signal \N__20071\ : std_logic;
signal \N__20070\ : std_logic;
signal \N__20067\ : std_logic;
signal \N__20064\ : std_logic;
signal \N__20061\ : std_logic;
signal \N__20056\ : std_logic;
signal \N__20053\ : std_logic;
signal \N__20050\ : std_logic;
signal \N__20045\ : std_logic;
signal \N__20042\ : std_logic;
signal \N__20039\ : std_logic;
signal \N__20036\ : std_logic;
signal \N__20033\ : std_logic;
signal \N__20030\ : std_logic;
signal \N__20027\ : std_logic;
signal \N__20024\ : std_logic;
signal \N__20023\ : std_logic;
signal \N__20022\ : std_logic;
signal \N__20019\ : std_logic;
signal \N__20016\ : std_logic;
signal \N__20013\ : std_logic;
signal \N__20006\ : std_logic;
signal \N__20003\ : std_logic;
signal \N__20000\ : std_logic;
signal \N__19997\ : std_logic;
signal \N__19996\ : std_logic;
signal \N__19993\ : std_logic;
signal \N__19990\ : std_logic;
signal \N__19987\ : std_logic;
signal \N__19984\ : std_logic;
signal \N__19983\ : std_logic;
signal \N__19980\ : std_logic;
signal \N__19977\ : std_logic;
signal \N__19974\ : std_logic;
signal \N__19967\ : std_logic;
signal \N__19966\ : std_logic;
signal \N__19965\ : std_logic;
signal \N__19964\ : std_logic;
signal \N__19963\ : std_logic;
signal \N__19960\ : std_logic;
signal \N__19959\ : std_logic;
signal \N__19958\ : std_logic;
signal \N__19955\ : std_logic;
signal \N__19954\ : std_logic;
signal \N__19953\ : std_logic;
signal \N__19952\ : std_logic;
signal \N__19949\ : std_logic;
signal \N__19948\ : std_logic;
signal \N__19945\ : std_logic;
signal \N__19944\ : std_logic;
signal \N__19943\ : std_logic;
signal \N__19936\ : std_logic;
signal \N__19935\ : std_logic;
signal \N__19934\ : std_logic;
signal \N__19931\ : std_logic;
signal \N__19930\ : std_logic;
signal \N__19925\ : std_logic;
signal \N__19920\ : std_logic;
signal \N__19915\ : std_logic;
signal \N__19908\ : std_logic;
signal \N__19905\ : std_logic;
signal \N__19902\ : std_logic;
signal \N__19895\ : std_logic;
signal \N__19892\ : std_logic;
signal \N__19877\ : std_logic;
signal \N__19874\ : std_logic;
signal \N__19873\ : std_logic;
signal \N__19870\ : std_logic;
signal \N__19869\ : std_logic;
signal \N__19866\ : std_logic;
signal \N__19863\ : std_logic;
signal \N__19860\ : std_logic;
signal \N__19853\ : std_logic;
signal \N__19850\ : std_logic;
signal \N__19847\ : std_logic;
signal \N__19844\ : std_logic;
signal \N__19843\ : std_logic;
signal \N__19842\ : std_logic;
signal \N__19839\ : std_logic;
signal \N__19836\ : std_logic;
signal \N__19833\ : std_logic;
signal \N__19826\ : std_logic;
signal \N__19823\ : std_logic;
signal \N__19820\ : std_logic;
signal \N__19817\ : std_logic;
signal \N__19814\ : std_logic;
signal \N__19811\ : std_logic;
signal \N__19808\ : std_logic;
signal \N__19805\ : std_logic;
signal \N__19802\ : std_logic;
signal \N__19801\ : std_logic;
signal \N__19798\ : std_logic;
signal \N__19795\ : std_logic;
signal \N__19792\ : std_logic;
signal \N__19787\ : std_logic;
signal \N__19784\ : std_logic;
signal \N__19783\ : std_logic;
signal \N__19780\ : std_logic;
signal \N__19777\ : std_logic;
signal \N__19774\ : std_logic;
signal \N__19769\ : std_logic;
signal \N__19766\ : std_logic;
signal \N__19763\ : std_logic;
signal \N__19760\ : std_logic;
signal \N__19757\ : std_logic;
signal \N__19754\ : std_logic;
signal \N__19751\ : std_logic;
signal \N__19748\ : std_logic;
signal \N__19747\ : std_logic;
signal \N__19744\ : std_logic;
signal \N__19741\ : std_logic;
signal \N__19736\ : std_logic;
signal \N__19733\ : std_logic;
signal \N__19732\ : std_logic;
signal \N__19731\ : std_logic;
signal \N__19728\ : std_logic;
signal \N__19725\ : std_logic;
signal \N__19722\ : std_logic;
signal \N__19719\ : std_logic;
signal \N__19712\ : std_logic;
signal \N__19709\ : std_logic;
signal \N__19706\ : std_logic;
signal \N__19703\ : std_logic;
signal \N__19702\ : std_logic;
signal \N__19701\ : std_logic;
signal \N__19698\ : std_logic;
signal \N__19693\ : std_logic;
signal \N__19690\ : std_logic;
signal \N__19685\ : std_logic;
signal \N__19682\ : std_logic;
signal \N__19679\ : std_logic;
signal \N__19676\ : std_logic;
signal \N__19673\ : std_logic;
signal \N__19670\ : std_logic;
signal \N__19669\ : std_logic;
signal \N__19668\ : std_logic;
signal \N__19665\ : std_logic;
signal \N__19662\ : std_logic;
signal \N__19659\ : std_logic;
signal \N__19656\ : std_logic;
signal \N__19651\ : std_logic;
signal \N__19646\ : std_logic;
signal \N__19643\ : std_logic;
signal \N__19640\ : std_logic;
signal \N__19637\ : std_logic;
signal \N__19634\ : std_logic;
signal \N__19633\ : std_logic;
signal \N__19630\ : std_logic;
signal \N__19627\ : std_logic;
signal \N__19624\ : std_logic;
signal \N__19621\ : std_logic;
signal \N__19616\ : std_logic;
signal \N__19615\ : std_logic;
signal \N__19612\ : std_logic;
signal \N__19609\ : std_logic;
signal \N__19604\ : std_logic;
signal \N__19603\ : std_logic;
signal \N__19600\ : std_logic;
signal \N__19597\ : std_logic;
signal \N__19594\ : std_logic;
signal \N__19589\ : std_logic;
signal \N__19586\ : std_logic;
signal \N__19583\ : std_logic;
signal \N__19580\ : std_logic;
signal \N__19577\ : std_logic;
signal \N__19574\ : std_logic;
signal \N__19571\ : std_logic;
signal \N__19568\ : std_logic;
signal \N__19565\ : std_logic;
signal \N__19562\ : std_logic;
signal \N__19559\ : std_logic;
signal \N__19556\ : std_logic;
signal \N__19553\ : std_logic;
signal \N__19550\ : std_logic;
signal \N__19549\ : std_logic;
signal \N__19546\ : std_logic;
signal \N__19543\ : std_logic;
signal \N__19540\ : std_logic;
signal \N__19539\ : std_logic;
signal \N__19536\ : std_logic;
signal \N__19533\ : std_logic;
signal \N__19530\ : std_logic;
signal \N__19523\ : std_logic;
signal \N__19520\ : std_logic;
signal \N__19519\ : std_logic;
signal \N__19516\ : std_logic;
signal \N__19513\ : std_logic;
signal \N__19512\ : std_logic;
signal \N__19509\ : std_logic;
signal \N__19506\ : std_logic;
signal \N__19503\ : std_logic;
signal \N__19500\ : std_logic;
signal \N__19497\ : std_logic;
signal \N__19494\ : std_logic;
signal \N__19487\ : std_logic;
signal \N__19484\ : std_logic;
signal \N__19483\ : std_logic;
signal \N__19480\ : std_logic;
signal \N__19477\ : std_logic;
signal \N__19474\ : std_logic;
signal \N__19471\ : std_logic;
signal \N__19466\ : std_logic;
signal \N__19463\ : std_logic;
signal \N__19460\ : std_logic;
signal \N__19457\ : std_logic;
signal \N__19454\ : std_logic;
signal \N__19451\ : std_logic;
signal \N__19448\ : std_logic;
signal \N__19445\ : std_logic;
signal \N__19442\ : std_logic;
signal \N__19439\ : std_logic;
signal \N__19438\ : std_logic;
signal \N__19435\ : std_logic;
signal \N__19432\ : std_logic;
signal \N__19431\ : std_logic;
signal \N__19428\ : std_logic;
signal \N__19425\ : std_logic;
signal \N__19422\ : std_logic;
signal \N__19419\ : std_logic;
signal \N__19416\ : std_logic;
signal \N__19409\ : std_logic;
signal \N__19406\ : std_logic;
signal \N__19403\ : std_logic;
signal \N__19400\ : std_logic;
signal \N__19399\ : std_logic;
signal \N__19396\ : std_logic;
signal \N__19395\ : std_logic;
signal \N__19392\ : std_logic;
signal \N__19389\ : std_logic;
signal \N__19386\ : std_logic;
signal \N__19383\ : std_logic;
signal \N__19378\ : std_logic;
signal \N__19373\ : std_logic;
signal \N__19370\ : std_logic;
signal \N__19367\ : std_logic;
signal \N__19364\ : std_logic;
signal \N__19361\ : std_logic;
signal \N__19360\ : std_logic;
signal \N__19357\ : std_logic;
signal \N__19354\ : std_logic;
signal \N__19353\ : std_logic;
signal \N__19350\ : std_logic;
signal \N__19347\ : std_logic;
signal \N__19344\ : std_logic;
signal \N__19337\ : std_logic;
signal \N__19336\ : std_logic;
signal \N__19333\ : std_logic;
signal \N__19330\ : std_logic;
signal \N__19327\ : std_logic;
signal \N__19324\ : std_logic;
signal \N__19321\ : std_logic;
signal \N__19316\ : std_logic;
signal \N__19313\ : std_logic;
signal \N__19310\ : std_logic;
signal \N__19309\ : std_logic;
signal \N__19308\ : std_logic;
signal \N__19305\ : std_logic;
signal \N__19302\ : std_logic;
signal \N__19297\ : std_logic;
signal \N__19292\ : std_logic;
signal \N__19289\ : std_logic;
signal \N__19286\ : std_logic;
signal \N__19283\ : std_logic;
signal \N__19280\ : std_logic;
signal \N__19277\ : std_logic;
signal \N__19274\ : std_logic;
signal \N__19271\ : std_logic;
signal \N__19268\ : std_logic;
signal \N__19267\ : std_logic;
signal \N__19266\ : std_logic;
signal \N__19263\ : std_logic;
signal \N__19262\ : std_logic;
signal \N__19261\ : std_logic;
signal \N__19260\ : std_logic;
signal \N__19259\ : std_logic;
signal \N__19258\ : std_logic;
signal \N__19257\ : std_logic;
signal \N__19256\ : std_logic;
signal \N__19255\ : std_logic;
signal \N__19254\ : std_logic;
signal \N__19253\ : std_logic;
signal \N__19250\ : std_logic;
signal \N__19247\ : std_logic;
signal \N__19244\ : std_logic;
signal \N__19241\ : std_logic;
signal \N__19240\ : std_logic;
signal \N__19239\ : std_logic;
signal \N__19236\ : std_logic;
signal \N__19233\ : std_logic;
signal \N__19230\ : std_logic;
signal \N__19227\ : std_logic;
signal \N__19226\ : std_logic;
signal \N__19225\ : std_logic;
signal \N__19224\ : std_logic;
signal \N__19221\ : std_logic;
signal \N__19218\ : std_logic;
signal \N__19215\ : std_logic;
signal \N__19212\ : std_logic;
signal \N__19211\ : std_logic;
signal \N__19208\ : std_logic;
signal \N__19201\ : std_logic;
signal \N__19194\ : std_logic;
signal \N__19193\ : std_logic;
signal \N__19188\ : std_logic;
signal \N__19179\ : std_logic;
signal \N__19168\ : std_logic;
signal \N__19165\ : std_logic;
signal \N__19162\ : std_logic;
signal \N__19157\ : std_logic;
signal \N__19154\ : std_logic;
signal \N__19139\ : std_logic;
signal \N__19136\ : std_logic;
signal \N__19135\ : std_logic;
signal \N__19132\ : std_logic;
signal \N__19131\ : std_logic;
signal \N__19128\ : std_logic;
signal \N__19125\ : std_logic;
signal \N__19122\ : std_logic;
signal \N__19115\ : std_logic;
signal \N__19112\ : std_logic;
signal \N__19111\ : std_logic;
signal \N__19110\ : std_logic;
signal \N__19107\ : std_logic;
signal \N__19102\ : std_logic;
signal \N__19099\ : std_logic;
signal \N__19094\ : std_logic;
signal \N__19091\ : std_logic;
signal \N__19090\ : std_logic;
signal \N__19089\ : std_logic;
signal \N__19086\ : std_logic;
signal \N__19083\ : std_logic;
signal \N__19080\ : std_logic;
signal \N__19073\ : std_logic;
signal \N__19070\ : std_logic;
signal \N__19067\ : std_logic;
signal \N__19064\ : std_logic;
signal \N__19063\ : std_logic;
signal \N__19062\ : std_logic;
signal \N__19059\ : std_logic;
signal \N__19056\ : std_logic;
signal \N__19053\ : std_logic;
signal \N__19050\ : std_logic;
signal \N__19043\ : std_logic;
signal \N__19040\ : std_logic;
signal \N__19037\ : std_logic;
signal \N__19034\ : std_logic;
signal \N__19031\ : std_logic;
signal \N__19028\ : std_logic;
signal \N__19025\ : std_logic;
signal \N__19022\ : std_logic;
signal \N__19021\ : std_logic;
signal \N__19018\ : std_logic;
signal \N__19017\ : std_logic;
signal \N__19014\ : std_logic;
signal \N__19011\ : std_logic;
signal \N__19008\ : std_logic;
signal \N__19005\ : std_logic;
signal \N__18998\ : std_logic;
signal \N__18995\ : std_logic;
signal \N__18992\ : std_logic;
signal \N__18989\ : std_logic;
signal \N__18986\ : std_logic;
signal \N__18983\ : std_logic;
signal \N__18980\ : std_logic;
signal \N__18979\ : std_logic;
signal \N__18976\ : std_logic;
signal \N__18975\ : std_logic;
signal \N__18972\ : std_logic;
signal \N__18969\ : std_logic;
signal \N__18964\ : std_logic;
signal \N__18959\ : std_logic;
signal \N__18956\ : std_logic;
signal \N__18953\ : std_logic;
signal \N__18950\ : std_logic;
signal \N__18947\ : std_logic;
signal \N__18946\ : std_logic;
signal \N__18945\ : std_logic;
signal \N__18942\ : std_logic;
signal \N__18937\ : std_logic;
signal \N__18934\ : std_logic;
signal \N__18929\ : std_logic;
signal \N__18926\ : std_logic;
signal \N__18923\ : std_logic;
signal \N__18920\ : std_logic;
signal \N__18917\ : std_logic;
signal \N__18914\ : std_logic;
signal \N__18911\ : std_logic;
signal \N__18910\ : std_logic;
signal \N__18907\ : std_logic;
signal \N__18906\ : std_logic;
signal \N__18903\ : std_logic;
signal \N__18900\ : std_logic;
signal \N__18897\ : std_logic;
signal \N__18894\ : std_logic;
signal \N__18887\ : std_logic;
signal \N__18884\ : std_logic;
signal \N__18881\ : std_logic;
signal \N__18878\ : std_logic;
signal \N__18875\ : std_logic;
signal \N__18872\ : std_logic;
signal \N__18869\ : std_logic;
signal \N__18866\ : std_logic;
signal \N__18863\ : std_logic;
signal \N__18862\ : std_logic;
signal \N__18859\ : std_logic;
signal \N__18856\ : std_logic;
signal \N__18855\ : std_logic;
signal \N__18852\ : std_logic;
signal \N__18849\ : std_logic;
signal \N__18846\ : std_logic;
signal \N__18839\ : std_logic;
signal \N__18836\ : std_logic;
signal \N__18833\ : std_logic;
signal \N__18830\ : std_logic;
signal \N__18827\ : std_logic;
signal \N__18824\ : std_logic;
signal \N__18821\ : std_logic;
signal \N__18818\ : std_logic;
signal \N__18815\ : std_logic;
signal \N__18812\ : std_logic;
signal \N__18809\ : std_logic;
signal \N__18806\ : std_logic;
signal \N__18805\ : std_logic;
signal \N__18804\ : std_logic;
signal \N__18801\ : std_logic;
signal \N__18796\ : std_logic;
signal \N__18791\ : std_logic;
signal \N__18788\ : std_logic;
signal \N__18785\ : std_logic;
signal \N__18782\ : std_logic;
signal \N__18781\ : std_logic;
signal \N__18778\ : std_logic;
signal \N__18777\ : std_logic;
signal \N__18774\ : std_logic;
signal \N__18771\ : std_logic;
signal \N__18768\ : std_logic;
signal \N__18761\ : std_logic;
signal \N__18758\ : std_logic;
signal \N__18757\ : std_logic;
signal \N__18756\ : std_logic;
signal \N__18753\ : std_logic;
signal \N__18750\ : std_logic;
signal \N__18747\ : std_logic;
signal \N__18744\ : std_logic;
signal \N__18739\ : std_logic;
signal \N__18736\ : std_logic;
signal \N__18731\ : std_logic;
signal \N__18728\ : std_logic;
signal \N__18725\ : std_logic;
signal \N__18722\ : std_logic;
signal \N__18719\ : std_logic;
signal \N__18718\ : std_logic;
signal \N__18717\ : std_logic;
signal \N__18714\ : std_logic;
signal \N__18709\ : std_logic;
signal \N__18706\ : std_logic;
signal \N__18701\ : std_logic;
signal \N__18698\ : std_logic;
signal \N__18695\ : std_logic;
signal \N__18694\ : std_logic;
signal \N__18693\ : std_logic;
signal \N__18690\ : std_logic;
signal \N__18687\ : std_logic;
signal \N__18684\ : std_logic;
signal \N__18677\ : std_logic;
signal \N__18674\ : std_logic;
signal \N__18671\ : std_logic;
signal \N__18668\ : std_logic;
signal \N__18665\ : std_logic;
signal \N__18662\ : std_logic;
signal \N__18659\ : std_logic;
signal \N__18656\ : std_logic;
signal \N__18655\ : std_logic;
signal \N__18654\ : std_logic;
signal \N__18649\ : std_logic;
signal \N__18646\ : std_logic;
signal \N__18643\ : std_logic;
signal \N__18640\ : std_logic;
signal \N__18635\ : std_logic;
signal \N__18632\ : std_logic;
signal \N__18629\ : std_logic;
signal \N__18626\ : std_logic;
signal \N__18623\ : std_logic;
signal \N__18622\ : std_logic;
signal \N__18621\ : std_logic;
signal \N__18616\ : std_logic;
signal \N__18613\ : std_logic;
signal \N__18610\ : std_logic;
signal \N__18607\ : std_logic;
signal \N__18604\ : std_logic;
signal \N__18601\ : std_logic;
signal \N__18596\ : std_logic;
signal \N__18593\ : std_logic;
signal \N__18590\ : std_logic;
signal \N__18587\ : std_logic;
signal \N__18586\ : std_logic;
signal \N__18583\ : std_logic;
signal \N__18580\ : std_logic;
signal \N__18577\ : std_logic;
signal \N__18572\ : std_logic;
signal \N__18569\ : std_logic;
signal \N__18566\ : std_logic;
signal \N__18563\ : std_logic;
signal \N__18560\ : std_logic;
signal \N__18557\ : std_logic;
signal \N__18554\ : std_logic;
signal \N__18551\ : std_logic;
signal \N__18550\ : std_logic;
signal \N__18547\ : std_logic;
signal \N__18546\ : std_logic;
signal \N__18543\ : std_logic;
signal \N__18540\ : std_logic;
signal \N__18537\ : std_logic;
signal \N__18534\ : std_logic;
signal \N__18527\ : std_logic;
signal \N__18524\ : std_logic;
signal \N__18521\ : std_logic;
signal \N__18518\ : std_logic;
signal \N__18515\ : std_logic;
signal \N__18512\ : std_logic;
signal \N__18511\ : std_logic;
signal \N__18508\ : std_logic;
signal \N__18505\ : std_logic;
signal \N__18504\ : std_logic;
signal \N__18501\ : std_logic;
signal \N__18498\ : std_logic;
signal \N__18495\ : std_logic;
signal \N__18490\ : std_logic;
signal \N__18485\ : std_logic;
signal \N__18482\ : std_logic;
signal \N__18479\ : std_logic;
signal \N__18476\ : std_logic;
signal \N__18473\ : std_logic;
signal \N__18472\ : std_logic;
signal \N__18469\ : std_logic;
signal \N__18466\ : std_logic;
signal \N__18463\ : std_logic;
signal \N__18460\ : std_logic;
signal \N__18459\ : std_logic;
signal \N__18454\ : std_logic;
signal \N__18451\ : std_logic;
signal \N__18446\ : std_logic;
signal \N__18443\ : std_logic;
signal \N__18440\ : std_logic;
signal \N__18437\ : std_logic;
signal \N__18434\ : std_logic;
signal \N__18433\ : std_logic;
signal \N__18430\ : std_logic;
signal \N__18427\ : std_logic;
signal \N__18424\ : std_logic;
signal \N__18421\ : std_logic;
signal \N__18416\ : std_logic;
signal \N__18413\ : std_logic;
signal \N__18410\ : std_logic;
signal \N__18409\ : std_logic;
signal \N__18406\ : std_logic;
signal \N__18403\ : std_logic;
signal \N__18402\ : std_logic;
signal \N__18397\ : std_logic;
signal \N__18394\ : std_logic;
signal \N__18389\ : std_logic;
signal \N__18386\ : std_logic;
signal \N__18383\ : std_logic;
signal \N__18382\ : std_logic;
signal \N__18379\ : std_logic;
signal \N__18376\ : std_logic;
signal \N__18373\ : std_logic;
signal \N__18370\ : std_logic;
signal \N__18369\ : std_logic;
signal \N__18366\ : std_logic;
signal \N__18363\ : std_logic;
signal \N__18360\ : std_logic;
signal \N__18353\ : std_logic;
signal \N__18350\ : std_logic;
signal \N__18347\ : std_logic;
signal \N__18344\ : std_logic;
signal \N__18341\ : std_logic;
signal \N__18340\ : std_logic;
signal \N__18339\ : std_logic;
signal \N__18338\ : std_logic;
signal \N__18337\ : std_logic;
signal \N__18336\ : std_logic;
signal \N__18333\ : std_logic;
signal \N__18332\ : std_logic;
signal \N__18331\ : std_logic;
signal \N__18328\ : std_logic;
signal \N__18327\ : std_logic;
signal \N__18326\ : std_logic;
signal \N__18323\ : std_logic;
signal \N__18320\ : std_logic;
signal \N__18319\ : std_logic;
signal \N__18316\ : std_logic;
signal \N__18315\ : std_logic;
signal \N__18314\ : std_logic;
signal \N__18313\ : std_logic;
signal \N__18304\ : std_logic;
signal \N__18299\ : std_logic;
signal \N__18296\ : std_logic;
signal \N__18285\ : std_logic;
signal \N__18282\ : std_logic;
signal \N__18279\ : std_logic;
signal \N__18278\ : std_logic;
signal \N__18273\ : std_logic;
signal \N__18268\ : std_logic;
signal \N__18261\ : std_logic;
signal \N__18258\ : std_logic;
signal \N__18251\ : std_logic;
signal \N__18248\ : std_logic;
signal \N__18247\ : std_logic;
signal \N__18244\ : std_logic;
signal \N__18241\ : std_logic;
signal \N__18236\ : std_logic;
signal \N__18233\ : std_logic;
signal \N__18230\ : std_logic;
signal \N__18227\ : std_logic;
signal \N__18224\ : std_logic;
signal \N__18221\ : std_logic;
signal \N__18218\ : std_logic;
signal \N__18215\ : std_logic;
signal \N__18212\ : std_logic;
signal \N__18209\ : std_logic;
signal \N__18206\ : std_logic;
signal \N__18203\ : std_logic;
signal \N__18202\ : std_logic;
signal \N__18199\ : std_logic;
signal \N__18196\ : std_logic;
signal \N__18193\ : std_logic;
signal \N__18190\ : std_logic;
signal \N__18185\ : std_logic;
signal \N__18182\ : std_logic;
signal \N__18179\ : std_logic;
signal \N__18176\ : std_logic;
signal \N__18173\ : std_logic;
signal \N__18170\ : std_logic;
signal \N__18167\ : std_logic;
signal \N__18164\ : std_logic;
signal \N__18161\ : std_logic;
signal \N__18158\ : std_logic;
signal \N__18155\ : std_logic;
signal \N__18152\ : std_logic;
signal \N__18149\ : std_logic;
signal \N__18146\ : std_logic;
signal \N__18143\ : std_logic;
signal \N__18140\ : std_logic;
signal \N__18139\ : std_logic;
signal \N__18136\ : std_logic;
signal \N__18133\ : std_logic;
signal \N__18132\ : std_logic;
signal \N__18129\ : std_logic;
signal \N__18126\ : std_logic;
signal \N__18123\ : std_logic;
signal \N__18116\ : std_logic;
signal \N__18113\ : std_logic;
signal \N__18110\ : std_logic;
signal \N__18107\ : std_logic;
signal \N__18104\ : std_logic;
signal \N__18101\ : std_logic;
signal \N__18098\ : std_logic;
signal \N__18095\ : std_logic;
signal \N__18094\ : std_logic;
signal \N__18091\ : std_logic;
signal \N__18088\ : std_logic;
signal \N__18085\ : std_logic;
signal \N__18082\ : std_logic;
signal \N__18077\ : std_logic;
signal \N__18074\ : std_logic;
signal \N__18071\ : std_logic;
signal \N__18068\ : std_logic;
signal \N__18065\ : std_logic;
signal \N__18062\ : std_logic;
signal \N__18059\ : std_logic;
signal \N__18056\ : std_logic;
signal \N__18053\ : std_logic;
signal \N__18050\ : std_logic;
signal \N__18047\ : std_logic;
signal \N__18044\ : std_logic;
signal \N__18041\ : std_logic;
signal \N__18038\ : std_logic;
signal \N__18035\ : std_logic;
signal \N__18034\ : std_logic;
signal \N__18033\ : std_logic;
signal \N__18030\ : std_logic;
signal \N__18025\ : std_logic;
signal \N__18020\ : std_logic;
signal \N__18017\ : std_logic;
signal \N__18014\ : std_logic;
signal \N__18011\ : std_logic;
signal \N__18008\ : std_logic;
signal \N__18005\ : std_logic;
signal \N__18002\ : std_logic;
signal \N__17999\ : std_logic;
signal \N__17996\ : std_logic;
signal \N__17993\ : std_logic;
signal \N__17990\ : std_logic;
signal \N__17987\ : std_logic;
signal \N__17984\ : std_logic;
signal \N__17981\ : std_logic;
signal \N__17978\ : std_logic;
signal \N__17975\ : std_logic;
signal \N__17972\ : std_logic;
signal \N__17969\ : std_logic;
signal \N__17966\ : std_logic;
signal \N__17963\ : std_logic;
signal \N__17960\ : std_logic;
signal \N__17957\ : std_logic;
signal \N__17954\ : std_logic;
signal \N__17951\ : std_logic;
signal \N__17950\ : std_logic;
signal \N__17947\ : std_logic;
signal \N__17944\ : std_logic;
signal \N__17941\ : std_logic;
signal \N__17938\ : std_logic;
signal \N__17933\ : std_logic;
signal \N__17930\ : std_logic;
signal \N__17927\ : std_logic;
signal \N__17924\ : std_logic;
signal \N__17921\ : std_logic;
signal \N__17918\ : std_logic;
signal \N__17915\ : std_logic;
signal \N__17914\ : std_logic;
signal \N__17911\ : std_logic;
signal \N__17908\ : std_logic;
signal \N__17905\ : std_logic;
signal \N__17900\ : std_logic;
signal \N__17897\ : std_logic;
signal \N__17894\ : std_logic;
signal \N__17891\ : std_logic;
signal \N__17888\ : std_logic;
signal \N__17885\ : std_logic;
signal \N__17882\ : std_logic;
signal \N__17879\ : std_logic;
signal \N__17876\ : std_logic;
signal \N__17873\ : std_logic;
signal \N__17870\ : std_logic;
signal \N__17867\ : std_logic;
signal \N__17864\ : std_logic;
signal \N__17861\ : std_logic;
signal \N__17858\ : std_logic;
signal \N__17855\ : std_logic;
signal \N__17852\ : std_logic;
signal \N__17849\ : std_logic;
signal \N__17846\ : std_logic;
signal \N__17843\ : std_logic;
signal \N__17840\ : std_logic;
signal \N__17837\ : std_logic;
signal \N__17834\ : std_logic;
signal \N__17831\ : std_logic;
signal \N__17828\ : std_logic;
signal \N__17825\ : std_logic;
signal \N__17822\ : std_logic;
signal \N__17819\ : std_logic;
signal \N__17816\ : std_logic;
signal \N__17813\ : std_logic;
signal \N__17810\ : std_logic;
signal \N__17807\ : std_logic;
signal \N__17804\ : std_logic;
signal \N__17801\ : std_logic;
signal \N__17798\ : std_logic;
signal \N__17795\ : std_logic;
signal \N__17792\ : std_logic;
signal \N__17789\ : std_logic;
signal \N__17786\ : std_logic;
signal \N__17783\ : std_logic;
signal \N__17780\ : std_logic;
signal \N__17777\ : std_logic;
signal \N__17774\ : std_logic;
signal \N__17771\ : std_logic;
signal \N__17768\ : std_logic;
signal \N__17765\ : std_logic;
signal \N__17762\ : std_logic;
signal \N__17759\ : std_logic;
signal \N__17756\ : std_logic;
signal \N__17753\ : std_logic;
signal \N__17750\ : std_logic;
signal \N__17747\ : std_logic;
signal \N__17744\ : std_logic;
signal \N__17741\ : std_logic;
signal \N__17738\ : std_logic;
signal \N__17735\ : std_logic;
signal \N__17732\ : std_logic;
signal \N__17729\ : std_logic;
signal \N__17726\ : std_logic;
signal \N__17723\ : std_logic;
signal \N__17720\ : std_logic;
signal \N__17717\ : std_logic;
signal \N__17714\ : std_logic;
signal \N__17713\ : std_logic;
signal \N__17710\ : std_logic;
signal \N__17707\ : std_logic;
signal \N__17706\ : std_logic;
signal \N__17703\ : std_logic;
signal \N__17700\ : std_logic;
signal \N__17697\ : std_logic;
signal \N__17690\ : std_logic;
signal \N__17687\ : std_logic;
signal \N__17684\ : std_logic;
signal \N__17681\ : std_logic;
signal \N__17680\ : std_logic;
signal \N__17677\ : std_logic;
signal \N__17674\ : std_logic;
signal \N__17671\ : std_logic;
signal \N__17668\ : std_logic;
signal \N__17665\ : std_logic;
signal \N__17662\ : std_logic;
signal \N__17657\ : std_logic;
signal \N__17654\ : std_logic;
signal \N__17651\ : std_logic;
signal \N__17648\ : std_logic;
signal \N__17645\ : std_logic;
signal \N__17642\ : std_logic;
signal \N__17639\ : std_logic;
signal \N__17636\ : std_logic;
signal \N__17633\ : std_logic;
signal \N__17630\ : std_logic;
signal \N__17627\ : std_logic;
signal \N__17624\ : std_logic;
signal \N__17621\ : std_logic;
signal \N__17618\ : std_logic;
signal \N__17615\ : std_logic;
signal \N__17612\ : std_logic;
signal \N__17609\ : std_logic;
signal \N__17606\ : std_logic;
signal \N__17603\ : std_logic;
signal \N__17600\ : std_logic;
signal \N__17597\ : std_logic;
signal \N__17594\ : std_logic;
signal \N__17591\ : std_logic;
signal \N__17588\ : std_logic;
signal \N__17585\ : std_logic;
signal \N__17582\ : std_logic;
signal \N__17579\ : std_logic;
signal \N__17576\ : std_logic;
signal \N__17573\ : std_logic;
signal \N__17570\ : std_logic;
signal \N__17567\ : std_logic;
signal \N__17564\ : std_logic;
signal \N__17561\ : std_logic;
signal \N__17558\ : std_logic;
signal \N__17555\ : std_logic;
signal \N__17552\ : std_logic;
signal \N__17549\ : std_logic;
signal \N__17546\ : std_logic;
signal \N__17543\ : std_logic;
signal \N__17540\ : std_logic;
signal \N__17537\ : std_logic;
signal \N__17534\ : std_logic;
signal \N__17531\ : std_logic;
signal \N__17528\ : std_logic;
signal \N__17525\ : std_logic;
signal \N__17522\ : std_logic;
signal \N__17519\ : std_logic;
signal \N__17518\ : std_logic;
signal \N__17515\ : std_logic;
signal \N__17512\ : std_logic;
signal \N__17509\ : std_logic;
signal \N__17506\ : std_logic;
signal \N__17501\ : std_logic;
signal \N__17498\ : std_logic;
signal \N__17495\ : std_logic;
signal \N__17492\ : std_logic;
signal \N__17491\ : std_logic;
signal \N__17488\ : std_logic;
signal \N__17487\ : std_logic;
signal \N__17484\ : std_logic;
signal \N__17481\ : std_logic;
signal \N__17478\ : std_logic;
signal \N__17473\ : std_logic;
signal \N__17470\ : std_logic;
signal \N__17465\ : std_logic;
signal \N__17462\ : std_logic;
signal \N__17459\ : std_logic;
signal \N__17458\ : std_logic;
signal \N__17457\ : std_logic;
signal \N__17454\ : std_logic;
signal \N__17451\ : std_logic;
signal \N__17448\ : std_logic;
signal \N__17441\ : std_logic;
signal \N__17438\ : std_logic;
signal \N__17437\ : std_logic;
signal \N__17434\ : std_logic;
signal \N__17431\ : std_logic;
signal \N__17430\ : std_logic;
signal \N__17427\ : std_logic;
signal \N__17424\ : std_logic;
signal \N__17421\ : std_logic;
signal \N__17416\ : std_logic;
signal \N__17411\ : std_logic;
signal \N__17408\ : std_logic;
signal \N__17405\ : std_logic;
signal \N__17402\ : std_logic;
signal \N__17399\ : std_logic;
signal \N__17396\ : std_logic;
signal \N__17393\ : std_logic;
signal \N__17390\ : std_logic;
signal \N__17389\ : std_logic;
signal \N__17386\ : std_logic;
signal \N__17383\ : std_logic;
signal \N__17380\ : std_logic;
signal \N__17377\ : std_logic;
signal \N__17376\ : std_logic;
signal \N__17371\ : std_logic;
signal \N__17368\ : std_logic;
signal \N__17363\ : std_logic;
signal \N__17362\ : std_logic;
signal \N__17359\ : std_logic;
signal \N__17356\ : std_logic;
signal \N__17353\ : std_logic;
signal \N__17350\ : std_logic;
signal \N__17345\ : std_logic;
signal \N__17342\ : std_logic;
signal \N__17339\ : std_logic;
signal \N__17336\ : std_logic;
signal \N__17333\ : std_logic;
signal \N__17330\ : std_logic;
signal \N__17327\ : std_logic;
signal \N__17324\ : std_logic;
signal \N__17323\ : std_logic;
signal \N__17320\ : std_logic;
signal \N__17319\ : std_logic;
signal \N__17316\ : std_logic;
signal \N__17313\ : std_logic;
signal \N__17310\ : std_logic;
signal \N__17303\ : std_logic;
signal \N__17300\ : std_logic;
signal \N__17297\ : std_logic;
signal \N__17294\ : std_logic;
signal \N__17291\ : std_logic;
signal \N__17288\ : std_logic;
signal \N__17285\ : std_logic;
signal \N__17282\ : std_logic;
signal \N__17279\ : std_logic;
signal \N__17276\ : std_logic;
signal \N__17273\ : std_logic;
signal \N__17270\ : std_logic;
signal \N__17267\ : std_logic;
signal \N__17264\ : std_logic;
signal \N__17261\ : std_logic;
signal \N__17258\ : std_logic;
signal \N__17255\ : std_logic;
signal \N__17254\ : std_logic;
signal \N__17251\ : std_logic;
signal \N__17248\ : std_logic;
signal \N__17247\ : std_logic;
signal \N__17244\ : std_logic;
signal \N__17241\ : std_logic;
signal \N__17238\ : std_logic;
signal \N__17231\ : std_logic;
signal \N__17228\ : std_logic;
signal \N__17225\ : std_logic;
signal \N__17222\ : std_logic;
signal \N__17221\ : std_logic;
signal \N__17220\ : std_logic;
signal \N__17219\ : std_logic;
signal \N__17218\ : std_logic;
signal \N__17217\ : std_logic;
signal \N__17214\ : std_logic;
signal \N__17213\ : std_logic;
signal \N__17212\ : std_logic;
signal \N__17211\ : std_logic;
signal \N__17210\ : std_logic;
signal \N__17207\ : std_logic;
signal \N__17204\ : std_logic;
signal \N__17203\ : std_logic;
signal \N__17202\ : std_logic;
signal \N__17199\ : std_logic;
signal \N__17198\ : std_logic;
signal \N__17195\ : std_logic;
signal \N__17194\ : std_logic;
signal \N__17191\ : std_logic;
signal \N__17188\ : std_logic;
signal \N__17185\ : std_logic;
signal \N__17180\ : std_logic;
signal \N__17171\ : std_logic;
signal \N__17160\ : std_logic;
signal \N__17147\ : std_logic;
signal \N__17144\ : std_logic;
signal \N__17141\ : std_logic;
signal \N__17138\ : std_logic;
signal \N__17135\ : std_logic;
signal \N__17132\ : std_logic;
signal \N__17129\ : std_logic;
signal \N__17126\ : std_logic;
signal \N__17123\ : std_logic;
signal \N__17122\ : std_logic;
signal \N__17121\ : std_logic;
signal \N__17118\ : std_logic;
signal \N__17115\ : std_logic;
signal \N__17112\ : std_logic;
signal \N__17109\ : std_logic;
signal \N__17104\ : std_logic;
signal \N__17101\ : std_logic;
signal \N__17098\ : std_logic;
signal \N__17093\ : std_logic;
signal \N__17090\ : std_logic;
signal \N__17087\ : std_logic;
signal \N__17084\ : std_logic;
signal \N__17081\ : std_logic;
signal \N__17080\ : std_logic;
signal \N__17077\ : std_logic;
signal \N__17074\ : std_logic;
signal \N__17071\ : std_logic;
signal \N__17066\ : std_logic;
signal \N__17063\ : std_logic;
signal \N__17060\ : std_logic;
signal \N__17057\ : std_logic;
signal \N__17054\ : std_logic;
signal \N__17051\ : std_logic;
signal \N__17050\ : std_logic;
signal \N__17047\ : std_logic;
signal \N__17046\ : std_logic;
signal \N__17043\ : std_logic;
signal \N__17040\ : std_logic;
signal \N__17037\ : std_logic;
signal \N__17030\ : std_logic;
signal \N__17027\ : std_logic;
signal \N__17024\ : std_logic;
signal \N__17021\ : std_logic;
signal \N__17018\ : std_logic;
signal \N__17015\ : std_logic;
signal \N__17012\ : std_logic;
signal \N__17009\ : std_logic;
signal \N__17006\ : std_logic;
signal \N__17003\ : std_logic;
signal \N__17002\ : std_logic;
signal \N__16999\ : std_logic;
signal \N__16996\ : std_logic;
signal \N__16993\ : std_logic;
signal \N__16990\ : std_logic;
signal \N__16985\ : std_logic;
signal \N__16982\ : std_logic;
signal \N__16981\ : std_logic;
signal \N__16980\ : std_logic;
signal \N__16977\ : std_logic;
signal \N__16972\ : std_logic;
signal \N__16967\ : std_logic;
signal \N__16964\ : std_logic;
signal \N__16961\ : std_logic;
signal \N__16958\ : std_logic;
signal \N__16957\ : std_logic;
signal \N__16954\ : std_logic;
signal \N__16953\ : std_logic;
signal \N__16950\ : std_logic;
signal \N__16947\ : std_logic;
signal \N__16942\ : std_logic;
signal \N__16937\ : std_logic;
signal \N__16934\ : std_logic;
signal \N__16931\ : std_logic;
signal \N__16928\ : std_logic;
signal \N__16925\ : std_logic;
signal \N__16922\ : std_logic;
signal \N__16919\ : std_logic;
signal \N__16916\ : std_logic;
signal \N__16915\ : std_logic;
signal \N__16912\ : std_logic;
signal \N__16909\ : std_logic;
signal \N__16908\ : std_logic;
signal \N__16905\ : std_logic;
signal \N__16902\ : std_logic;
signal \N__16899\ : std_logic;
signal \N__16892\ : std_logic;
signal \N__16891\ : std_logic;
signal \N__16888\ : std_logic;
signal \N__16885\ : std_logic;
signal \N__16884\ : std_logic;
signal \N__16881\ : std_logic;
signal \N__16878\ : std_logic;
signal \N__16875\ : std_logic;
signal \N__16868\ : std_logic;
signal \N__16865\ : std_logic;
signal \N__16862\ : std_logic;
signal \N__16859\ : std_logic;
signal \N__16856\ : std_logic;
signal \N__16855\ : std_logic;
signal \N__16852\ : std_logic;
signal \N__16849\ : std_logic;
signal \N__16846\ : std_logic;
signal \N__16843\ : std_logic;
signal \N__16842\ : std_logic;
signal \N__16839\ : std_logic;
signal \N__16836\ : std_logic;
signal \N__16833\ : std_logic;
signal \N__16826\ : std_logic;
signal \N__16823\ : std_logic;
signal \N__16820\ : std_logic;
signal \N__16817\ : std_logic;
signal \N__16814\ : std_logic;
signal \N__16811\ : std_logic;
signal \N__16810\ : std_logic;
signal \N__16809\ : std_logic;
signal \N__16806\ : std_logic;
signal \N__16803\ : std_logic;
signal \N__16800\ : std_logic;
signal \N__16797\ : std_logic;
signal \N__16790\ : std_logic;
signal \N__16787\ : std_logic;
signal \N__16784\ : std_logic;
signal \N__16781\ : std_logic;
signal \N__16778\ : std_logic;
signal \N__16775\ : std_logic;
signal \N__16772\ : std_logic;
signal \N__16769\ : std_logic;
signal \N__16766\ : std_logic;
signal \N__16763\ : std_logic;
signal \N__16762\ : std_logic;
signal \N__16761\ : std_logic;
signal \N__16758\ : std_logic;
signal \N__16755\ : std_logic;
signal \N__16752\ : std_logic;
signal \N__16747\ : std_logic;
signal \N__16744\ : std_logic;
signal \N__16741\ : std_logic;
signal \N__16736\ : std_logic;
signal \N__16733\ : std_logic;
signal \N__16730\ : std_logic;
signal \N__16727\ : std_logic;
signal \N__16724\ : std_logic;
signal \N__16721\ : std_logic;
signal \N__16718\ : std_logic;
signal \N__16715\ : std_logic;
signal \N__16712\ : std_logic;
signal \N__16709\ : std_logic;
signal \N__16708\ : std_logic;
signal \N__16707\ : std_logic;
signal \N__16704\ : std_logic;
signal \N__16701\ : std_logic;
signal \N__16698\ : std_logic;
signal \N__16695\ : std_logic;
signal \N__16692\ : std_logic;
signal \N__16685\ : std_logic;
signal \N__16682\ : std_logic;
signal \N__16679\ : std_logic;
signal \N__16676\ : std_logic;
signal \N__16675\ : std_logic;
signal \N__16674\ : std_logic;
signal \N__16671\ : std_logic;
signal \N__16666\ : std_logic;
signal \N__16663\ : std_logic;
signal \N__16660\ : std_logic;
signal \N__16655\ : std_logic;
signal \N__16652\ : std_logic;
signal \N__16649\ : std_logic;
signal \N__16646\ : std_logic;
signal \N__16643\ : std_logic;
signal \N__16640\ : std_logic;
signal \N__16637\ : std_logic;
signal \N__16636\ : std_logic;
signal \N__16633\ : std_logic;
signal \N__16630\ : std_logic;
signal \N__16629\ : std_logic;
signal \N__16626\ : std_logic;
signal \N__16621\ : std_logic;
signal \N__16616\ : std_logic;
signal \N__16613\ : std_logic;
signal \N__16610\ : std_logic;
signal \N__16607\ : std_logic;
signal \N__16604\ : std_logic;
signal \N__16603\ : std_logic;
signal \N__16602\ : std_logic;
signal \N__16601\ : std_logic;
signal \N__16600\ : std_logic;
signal \N__16599\ : std_logic;
signal \N__16598\ : std_logic;
signal \N__16597\ : std_logic;
signal \N__16594\ : std_logic;
signal \N__16593\ : std_logic;
signal \N__16592\ : std_logic;
signal \N__16591\ : std_logic;
signal \N__16588\ : std_logic;
signal \N__16583\ : std_logic;
signal \N__16580\ : std_logic;
signal \N__16575\ : std_logic;
signal \N__16572\ : std_logic;
signal \N__16569\ : std_logic;
signal \N__16562\ : std_logic;
signal \N__16547\ : std_logic;
signal \N__16546\ : std_logic;
signal \N__16543\ : std_logic;
signal \N__16540\ : std_logic;
signal \N__16537\ : std_logic;
signal \N__16534\ : std_logic;
signal \N__16531\ : std_logic;
signal \N__16526\ : std_logic;
signal \N__16523\ : std_logic;
signal \N__16522\ : std_logic;
signal \N__16519\ : std_logic;
signal \N__16516\ : std_logic;
signal \N__16513\ : std_logic;
signal \N__16510\ : std_logic;
signal \N__16507\ : std_logic;
signal \N__16504\ : std_logic;
signal \N__16499\ : std_logic;
signal \N__16498\ : std_logic;
signal \N__16495\ : std_logic;
signal \N__16492\ : std_logic;
signal \N__16489\ : std_logic;
signal \N__16486\ : std_logic;
signal \N__16485\ : std_logic;
signal \N__16482\ : std_logic;
signal \N__16479\ : std_logic;
signal \N__16476\ : std_logic;
signal \N__16469\ : std_logic;
signal \N__16466\ : std_logic;
signal \N__16463\ : std_logic;
signal \N__16460\ : std_logic;
signal \N__16457\ : std_logic;
signal \N__16456\ : std_logic;
signal \N__16453\ : std_logic;
signal \N__16450\ : std_logic;
signal \N__16447\ : std_logic;
signal \N__16444\ : std_logic;
signal \N__16439\ : std_logic;
signal \N__16436\ : std_logic;
signal \N__16433\ : std_logic;
signal \N__16430\ : std_logic;
signal \N__16427\ : std_logic;
signal \N__16426\ : std_logic;
signal \N__16423\ : std_logic;
signal \N__16420\ : std_logic;
signal \N__16417\ : std_logic;
signal \N__16414\ : std_logic;
signal \N__16413\ : std_logic;
signal \N__16410\ : std_logic;
signal \N__16407\ : std_logic;
signal \N__16404\ : std_logic;
signal \N__16397\ : std_logic;
signal \N__16396\ : std_logic;
signal \N__16393\ : std_logic;
signal \N__16390\ : std_logic;
signal \N__16387\ : std_logic;
signal \N__16386\ : std_logic;
signal \N__16383\ : std_logic;
signal \N__16380\ : std_logic;
signal \N__16377\ : std_logic;
signal \N__16370\ : std_logic;
signal \N__16369\ : std_logic;
signal \N__16368\ : std_logic;
signal \N__16367\ : std_logic;
signal \N__16366\ : std_logic;
signal \N__16365\ : std_logic;
signal \N__16364\ : std_logic;
signal \N__16361\ : std_logic;
signal \N__16358\ : std_logic;
signal \N__16355\ : std_logic;
signal \N__16354\ : std_logic;
signal \N__16353\ : std_logic;
signal \N__16350\ : std_logic;
signal \N__16347\ : std_logic;
signal \N__16346\ : std_logic;
signal \N__16343\ : std_logic;
signal \N__16340\ : std_logic;
signal \N__16339\ : std_logic;
signal \N__16336\ : std_logic;
signal \N__16333\ : std_logic;
signal \N__16328\ : std_logic;
signal \N__16319\ : std_logic;
signal \N__16312\ : std_logic;
signal \N__16309\ : std_logic;
signal \N__16298\ : std_logic;
signal \N__16295\ : std_logic;
signal \N__16292\ : std_logic;
signal \N__16289\ : std_logic;
signal \N__16288\ : std_logic;
signal \N__16285\ : std_logic;
signal \N__16282\ : std_logic;
signal \N__16277\ : std_logic;
signal \N__16274\ : std_logic;
signal \N__16271\ : std_logic;
signal \N__16268\ : std_logic;
signal \N__16265\ : std_logic;
signal \N__16262\ : std_logic;
signal \N__16259\ : std_logic;
signal \N__16258\ : std_logic;
signal \N__16255\ : std_logic;
signal \N__16252\ : std_logic;
signal \N__16247\ : std_logic;
signal \N__16244\ : std_logic;
signal \N__16241\ : std_logic;
signal \N__16238\ : std_logic;
signal \N__16237\ : std_logic;
signal \N__16234\ : std_logic;
signal \N__16231\ : std_logic;
signal \N__16230\ : std_logic;
signal \N__16227\ : std_logic;
signal \N__16224\ : std_logic;
signal \N__16221\ : std_logic;
signal \N__16214\ : std_logic;
signal \N__16211\ : std_logic;
signal \N__16208\ : std_logic;
signal \N__16205\ : std_logic;
signal \N__16204\ : std_logic;
signal \N__16203\ : std_logic;
signal \N__16200\ : std_logic;
signal \N__16197\ : std_logic;
signal \N__16194\ : std_logic;
signal \N__16191\ : std_logic;
signal \N__16188\ : std_logic;
signal \N__16181\ : std_logic;
signal \N__16178\ : std_logic;
signal \N__16175\ : std_logic;
signal \N__16172\ : std_logic;
signal \N__16169\ : std_logic;
signal \N__16166\ : std_logic;
signal \N__16165\ : std_logic;
signal \N__16162\ : std_logic;
signal \N__16159\ : std_logic;
signal \N__16154\ : std_logic;
signal \N__16151\ : std_logic;
signal \N__16148\ : std_logic;
signal \N__16145\ : std_logic;
signal \N__16142\ : std_logic;
signal \N__16139\ : std_logic;
signal \N__16136\ : std_logic;
signal \N__16135\ : std_logic;
signal \N__16132\ : std_logic;
signal \N__16129\ : std_logic;
signal \N__16124\ : std_logic;
signal \N__16121\ : std_logic;
signal \N__16118\ : std_logic;
signal \N__16115\ : std_logic;
signal \N__16114\ : std_logic;
signal \N__16111\ : std_logic;
signal \N__16108\ : std_logic;
signal \N__16107\ : std_logic;
signal \N__16104\ : std_logic;
signal \N__16101\ : std_logic;
signal \N__16098\ : std_logic;
signal \N__16091\ : std_logic;
signal \N__16090\ : std_logic;
signal \N__16087\ : std_logic;
signal \N__16084\ : std_logic;
signal \N__16083\ : std_logic;
signal \N__16080\ : std_logic;
signal \N__16077\ : std_logic;
signal \N__16074\ : std_logic;
signal \N__16067\ : std_logic;
signal \N__16064\ : std_logic;
signal \N__16061\ : std_logic;
signal \N__16058\ : std_logic;
signal \N__16055\ : std_logic;
signal \N__16052\ : std_logic;
signal \N__16051\ : std_logic;
signal \N__16050\ : std_logic;
signal \N__16047\ : std_logic;
signal \N__16044\ : std_logic;
signal \N__16041\ : std_logic;
signal \N__16038\ : std_logic;
signal \N__16035\ : std_logic;
signal \N__16032\ : std_logic;
signal \N__16025\ : std_logic;
signal \N__16022\ : std_logic;
signal \N__16021\ : std_logic;
signal \N__16018\ : std_logic;
signal \N__16015\ : std_logic;
signal \N__16014\ : std_logic;
signal \N__16011\ : std_logic;
signal \N__16008\ : std_logic;
signal \N__16005\ : std_logic;
signal \N__15998\ : std_logic;
signal \N__15995\ : std_logic;
signal \N__15992\ : std_logic;
signal \N__15989\ : std_logic;
signal \N__15986\ : std_logic;
signal \N__15983\ : std_logic;
signal \N__15982\ : std_logic;
signal \N__15979\ : std_logic;
signal \N__15978\ : std_logic;
signal \N__15977\ : std_logic;
signal \N__15974\ : std_logic;
signal \N__15973\ : std_logic;
signal \N__15972\ : std_logic;
signal \N__15967\ : std_logic;
signal \N__15964\ : std_logic;
signal \N__15963\ : std_logic;
signal \N__15962\ : std_logic;
signal \N__15961\ : std_logic;
signal \N__15960\ : std_logic;
signal \N__15959\ : std_logic;
signal \N__15956\ : std_logic;
signal \N__15951\ : std_logic;
signal \N__15948\ : std_logic;
signal \N__15941\ : std_logic;
signal \N__15936\ : std_logic;
signal \N__15935\ : std_logic;
signal \N__15932\ : std_logic;
signal \N__15931\ : std_logic;
signal \N__15928\ : std_logic;
signal \N__15925\ : std_logic;
signal \N__15920\ : std_logic;
signal \N__15917\ : std_logic;
signal \N__15910\ : std_logic;
signal \N__15899\ : std_logic;
signal \N__15898\ : std_logic;
signal \N__15897\ : std_logic;
signal \N__15894\ : std_logic;
signal \N__15891\ : std_logic;
signal \N__15888\ : std_logic;
signal \N__15885\ : std_logic;
signal \N__15878\ : std_logic;
signal \N__15875\ : std_logic;
signal \N__15872\ : std_logic;
signal \N__15869\ : std_logic;
signal \N__15868\ : std_logic;
signal \N__15865\ : std_logic;
signal \N__15862\ : std_logic;
signal \N__15859\ : std_logic;
signal \N__15858\ : std_logic;
signal \N__15855\ : std_logic;
signal \N__15852\ : std_logic;
signal \N__15849\ : std_logic;
signal \N__15846\ : std_logic;
signal \N__15839\ : std_logic;
signal \N__15836\ : std_logic;
signal \N__15833\ : std_logic;
signal \N__15830\ : std_logic;
signal \N__15829\ : std_logic;
signal \N__15826\ : std_logic;
signal \N__15823\ : std_logic;
signal \N__15820\ : std_logic;
signal \N__15819\ : std_logic;
signal \N__15816\ : std_logic;
signal \N__15813\ : std_logic;
signal \N__15810\ : std_logic;
signal \N__15807\ : std_logic;
signal \N__15804\ : std_logic;
signal \N__15801\ : std_logic;
signal \N__15794\ : std_logic;
signal \N__15793\ : std_logic;
signal \N__15790\ : std_logic;
signal \N__15787\ : std_logic;
signal \N__15784\ : std_logic;
signal \N__15781\ : std_logic;
signal \N__15780\ : std_logic;
signal \N__15777\ : std_logic;
signal \N__15774\ : std_logic;
signal \N__15771\ : std_logic;
signal \N__15768\ : std_logic;
signal \N__15761\ : std_logic;
signal \N__15758\ : std_logic;
signal \N__15755\ : std_logic;
signal \N__15752\ : std_logic;
signal \N__15751\ : std_logic;
signal \N__15750\ : std_logic;
signal \N__15747\ : std_logic;
signal \N__15744\ : std_logic;
signal \N__15741\ : std_logic;
signal \N__15738\ : std_logic;
signal \N__15731\ : std_logic;
signal \N__15728\ : std_logic;
signal \N__15727\ : std_logic;
signal \N__15724\ : std_logic;
signal \N__15721\ : std_logic;
signal \N__15718\ : std_logic;
signal \N__15717\ : std_logic;
signal \N__15712\ : std_logic;
signal \N__15709\ : std_logic;
signal \N__15706\ : std_logic;
signal \N__15701\ : std_logic;
signal \N__15698\ : std_logic;
signal \N__15695\ : std_logic;
signal \N__15692\ : std_logic;
signal \N__15689\ : std_logic;
signal \N__15686\ : std_logic;
signal \N__15685\ : std_logic;
signal \N__15684\ : std_logic;
signal \N__15681\ : std_logic;
signal \N__15678\ : std_logic;
signal \N__15675\ : std_logic;
signal \N__15668\ : std_logic;
signal \N__15665\ : std_logic;
signal \N__15662\ : std_logic;
signal \N__15659\ : std_logic;
signal \N__15656\ : std_logic;
signal \N__15653\ : std_logic;
signal \N__15652\ : std_logic;
signal \N__15649\ : std_logic;
signal \N__15646\ : std_logic;
signal \N__15643\ : std_logic;
signal \N__15640\ : std_logic;
signal \N__15635\ : std_logic;
signal \N__15632\ : std_logic;
signal \N__15629\ : std_logic;
signal \N__15626\ : std_logic;
signal \N__15623\ : std_logic;
signal \N__15620\ : std_logic;
signal \N__15617\ : std_logic;
signal \N__15616\ : std_logic;
signal \N__15613\ : std_logic;
signal \N__15610\ : std_logic;
signal \N__15609\ : std_logic;
signal \N__15606\ : std_logic;
signal \N__15603\ : std_logic;
signal \N__15600\ : std_logic;
signal \N__15597\ : std_logic;
signal \N__15594\ : std_logic;
signal \N__15587\ : std_logic;
signal \N__15584\ : std_logic;
signal \N__15583\ : std_logic;
signal \N__15580\ : std_logic;
signal \N__15579\ : std_logic;
signal \N__15576\ : std_logic;
signal \N__15573\ : std_logic;
signal \N__15570\ : std_logic;
signal \N__15565\ : std_logic;
signal \N__15560\ : std_logic;
signal \N__15557\ : std_logic;
signal \N__15554\ : std_logic;
signal \N__15551\ : std_logic;
signal \N__15548\ : std_logic;
signal \N__15547\ : std_logic;
signal \N__15544\ : std_logic;
signal \N__15541\ : std_logic;
signal \N__15538\ : std_logic;
signal \N__15537\ : std_logic;
signal \N__15534\ : std_logic;
signal \N__15531\ : std_logic;
signal \N__15528\ : std_logic;
signal \N__15521\ : std_logic;
signal \N__15520\ : std_logic;
signal \N__15519\ : std_logic;
signal \N__15518\ : std_logic;
signal \N__15517\ : std_logic;
signal \N__15514\ : std_logic;
signal \N__15513\ : std_logic;
signal \N__15512\ : std_logic;
signal \N__15509\ : std_logic;
signal \N__15506\ : std_logic;
signal \N__15505\ : std_logic;
signal \N__15504\ : std_logic;
signal \N__15501\ : std_logic;
signal \N__15500\ : std_logic;
signal \N__15499\ : std_logic;
signal \N__15498\ : std_logic;
signal \N__15495\ : std_logic;
signal \N__15494\ : std_logic;
signal \N__15489\ : std_logic;
signal \N__15484\ : std_logic;
signal \N__15479\ : std_logic;
signal \N__15472\ : std_logic;
signal \N__15469\ : std_logic;
signal \N__15462\ : std_logic;
signal \N__15457\ : std_logic;
signal \N__15446\ : std_logic;
signal \N__15443\ : std_logic;
signal \N__15440\ : std_logic;
signal \N__15437\ : std_logic;
signal \N__15434\ : std_logic;
signal \N__15431\ : std_logic;
signal \N__15430\ : std_logic;
signal \N__15427\ : std_logic;
signal \N__15424\ : std_logic;
signal \N__15419\ : std_logic;
signal \N__15418\ : std_logic;
signal \N__15415\ : std_logic;
signal \N__15412\ : std_logic;
signal \N__15409\ : std_logic;
signal \N__15406\ : std_logic;
signal \N__15401\ : std_logic;
signal \N__15398\ : std_logic;
signal \N__15395\ : std_logic;
signal \N__15392\ : std_logic;
signal \N__15389\ : std_logic;
signal \N__15386\ : std_logic;
signal \N__15383\ : std_logic;
signal \N__15380\ : std_logic;
signal \N__15377\ : std_logic;
signal \N__15374\ : std_logic;
signal \N__15371\ : std_logic;
signal \N__15370\ : std_logic;
signal \N__15369\ : std_logic;
signal \N__15366\ : std_logic;
signal \N__15363\ : std_logic;
signal \N__15360\ : std_logic;
signal \N__15357\ : std_logic;
signal \N__15354\ : std_logic;
signal \N__15347\ : std_logic;
signal \N__15344\ : std_logic;
signal \N__15341\ : std_logic;
signal \N__15338\ : std_logic;
signal \N__15335\ : std_logic;
signal \N__15334\ : std_logic;
signal \N__15331\ : std_logic;
signal \N__15328\ : std_logic;
signal \N__15327\ : std_logic;
signal \N__15324\ : std_logic;
signal \N__15321\ : std_logic;
signal \N__15318\ : std_logic;
signal \N__15315\ : std_logic;
signal \N__15312\ : std_logic;
signal \N__15309\ : std_logic;
signal \N__15306\ : std_logic;
signal \N__15301\ : std_logic;
signal \N__15296\ : std_logic;
signal \N__15293\ : std_logic;
signal \N__15290\ : std_logic;
signal \N__15287\ : std_logic;
signal \N__15284\ : std_logic;
signal \N__15283\ : std_logic;
signal \N__15280\ : std_logic;
signal \N__15277\ : std_logic;
signal \N__15276\ : std_logic;
signal \N__15273\ : std_logic;
signal \N__15270\ : std_logic;
signal \N__15267\ : std_logic;
signal \N__15262\ : std_logic;
signal \N__15259\ : std_logic;
signal \N__15256\ : std_logic;
signal \N__15253\ : std_logic;
signal \N__15250\ : std_logic;
signal \N__15247\ : std_logic;
signal \N__15242\ : std_logic;
signal \N__15239\ : std_logic;
signal \N__15236\ : std_logic;
signal \N__15233\ : std_logic;
signal \N__15230\ : std_logic;
signal \N__15227\ : std_logic;
signal \N__15224\ : std_logic;
signal \N__15223\ : std_logic;
signal \N__15220\ : std_logic;
signal \N__15217\ : std_logic;
signal \N__15214\ : std_logic;
signal \N__15211\ : std_logic;
signal \N__15206\ : std_logic;
signal \N__15203\ : std_logic;
signal \N__15200\ : std_logic;
signal \N__15197\ : std_logic;
signal \N__15194\ : std_logic;
signal \N__15191\ : std_logic;
signal \N__15188\ : std_logic;
signal \N__15187\ : std_logic;
signal \N__15184\ : std_logic;
signal \N__15181\ : std_logic;
signal \N__15180\ : std_logic;
signal \N__15175\ : std_logic;
signal \N__15172\ : std_logic;
signal \N__15169\ : std_logic;
signal \N__15164\ : std_logic;
signal \N__15161\ : std_logic;
signal \N__15158\ : std_logic;
signal \N__15155\ : std_logic;
signal \N__15152\ : std_logic;
signal \N__15149\ : std_logic;
signal \N__15148\ : std_logic;
signal \N__15145\ : std_logic;
signal \N__15144\ : std_logic;
signal \N__15141\ : std_logic;
signal \N__15138\ : std_logic;
signal \N__15135\ : std_logic;
signal \N__15132\ : std_logic;
signal \N__15125\ : std_logic;
signal \N__15122\ : std_logic;
signal \N__15119\ : std_logic;
signal \N__15116\ : std_logic;
signal \N__15113\ : std_logic;
signal \N__15112\ : std_logic;
signal \N__15109\ : std_logic;
signal \N__15106\ : std_logic;
signal \N__15103\ : std_logic;
signal \N__15100\ : std_logic;
signal \N__15097\ : std_logic;
signal \N__15096\ : std_logic;
signal \N__15093\ : std_logic;
signal \N__15090\ : std_logic;
signal \N__15087\ : std_logic;
signal \N__15080\ : std_logic;
signal \N__15077\ : std_logic;
signal \N__15074\ : std_logic;
signal \N__15071\ : std_logic;
signal \N__15068\ : std_logic;
signal \N__15067\ : std_logic;
signal \N__15064\ : std_logic;
signal \N__15061\ : std_logic;
signal \N__15058\ : std_logic;
signal \N__15055\ : std_logic;
signal \N__15052\ : std_logic;
signal \N__15051\ : std_logic;
signal \N__15048\ : std_logic;
signal \N__15045\ : std_logic;
signal \N__15042\ : std_logic;
signal \N__15035\ : std_logic;
signal \N__15032\ : std_logic;
signal \N__15029\ : std_logic;
signal \N__15026\ : std_logic;
signal \N__15023\ : std_logic;
signal \N__15020\ : std_logic;
signal \N__15019\ : std_logic;
signal \N__15016\ : std_logic;
signal \N__15013\ : std_logic;
signal \N__15010\ : std_logic;
signal \N__15007\ : std_logic;
signal \N__15006\ : std_logic;
signal \N__15003\ : std_logic;
signal \N__15000\ : std_logic;
signal \N__14997\ : std_logic;
signal \N__14994\ : std_logic;
signal \N__14991\ : std_logic;
signal \N__14988\ : std_logic;
signal \N__14981\ : std_logic;
signal \N__14978\ : std_logic;
signal \N__14975\ : std_logic;
signal \N__14972\ : std_logic;
signal \N__14969\ : std_logic;
signal \N__14968\ : std_logic;
signal \N__14965\ : std_logic;
signal \N__14962\ : std_logic;
signal \N__14959\ : std_logic;
signal \N__14958\ : std_logic;
signal \N__14955\ : std_logic;
signal \N__14952\ : std_logic;
signal \N__14949\ : std_logic;
signal \N__14942\ : std_logic;
signal \N__14939\ : std_logic;
signal \N__14936\ : std_logic;
signal \N__14933\ : std_logic;
signal \N__14930\ : std_logic;
signal \N__14927\ : std_logic;
signal \N__14924\ : std_logic;
signal \N__14921\ : std_logic;
signal \N__14918\ : std_logic;
signal \N__14915\ : std_logic;
signal \N__14914\ : std_logic;
signal \N__14911\ : std_logic;
signal \N__14910\ : std_logic;
signal \N__14907\ : std_logic;
signal \N__14904\ : std_logic;
signal \N__14901\ : std_logic;
signal \N__14894\ : std_logic;
signal \N__14891\ : std_logic;
signal \N__14888\ : std_logic;
signal \N__14885\ : std_logic;
signal \N__14882\ : std_logic;
signal \N__14879\ : std_logic;
signal \N__14878\ : std_logic;
signal \N__14875\ : std_logic;
signal \N__14874\ : std_logic;
signal \N__14871\ : std_logic;
signal \N__14868\ : std_logic;
signal \N__14865\ : std_logic;
signal \N__14858\ : std_logic;
signal \N__14855\ : std_logic;
signal \N__14852\ : std_logic;
signal \N__14849\ : std_logic;
signal \N__14846\ : std_logic;
signal \N__14843\ : std_logic;
signal \N__14840\ : std_logic;
signal \N__14837\ : std_logic;
signal \N__14834\ : std_logic;
signal \N__14831\ : std_logic;
signal \N__14828\ : std_logic;
signal \N__14825\ : std_logic;
signal \N__14822\ : std_logic;
signal \N__14819\ : std_logic;
signal \N__14816\ : std_logic;
signal \N__14813\ : std_logic;
signal \N__14810\ : std_logic;
signal \N__14807\ : std_logic;
signal \N__14804\ : std_logic;
signal \N__14801\ : std_logic;
signal \N__14800\ : std_logic;
signal \N__14799\ : std_logic;
signal \N__14794\ : std_logic;
signal \N__14791\ : std_logic;
signal \N__14786\ : std_logic;
signal \N__14783\ : std_logic;
signal \N__14782\ : std_logic;
signal \N__14781\ : std_logic;
signal \N__14776\ : std_logic;
signal \N__14773\ : std_logic;
signal \N__14768\ : std_logic;
signal \N__14765\ : std_logic;
signal \N__14764\ : std_logic;
signal \N__14761\ : std_logic;
signal \N__14760\ : std_logic;
signal \N__14755\ : std_logic;
signal \N__14752\ : std_logic;
signal \N__14747\ : std_logic;
signal \N__14744\ : std_logic;
signal \N__14743\ : std_logic;
signal \N__14742\ : std_logic;
signal \N__14737\ : std_logic;
signal \N__14734\ : std_logic;
signal \N__14729\ : std_logic;
signal \N__14726\ : std_logic;
signal \N__14723\ : std_logic;
signal \N__14722\ : std_logic;
signal \N__14719\ : std_logic;
signal \N__14716\ : std_logic;
signal \N__14711\ : std_logic;
signal \N__14708\ : std_logic;
signal \N__14705\ : std_logic;
signal \N__14702\ : std_logic;
signal \N__14699\ : std_logic;
signal \N__14696\ : std_logic;
signal \N__14693\ : std_logic;
signal \N__14690\ : std_logic;
signal \N__14687\ : std_logic;
signal \N__14684\ : std_logic;
signal \N__14681\ : std_logic;
signal \N__14678\ : std_logic;
signal \N__14675\ : std_logic;
signal \N__14672\ : std_logic;
signal \N__14669\ : std_logic;
signal \N__14666\ : std_logic;
signal \N__14663\ : std_logic;
signal \N__14660\ : std_logic;
signal \N__14657\ : std_logic;
signal \N__14654\ : std_logic;
signal \N__14651\ : std_logic;
signal \N__14648\ : std_logic;
signal \N__14645\ : std_logic;
signal \N__14642\ : std_logic;
signal \N__14639\ : std_logic;
signal \N__14636\ : std_logic;
signal \N__14633\ : std_logic;
signal \N__14630\ : std_logic;
signal \N__14627\ : std_logic;
signal \N__14624\ : std_logic;
signal \N__14621\ : std_logic;
signal \N__14618\ : std_logic;
signal \N__14615\ : std_logic;
signal \N__14612\ : std_logic;
signal \N__14609\ : std_logic;
signal \N__14606\ : std_logic;
signal \N__14603\ : std_logic;
signal \N__14600\ : std_logic;
signal \N__14597\ : std_logic;
signal \N__14594\ : std_logic;
signal \N__14591\ : std_logic;
signal \N__14588\ : std_logic;
signal \N__14585\ : std_logic;
signal \N__14582\ : std_logic;
signal \N__14579\ : std_logic;
signal \N__14576\ : std_logic;
signal \N__14573\ : std_logic;
signal \N__14570\ : std_logic;
signal \N__14567\ : std_logic;
signal \N__14564\ : std_logic;
signal \N__14561\ : std_logic;
signal \N__14558\ : std_logic;
signal \N__14557\ : std_logic;
signal \N__14556\ : std_logic;
signal \N__14553\ : std_logic;
signal \N__14550\ : std_logic;
signal \N__14547\ : std_logic;
signal \N__14544\ : std_logic;
signal \N__14541\ : std_logic;
signal \N__14538\ : std_logic;
signal \N__14531\ : std_logic;
signal \N__14528\ : std_logic;
signal \N__14525\ : std_logic;
signal \N__14522\ : std_logic;
signal \N__14519\ : std_logic;
signal \N__14516\ : std_logic;
signal \N__14515\ : std_logic;
signal \N__14512\ : std_logic;
signal \N__14509\ : std_logic;
signal \N__14506\ : std_logic;
signal \N__14503\ : std_logic;
signal \N__14500\ : std_logic;
signal \N__14497\ : std_logic;
signal \N__14492\ : std_logic;
signal \N__14489\ : std_logic;
signal \N__14486\ : std_logic;
signal \N__14483\ : std_logic;
signal \N__14480\ : std_logic;
signal \N__14479\ : std_logic;
signal \N__14478\ : std_logic;
signal \N__14475\ : std_logic;
signal \N__14470\ : std_logic;
signal \N__14467\ : std_logic;
signal \N__14462\ : std_logic;
signal \N__14459\ : std_logic;
signal \N__14456\ : std_logic;
signal \N__14453\ : std_logic;
signal \N__14450\ : std_logic;
signal \N__14447\ : std_logic;
signal \N__14444\ : std_logic;
signal \N__14441\ : std_logic;
signal \N__14440\ : std_logic;
signal \N__14437\ : std_logic;
signal \N__14436\ : std_logic;
signal \N__14433\ : std_logic;
signal \N__14430\ : std_logic;
signal \N__14427\ : std_logic;
signal \N__14424\ : std_logic;
signal \N__14419\ : std_logic;
signal \N__14414\ : std_logic;
signal \N__14411\ : std_logic;
signal \N__14408\ : std_logic;
signal \N__14405\ : std_logic;
signal \N__14402\ : std_logic;
signal \N__14399\ : std_logic;
signal \N__14398\ : std_logic;
signal \N__14395\ : std_logic;
signal \N__14392\ : std_logic;
signal \N__14387\ : std_logic;
signal \N__14384\ : std_logic;
signal \N__14381\ : std_logic;
signal \N__14378\ : std_logic;
signal \N__14375\ : std_logic;
signal \N__14372\ : std_logic;
signal \N__14369\ : std_logic;
signal \N__14366\ : std_logic;
signal \N__14363\ : std_logic;
signal \N__14360\ : std_logic;
signal \N__14357\ : std_logic;
signal \N__14354\ : std_logic;
signal \N__14351\ : std_logic;
signal \N__14348\ : std_logic;
signal \N__14345\ : std_logic;
signal \N__14344\ : std_logic;
signal \N__14343\ : std_logic;
signal \N__14340\ : std_logic;
signal \N__14335\ : std_logic;
signal \N__14332\ : std_logic;
signal \N__14327\ : std_logic;
signal \N__14324\ : std_logic;
signal \N__14321\ : std_logic;
signal \N__14318\ : std_logic;
signal \N__14315\ : std_logic;
signal \N__14314\ : std_logic;
signal \N__14311\ : std_logic;
signal \N__14308\ : std_logic;
signal \N__14305\ : std_logic;
signal \N__14302\ : std_logic;
signal \N__14299\ : std_logic;
signal \N__14296\ : std_logic;
signal \N__14295\ : std_logic;
signal \N__14290\ : std_logic;
signal \N__14287\ : std_logic;
signal \N__14282\ : std_logic;
signal \N__14279\ : std_logic;
signal \N__14276\ : std_logic;
signal \N__14273\ : std_logic;
signal \N__14272\ : std_logic;
signal \N__14269\ : std_logic;
signal \N__14266\ : std_logic;
signal \N__14263\ : std_logic;
signal \N__14262\ : std_logic;
signal \N__14257\ : std_logic;
signal \N__14254\ : std_logic;
signal \N__14249\ : std_logic;
signal \N__14246\ : std_logic;
signal \N__14245\ : std_logic;
signal \N__14242\ : std_logic;
signal \N__14239\ : std_logic;
signal \N__14234\ : std_logic;
signal \N__14231\ : std_logic;
signal \N__14228\ : std_logic;
signal \N__14225\ : std_logic;
signal \N__14224\ : std_logic;
signal \N__14221\ : std_logic;
signal \N__14218\ : std_logic;
signal \N__14215\ : std_logic;
signal \N__14210\ : std_logic;
signal \N__14207\ : std_logic;
signal \N__14204\ : std_logic;
signal \N__14201\ : std_logic;
signal \N__14198\ : std_logic;
signal \N__14195\ : std_logic;
signal \N__14192\ : std_logic;
signal \N__14189\ : std_logic;
signal \N__14186\ : std_logic;
signal \N__14185\ : std_logic;
signal \N__14182\ : std_logic;
signal \N__14179\ : std_logic;
signal \N__14178\ : std_logic;
signal \N__14175\ : std_logic;
signal \N__14172\ : std_logic;
signal \N__14169\ : std_logic;
signal \N__14164\ : std_logic;
signal \N__14159\ : std_logic;
signal \N__14156\ : std_logic;
signal \N__14155\ : std_logic;
signal \N__14152\ : std_logic;
signal \N__14149\ : std_logic;
signal \N__14146\ : std_logic;
signal \N__14145\ : std_logic;
signal \N__14142\ : std_logic;
signal \N__14139\ : std_logic;
signal \N__14136\ : std_logic;
signal \N__14129\ : std_logic;
signal \N__14128\ : std_logic;
signal \N__14127\ : std_logic;
signal \N__14124\ : std_logic;
signal \N__14121\ : std_logic;
signal \N__14118\ : std_logic;
signal \N__14115\ : std_logic;
signal \N__14112\ : std_logic;
signal \N__14109\ : std_logic;
signal \N__14104\ : std_logic;
signal \N__14099\ : std_logic;
signal \N__14096\ : std_logic;
signal \N__14093\ : std_logic;
signal \N__14090\ : std_logic;
signal \N__14087\ : std_logic;
signal \N__14084\ : std_logic;
signal \N__14081\ : std_logic;
signal \N__14078\ : std_logic;
signal \N__14075\ : std_logic;
signal \N__14072\ : std_logic;
signal \N__14069\ : std_logic;
signal \N__14068\ : std_logic;
signal \N__14065\ : std_logic;
signal \N__14064\ : std_logic;
signal \N__14061\ : std_logic;
signal \N__14058\ : std_logic;
signal \N__14055\ : std_logic;
signal \N__14052\ : std_logic;
signal \N__14045\ : std_logic;
signal \N__14042\ : std_logic;
signal \N__14039\ : std_logic;
signal \N__14036\ : std_logic;
signal \N__14035\ : std_logic;
signal \N__14034\ : std_logic;
signal \N__14031\ : std_logic;
signal \N__14028\ : std_logic;
signal \N__14025\ : std_logic;
signal \N__14022\ : std_logic;
signal \N__14019\ : std_logic;
signal \N__14012\ : std_logic;
signal \N__14011\ : std_logic;
signal \N__14008\ : std_logic;
signal \N__14005\ : std_logic;
signal \N__14004\ : std_logic;
signal \N__14001\ : std_logic;
signal \N__13998\ : std_logic;
signal \N__13995\ : std_logic;
signal \N__13988\ : std_logic;
signal \N__13985\ : std_logic;
signal \N__13982\ : std_logic;
signal \N__13979\ : std_logic;
signal \N__13978\ : std_logic;
signal \N__13975\ : std_logic;
signal \N__13974\ : std_logic;
signal \N__13971\ : std_logic;
signal \N__13968\ : std_logic;
signal \N__13965\ : std_logic;
signal \N__13958\ : std_logic;
signal \N__13955\ : std_logic;
signal \N__13952\ : std_logic;
signal \N__13951\ : std_logic;
signal \N__13950\ : std_logic;
signal \N__13949\ : std_logic;
signal \N__13946\ : std_logic;
signal \N__13943\ : std_logic;
signal \N__13940\ : std_logic;
signal \N__13939\ : std_logic;
signal \N__13938\ : std_logic;
signal \N__13937\ : std_logic;
signal \N__13936\ : std_logic;
signal \N__13935\ : std_logic;
signal \N__13932\ : std_logic;
signal \N__13931\ : std_logic;
signal \N__13928\ : std_logic;
signal \N__13917\ : std_logic;
signal \N__13908\ : std_logic;
signal \N__13901\ : std_logic;
signal \N__13898\ : std_logic;
signal \N__13897\ : std_logic;
signal \N__13894\ : std_logic;
signal \N__13891\ : std_logic;
signal \N__13886\ : std_logic;
signal \N__13885\ : std_logic;
signal \N__13884\ : std_logic;
signal \N__13881\ : std_logic;
signal \N__13878\ : std_logic;
signal \N__13875\ : std_logic;
signal \N__13872\ : std_logic;
signal \N__13869\ : std_logic;
signal \N__13862\ : std_logic;
signal \N__13859\ : std_logic;
signal \N__13856\ : std_logic;
signal \N__13853\ : std_logic;
signal \N__13850\ : std_logic;
signal \N__13847\ : std_logic;
signal \N__13844\ : std_logic;
signal \N__13843\ : std_logic;
signal \N__13840\ : std_logic;
signal \N__13837\ : std_logic;
signal \N__13834\ : std_logic;
signal \N__13831\ : std_logic;
signal \N__13826\ : std_logic;
signal \N__13823\ : std_logic;
signal \N__13820\ : std_logic;
signal \N__13817\ : std_logic;
signal \N__13814\ : std_logic;
signal \N__13813\ : std_logic;
signal \N__13810\ : std_logic;
signal \N__13807\ : std_logic;
signal \N__13804\ : std_logic;
signal \N__13801\ : std_logic;
signal \N__13796\ : std_logic;
signal \N__13793\ : std_logic;
signal \N__13792\ : std_logic;
signal \N__13791\ : std_logic;
signal \N__13788\ : std_logic;
signal \N__13785\ : std_logic;
signal \N__13782\ : std_logic;
signal \N__13777\ : std_logic;
signal \N__13772\ : std_logic;
signal \N__13769\ : std_logic;
signal \N__13766\ : std_logic;
signal \N__13763\ : std_logic;
signal \N__13760\ : std_logic;
signal \N__13757\ : std_logic;
signal \N__13756\ : std_logic;
signal \N__13753\ : std_logic;
signal \N__13750\ : std_logic;
signal \N__13747\ : std_logic;
signal \N__13744\ : std_logic;
signal \N__13743\ : std_logic;
signal \N__13738\ : std_logic;
signal \N__13735\ : std_logic;
signal \N__13730\ : std_logic;
signal \N__13727\ : std_logic;
signal \N__13724\ : std_logic;
signal \N__13721\ : std_logic;
signal \N__13720\ : std_logic;
signal \N__13719\ : std_logic;
signal \N__13716\ : std_logic;
signal \N__13713\ : std_logic;
signal \N__13710\ : std_logic;
signal \N__13705\ : std_logic;
signal \N__13702\ : std_logic;
signal \N__13699\ : std_logic;
signal \N__13694\ : std_logic;
signal \N__13691\ : std_logic;
signal \N__13688\ : std_logic;
signal \N__13685\ : std_logic;
signal \N__13682\ : std_logic;
signal \N__13679\ : std_logic;
signal \N__13678\ : std_logic;
signal \N__13675\ : std_logic;
signal \N__13674\ : std_logic;
signal \N__13671\ : std_logic;
signal \N__13668\ : std_logic;
signal \N__13665\ : std_logic;
signal \N__13658\ : std_logic;
signal \N__13655\ : std_logic;
signal \N__13652\ : std_logic;
signal \N__13649\ : std_logic;
signal \N__13646\ : std_logic;
signal \N__13643\ : std_logic;
signal \N__13640\ : std_logic;
signal \N__13637\ : std_logic;
signal \N__13636\ : std_logic;
signal \N__13633\ : std_logic;
signal \N__13632\ : std_logic;
signal \N__13629\ : std_logic;
signal \N__13626\ : std_logic;
signal \N__13623\ : std_logic;
signal \N__13616\ : std_logic;
signal \N__13613\ : std_logic;
signal \N__13610\ : std_logic;
signal \N__13607\ : std_logic;
signal \N__13604\ : std_logic;
signal \N__13601\ : std_logic;
signal \N__13598\ : std_logic;
signal \N__13595\ : std_logic;
signal \N__13592\ : std_logic;
signal \N__13589\ : std_logic;
signal \N__13586\ : std_logic;
signal \N__13585\ : std_logic;
signal \N__13584\ : std_logic;
signal \N__13581\ : std_logic;
signal \N__13578\ : std_logic;
signal \N__13575\ : std_logic;
signal \N__13570\ : std_logic;
signal \N__13565\ : std_logic;
signal \N__13562\ : std_logic;
signal \N__13559\ : std_logic;
signal \N__13556\ : std_logic;
signal \N__13553\ : std_logic;
signal \N__13550\ : std_logic;
signal \N__13547\ : std_logic;
signal \N__13544\ : std_logic;
signal \N__13541\ : std_logic;
signal \N__13538\ : std_logic;
signal \N__13535\ : std_logic;
signal \N__13532\ : std_logic;
signal \N__13531\ : std_logic;
signal \N__13528\ : std_logic;
signal \N__13525\ : std_logic;
signal \N__13520\ : std_logic;
signal \N__13517\ : std_logic;
signal \N__13514\ : std_logic;
signal \N__13511\ : std_logic;
signal \N__13508\ : std_logic;
signal \N__13505\ : std_logic;
signal \N__13502\ : std_logic;
signal \N__13499\ : std_logic;
signal \N__13496\ : std_logic;
signal \N__13493\ : std_logic;
signal \N__13490\ : std_logic;
signal \N__13487\ : std_logic;
signal \N__13484\ : std_logic;
signal \N__13481\ : std_logic;
signal \N__13478\ : std_logic;
signal \N__13475\ : std_logic;
signal \N__13474\ : std_logic;
signal \N__13471\ : std_logic;
signal \N__13470\ : std_logic;
signal \N__13467\ : std_logic;
signal \N__13464\ : std_logic;
signal \N__13461\ : std_logic;
signal \N__13454\ : std_logic;
signal \N__13451\ : std_logic;
signal \N__13448\ : std_logic;
signal \N__13445\ : std_logic;
signal \N__13442\ : std_logic;
signal \N__13439\ : std_logic;
signal \N__13436\ : std_logic;
signal \N__13433\ : std_logic;
signal \N__13430\ : std_logic;
signal \N__13429\ : std_logic;
signal \N__13426\ : std_logic;
signal \N__13423\ : std_logic;
signal \N__13418\ : std_logic;
signal \N__13415\ : std_logic;
signal \N__13414\ : std_logic;
signal \N__13413\ : std_logic;
signal \N__13408\ : std_logic;
signal \N__13405\ : std_logic;
signal \N__13400\ : std_logic;
signal \N__13397\ : std_logic;
signal \N__13394\ : std_logic;
signal \N__13391\ : std_logic;
signal \N__13388\ : std_logic;
signal \N__13385\ : std_logic;
signal \N__13382\ : std_logic;
signal \N__13381\ : std_logic;
signal \N__13376\ : std_logic;
signal \N__13375\ : std_logic;
signal \N__13372\ : std_logic;
signal \N__13369\ : std_logic;
signal \N__13364\ : std_logic;
signal \N__13361\ : std_logic;
signal \N__13360\ : std_logic;
signal \N__13359\ : std_logic;
signal \N__13356\ : std_logic;
signal \N__13351\ : std_logic;
signal \N__13348\ : std_logic;
signal \N__13343\ : std_logic;
signal \N__13340\ : std_logic;
signal \N__13337\ : std_logic;
signal \N__13334\ : std_logic;
signal \N__13331\ : std_logic;
signal \N__13328\ : std_logic;
signal \N__13325\ : std_logic;
signal \N__13324\ : std_logic;
signal \N__13321\ : std_logic;
signal \N__13320\ : std_logic;
signal \N__13317\ : std_logic;
signal \N__13314\ : std_logic;
signal \N__13311\ : std_logic;
signal \N__13304\ : std_logic;
signal \N__13301\ : std_logic;
signal \N__13298\ : std_logic;
signal \N__13295\ : std_logic;
signal \N__13292\ : std_logic;
signal \N__13289\ : std_logic;
signal \N__13288\ : std_logic;
signal \N__13285\ : std_logic;
signal \N__13284\ : std_logic;
signal \N__13281\ : std_logic;
signal \N__13278\ : std_logic;
signal \N__13273\ : std_logic;
signal \N__13268\ : std_logic;
signal \N__13265\ : std_logic;
signal \N__13262\ : std_logic;
signal \N__13259\ : std_logic;
signal \N__13256\ : std_logic;
signal \N__13255\ : std_logic;
signal \N__13254\ : std_logic;
signal \N__13251\ : std_logic;
signal \N__13248\ : std_logic;
signal \N__13245\ : std_logic;
signal \N__13242\ : std_logic;
signal \N__13239\ : std_logic;
signal \N__13232\ : std_logic;
signal \N__13229\ : std_logic;
signal \N__13226\ : std_logic;
signal \N__13223\ : std_logic;
signal \N__13220\ : std_logic;
signal \N__13217\ : std_logic;
signal \N__13216\ : std_logic;
signal \N__13213\ : std_logic;
signal \N__13210\ : std_logic;
signal \N__13209\ : std_logic;
signal \N__13206\ : std_logic;
signal \N__13201\ : std_logic;
signal \N__13196\ : std_logic;
signal \N__13193\ : std_logic;
signal \N__13190\ : std_logic;
signal \N__13187\ : std_logic;
signal \N__13184\ : std_logic;
signal \N__13181\ : std_logic;
signal \N__13178\ : std_logic;
signal \N__13175\ : std_logic;
signal \N__13172\ : std_logic;
signal \N__13171\ : std_logic;
signal \N__13168\ : std_logic;
signal \N__13165\ : std_logic;
signal \N__13160\ : std_logic;
signal \N__13157\ : std_logic;
signal \N__13154\ : std_logic;
signal \N__13151\ : std_logic;
signal \N__13148\ : std_logic;
signal \N__13145\ : std_logic;
signal \N__13142\ : std_logic;
signal \N__13139\ : std_logic;
signal \N__13136\ : std_logic;
signal \N__13133\ : std_logic;
signal \N__13130\ : std_logic;
signal \N__13127\ : std_logic;
signal \N__13124\ : std_logic;
signal \N__13121\ : std_logic;
signal \N__13118\ : std_logic;
signal \N__13117\ : std_logic;
signal \N__13116\ : std_logic;
signal \N__13115\ : std_logic;
signal \N__13114\ : std_logic;
signal \N__13113\ : std_logic;
signal \N__13110\ : std_logic;
signal \N__13107\ : std_logic;
signal \N__13104\ : std_logic;
signal \N__13103\ : std_logic;
signal \N__13102\ : std_logic;
signal \N__13101\ : std_logic;
signal \N__13100\ : std_logic;
signal \N__13097\ : std_logic;
signal \N__13094\ : std_logic;
signal \N__13091\ : std_logic;
signal \N__13090\ : std_logic;
signal \N__13087\ : std_logic;
signal \N__13076\ : std_logic;
signal \N__13073\ : std_logic;
signal \N__13064\ : std_logic;
signal \N__13055\ : std_logic;
signal \N__13052\ : std_logic;
signal \N__13051\ : std_logic;
signal \N__13050\ : std_logic;
signal \N__13047\ : std_logic;
signal \N__13044\ : std_logic;
signal \N__13041\ : std_logic;
signal \N__13036\ : std_logic;
signal \N__13031\ : std_logic;
signal \N__13028\ : std_logic;
signal \N__13025\ : std_logic;
signal \N__13022\ : std_logic;
signal \N__13019\ : std_logic;
signal \N__13016\ : std_logic;
signal \N__13013\ : std_logic;
signal \N__13010\ : std_logic;
signal \N__13009\ : std_logic;
signal \N__13006\ : std_logic;
signal \N__13003\ : std_logic;
signal \N__12998\ : std_logic;
signal \N__12995\ : std_logic;
signal \N__12992\ : std_logic;
signal \N__12989\ : std_logic;
signal \N__12986\ : std_logic;
signal \N__12983\ : std_logic;
signal \N__12980\ : std_logic;
signal \N__12977\ : std_logic;
signal \N__12976\ : std_logic;
signal \N__12975\ : std_logic;
signal \N__12972\ : std_logic;
signal \N__12969\ : std_logic;
signal \N__12966\ : std_logic;
signal \N__12959\ : std_logic;
signal \N__12956\ : std_logic;
signal \N__12953\ : std_logic;
signal \N__12950\ : std_logic;
signal \N__12947\ : std_logic;
signal \N__12946\ : std_logic;
signal \N__12943\ : std_logic;
signal \N__12940\ : std_logic;
signal \N__12937\ : std_logic;
signal \N__12934\ : std_logic;
signal \N__12929\ : std_logic;
signal \N__12928\ : std_logic;
signal \N__12927\ : std_logic;
signal \N__12926\ : std_logic;
signal \N__12923\ : std_logic;
signal \N__12920\ : std_logic;
signal \N__12917\ : std_logic;
signal \N__12916\ : std_logic;
signal \N__12915\ : std_logic;
signal \N__12912\ : std_logic;
signal \N__12911\ : std_logic;
signal \N__12908\ : std_logic;
signal \N__12899\ : std_logic;
signal \N__12894\ : std_logic;
signal \N__12887\ : std_logic;
signal \N__12884\ : std_logic;
signal \N__12881\ : std_logic;
signal \N__12878\ : std_logic;
signal \N__12875\ : std_logic;
signal \N__12872\ : std_logic;
signal \N__12869\ : std_logic;
signal \N__12866\ : std_logic;
signal \N__12863\ : std_logic;
signal \N__12860\ : std_logic;
signal \N__12857\ : std_logic;
signal \N__12854\ : std_logic;
signal \N__12851\ : std_logic;
signal \N__12848\ : std_logic;
signal \N__12845\ : std_logic;
signal \N__12842\ : std_logic;
signal \N__12839\ : std_logic;
signal \N__12836\ : std_logic;
signal \N__12833\ : std_logic;
signal \N__12832\ : std_logic;
signal \N__12829\ : std_logic;
signal \N__12828\ : std_logic;
signal \N__12825\ : std_logic;
signal \N__12822\ : std_logic;
signal \N__12819\ : std_logic;
signal \N__12812\ : std_logic;
signal \N__12809\ : std_logic;
signal \N__12806\ : std_logic;
signal \N__12803\ : std_logic;
signal \N__12800\ : std_logic;
signal \N__12797\ : std_logic;
signal \N__12794\ : std_logic;
signal \N__12793\ : std_logic;
signal \N__12792\ : std_logic;
signal \N__12789\ : std_logic;
signal \N__12784\ : std_logic;
signal \N__12781\ : std_logic;
signal \N__12776\ : std_logic;
signal \N__12773\ : std_logic;
signal \N__12770\ : std_logic;
signal \N__12767\ : std_logic;
signal \N__12766\ : std_logic;
signal \N__12765\ : std_logic;
signal \N__12762\ : std_logic;
signal \N__12759\ : std_logic;
signal \N__12756\ : std_logic;
signal \N__12753\ : std_logic;
signal \N__12746\ : std_logic;
signal \N__12743\ : std_logic;
signal \N__12742\ : std_logic;
signal \N__12739\ : std_logic;
signal \N__12736\ : std_logic;
signal \N__12733\ : std_logic;
signal \N__12728\ : std_logic;
signal \N__12727\ : std_logic;
signal \N__12726\ : std_logic;
signal \N__12723\ : std_logic;
signal \N__12720\ : std_logic;
signal \N__12715\ : std_logic;
signal \N__12712\ : std_logic;
signal \N__12709\ : std_logic;
signal \N__12704\ : std_logic;
signal \N__12701\ : std_logic;
signal \N__12698\ : std_logic;
signal \N__12695\ : std_logic;
signal \N__12692\ : std_logic;
signal \N__12689\ : std_logic;
signal \N__12686\ : std_logic;
signal \N__12685\ : std_logic;
signal \N__12682\ : std_logic;
signal \N__12681\ : std_logic;
signal \N__12678\ : std_logic;
signal \N__12675\ : std_logic;
signal \N__12672\ : std_logic;
signal \N__12665\ : std_logic;
signal \N__12662\ : std_logic;
signal \N__12661\ : std_logic;
signal \N__12660\ : std_logic;
signal \N__12657\ : std_logic;
signal \N__12654\ : std_logic;
signal \N__12651\ : std_logic;
signal \N__12648\ : std_logic;
signal \N__12645\ : std_logic;
signal \N__12638\ : std_logic;
signal \N__12635\ : std_logic;
signal \N__12632\ : std_logic;
signal \N__12629\ : std_logic;
signal \N__12626\ : std_logic;
signal \N__12623\ : std_logic;
signal \N__12620\ : std_logic;
signal \N__12617\ : std_logic;
signal \N__12616\ : std_logic;
signal \N__12611\ : std_logic;
signal \N__12608\ : std_logic;
signal \N__12607\ : std_logic;
signal \N__12606\ : std_logic;
signal \N__12605\ : std_logic;
signal \N__12602\ : std_logic;
signal \N__12601\ : std_logic;
signal \N__12600\ : std_logic;
signal \N__12599\ : std_logic;
signal \N__12598\ : std_logic;
signal \N__12595\ : std_logic;
signal \N__12590\ : std_logic;
signal \N__12587\ : std_logic;
signal \N__12578\ : std_logic;
signal \N__12575\ : std_logic;
signal \N__12566\ : std_logic;
signal \N__12563\ : std_logic;
signal \N__12560\ : std_logic;
signal \N__12557\ : std_logic;
signal \N__12554\ : std_logic;
signal \N__12551\ : std_logic;
signal \N__12548\ : std_logic;
signal \N__12545\ : std_logic;
signal \N__12542\ : std_logic;
signal \N__12539\ : std_logic;
signal \N__12536\ : std_logic;
signal \N__12533\ : std_logic;
signal \N__12530\ : std_logic;
signal \N__12527\ : std_logic;
signal \N__12524\ : std_logic;
signal \N__12521\ : std_logic;
signal \N__12518\ : std_logic;
signal \N__12515\ : std_logic;
signal \N__12512\ : std_logic;
signal \N__12511\ : std_logic;
signal \N__12508\ : std_logic;
signal \N__12507\ : std_logic;
signal \N__12504\ : std_logic;
signal \N__12501\ : std_logic;
signal \N__12498\ : std_logic;
signal \N__12491\ : std_logic;
signal \N__12488\ : std_logic;
signal \N__12487\ : std_logic;
signal \N__12484\ : std_logic;
signal \N__12481\ : std_logic;
signal \N__12478\ : std_logic;
signal \N__12473\ : std_logic;
signal \N__12472\ : std_logic;
signal \N__12471\ : std_logic;
signal \N__12470\ : std_logic;
signal \N__12467\ : std_logic;
signal \N__12466\ : std_logic;
signal \N__12463\ : std_logic;
signal \N__12460\ : std_logic;
signal \N__12459\ : std_logic;
signal \N__12456\ : std_logic;
signal \N__12453\ : std_logic;
signal \N__12450\ : std_logic;
signal \N__12443\ : std_logic;
signal \N__12434\ : std_logic;
signal \N__12431\ : std_logic;
signal \N__12428\ : std_logic;
signal \N__12425\ : std_logic;
signal \N__12422\ : std_logic;
signal \N__12419\ : std_logic;
signal \N__12416\ : std_logic;
signal \N__12413\ : std_logic;
signal \N__12410\ : std_logic;
signal \N__12407\ : std_logic;
signal \N__12404\ : std_logic;
signal \N__12401\ : std_logic;
signal \N__12398\ : std_logic;
signal \N__12397\ : std_logic;
signal \N__12394\ : std_logic;
signal \N__12393\ : std_logic;
signal \N__12390\ : std_logic;
signal \N__12387\ : std_logic;
signal \N__12384\ : std_logic;
signal \N__12377\ : std_logic;
signal \N__12374\ : std_logic;
signal \N__12371\ : std_logic;
signal \N__12368\ : std_logic;
signal \N__12365\ : std_logic;
signal \N__12362\ : std_logic;
signal \N__12359\ : std_logic;
signal \N__12356\ : std_logic;
signal \N__12353\ : std_logic;
signal \N__12350\ : std_logic;
signal \N__12347\ : std_logic;
signal \N__12344\ : std_logic;
signal \N__12341\ : std_logic;
signal \N__12338\ : std_logic;
signal \N__12335\ : std_logic;
signal \N__12334\ : std_logic;
signal \N__12331\ : std_logic;
signal \N__12330\ : std_logic;
signal \N__12327\ : std_logic;
signal \N__12324\ : std_logic;
signal \N__12321\ : std_logic;
signal \N__12314\ : std_logic;
signal \N__12311\ : std_logic;
signal \N__12308\ : std_logic;
signal \N__12307\ : std_logic;
signal \N__12306\ : std_logic;
signal \N__12303\ : std_logic;
signal \N__12300\ : std_logic;
signal \N__12297\ : std_logic;
signal \N__12292\ : std_logic;
signal \N__12287\ : std_logic;
signal \N__12284\ : std_logic;
signal \N__12281\ : std_logic;
signal \N__12278\ : std_logic;
signal \N__12275\ : std_logic;
signal \N__12272\ : std_logic;
signal \N__12271\ : std_logic;
signal \N__12268\ : std_logic;
signal \N__12267\ : std_logic;
signal \N__12264\ : std_logic;
signal \N__12261\ : std_logic;
signal \N__12258\ : std_logic;
signal \N__12251\ : std_logic;
signal \N__12248\ : std_logic;
signal \N__12245\ : std_logic;
signal \N__12242\ : std_logic;
signal \N__12239\ : std_logic;
signal \N__12236\ : std_logic;
signal \N__12233\ : std_logic;
signal \N__12230\ : std_logic;
signal \N__12229\ : std_logic;
signal \N__12228\ : std_logic;
signal \N__12225\ : std_logic;
signal \N__12222\ : std_logic;
signal \N__12219\ : std_logic;
signal \N__12216\ : std_logic;
signal \N__12209\ : std_logic;
signal \N__12206\ : std_logic;
signal \N__12205\ : std_logic;
signal \N__12202\ : std_logic;
signal \N__12199\ : std_logic;
signal \N__12194\ : std_logic;
signal \N__12191\ : std_logic;
signal \N__12188\ : std_logic;
signal \N__12187\ : std_logic;
signal \N__12184\ : std_logic;
signal \N__12181\ : std_logic;
signal \N__12178\ : std_logic;
signal \N__12175\ : std_logic;
signal \N__12172\ : std_logic;
signal \N__12167\ : std_logic;
signal \N__12166\ : std_logic;
signal \N__12165\ : std_logic;
signal \N__12162\ : std_logic;
signal \N__12159\ : std_logic;
signal \N__12156\ : std_logic;
signal \N__12149\ : std_logic;
signal \N__12146\ : std_logic;
signal \N__12143\ : std_logic;
signal \N__12140\ : std_logic;
signal \N__12137\ : std_logic;
signal \N__12134\ : std_logic;
signal \N__12131\ : std_logic;
signal \N__12130\ : std_logic;
signal \N__12127\ : std_logic;
signal \N__12124\ : std_logic;
signal \N__12119\ : std_logic;
signal \N__12116\ : std_logic;
signal \N__12113\ : std_logic;
signal \N__12110\ : std_logic;
signal \N__12107\ : std_logic;
signal \N__12104\ : std_logic;
signal \N__12101\ : std_logic;
signal \N__12098\ : std_logic;
signal \N__12095\ : std_logic;
signal \N__12094\ : std_logic;
signal \N__12091\ : std_logic;
signal \N__12090\ : std_logic;
signal \N__12087\ : std_logic;
signal \N__12084\ : std_logic;
signal \N__12081\ : std_logic;
signal \N__12074\ : std_logic;
signal \N__12071\ : std_logic;
signal \N__12068\ : std_logic;
signal \N__12065\ : std_logic;
signal \N__12062\ : std_logic;
signal \N__12059\ : std_logic;
signal \N__12056\ : std_logic;
signal \N__12053\ : std_logic;
signal \N__12050\ : std_logic;
signal \N__12047\ : std_logic;
signal \N__12044\ : std_logic;
signal \N__12043\ : std_logic;
signal \N__12040\ : std_logic;
signal \N__12037\ : std_logic;
signal \N__12034\ : std_logic;
signal \N__12031\ : std_logic;
signal \N__12028\ : std_logic;
signal \N__12025\ : std_logic;
signal \N__12020\ : std_logic;
signal \N__12017\ : std_logic;
signal \N__12014\ : std_logic;
signal \N__12011\ : std_logic;
signal \N__12008\ : std_logic;
signal \N__12005\ : std_logic;
signal \N__12004\ : std_logic;
signal \N__12001\ : std_logic;
signal \N__11998\ : std_logic;
signal \N__11995\ : std_logic;
signal \N__11990\ : std_logic;
signal \N__11987\ : std_logic;
signal \N__11984\ : std_logic;
signal \N__11983\ : std_logic;
signal \N__11982\ : std_logic;
signal \N__11979\ : std_logic;
signal \N__11976\ : std_logic;
signal \N__11973\ : std_logic;
signal \N__11970\ : std_logic;
signal \N__11967\ : std_logic;
signal \N__11960\ : std_logic;
signal \N__11957\ : std_logic;
signal \N__11954\ : std_logic;
signal \N__11951\ : std_logic;
signal \N__11948\ : std_logic;
signal \N__11945\ : std_logic;
signal \N__11942\ : std_logic;
signal \N__11939\ : std_logic;
signal \N__11936\ : std_logic;
signal \N__11935\ : std_logic;
signal \N__11930\ : std_logic;
signal \N__11927\ : std_logic;
signal \N__11924\ : std_logic;
signal \N__11921\ : std_logic;
signal \N__11920\ : std_logic;
signal \N__11919\ : std_logic;
signal \N__11916\ : std_logic;
signal \N__11913\ : std_logic;
signal \N__11910\ : std_logic;
signal \N__11903\ : std_logic;
signal \N__11902\ : std_logic;
signal \N__11899\ : std_logic;
signal \N__11896\ : std_logic;
signal \N__11893\ : std_logic;
signal \N__11888\ : std_logic;
signal \N__11885\ : std_logic;
signal \N__11882\ : std_logic;
signal \N__11879\ : std_logic;
signal \N__11876\ : std_logic;
signal \N__11873\ : std_logic;
signal \N__11870\ : std_logic;
signal \N__11867\ : std_logic;
signal \N__11864\ : std_logic;
signal \N__11863\ : std_logic;
signal \N__11862\ : std_logic;
signal \N__11859\ : std_logic;
signal \N__11856\ : std_logic;
signal \N__11851\ : std_logic;
signal \N__11846\ : std_logic;
signal \N__11843\ : std_logic;
signal \N__11840\ : std_logic;
signal \N__11837\ : std_logic;
signal \N__11834\ : std_logic;
signal \N__11831\ : std_logic;
signal \N__11828\ : std_logic;
signal \N__11825\ : std_logic;
signal \N__11822\ : std_logic;
signal \N__11819\ : std_logic;
signal \N__11816\ : std_logic;
signal \N__11813\ : std_logic;
signal \N__11812\ : std_logic;
signal \N__11809\ : std_logic;
signal \N__11808\ : std_logic;
signal \N__11805\ : std_logic;
signal \N__11802\ : std_logic;
signal \N__11799\ : std_logic;
signal \N__11792\ : std_logic;
signal \N__11789\ : std_logic;
signal \N__11786\ : std_logic;
signal \N__11783\ : std_logic;
signal \N__11780\ : std_logic;
signal \N__11777\ : std_logic;
signal \N__11774\ : std_logic;
signal \N__11771\ : std_logic;
signal \N__11768\ : std_logic;
signal \N__11765\ : std_logic;
signal \N__11762\ : std_logic;
signal \N__11759\ : std_logic;
signal \N__11756\ : std_logic;
signal \N__11753\ : std_logic;
signal \N__11750\ : std_logic;
signal \N__11747\ : std_logic;
signal \N__11744\ : std_logic;
signal \N__11741\ : std_logic;
signal \N__11738\ : std_logic;
signal \N__11735\ : std_logic;
signal \N__11732\ : std_logic;
signal \N__11731\ : std_logic;
signal \N__11728\ : std_logic;
signal \N__11727\ : std_logic;
signal \N__11724\ : std_logic;
signal \N__11721\ : std_logic;
signal \N__11718\ : std_logic;
signal \N__11711\ : std_logic;
signal \N__11708\ : std_logic;
signal \N__11705\ : std_logic;
signal \N__11702\ : std_logic;
signal \N__11699\ : std_logic;
signal \N__11696\ : std_logic;
signal \N__11693\ : std_logic;
signal \N__11690\ : std_logic;
signal \N__11687\ : std_logic;
signal \N__11684\ : std_logic;
signal \N__11681\ : std_logic;
signal \N__11678\ : std_logic;
signal \N__11675\ : std_logic;
signal \N__11672\ : std_logic;
signal \N__11669\ : std_logic;
signal \N__11666\ : std_logic;
signal \N__11663\ : std_logic;
signal \N__11660\ : std_logic;
signal \N__11657\ : std_logic;
signal \N__11654\ : std_logic;
signal \N__11651\ : std_logic;
signal \N__11648\ : std_logic;
signal \N__11645\ : std_logic;
signal \N__11642\ : std_logic;
signal \N__11639\ : std_logic;
signal \N__11636\ : std_logic;
signal \N__11633\ : std_logic;
signal \N__11630\ : std_logic;
signal \N__11627\ : std_logic;
signal \N__11624\ : std_logic;
signal \N__11621\ : std_logic;
signal \N__11618\ : std_logic;
signal \N__11615\ : std_logic;
signal \N__11612\ : std_logic;
signal \N__11609\ : std_logic;
signal \N__11606\ : std_logic;
signal \N__11603\ : std_logic;
signal \N__11600\ : std_logic;
signal \N__11597\ : std_logic;
signal \N__11594\ : std_logic;
signal \N__11591\ : std_logic;
signal \N__11588\ : std_logic;
signal \N__11585\ : std_logic;
signal \N__11582\ : std_logic;
signal \N__11579\ : std_logic;
signal \N__11576\ : std_logic;
signal \N__11573\ : std_logic;
signal \N__11570\ : std_logic;
signal \N__11567\ : std_logic;
signal \N__11564\ : std_logic;
signal \N__11561\ : std_logic;
signal \N__11558\ : std_logic;
signal \N__11555\ : std_logic;
signal \N__11552\ : std_logic;
signal \N__11549\ : std_logic;
signal \N__11546\ : std_logic;
signal \N__11543\ : std_logic;
signal \N__11540\ : std_logic;
signal \N__11537\ : std_logic;
signal \N__11536\ : std_logic;
signal \N__11535\ : std_logic;
signal \N__11532\ : std_logic;
signal \N__11529\ : std_logic;
signal \N__11526\ : std_logic;
signal \N__11521\ : std_logic;
signal \N__11516\ : std_logic;
signal \N__11513\ : std_logic;
signal \N__11510\ : std_logic;
signal \N__11507\ : std_logic;
signal \N__11504\ : std_logic;
signal \N__11501\ : std_logic;
signal \N__11498\ : std_logic;
signal \N__11495\ : std_logic;
signal \N__11492\ : std_logic;
signal \N__11489\ : std_logic;
signal \N__11486\ : std_logic;
signal \N__11483\ : std_logic;
signal \N__11480\ : std_logic;
signal \N__11477\ : std_logic;
signal \N__11474\ : std_logic;
signal \N__11471\ : std_logic;
signal \N__11468\ : std_logic;
signal \N__11465\ : std_logic;
signal \N__11462\ : std_logic;
signal \N__11459\ : std_logic;
signal \N__11456\ : std_logic;
signal \N__11453\ : std_logic;
signal \N__11450\ : std_logic;
signal \N__11447\ : std_logic;
signal \N__11444\ : std_logic;
signal \N__11441\ : std_logic;
signal \N__11438\ : std_logic;
signal \N__11435\ : std_logic;
signal \N__11432\ : std_logic;
signal \N__11429\ : std_logic;
signal \N__11426\ : std_logic;
signal \N__11423\ : std_logic;
signal \N__11420\ : std_logic;
signal \N__11417\ : std_logic;
signal \N__11414\ : std_logic;
signal \N__11411\ : std_logic;
signal \N__11408\ : std_logic;
signal \N__11405\ : std_logic;
signal \N__11402\ : std_logic;
signal \N__11399\ : std_logic;
signal \N__11396\ : std_logic;
signal \N__11393\ : std_logic;
signal \N__11390\ : std_logic;
signal \N__11387\ : std_logic;
signal \N__11384\ : std_logic;
signal \N__11381\ : std_logic;
signal \N__11378\ : std_logic;
signal \N__11375\ : std_logic;
signal \N__11372\ : std_logic;
signal \N__11369\ : std_logic;
signal \N__11366\ : std_logic;
signal \N__11363\ : std_logic;
signal \N__11360\ : std_logic;
signal \N__11357\ : std_logic;
signal \N__11354\ : std_logic;
signal \N__11351\ : std_logic;
signal \N__11348\ : std_logic;
signal \N__11345\ : std_logic;
signal \N__11342\ : std_logic;
signal \N__11339\ : std_logic;
signal \N__11336\ : std_logic;
signal \N__11333\ : std_logic;
signal \N__11330\ : std_logic;
signal \N__11327\ : std_logic;
signal \N__11324\ : std_logic;
signal \N__11321\ : std_logic;
signal \N__11318\ : std_logic;
signal \N__11315\ : std_logic;
signal \N__11312\ : std_logic;
signal \N__11309\ : std_logic;
signal \N__11306\ : std_logic;
signal \N__11303\ : std_logic;
signal \N__11300\ : std_logic;
signal \N__11297\ : std_logic;
signal \N__11294\ : std_logic;
signal \N__11291\ : std_logic;
signal \N__11288\ : std_logic;
signal \N__11285\ : std_logic;
signal \N__11282\ : std_logic;
signal \N__11279\ : std_logic;
signal \N__11276\ : std_logic;
signal \N__11273\ : std_logic;
signal \N__11270\ : std_logic;
signal \N__11267\ : std_logic;
signal \N__11264\ : std_logic;
signal \N__11261\ : std_logic;
signal \N__11258\ : std_logic;
signal \N__11255\ : std_logic;
signal \N__11252\ : std_logic;
signal \N__11249\ : std_logic;
signal \N__11246\ : std_logic;
signal \N__11243\ : std_logic;
signal \N__11240\ : std_logic;
signal \N__11237\ : std_logic;
signal \N__11234\ : std_logic;
signal \N__11231\ : std_logic;
signal \N__11230\ : std_logic;
signal \N__11227\ : std_logic;
signal \N__11226\ : std_logic;
signal \N__11223\ : std_logic;
signal \N__11220\ : std_logic;
signal \N__11217\ : std_logic;
signal \N__11212\ : std_logic;
signal \N__11207\ : std_logic;
signal \N__11204\ : std_logic;
signal \N__11201\ : std_logic;
signal \N__11198\ : std_logic;
signal \N__11197\ : std_logic;
signal \N__11192\ : std_logic;
signal \N__11191\ : std_logic;
signal \N__11188\ : std_logic;
signal \N__11185\ : std_logic;
signal \N__11182\ : std_logic;
signal \N__11177\ : std_logic;
signal \N__11174\ : std_logic;
signal \N__11171\ : std_logic;
signal \N__11168\ : std_logic;
signal \N__11165\ : std_logic;
signal \N__11162\ : std_logic;
signal \N__11159\ : std_logic;
signal \N__11156\ : std_logic;
signal \N__11153\ : std_logic;
signal \N__11150\ : std_logic;
signal \N__11147\ : std_logic;
signal \N__11144\ : std_logic;
signal \N__11141\ : std_logic;
signal \N__11138\ : std_logic;
signal \N__11137\ : std_logic;
signal \N__11136\ : std_logic;
signal \N__11133\ : std_logic;
signal \N__11128\ : std_logic;
signal \N__11123\ : std_logic;
signal \N__11120\ : std_logic;
signal \N__11117\ : std_logic;
signal \N__11114\ : std_logic;
signal \N__11111\ : std_logic;
signal \N__11108\ : std_logic;
signal \N__11105\ : std_logic;
signal \N__11102\ : std_logic;
signal \N__11099\ : std_logic;
signal \N__11096\ : std_logic;
signal \CLK_pad_gb_input\ : std_logic;
signal \VCCG0\ : std_logic;
signal \GNDG0\ : std_logic;
signal \bfn_2_17_0_\ : std_logic;
signal \eeprom.n3454\ : std_logic;
signal \eeprom.n3455\ : std_logic;
signal \eeprom.n3456\ : std_logic;
signal \eeprom.n3457\ : std_logic;
signal \eeprom.n3458\ : std_logic;
signal \eeprom.n3459\ : std_logic;
signal \eeprom.n3460\ : std_logic;
signal \eeprom.n3461\ : std_logic;
signal \bfn_2_18_0_\ : std_logic;
signal \eeprom.n3462\ : std_logic;
signal \eeprom.n3463\ : std_logic;
signal \eeprom.delay_counter_11\ : std_logic;
signal \eeprom.n3464\ : std_logic;
signal \eeprom.n3465\ : std_logic;
signal \eeprom.delay_counter_13\ : std_logic;
signal \eeprom.n3466\ : std_logic;
signal \eeprom.n3467\ : std_logic;
signal \eeprom.n3468\ : std_logic;
signal \eeprom.n3469\ : std_logic;
signal \eeprom.delay_counter_16\ : std_logic;
signal \bfn_2_19_0_\ : std_logic;
signal \eeprom.n3470\ : std_logic;
signal \eeprom.n3471\ : std_logic;
signal \eeprom.n3472\ : std_logic;
signal \eeprom.n3473\ : std_logic;
signal \eeprom.n3474\ : std_logic;
signal \eeprom.n3475\ : std_logic;
signal \eeprom.n3476\ : std_logic;
signal \eeprom.n3477\ : std_logic;
signal \bfn_2_20_0_\ : std_logic;
signal \eeprom.n3478\ : std_logic;
signal \eeprom.n3479\ : std_logic;
signal \eeprom.n3480\ : std_logic;
signal \eeprom.n3481\ : std_logic;
signal \eeprom.n3482\ : std_logic;
signal \eeprom.n3483\ : std_logic;
signal \eeprom.n3484\ : std_logic;
signal \bfn_2_21_0_\ : std_logic;
signal \eeprom.n3786\ : std_logic;
signal \eeprom.n31_adj_457\ : std_logic;
signal \eeprom.n3787\ : std_logic;
signal \eeprom.n3788\ : std_logic;
signal \eeprom.n3789\ : std_logic;
signal \eeprom.n28_adj_461\ : std_logic;
signal \eeprom.n3790\ : std_logic;
signal \eeprom.n27_adj_462\ : std_logic;
signal \eeprom.n3791\ : std_logic;
signal \eeprom.n3792\ : std_logic;
signal \eeprom.n3793\ : std_logic;
signal \bfn_2_22_0_\ : std_logic;
signal \eeprom.n24_adj_463\ : std_logic;
signal \eeprom.n3794\ : std_logic;
signal \eeprom.n23\ : std_logic;
signal \eeprom.n3795\ : std_logic;
signal \eeprom.n22_adj_448\ : std_logic;
signal \eeprom.n22_adj_447\ : std_logic;
signal \eeprom.n3796\ : std_logic;
signal \eeprom.n21_adj_440\ : std_logic;
signal \eeprom.n3797\ : std_logic;
signal \eeprom.n20_adj_431\ : std_logic;
signal \eeprom.n20_adj_430\ : std_logic;
signal \eeprom.n3798\ : std_logic;
signal \eeprom.n3799\ : std_logic;
signal \eeprom.n18_adj_427\ : std_logic;
signal \eeprom.n3800\ : std_logic;
signal \eeprom.n3801\ : std_logic;
signal \eeprom.n17_adj_425\ : std_logic;
signal \eeprom.n17\ : std_logic;
signal \bfn_2_23_0_\ : std_logic;
signal \eeprom.n16_adj_424\ : std_logic;
signal \eeprom.n3802\ : std_logic;
signal \eeprom.n3803\ : std_logic;
signal \eeprom.n14_adj_413\ : std_logic;
signal \eeprom.n3804\ : std_logic;
signal \eeprom.n3805\ : std_logic;
signal \eeprom.n3806\ : std_logic;
signal \eeprom.n3807\ : std_logic;
signal \eeprom.n3808\ : std_logic;
signal \eeprom.n3809\ : std_logic;
signal \bfn_2_24_0_\ : std_logic;
signal \eeprom.n8_adj_407\ : std_logic;
signal \eeprom.n3810\ : std_logic;
signal \eeprom.n7_adj_405\ : std_logic;
signal \eeprom.n3811\ : std_logic;
signal \eeprom.n6_adj_403\ : std_logic;
signal \eeprom.n3812\ : std_logic;
signal \eeprom.n3813\ : std_logic;
signal \eeprom.n4_adj_397\ : std_logic;
signal \eeprom.n3814\ : std_logic;
signal \eeprom.n3_adj_396\ : std_logic;
signal \eeprom.n3815\ : std_logic;
signal \eeprom.n3816\ : std_logic;
signal \eeprom.n14\ : std_logic;
signal \eeprom.delay_counter_19\ : std_logic;
signal \eeprom.n11_adj_410\ : std_logic;
signal \bfn_3_17_0_\ : std_logic;
signal \eeprom.n3448\ : std_logic;
signal \eeprom.n3449\ : std_logic;
signal \eeprom.n3450\ : std_logic;
signal \eeprom.n3451\ : std_logic;
signal \eeprom.n3452\ : std_logic;
signal \eeprom.n3453\ : std_logic;
signal \eeprom.n30_adj_458\ : std_logic;
signal \eeprom.n26\ : std_logic;
signal \eeprom.delay_counter_30\ : std_logic;
signal \eeprom.n3\ : std_logic;
signal \eeprom.n1341\ : std_logic;
signal \eeprom.n1256_cascade_\ : std_logic;
signal \eeprom.n5_adj_400\ : std_logic;
signal \eeprom.n15_adj_415\ : std_logic;
signal \eeprom.n33\ : std_logic;
signal \eeprom.delay_counter_25\ : std_logic;
signal \eeprom.n8\ : std_logic;
signal \eeprom.n1141_cascade_\ : std_logic;
signal \eeprom.n2_adj_395\ : std_logic;
signal \eeprom.n4399_cascade_\ : std_logic;
signal \eeprom.n1343\ : std_logic;
signal \eeprom.n1141\ : std_logic;
signal \eeprom.n4405_cascade_\ : std_logic;
signal \eeprom.delay_counter_28\ : std_logic;
signal \eeprom.n5\ : std_logic;
signal \eeprom.n1342\ : std_logic;
signal \eeprom.n6_adj_402\ : std_logic;
signal \eeprom.delay_counter_27\ : std_logic;
signal \eeprom.n1139\ : std_logic;
signal \eeprom.n25\ : std_logic;
signal \eeprom.n9\ : std_logic;
signal \eeprom.delay_counter_24\ : std_logic;
signal \eeprom.n9_adj_408\ : std_logic;
signal \eeprom.n32\ : std_logic;
signal \eeprom.delay_counter_26\ : std_logic;
signal \eeprom.n7\ : std_logic;
signal \eeprom.n1140\ : std_logic;
signal \eeprom.delay_counter_29\ : std_logic;
signal \eeprom.n4\ : std_logic;
signal \eeprom.n1137\ : std_logic;
signal \eeprom.n1339\ : std_logic;
signal \eeprom.n1137_cascade_\ : std_logic;
signal \eeprom.n24_adj_467\ : std_logic;
signal \eeprom.delay_counter_9\ : std_logic;
signal \eeprom.n33_adj_483\ : std_logic;
signal \eeprom.n13_adj_412\ : std_logic;
signal \eeprom.n10_adj_409\ : std_logic;
signal \eeprom.n19_adj_428\ : std_logic;
signal \eeprom.delay_counter_18\ : std_logic;
signal \eeprom.n15_adj_414\ : std_logic;
signal \eeprom.delay_counter_23\ : std_logic;
signal \eeprom.n10\ : std_logic;
signal \eeprom.n18_adj_426\ : std_logic;
signal \eeprom.delay_counter_15\ : std_logic;
signal \bfn_3_23_0_\ : std_logic;
signal \eeprom.n3551\ : std_logic;
signal \eeprom.n3552\ : std_logic;
signal \eeprom.n2383\ : std_logic;
signal \eeprom.n3553\ : std_logic;
signal \eeprom.n3554\ : std_logic;
signal \eeprom.n3555\ : std_logic;
signal \eeprom.n3556\ : std_logic;
signal \eeprom.n3557\ : std_logic;
signal \eeprom.n3558\ : std_logic;
signal \bfn_3_24_0_\ : std_logic;
signal \eeprom.n3559\ : std_logic;
signal \eeprom.n3560\ : std_logic;
signal \eeprom.n3561\ : std_logic;
signal \eeprom.n2386\ : std_logic;
signal \eeprom.n2381\ : std_logic;
signal \eeprom.n2384\ : std_logic;
signal \eeprom.n2378\ : std_logic;
signal \eeprom.n4733\ : std_logic;
signal \eeprom.n1340\ : std_logic;
signal \eeprom.n1138\ : std_logic;
signal \eeprom.n1915_cascade_\ : std_logic;
signal \eeprom.n1135\ : std_logic;
signal \eeprom.n4405\ : std_logic;
signal \eeprom.n1337\ : std_logic;
signal \eeprom.n12_adj_411\ : std_logic;
signal \eeprom.n25_adj_471\ : std_logic;
signal \eeprom.delay_counter_8\ : std_logic;
signal \eeprom.delay_counter_17\ : std_logic;
signal \eeprom.n16_adj_377\ : std_logic;
signal \eeprom.n4734\ : std_logic;
signal \eeprom.n1256\ : std_logic;
signal \bfn_4_19_0_\ : std_logic;
signal \eeprom.n3517\ : std_logic;
signal \eeprom.n3518\ : std_logic;
signal \eeprom.n3519\ : std_logic;
signal \eeprom.n3520\ : std_logic;
signal \eeprom.n3521\ : std_logic;
signal \eeprom.n3522\ : std_logic;
signal \eeprom.n3523\ : std_logic;
signal \eeprom.n26_adj_469\ : std_logic;
signal \eeprom.delay_counter_7\ : std_logic;
signal \eeprom.n1984\ : std_logic;
signal \eeprom.n1985\ : std_logic;
signal \eeprom.n2017_cascade_\ : std_logic;
signal \eeprom.n1917\ : std_logic;
signal \eeprom.n4437\ : std_logic;
signal \eeprom.n1918\ : std_logic;
signal \eeprom.n4441_cascade_\ : std_logic;
signal \eeprom.n1912\ : std_logic;
signal \eeprom.n1916\ : std_logic;
signal \eeprom.n1945_cascade_\ : std_logic;
signal \eeprom.n1983\ : std_logic;
signal \eeprom.n1981\ : std_logic;
signal \eeprom.n1914\ : std_logic;
signal \eeprom.n1915\ : std_logic;
signal \eeprom.n1982\ : std_logic;
signal \eeprom.n2014_cascade_\ : std_logic;
signal \eeprom.n4415\ : std_logic;
signal \eeprom.n1919\ : std_logic;
signal \eeprom.n1986\ : std_logic;
signal \eeprom.n1913\ : std_logic;
signal \eeprom.n1945\ : std_logic;
signal \eeprom.n1980\ : std_logic;
signal \eeprom.n4419\ : std_logic;
signal \eeprom.n4575_cascade_\ : std_logic;
signal \eeprom.n4579\ : std_logic;
signal \eeprom.n13\ : std_logic;
signal \eeprom.delay_counter_20\ : std_logic;
signal \eeprom.n4479_cascade_\ : std_logic;
signal \eeprom.n4477\ : std_logic;
signal \eeprom.n2385\ : std_logic;
signal \eeprom.n2341_cascade_\ : std_logic;
signal \eeprom.n2376\ : std_logic;
signal \eeprom.n2312\ : std_logic;
signal \eeprom.n2312_cascade_\ : std_logic;
signal \eeprom.n2379\ : std_logic;
signal \eeprom.n2411_cascade_\ : std_logic;
signal \eeprom.n4133\ : std_logic;
signal \eeprom.n12_adj_472_cascade_\ : std_logic;
signal \eeprom.n2382\ : std_logic;
signal \eeprom.n2377\ : std_logic;
signal \eeprom.n2380\ : std_logic;
signal \eeprom.n2341\ : std_logic;
signal \bfn_4_25_0_\ : std_logic;
signal \eeprom.n2418\ : std_logic;
signal \eeprom.n2485\ : std_logic;
signal \eeprom.n3562\ : std_logic;
signal \eeprom.n2417\ : std_logic;
signal \eeprom.n2484\ : std_logic;
signal \eeprom.n3563\ : std_logic;
signal \eeprom.n2416\ : std_logic;
signal \eeprom.n2483\ : std_logic;
signal \eeprom.n3564\ : std_logic;
signal \eeprom.n2415\ : std_logic;
signal \eeprom.n2482\ : std_logic;
signal \eeprom.n3565\ : std_logic;
signal \eeprom.n2414\ : std_logic;
signal \eeprom.n2481\ : std_logic;
signal \eeprom.n3566\ : std_logic;
signal \eeprom.n3567\ : std_logic;
signal \eeprom.n3568\ : std_logic;
signal \eeprom.n3569\ : std_logic;
signal \bfn_4_26_0_\ : std_logic;
signal \eeprom.n3570\ : std_logic;
signal \eeprom.n3571\ : std_logic;
signal \eeprom.n3572\ : std_logic;
signal \eeprom.n2407\ : std_logic;
signal \eeprom.n3573\ : std_logic;
signal \eeprom.n2410\ : std_logic;
signal \eeprom.n2477\ : std_logic;
signal \eeprom.n2476\ : std_logic;
signal \eeprom.n2409\ : std_logic;
signal n4826 : std_logic;
signal \n4825_cascade_\ : std_logic;
signal \LED_c\ : std_logic;
signal \eeprom.n23_adj_464\ : std_logic;
signal \eeprom.delay_counter_10\ : std_logic;
signal \eeprom.n2615_cascade_\ : std_logic;
signal \eeprom.n4497_cascade_\ : std_logic;
signal \eeprom.n4501_cascade_\ : std_logic;
signal \eeprom.n13_adj_474_cascade_\ : std_logic;
signal \eeprom.n11_adj_473\ : std_logic;
signal \eeprom.n2539_cascade_\ : std_logic;
signal \eeprom.delay_counter_14\ : std_logic;
signal \eeprom.n19_adj_429\ : std_logic;
signal \eeprom.n30\ : std_logic;
signal \eeprom.n2114_cascade_\ : std_logic;
signal \eeprom.n2411\ : std_logic;
signal \eeprom.n2478\ : std_logic;
signal \eeprom.n2419\ : std_logic;
signal \eeprom.n2486\ : std_logic;
signal \bfn_5_22_0_\ : std_logic;
signal \eeprom.n2018\ : std_logic;
signal \eeprom.n2085\ : std_logic;
signal \eeprom.n3524\ : std_logic;
signal \eeprom.n3525\ : std_logic;
signal \eeprom.n3526\ : std_logic;
signal \eeprom.n2015\ : std_logic;
signal \eeprom.n2082\ : std_logic;
signal \eeprom.n3527\ : std_logic;
signal \eeprom.n3528\ : std_logic;
signal \eeprom.n2013\ : std_logic;
signal \eeprom.n2080\ : std_logic;
signal \eeprom.n3529\ : std_logic;
signal \eeprom.n3530\ : std_logic;
signal \eeprom.n3531\ : std_logic;
signal \eeprom.n2011\ : std_logic;
signal \bfn_5_23_0_\ : std_logic;
signal \eeprom.n2081\ : std_logic;
signal \eeprom.n2014\ : std_logic;
signal \eeprom.n2012\ : std_logic;
signal \eeprom.n2079\ : std_logic;
signal \eeprom.n2083\ : std_logic;
signal \eeprom.n2016\ : std_logic;
signal \eeprom.n7_adj_470\ : std_logic;
signal \eeprom.n2019\ : std_logic;
signal \eeprom.n2086\ : std_logic;
signal \eeprom.n2309\ : std_logic;
signal \eeprom.n2319\ : std_logic;
signal \eeprom.n4509_cascade_\ : std_logic;
signal \eeprom.n8_adj_468\ : std_logic;
signal \eeprom.n2310\ : std_logic;
signal \eeprom.n6_cascade_\ : std_logic;
signal \eeprom.n2242_cascade_\ : std_logic;
signal \eeprom.n2044\ : std_logic;
signal \eeprom.n2084\ : std_logic;
signal \eeprom.n2214_cascade_\ : std_logic;
signal \eeprom.n2313\ : std_logic;
signal \eeprom.n2313_cascade_\ : std_logic;
signal \eeprom.n4505\ : std_logic;
signal \eeprom.n11\ : std_logic;
signal \eeprom.delay_counter_22\ : std_logic;
signal \eeprom.n2315\ : std_logic;
signal \eeprom.n2311\ : std_logic;
signal \eeprom.n4461\ : std_logic;
signal \eeprom.n4463\ : std_logic;
signal \eeprom.n4225_cascade_\ : std_logic;
signal \eeprom.n2143_cascade_\ : std_logic;
signal \bfn_5_27_0_\ : std_logic;
signal \eeprom.n2118\ : std_logic;
signal \eeprom.n2185\ : std_logic;
signal \eeprom.n3532\ : std_logic;
signal \eeprom.n2117\ : std_logic;
signal \eeprom.n2184\ : std_logic;
signal \eeprom.n3533\ : std_logic;
signal \eeprom.n2116\ : std_logic;
signal \eeprom.n2183\ : std_logic;
signal \eeprom.n3534\ : std_logic;
signal \eeprom.n2115\ : std_logic;
signal \eeprom.n2182\ : std_logic;
signal \eeprom.n3535\ : std_logic;
signal \eeprom.n2114\ : std_logic;
signal \eeprom.n2181\ : std_logic;
signal \eeprom.n3536\ : std_logic;
signal \eeprom.n3537\ : std_logic;
signal \eeprom.n2112\ : std_logic;
signal \eeprom.n2179\ : std_logic;
signal \eeprom.n3538\ : std_logic;
signal \eeprom.n3539\ : std_logic;
signal \eeprom.n2111\ : std_logic;
signal \eeprom.n2178\ : std_logic;
signal \bfn_5_28_0_\ : std_logic;
signal \eeprom.n2110\ : std_logic;
signal \eeprom.n3540\ : std_logic;
signal n26 : std_logic;
signal \bfn_5_29_0_\ : std_logic;
signal n25 : std_logic;
signal n3485 : std_logic;
signal n24 : std_logic;
signal n3486 : std_logic;
signal n23 : std_logic;
signal n3487 : std_logic;
signal n22 : std_logic;
signal n3488 : std_logic;
signal n21 : std_logic;
signal n3489 : std_logic;
signal n20 : std_logic;
signal n3490 : std_logic;
signal n19 : std_logic;
signal n3491 : std_logic;
signal n3492 : std_logic;
signal n18 : std_logic;
signal \bfn_5_30_0_\ : std_logic;
signal n17 : std_logic;
signal n3493 : std_logic;
signal n16 : std_logic;
signal n3494 : std_logic;
signal n15 : std_logic;
signal n3495 : std_logic;
signal n14 : std_logic;
signal n3496 : std_logic;
signal n13 : std_logic;
signal n3497 : std_logic;
signal n12 : std_logic;
signal n3498 : std_logic;
signal n11 : std_logic;
signal n3499 : std_logic;
signal n3500 : std_logic;
signal n10 : std_logic;
signal \bfn_5_31_0_\ : std_logic;
signal n9 : std_logic;
signal n3501 : std_logic;
signal n8 : std_logic;
signal n3502 : std_logic;
signal n7 : std_logic;
signal n3503 : std_logic;
signal n6 : std_logic;
signal n3504 : std_logic;
signal blink_counter_21 : std_logic;
signal n3505 : std_logic;
signal blink_counter_22 : std_logic;
signal n3506 : std_logic;
signal blink_counter_23 : std_logic;
signal n3507 : std_logic;
signal n3508 : std_logic;
signal blink_counter_24 : std_logic;
signal \bfn_5_32_0_\ : std_logic;
signal n3509 : std_logic;
signal blink_counter_25 : std_logic;
signal \bfn_6_18_0_\ : std_logic;
signal \eeprom.n3587\ : std_logic;
signal \eeprom.n3588\ : std_logic;
signal \eeprom.n3589\ : std_logic;
signal \eeprom.n3590\ : std_logic;
signal \eeprom.n3591\ : std_logic;
signal \eeprom.n3592\ : std_logic;
signal \eeprom.n3593\ : std_logic;
signal \eeprom.n3594\ : std_logic;
signal \bfn_6_19_0_\ : std_logic;
signal \eeprom.n3595\ : std_logic;
signal \eeprom.n3596\ : std_logic;
signal \eeprom.n3597\ : std_logic;
signal \eeprom.n3598\ : std_logic;
signal \eeprom.n3599\ : std_logic;
signal \eeprom.n3600\ : std_logic;
signal \eeprom.n21\ : std_logic;
signal \eeprom.delay_counter_12\ : std_logic;
signal \eeprom.n29_adj_460\ : std_logic;
signal \eeprom.n2609\ : std_logic;
signal \eeprom.n2676\ : std_logic;
signal \eeprom.n2678\ : std_logic;
signal \eeprom.n2611_cascade_\ : std_logic;
signal \eeprom.n2519\ : std_logic;
signal \eeprom.n2586\ : std_logic;
signal \bfn_6_21_0_\ : std_logic;
signal \eeprom.n2518\ : std_logic;
signal \eeprom.n2585\ : std_logic;
signal \eeprom.n3574\ : std_logic;
signal \eeprom.n2517\ : std_logic;
signal \eeprom.n2584\ : std_logic;
signal \eeprom.n3575\ : std_logic;
signal \eeprom.n2516\ : std_logic;
signal \eeprom.n2583\ : std_logic;
signal \eeprom.n3576\ : std_logic;
signal \eeprom.n2515\ : std_logic;
signal \eeprom.n2582\ : std_logic;
signal \eeprom.n3577\ : std_logic;
signal \eeprom.n2514\ : std_logic;
signal \eeprom.n2581\ : std_logic;
signal \eeprom.n3578\ : std_logic;
signal \eeprom.n3579\ : std_logic;
signal \eeprom.n2579\ : std_logic;
signal \eeprom.n3580\ : std_logic;
signal \eeprom.n3581\ : std_logic;
signal \bfn_6_22_0_\ : std_logic;
signal \eeprom.n2510\ : std_logic;
signal \eeprom.n2577\ : std_logic;
signal \eeprom.n3582\ : std_logic;
signal \eeprom.n2509\ : std_logic;
signal \eeprom.n2576\ : std_logic;
signal \eeprom.n3583\ : std_logic;
signal \eeprom.n2508\ : std_logic;
signal \eeprom.n2575\ : std_logic;
signal \eeprom.n3584\ : std_logic;
signal \eeprom.n3585\ : std_logic;
signal \eeprom.n2506\ : std_logic;
signal \eeprom.n3586\ : std_logic;
signal \eeprom.n2412\ : std_logic;
signal \eeprom.n2479\ : std_logic;
signal \eeprom.n2511\ : std_logic;
signal \eeprom.n2578\ : std_logic;
signal \eeprom.n2511_cascade_\ : std_logic;
signal \eeprom.n12_adj_351\ : std_logic;
signal \eeprom.delay_counter_21\ : std_logic;
signal \eeprom.n2219_cascade_\ : std_logic;
signal \eeprom.n2318\ : std_logic;
signal \eeprom.n2580\ : std_logic;
signal \eeprom.n2513\ : std_logic;
signal \eeprom.n2539\ : std_logic;
signal \eeprom.n2574\ : std_logic;
signal \eeprom.n2606_cascade_\ : std_logic;
signal \eeprom.n2605\ : std_logic;
signal \eeprom.n2611\ : std_logic;
signal \eeprom.n10_adj_475_cascade_\ : std_logic;
signal \eeprom.n2413\ : std_logic;
signal \eeprom.n2480\ : std_logic;
signal \eeprom.n2512\ : std_logic;
signal \eeprom.n2408\ : std_logic;
signal \eeprom.n2475\ : std_logic;
signal \eeprom.n2440\ : std_logic;
signal \eeprom.n2507\ : std_logic;
signal \eeprom.n4801\ : std_logic;
signal \eeprom.n2017\ : std_logic;
signal \eeprom.n4799_cascade_\ : std_logic;
signal \eeprom.n4872\ : std_logic;
signal \eeprom.n2314\ : std_logic;
signal \eeprom.n2316\ : std_logic;
signal \eeprom.n2186\ : std_logic;
signal \eeprom.n2119\ : std_logic;
signal \eeprom.n2218_cascade_\ : std_logic;
signal \eeprom.n2317\ : std_logic;
signal \eeprom.n4447_cascade_\ : std_logic;
signal \eeprom.n4218\ : std_logic;
signal \eeprom.n2113\ : std_logic;
signal \eeprom.n2143\ : std_logic;
signal \eeprom.n2180\ : std_logic;
signal \eeprom.n2219\ : std_logic;
signal \eeprom.n2286\ : std_logic;
signal \bfn_6_26_0_\ : std_logic;
signal \eeprom.n2218\ : std_logic;
signal \eeprom.n2285\ : std_logic;
signal \eeprom.n3541\ : std_logic;
signal \eeprom.n2217\ : std_logic;
signal \eeprom.n2284\ : std_logic;
signal \eeprom.n3542\ : std_logic;
signal \eeprom.n2216\ : std_logic;
signal \eeprom.n2283\ : std_logic;
signal \eeprom.n3543\ : std_logic;
signal \eeprom.n2215\ : std_logic;
signal \eeprom.n2282\ : std_logic;
signal \eeprom.n3544\ : std_logic;
signal \eeprom.n2214\ : std_logic;
signal \eeprom.n2281\ : std_logic;
signal \eeprom.n3545\ : std_logic;
signal \eeprom.n2213\ : std_logic;
signal \eeprom.n2280\ : std_logic;
signal \eeprom.n3546\ : std_logic;
signal \eeprom.n2212\ : std_logic;
signal \eeprom.n2279\ : std_logic;
signal \eeprom.n3547\ : std_logic;
signal \eeprom.n3548\ : std_logic;
signal \eeprom.n2211\ : std_logic;
signal \eeprom.n2278\ : std_logic;
signal \bfn_6_27_0_\ : std_logic;
signal \eeprom.n2210\ : std_logic;
signal \eeprom.n2277\ : std_logic;
signal \eeprom.n3549\ : std_logic;
signal \eeprom.n2242\ : std_logic;
signal \eeprom.n2209\ : std_logic;
signal \eeprom.n3550\ : std_logic;
signal \eeprom.n2308\ : std_logic;
signal \eeprom.n2612\ : std_logic;
signal \eeprom.n2679\ : std_logic;
signal \eeprom.n2606\ : std_logic;
signal \eeprom.n2673\ : std_logic;
signal \eeprom.n2680\ : std_logic;
signal \eeprom.n2613\ : std_logic;
signal \eeprom.n2614\ : std_logic;
signal \eeprom.n2681\ : std_logic;
signal \eeprom.n2713_cascade_\ : std_logic;
signal \eeprom.n4695_cascade_\ : std_logic;
signal \eeprom.n16_adj_416_cascade_\ : std_logic;
signal \eeprom.n2618\ : std_logic;
signal \eeprom.n2685\ : std_logic;
signal \eeprom.n2674\ : std_logic;
signal \eeprom.n2686\ : std_logic;
signal \eeprom.n2619\ : std_logic;
signal \eeprom.n2718_cascade_\ : std_logic;
signal \eeprom.n4699\ : std_logic;
signal \eeprom.n2675\ : std_logic;
signal \eeprom.n2682\ : std_logic;
signal \eeprom.n2615\ : std_logic;
signal \eeprom.n2608\ : std_logic;
signal \eeprom.n12\ : std_logic;
signal \eeprom.n2607\ : std_logic;
signal \eeprom.n16\ : std_logic;
signal \eeprom.n2683\ : std_logic;
signal \eeprom.n2638_cascade_\ : std_logic;
signal \eeprom.n2616\ : std_logic;
signal \eeprom.n2617\ : std_logic;
signal \eeprom.n2684\ : std_logic;
signal \eeprom.n2815_cascade_\ : std_logic;
signal \eeprom.n28\ : std_logic;
signal \eeprom.n2610\ : std_logic;
signal \eeprom.n2677\ : std_logic;
signal \eeprom.n2638\ : std_logic;
signal \eeprom.n18\ : std_logic;
signal \eeprom.n2709_cascade_\ : std_logic;
signal \eeprom.n13_adj_417\ : std_logic;
signal \eeprom.n2737_cascade_\ : std_logic;
signal \eeprom.n2719\ : std_logic;
signal \eeprom.n2786\ : std_logic;
signal \bfn_7_21_0_\ : std_logic;
signal \eeprom.n2718\ : std_logic;
signal \eeprom.n2785\ : std_logic;
signal \eeprom.n3601\ : std_logic;
signal \eeprom.n3602\ : std_logic;
signal \eeprom.n2716\ : std_logic;
signal \eeprom.n2783\ : std_logic;
signal \eeprom.n3603\ : std_logic;
signal \eeprom.n3604\ : std_logic;
signal \eeprom.n2714\ : std_logic;
signal \eeprom.n2781\ : std_logic;
signal \eeprom.n3605\ : std_logic;
signal \eeprom.n3606\ : std_logic;
signal \eeprom.n3607\ : std_logic;
signal \eeprom.n3608\ : std_logic;
signal \bfn_7_22_0_\ : std_logic;
signal \eeprom.n3609\ : std_logic;
signal \eeprom.n3610\ : std_logic;
signal \eeprom.n3611\ : std_logic;
signal \eeprom.n3612\ : std_logic;
signal \eeprom.n3613\ : std_logic;
signal \eeprom.n3614\ : std_logic;
signal \eeprom.n2704\ : std_logic;
signal \eeprom.n3615\ : std_logic;
signal \eeprom.n2777\ : std_logic;
signal \eeprom.n2710\ : std_logic;
signal \eeprom.n2778\ : std_logic;
signal \eeprom.n2711\ : std_logic;
signal \eeprom.n2717\ : std_logic;
signal \eeprom.n2784\ : std_logic;
signal \eeprom.n2782\ : std_logic;
signal \eeprom.n2715\ : std_logic;
signal \eeprom.n2713\ : std_logic;
signal \eeprom.n2780\ : std_logic;
signal \bfn_9_17_0_\ : std_logic;
signal \eeprom.n3706\ : std_logic;
signal \eeprom.n3707\ : std_logic;
signal \eeprom.n3708\ : std_logic;
signal \eeprom.n3709\ : std_logic;
signal \eeprom.n3710\ : std_logic;
signal \eeprom.n3711\ : std_logic;
signal \eeprom.n3712\ : std_logic;
signal \eeprom.n3713\ : std_logic;
signal \bfn_9_18_0_\ : std_logic;
signal \eeprom.n3714\ : std_logic;
signal \eeprom.n3715\ : std_logic;
signal \eeprom.n3716\ : std_logic;
signal \eeprom.n3717\ : std_logic;
signal \eeprom.n3718\ : std_logic;
signal \eeprom.n3719\ : std_logic;
signal \eeprom.n3720\ : std_logic;
signal \eeprom.n3721\ : std_logic;
signal \bfn_9_19_0_\ : std_logic;
signal \eeprom.n3722\ : std_logic;
signal \eeprom.n3723\ : std_logic;
signal \eeprom.n3724\ : std_logic;
signal \eeprom.n3725\ : std_logic;
signal \eeprom.n3726\ : std_logic;
signal \bfn_9_20_0_\ : std_logic;
signal \eeprom.n3686\ : std_logic;
signal \eeprom.n3687\ : std_logic;
signal \eeprom.n3688\ : std_logic;
signal \eeprom.n3689\ : std_logic;
signal \eeprom.n3281\ : std_logic;
signal \eeprom.n3690\ : std_logic;
signal \eeprom.n3691\ : std_logic;
signal \eeprom.n3692\ : std_logic;
signal \eeprom.n3693\ : std_logic;
signal \bfn_9_21_0_\ : std_logic;
signal \eeprom.n3694\ : std_logic;
signal \eeprom.n3695\ : std_logic;
signal \eeprom.n3696\ : std_logic;
signal \eeprom.n3697\ : std_logic;
signal \eeprom.n3698\ : std_logic;
signal \eeprom.n3699\ : std_logic;
signal \eeprom.n3700\ : std_logic;
signal \eeprom.n3701\ : std_logic;
signal \bfn_9_22_0_\ : std_logic;
signal \eeprom.n3702\ : std_logic;
signal \eeprom.n3703\ : std_logic;
signal \eeprom.n3704\ : std_logic;
signal \eeprom.n3705\ : std_logic;
signal \eeprom.n2706\ : std_logic;
signal \eeprom.n2773\ : std_logic;
signal \eeprom.n2709\ : std_logic;
signal \eeprom.n2776\ : std_logic;
signal \bfn_9_23_0_\ : std_logic;
signal \eeprom.n3616\ : std_logic;
signal \eeprom.n3617\ : std_logic;
signal \eeprom.n3618\ : std_logic;
signal \eeprom.n3619\ : std_logic;
signal \eeprom.n3620\ : std_logic;
signal \eeprom.n3621\ : std_logic;
signal \eeprom.n3622\ : std_logic;
signal \eeprom.n3623\ : std_logic;
signal \bfn_9_24_0_\ : std_logic;
signal \eeprom.n3624\ : std_logic;
signal \eeprom.n3625\ : std_logic;
signal \eeprom.n3626\ : std_logic;
signal \eeprom.n3627\ : std_logic;
signal \eeprom.n3628\ : std_logic;
signal \eeprom.n3629\ : std_logic;
signal \eeprom.n3630\ : std_logic;
signal \eeprom.n3631\ : std_logic;
signal \bfn_9_25_0_\ : std_logic;
signal \eeprom.n2873\ : std_logic;
signal \eeprom.n2872\ : std_logic;
signal \eeprom.n2904_cascade_\ : std_logic;
signal \eeprom.n3286\ : std_logic;
signal \eeprom.n3285\ : std_logic;
signal \eeprom.n3371\ : std_logic;
signal \eeprom.n3282\ : std_logic;
signal \eeprom.n3314_cascade_\ : std_logic;
signal \eeprom.n3272\ : std_logic;
signal \eeprom.n3274\ : std_logic;
signal \eeprom.n3273\ : std_logic;
signal \eeprom.n3280\ : std_logic;
signal \eeprom.n3312\ : std_logic;
signal \eeprom.n3379\ : std_logic;
signal \eeprom.n3312_cascade_\ : std_logic;
signal \eeprom.n3275\ : std_logic;
signal \eeprom.n3307\ : std_logic;
signal \eeprom.n3374\ : std_logic;
signal \eeprom.n3307_cascade_\ : std_logic;
signal \eeprom.n28_adj_482_cascade_\ : std_logic;
signal \eeprom.n3278\ : std_logic;
signal \eeprom.n3232_cascade_\ : std_logic;
signal \eeprom.n3367\ : std_logic;
signal \eeprom.n3276\ : std_logic;
signal \eeprom.n3279\ : std_logic;
signal \eeprom.n3271\ : std_logic;
signal \eeprom.n3277\ : std_logic;
signal \eeprom.n3209\ : std_logic;
signal \eeprom.n3369\ : std_logic;
signal \eeprom.n27\ : std_logic;
signal \eeprom.n3268\ : std_logic;
signal \eeprom.n32_adj_480\ : std_logic;
signal \eeprom.n3269\ : std_logic;
signal \eeprom.n2815\ : std_logic;
signal \eeprom.n2882\ : std_logic;
signal \eeprom.n2886\ : std_logic;
signal \eeprom.n2918_cascade_\ : std_logic;
signal \eeprom.n3267\ : std_logic;
signal \eeprom.n2705\ : std_logic;
signal \eeprom.n2772\ : std_logic;
signal \eeprom.n2803\ : std_logic;
signal \eeprom.n2804_cascade_\ : std_logic;
signal \eeprom.n3270\ : std_logic;
signal \eeprom.n2712\ : std_logic;
signal \eeprom.n2779\ : std_logic;
signal \eeprom.n2707\ : std_logic;
signal \eeprom.n2774\ : std_logic;
signal \eeprom.n2806\ : std_logic;
signal \eeprom.n2806_cascade_\ : std_logic;
signal \eeprom.n2805\ : std_logic;
signal \eeprom.n18_adj_418\ : std_logic;
signal \eeprom.n2708\ : std_logic;
signal \eeprom.n2775\ : std_logic;
signal \eeprom.n2737\ : std_logic;
signal \eeprom.n2807\ : std_logic;
signal \eeprom.n2874\ : std_logic;
signal \eeprom.n2807_cascade_\ : std_logic;
signal \eeprom.n2881\ : std_logic;
signal \eeprom.n2913_cascade_\ : std_logic;
signal \eeprom.n4529\ : std_logic;
signal \eeprom.n2814\ : std_logic;
signal \eeprom.n2819\ : std_logic;
signal \eeprom.n4533_cascade_\ : std_logic;
signal \eeprom.n20\ : std_logic;
signal \eeprom.n15_cascade_\ : std_logic;
signal \eeprom.n2816\ : std_logic;
signal \eeprom.n2836_cascade_\ : std_logic;
signal \eeprom.n2883\ : std_logic;
signal \eeprom.n2809\ : std_logic;
signal \eeprom.n2876\ : std_logic;
signal \eeprom.n2804\ : std_logic;
signal \eeprom.n2871\ : std_logic;
signal \eeprom.n19\ : std_logic;
signal \eeprom.n22_cascade_\ : std_logic;
signal \eeprom.n2885\ : std_logic;
signal \eeprom.n2818\ : std_logic;
signal \eeprom.n4703\ : std_logic;
signal \eeprom.n2917_cascade_\ : std_logic;
signal \eeprom.n4707_cascade_\ : std_logic;
signal \eeprom.n15_adj_419\ : std_logic;
signal \eeprom.n2875\ : std_logic;
signal \eeprom.n2808\ : std_logic;
signal \eeprom.n3385\ : std_logic;
signal \eeprom.n3283\ : std_logic;
signal \eeprom.n3315_cascade_\ : std_logic;
signal \eeprom.n3318\ : std_logic;
signal \eeprom.n4719_cascade_\ : std_logic;
signal \eeprom.n4721\ : std_logic;
signal \eeprom.n3304\ : std_logic;
signal \eeprom.n4151_cascade_\ : std_logic;
signal \eeprom.n3302\ : std_logic;
signal \eeprom.n3317\ : std_logic;
signal \eeprom.n3384\ : std_logic;
signal \eeprom.n3375\ : std_logic;
signal \eeprom.n3308\ : std_logic;
signal \eeprom.n3407_cascade_\ : std_logic;
signal \eeprom.n28_adj_484\ : std_logic;
signal \eeprom.n27_adj_486_cascade_\ : std_logic;
signal \eeprom.n26_adj_485\ : std_logic;
signal \eeprom.n3306\ : std_logic;
signal \eeprom.n3331_cascade_\ : std_logic;
signal \eeprom.n3373\ : std_logic;
signal \eeprom.n3305\ : std_logic;
signal \eeprom.n3372\ : std_logic;
signal \eeprom.n3376\ : std_logic;
signal \eeprom.n3309\ : std_logic;
signal \eeprom.n3219\ : std_logic;
signal \eeprom.n4615_cascade_\ : std_logic;
signal \eeprom.n3218\ : std_logic;
signal \eeprom.n21_adj_477\ : std_logic;
signal \eeprom.n4611\ : std_logic;
signal \eeprom.n3300\ : std_logic;
signal \eeprom.n3298\ : std_logic;
signal \eeprom.n25_adj_487\ : std_logic;
signal \eeprom.n3301\ : std_logic;
signal \eeprom.n3368\ : std_logic;
signal \eeprom.n3284\ : std_logic;
signal \eeprom.n3232\ : std_logic;
signal \eeprom.n3210\ : std_logic;
signal \eeprom.n3113_cascade_\ : std_logic;
signal \eeprom.n3212\ : std_logic;
signal \eeprom.n3208\ : std_logic;
signal \eeprom.n25_adj_478\ : std_logic;
signal \eeprom.n3213\ : std_logic;
signal \eeprom.n3116_cascade_\ : std_logic;
signal \eeprom.n3215\ : std_logic;
signal \bfn_11_21_0_\ : std_logic;
signal \eeprom.n2918\ : std_logic;
signal \eeprom.n2985\ : std_logic;
signal \eeprom.n3632\ : std_logic;
signal \eeprom.n3633\ : std_logic;
signal \eeprom.n3634\ : std_logic;
signal \eeprom.n3635\ : std_logic;
signal \eeprom.n3636\ : std_logic;
signal \eeprom.n3637\ : std_logic;
signal \eeprom.n3638\ : std_logic;
signal \eeprom.n3639\ : std_logic;
signal \bfn_11_22_0_\ : std_logic;
signal \eeprom.n3640\ : std_logic;
signal \eeprom.n3641\ : std_logic;
signal \eeprom.n3642\ : std_logic;
signal \eeprom.n3643\ : std_logic;
signal \eeprom.n3644\ : std_logic;
signal \eeprom.n3645\ : std_logic;
signal \eeprom.n3646\ : std_logic;
signal \eeprom.n3647\ : std_logic;
signal \bfn_11_23_0_\ : std_logic;
signal \eeprom.n2902\ : std_logic;
signal \eeprom.n3648\ : std_logic;
signal \eeprom.n2906\ : std_logic;
signal \eeprom.n2973\ : std_logic;
signal \eeprom.n2903\ : std_logic;
signal \eeprom.n2970\ : std_logic;
signal \eeprom.n2879\ : std_logic;
signal \eeprom.n2812\ : std_logic;
signal \eeprom.n2880\ : std_logic;
signal \eeprom.n2813\ : std_logic;
signal \eeprom.n2913\ : std_logic;
signal \eeprom.n2980\ : std_logic;
signal \eeprom.n2817\ : std_logic;
signal \eeprom.n2884\ : std_logic;
signal \eeprom.n2877\ : std_logic;
signal \eeprom.n2810\ : std_logic;
signal \eeprom.n2909_cascade_\ : std_logic;
signal \eeprom.n18_adj_420\ : std_logic;
signal \eeprom.n2975\ : std_logic;
signal \eeprom.n2908\ : std_logic;
signal \eeprom.n2878\ : std_logic;
signal \eeprom.n2811\ : std_logic;
signal \eeprom.n2836\ : std_logic;
signal \eeprom.n2915\ : std_logic;
signal \eeprom.n2982\ : std_logic;
signal \eeprom.n2911\ : std_logic;
signal \eeprom.n2978\ : std_logic;
signal \eeprom.n2984\ : std_logic;
signal \eeprom.n2917\ : std_logic;
signal \eeprom.n3315\ : std_logic;
signal \eeprom.n3382\ : std_logic;
signal \eeprom.n3414_cascade_\ : std_logic;
signal \eeprom.n4689_cascade_\ : std_logic;
signal \eeprom.n4144_cascade_\ : std_logic;
signal \eeprom.n3386\ : std_logic;
signal \eeprom.n3319\ : std_logic;
signal \eeprom.n3316\ : std_logic;
signal \eeprom.n3383\ : std_logic;
signal \eeprom.n3314\ : std_logic;
signal \eeprom.n3381\ : std_logic;
signal \eeprom.n3413_cascade_\ : std_logic;
signal \eeprom.n4687\ : std_logic;
signal \eeprom.n3378\ : std_logic;
signal \eeprom.n3311\ : std_logic;
signal \eeprom.n3410_cascade_\ : std_logic;
signal \eeprom.n3505_cascade_\ : std_logic;
signal \eeprom.n3310\ : std_logic;
signal \eeprom.n3377\ : std_logic;
signal \eeprom.n3608_adj_451_cascade_\ : std_logic;
signal \eeprom.n3313\ : std_logic;
signal \eeprom.n3380\ : std_logic;
signal \eeprom.n3412_cascade_\ : std_logic;
signal \eeprom.n3303\ : std_logic;
signal \eeprom.n3370\ : std_logic;
signal \eeprom.n3366\ : std_logic;
signal \eeprom.n3299\ : std_logic;
signal \eeprom.n3331\ : std_logic;
signal \eeprom.n3500_cascade_\ : std_logic;
signal \eeprom.n3216\ : std_logic;
signal \eeprom.n3203\ : std_logic;
signal \eeprom.n3217\ : std_logic;
signal \eeprom.n18_adj_432_cascade_\ : std_logic;
signal \eeprom.n26_adj_466_cascade_\ : std_logic;
signal \eeprom.n4711_cascade_\ : std_logic;
signal \eeprom.n4715\ : std_logic;
signal \eeprom.n3206\ : std_logic;
signal \eeprom.n3214\ : std_logic;
signal \eeprom.n3119\ : std_logic;
signal \eeprom.n3186\ : std_logic;
signal \bfn_12_22_0_\ : std_logic;
signal \eeprom.n3185\ : std_logic;
signal \eeprom.n3667\ : std_logic;
signal \eeprom.n3184\ : std_logic;
signal \eeprom.n3668\ : std_logic;
signal \eeprom.n3116\ : std_logic;
signal \eeprom.n3183\ : std_logic;
signal \eeprom.n3669\ : std_logic;
signal \eeprom.n3182\ : std_logic;
signal \eeprom.n3670\ : std_logic;
signal \eeprom.n3181\ : std_logic;
signal \eeprom.n3671\ : std_logic;
signal \eeprom.n3113\ : std_logic;
signal \eeprom.n3180\ : std_logic;
signal \eeprom.n3672\ : std_logic;
signal \eeprom.n3673\ : std_logic;
signal \eeprom.n3674\ : std_logic;
signal \eeprom.n3178\ : std_logic;
signal \bfn_12_23_0_\ : std_logic;
signal \eeprom.n3177\ : std_logic;
signal \eeprom.n3675\ : std_logic;
signal \eeprom.n3176\ : std_logic;
signal \eeprom.n3676\ : std_logic;
signal \eeprom.n3677\ : std_logic;
signal \eeprom.n3174\ : std_logic;
signal \eeprom.n3678\ : std_logic;
signal \eeprom.n3679\ : std_logic;
signal \eeprom.n3680\ : std_logic;
signal \eeprom.n3171\ : std_logic;
signal \eeprom.n3681\ : std_logic;
signal \eeprom.n3682\ : std_logic;
signal \bfn_12_24_0_\ : std_logic;
signal \eeprom.n3683\ : std_logic;
signal \eeprom.n3684\ : std_logic;
signal \eeprom.n3685\ : std_logic;
signal \eeprom.n2971\ : std_logic;
signal \eeprom.n2904\ : std_logic;
signal \eeprom.n2977\ : std_logic;
signal \eeprom.n2910\ : std_logic;
signal \eeprom.n3497_cascade_\ : std_logic;
signal \eeprom.n28_adj_493_cascade_\ : std_logic;
signal \eeprom.n18_adj_488_cascade_\ : std_logic;
signal \eeprom.n29_adj_491\ : std_logic;
signal \eeprom.n28_adj_490\ : std_logic;
signal \eeprom.n30_adj_489_cascade_\ : std_logic;
signal \eeprom.n27_adj_492\ : std_logic;
signal \eeprom.n3430_cascade_\ : std_logic;
signal \eeprom.n3609_adj_445\ : std_logic;
signal \eeprom.n3508_cascade_\ : std_logic;
signal \eeprom.n31_adj_496\ : std_logic;
signal \eeprom.n29_adj_497\ : std_logic;
signal \eeprom.n30_adj_495_cascade_\ : std_logic;
signal \eeprom.n32_adj_494\ : std_logic;
signal \eeprom.n3606_adj_446_cascade_\ : std_logic;
signal \eeprom.n4451_cascade_\ : std_logic;
signal \eeprom.n4453\ : std_logic;
signal \eeprom.n3599_adj_450_cascade_\ : std_logic;
signal \eeprom.n4429\ : std_logic;
signal \eeprom.n29\ : std_logic;
signal \eeprom.n3600_adj_449\ : std_logic;
signal \eeprom.n4581\ : std_logic;
signal \eeprom.n3117\ : std_logic;
signal \eeprom.n3108\ : std_logic;
signal \eeprom.n3175\ : std_logic;
signal \eeprom.n3108_cascade_\ : std_logic;
signal \eeprom.n3105\ : std_logic;
signal \eeprom.n3172\ : std_logic;
signal \eeprom.n3105_cascade_\ : std_logic;
signal \eeprom.n3204\ : std_logic;
signal \eeprom.n3179\ : std_logic;
signal \eeprom.n3211\ : std_logic;
signal \eeprom.n3115\ : std_logic;
signal \eeprom.n3169\ : std_logic;
signal \eeprom.n3201\ : std_logic;
signal \eeprom.n3207\ : std_logic;
signal \eeprom.n3201_cascade_\ : std_logic;
signal \eeprom.n24_adj_481\ : std_logic;
signal \eeprom.n3114\ : std_logic;
signal \eeprom.n2905\ : std_logic;
signal \eeprom.n2972\ : std_logic;
signal \eeprom.n3118\ : std_logic;
signal \eeprom.n3102\ : std_logic;
signal \eeprom.n3102_cascade_\ : std_logic;
signal \eeprom.n22_adj_465\ : std_logic;
signal \eeprom.n3104\ : std_logic;
signal \eeprom.n3170\ : std_logic;
signal \eeprom.n3202\ : std_logic;
signal \eeprom.n3168\ : std_logic;
signal \eeprom.n3200\ : std_logic;
signal \eeprom.n2983\ : std_logic;
signal \eeprom.n2916\ : std_logic;
signal \eeprom.n3106\ : std_logic;
signal \eeprom.n3173\ : std_logic;
signal \eeprom.n3106_cascade_\ : std_logic;
signal \eeprom.n3133\ : std_logic;
signal \eeprom.n3205\ : std_logic;
signal \eeprom.n3205_cascade_\ : std_logic;
signal \eeprom.n3199\ : std_logic;
signal \eeprom.n16_adj_479\ : std_logic;
signal \eeprom.n2907\ : std_logic;
signal \eeprom.n2974\ : std_logic;
signal \eeprom.n2914\ : std_logic;
signal \eeprom.n2981\ : std_logic;
signal \eeprom.n3101\ : std_logic;
signal \bfn_14_17_0_\ : std_logic;
signal \eeprom.n3727\ : std_logic;
signal \eeprom.n3728\ : std_logic;
signal \eeprom.n3729\ : std_logic;
signal \eeprom.n3415\ : std_logic;
signal \eeprom.n3482_adj_401\ : std_logic;
signal \eeprom.n3730\ : std_logic;
signal \eeprom.n3414\ : std_logic;
signal \eeprom.n3481_adj_399\ : std_logic;
signal \eeprom.n3731\ : std_logic;
signal \eeprom.n3413\ : std_logic;
signal \eeprom.n3480_adj_398\ : std_logic;
signal \eeprom.n3732\ : std_logic;
signal \eeprom.n3412\ : std_logic;
signal \eeprom.n3479_adj_394\ : std_logic;
signal \eeprom.n3733\ : std_logic;
signal \eeprom.n3734\ : std_logic;
signal \eeprom.n3411\ : std_logic;
signal \eeprom.n3478_adj_393\ : std_logic;
signal \bfn_14_18_0_\ : std_logic;
signal \eeprom.n3410\ : std_logic;
signal \eeprom.n3477_adj_392\ : std_logic;
signal \eeprom.n3735\ : std_logic;
signal \eeprom.n3409\ : std_logic;
signal \eeprom.n3476_adj_391\ : std_logic;
signal \eeprom.n3736\ : std_logic;
signal \eeprom.n3408\ : std_logic;
signal \eeprom.n3475_adj_390\ : std_logic;
signal \eeprom.n3737\ : std_logic;
signal \eeprom.n3407\ : std_logic;
signal \eeprom.n3474_adj_389\ : std_logic;
signal \eeprom.n3738\ : std_logic;
signal \eeprom.n3406\ : std_logic;
signal \eeprom.n3473_adj_388\ : std_logic;
signal \eeprom.n3739\ : std_logic;
signal \eeprom.n3405\ : std_logic;
signal \eeprom.n3472_adj_387\ : std_logic;
signal \eeprom.n3740\ : std_logic;
signal \eeprom.n3741\ : std_logic;
signal \eeprom.n3742\ : std_logic;
signal \eeprom.n3403\ : std_logic;
signal \eeprom.n3470_adj_385\ : std_logic;
signal \bfn_14_19_0_\ : std_logic;
signal \eeprom.n3402\ : std_logic;
signal \eeprom.n3469_adj_384\ : std_logic;
signal \eeprom.n3743\ : std_logic;
signal \eeprom.n3401\ : std_logic;
signal \eeprom.n3468_adj_383\ : std_logic;
signal \eeprom.n3744\ : std_logic;
signal \eeprom.n3400\ : std_logic;
signal \eeprom.n3467_adj_382\ : std_logic;
signal \eeprom.n3745\ : std_logic;
signal \eeprom.n3399\ : std_logic;
signal \eeprom.n3466_adj_381\ : std_logic;
signal \eeprom.n3746\ : std_logic;
signal \eeprom.n3398\ : std_logic;
signal \eeprom.n3465_adj_380\ : std_logic;
signal \eeprom.n3747\ : std_logic;
signal \eeprom.n3397\ : std_logic;
signal \eeprom.n3748\ : std_logic;
signal \eeprom.n4583\ : std_logic;
signal \eeprom.n31_cascade_\ : std_logic;
signal \eeprom.n4433\ : std_logic;
signal \eeprom.n3598_adj_452\ : std_logic;
signal \eeprom.n31_adj_476\ : std_logic;
signal \eeprom.delay_counter_31\ : std_logic;
signal \eeprom.n24_adj_459\ : std_logic;
signal \eeprom.n4559_cascade_\ : std_logic;
signal \eeprom.n4563_cascade_\ : std_logic;
signal \eeprom.n21_adj_422\ : std_logic;
signal \eeprom.n17_adj_421_cascade_\ : std_logic;
signal \eeprom.n24_cascade_\ : std_logic;
signal \eeprom.n20_adj_423\ : std_logic;
signal \eeprom.n3034_cascade_\ : std_logic;
signal \eeprom.n3112\ : std_logic;
signal \eeprom.n2912\ : std_logic;
signal \eeprom.n2979\ : std_logic;
signal \eeprom.n3103\ : std_logic;
signal \eeprom.n4137\ : std_logic;
signal \eeprom.n3417\ : std_logic;
signal \eeprom.n3484_adj_406\ : std_logic;
signal \eeprom.n3418\ : std_logic;
signal \eeprom.n3485\ : std_logic;
signal \eeprom.n3517_adj_374_cascade_\ : std_logic;
signal \eeprom.n4729\ : std_logic;
signal \eeprom.n3416\ : std_logic;
signal \eeprom.n3483_adj_404\ : std_logic;
signal \eeprom.n3515_adj_370_cascade_\ : std_logic;
signal \eeprom.n4727\ : std_logic;
signal \eeprom.n3419\ : std_logic;
signal \eeprom.n3486\ : std_logic;
signal \eeprom.n3471_adj_386\ : std_logic;
signal \eeprom.n3430\ : std_logic;
signal \eeprom.n3404\ : std_logic;
signal \eeprom.n3615_adj_344_cascade_\ : std_logic;
signal \eeprom.n3714_adj_442_cascade_\ : std_logic;
signal \eeprom.n3617_adj_346_cascade_\ : std_logic;
signal \eeprom.n4619\ : std_logic;
signal \eeprom.n4427_cascade_\ : std_logic;
signal \eeprom.n3596_adj_454\ : std_logic;
signal \eeprom.n28_adj_455_cascade_\ : std_logic;
signal \eeprom.n4567\ : std_logic;
signal \eeprom.n3628_adj_437_cascade_\ : std_logic;
signal \eeprom.n3716_adj_439_cascade_\ : std_logic;
signal \eeprom.n3605_adj_453\ : std_logic;
signal \eeprom.n3618_adj_350_cascade_\ : std_logic;
signal \eeprom.n4623\ : std_logic;
signal \eeprom.n4425\ : std_logic;
signal \eeprom.delay_counter_0\ : std_logic;
signal \eeprom.n1166\ : std_logic;
signal \bfn_15_20_0_\ : std_logic;
signal \eeprom.delay_counter_1\ : std_logic;
signal \eeprom.n3724_adj_335\ : std_logic;
signal \eeprom.n3772\ : std_logic;
signal \eeprom.delay_counter_2\ : std_logic;
signal \eeprom.n3723_adj_334\ : std_logic;
signal \eeprom.n3773\ : std_logic;
signal \eeprom.delay_counter_3\ : std_logic;
signal \eeprom.n3722_adj_433\ : std_logic;
signal \eeprom.n3774\ : std_logic;
signal \eeprom.delay_counter_4\ : std_logic;
signal \eeprom.n3721_adj_434\ : std_logic;
signal \eeprom.n3775\ : std_logic;
signal \eeprom.delay_counter_5\ : std_logic;
signal \eeprom.n3720_adj_435\ : std_logic;
signal \eeprom.n3776\ : std_logic;
signal \eeprom.delay_counter_6\ : std_logic;
signal \eeprom.n3719_adj_436\ : std_logic;
signal \eeprom.n3777\ : std_logic;
signal \eeprom.n3778\ : std_logic;
signal \eeprom.n3779\ : std_logic;
signal \bfn_15_21_0_\ : std_logic;
signal \eeprom.n4909\ : std_logic;
signal \eeprom.n3716_adj_439\ : std_logic;
signal \eeprom.n3780\ : std_logic;
signal \eeprom.n3781\ : std_logic;
signal \eeprom.n4915\ : std_logic;
signal \eeprom.n3714_adj_442\ : std_logic;
signal \eeprom.n3782\ : std_logic;
signal \eeprom.n3783\ : std_logic;
signal \eeprom.n4921\ : std_logic;
signal \eeprom.n3712_adj_444\ : std_logic;
signal \eeprom.n3784\ : std_logic;
signal \eeprom.n2\ : std_logic;
signal \eeprom.n4924\ : std_logic;
signal \eeprom.n3785\ : std_logic;
signal \eeprom.n3713_adj_443\ : std_logic;
signal \eeprom.n4918\ : std_logic;
signal \eeprom.number_of_bytes_7_N_68_5\ : std_logic;
signal \eeprom.number_of_bytes_7_N_68_4\ : std_logic;
signal \eeprom.number_of_bytes_7_N_68_3\ : std_logic;
signal \eeprom.number_of_bytes_7_N_68_6\ : std_logic;
signal \eeprom.number_of_bytes_7_N_68_8\ : std_logic;
signal \eeprom.n4301_cascade_\ : std_logic;
signal \eeprom.number_of_bytes_7_N_68_7\ : std_logic;
signal \eeprom.number_of_bytes_7_N_68_9\ : std_logic;
signal \eeprom.number_of_bytes_7_N_68_10\ : std_logic;
signal \eeprom.n4307_cascade_\ : std_logic;
signal \eeprom.number_of_bytes_7_N_68_11\ : std_logic;
signal \eeprom.number_of_bytes_7_N_68_12\ : std_logic;
signal \eeprom.number_of_bytes_7_N_68_13\ : std_logic;
signal \eeprom.n4313_cascade_\ : std_logic;
signal \eeprom.number_of_bytes_7_N_68_14\ : std_logic;
signal sda_enable : std_logic;
signal \CLK_N\ : std_logic;
signal \eeprom.number_of_bytes_7_N_68_2\ : std_logic;
signal \eeprom.number_of_bytes_7_N_68_0\ : std_logic;
signal \eeprom.number_of_bytes_7_N_68_1\ : std_logic;
signal \eeprom.n4295\ : std_logic;
signal \eeprom.n3111\ : std_logic;
signal \eeprom.n3109\ : std_logic;
signal \eeprom.n3110\ : std_logic;
signal \eeprom.n3107\ : std_logic;
signal \eeprom.n2986\ : std_logic;
signal \eeprom.n2919\ : std_logic;
signal \eeprom.n2909\ : std_logic;
signal \eeprom.n2976\ : std_logic;
signal \eeprom.n2935\ : std_logic;
signal \eeprom.n3519_adj_379\ : std_logic;
signal \eeprom.n3586_adj_378\ : std_logic;
signal \bfn_16_17_0_\ : std_logic;
signal \eeprom.n3518_adj_376\ : std_logic;
signal \eeprom.n3585_adj_375\ : std_logic;
signal \eeprom.n3749\ : std_logic;
signal \eeprom.n3517_adj_374\ : std_logic;
signal \eeprom.n3584_adj_373\ : std_logic;
signal \eeprom.n3750\ : std_logic;
signal \eeprom.n3516_adj_372\ : std_logic;
signal \eeprom.n3583_adj_371\ : std_logic;
signal \eeprom.n3751\ : std_logic;
signal \eeprom.n3515_adj_370\ : std_logic;
signal \eeprom.n3582_adj_369\ : std_logic;
signal \eeprom.n3752\ : std_logic;
signal \eeprom.n3514_adj_368\ : std_logic;
signal \eeprom.n3581_adj_367\ : std_logic;
signal \eeprom.n3753\ : std_logic;
signal \eeprom.n3513_adj_366\ : std_logic;
signal \eeprom.n3580_adj_365\ : std_logic;
signal \eeprom.n3754\ : std_logic;
signal \eeprom.n3512_adj_364\ : std_logic;
signal \eeprom.n3579_adj_363\ : std_logic;
signal \eeprom.n3755\ : std_logic;
signal \eeprom.n3756\ : std_logic;
signal \eeprom.n3511_adj_362\ : std_logic;
signal \eeprom.n3578_adj_361\ : std_logic;
signal \bfn_16_18_0_\ : std_logic;
signal \eeprom.n3510_adj_360\ : std_logic;
signal \eeprom.n3577_adj_359\ : std_logic;
signal \eeprom.n3757\ : std_logic;
signal \eeprom.n3509\ : std_logic;
signal \eeprom.n3576_adj_358\ : std_logic;
signal \eeprom.n3758\ : std_logic;
signal \eeprom.n3508\ : std_logic;
signal \eeprom.n3575_adj_357\ : std_logic;
signal \eeprom.n3759\ : std_logic;
signal \eeprom.n3507\ : std_logic;
signal \eeprom.n3574_adj_356\ : std_logic;
signal \eeprom.n3760\ : std_logic;
signal \eeprom.n3506\ : std_logic;
signal \eeprom.n3573_adj_355\ : std_logic;
signal \eeprom.n3761\ : std_logic;
signal \eeprom.n3505\ : std_logic;
signal \eeprom.n3572_adj_354\ : std_logic;
signal \eeprom.n3762\ : std_logic;
signal \eeprom.n3504\ : std_logic;
signal \eeprom.n3571_adj_353\ : std_logic;
signal \eeprom.n3763\ : std_logic;
signal \eeprom.n3764\ : std_logic;
signal \eeprom.n3503\ : std_logic;
signal \eeprom.n3570_adj_349\ : std_logic;
signal \bfn_16_19_0_\ : std_logic;
signal \eeprom.n3502\ : std_logic;
signal \eeprom.n3569_adj_348\ : std_logic;
signal \eeprom.n3765\ : std_logic;
signal \eeprom.n3501\ : std_logic;
signal \eeprom.n3568_adj_347\ : std_logic;
signal \eeprom.n3766\ : std_logic;
signal \eeprom.n3500\ : std_logic;
signal \eeprom.n3567_adj_341\ : std_logic;
signal \eeprom.n3767\ : std_logic;
signal \eeprom.n3499\ : std_logic;
signal \eeprom.n3566_adj_340\ : std_logic;
signal \eeprom.n3768\ : std_logic;
signal \eeprom.n3498\ : std_logic;
signal \eeprom.n3565_adj_338\ : std_logic;
signal \eeprom.n3769\ : std_logic;
signal \eeprom.n3497\ : std_logic;
signal \eeprom.n3564_adj_337\ : std_logic;
signal \eeprom.n3770\ : std_logic;
signal \eeprom.n3496\ : std_logic;
signal \eeprom.n3529_adj_336\ : std_logic;
signal \eeprom.n3771\ : std_logic;
signal \eeprom.n4765\ : std_logic;
signal \bfn_16_20_0_\ : std_logic;
signal \eeprom.n3510\ : std_logic;
signal \eeprom.n3617_adj_346\ : std_logic;
signal \eeprom.n1351\ : std_logic;
signal \eeprom.n3511\ : std_logic;
signal \eeprom.n3512\ : std_logic;
signal \eeprom.n3615_adj_344\ : std_logic;
signal \eeprom.n1349\ : std_logic;
signal \eeprom.n3513\ : std_logic;
signal \eeprom.n3614_adj_343\ : std_logic;
signal \eeprom.n1348\ : std_logic;
signal \eeprom.n3514\ : std_logic;
signal \eeprom.n3613_adj_342\ : std_logic;
signal \eeprom.n1347\ : std_logic;
signal \eeprom.n3515\ : std_logic;
signal \eeprom.n3612_adj_339\ : std_logic;
signal \eeprom.n3516\ : std_logic;
signal \eeprom.n1350\ : std_logic;
signal \eeprom.n3616_adj_345\ : std_logic;
signal \eeprom.n3715_adj_441\ : std_logic;
signal \eeprom.n3715_adj_441_cascade_\ : std_logic;
signal \eeprom.n4912\ : std_logic;
signal \eeprom.n1346\ : std_logic;
signal \eeprom.n3711_adj_456\ : std_logic;
signal \eeprom.n1352\ : std_logic;
signal \eeprom.n3618_adj_350\ : std_logic;
signal \eeprom.n3717_adj_438\ : std_logic;
signal \eeprom.n3717_adj_438_cascade_\ : std_logic;
signal \eeprom.n4906\ : std_logic;
signal \eeprom.n1353\ : std_logic;
signal \eeprom.n3619_adj_352\ : std_logic;
signal \eeprom.n3628_adj_437\ : std_logic;
signal \eeprom.n4766\ : std_logic;
signal \eeprom.n4766_cascade_\ : std_logic;
signal \eeprom.n4903\ : std_logic;
signal \eeprom.n3019\ : std_logic;
signal \eeprom.n3086\ : std_logic;
signal \bfn_16_23_0_\ : std_logic;
signal \eeprom.n3018\ : std_logic;
signal \eeprom.n3085\ : std_logic;
signal \eeprom.n3649\ : std_logic;
signal \eeprom.n3017\ : std_logic;
signal \eeprom.n3084\ : std_logic;
signal \eeprom.n3650\ : std_logic;
signal \eeprom.n3016\ : std_logic;
signal \eeprom.n3083\ : std_logic;
signal \eeprom.n3651\ : std_logic;
signal \eeprom.n3015\ : std_logic;
signal \eeprom.n3082\ : std_logic;
signal \eeprom.n3652\ : std_logic;
signal \eeprom.n3014\ : std_logic;
signal \eeprom.n3081\ : std_logic;
signal \eeprom.n3653\ : std_logic;
signal \eeprom.n3013\ : std_logic;
signal \eeprom.n3080\ : std_logic;
signal \eeprom.n3654\ : std_logic;
signal \eeprom.n3012\ : std_logic;
signal \eeprom.n3079\ : std_logic;
signal \eeprom.n3655\ : std_logic;
signal \eeprom.n3656\ : std_logic;
signal \eeprom.n3011\ : std_logic;
signal \eeprom.n3078\ : std_logic;
signal \bfn_16_24_0_\ : std_logic;
signal \eeprom.n3010\ : std_logic;
signal \eeprom.n3077\ : std_logic;
signal \eeprom.n3657\ : std_logic;
signal \eeprom.n3009\ : std_logic;
signal \eeprom.n3076\ : std_logic;
signal \eeprom.n3658\ : std_logic;
signal \eeprom.n3008\ : std_logic;
signal \eeprom.n3075\ : std_logic;
signal \eeprom.n3659\ : std_logic;
signal \eeprom.n3007\ : std_logic;
signal \eeprom.n3074\ : std_logic;
signal \eeprom.n3660\ : std_logic;
signal \eeprom.n3006\ : std_logic;
signal \eeprom.n3073\ : std_logic;
signal \eeprom.n3661\ : std_logic;
signal \eeprom.n3005\ : std_logic;
signal \eeprom.n3072\ : std_logic;
signal \eeprom.n3662\ : std_logic;
signal \eeprom.n3004\ : std_logic;
signal \eeprom.n3071\ : std_logic;
signal \eeprom.n3663\ : std_logic;
signal \eeprom.n3664\ : std_logic;
signal \eeprom.n3003\ : std_logic;
signal \eeprom.n3070\ : std_logic;
signal \bfn_16_25_0_\ : std_logic;
signal \eeprom.n3002\ : std_logic;
signal \eeprom.n3069\ : std_logic;
signal \eeprom.n3665\ : std_logic;
signal \eeprom.n3001\ : std_logic;
signal \eeprom.n3034\ : std_logic;
signal \eeprom.n3666\ : std_logic;
signal \eeprom.n3100\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \_gnd_net_\ : std_logic;

signal \CS_CLK_wire\ : std_logic;
signal \CS_wire\ : std_logic;
signal \DE_wire\ : std_logic;
signal \INHA_wire\ : std_logic;
signal \INHB_wire\ : std_logic;
signal \INHC_wire\ : std_logic;
signal \INLA_wire\ : std_logic;
signal \INLB_wire\ : std_logic;
signal \INLC_wire\ : std_logic;
signal \LED_wire\ : std_logic;
signal \NEOPXL_wire\ : std_logic;
signal \TX_wire\ : std_logic;
signal \USBPU_wire\ : std_logic;
signal \CLK_wire\ : std_logic;

begin
    CS_CLK <= \CS_CLK_wire\;
    CS <= \CS_wire\;
    DE <= \DE_wire\;
    INHA <= \INHA_wire\;
    INHB <= \INHB_wire\;
    INHC <= \INHC_wire\;
    INLA <= \INLA_wire\;
    INLB <= \INLB_wire\;
    INLC <= \INLC_wire\;
    LED <= \LED_wire\;
    NEOPXL <= \NEOPXL_wire\;
    TX <= \TX_wire\;
    USBPU <= \USBPU_wire\;
    \CLK_wire\ <= CLK;

    \CS_CLK_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__28245\,
            DIN => \N__28244\,
            DOUT => \N__28243\,
            PACKAGEPIN => \CS_CLK_wire\
        );

    \CS_CLK_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__28245\,
            PADOUT => \N__28244\,
            PADIN => \N__28243\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \CS_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__28236\,
            DIN => \N__28235\,
            DOUT => \N__28234\,
            PACKAGEPIN => \CS_wire\
        );

    \CS_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__28236\,
            PADOUT => \N__28235\,
            PADIN => \N__28234\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \DE_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__28227\,
            DIN => \N__28226\,
            DOUT => \N__28225\,
            PACKAGEPIN => \DE_wire\
        );

    \DE_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__28227\,
            PADOUT => \N__28226\,
            PADIN => \N__28225\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \INHA_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__28218\,
            DIN => \N__28217\,
            DOUT => \N__28216\,
            PACKAGEPIN => \INHA_wire\
        );

    \INHA_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__28218\,
            PADOUT => \N__28217\,
            PADIN => \N__28216\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \INHB_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__28209\,
            DIN => \N__28208\,
            DOUT => \N__28207\,
            PACKAGEPIN => \INHB_wire\
        );

    \INHB_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__28209\,
            PADOUT => \N__28208\,
            PADIN => \N__28207\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \INHC_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__28200\,
            DIN => \N__28199\,
            DOUT => \N__28198\,
            PACKAGEPIN => \INHC_wire\
        );

    \INHC_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__28200\,
            PADOUT => \N__28199\,
            PADIN => \N__28198\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \INLA_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__28191\,
            DIN => \N__28190\,
            DOUT => \N__28189\,
            PACKAGEPIN => \INLA_wire\
        );

    \INLA_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__28191\,
            PADOUT => \N__28190\,
            PADIN => \N__28189\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \INLB_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__28182\,
            DIN => \N__28181\,
            DOUT => \N__28180\,
            PACKAGEPIN => \INLB_wire\
        );

    \INLB_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__28182\,
            PADOUT => \N__28181\,
            PADIN => \N__28180\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \INLC_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__28173\,
            DIN => \N__28172\,
            DOUT => \N__28171\,
            PACKAGEPIN => \INLC_wire\
        );

    \INLC_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__28173\,
            PADOUT => \N__28172\,
            PADIN => \N__28171\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \LED_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__28164\,
            DIN => \N__28163\,
            DOUT => \N__28162\,
            PACKAGEPIN => \LED_wire\
        );

    \LED_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__28164\,
            PADOUT => \N__28163\,
            PADIN => \N__28162\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__13496\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \NEOPXL_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__28155\,
            DIN => \N__28154\,
            DOUT => \N__28153\,
            PACKAGEPIN => \NEOPXL_wire\
        );

    \NEOPXL_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__28155\,
            PADOUT => \N__28154\,
            PADIN => \N__28153\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \TX_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__28146\,
            DIN => \N__28145\,
            DOUT => \N__28144\,
            PACKAGEPIN => \TX_wire\
        );

    \TX_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__28146\,
            PADOUT => \N__28145\,
            PADIN => \N__28144\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \USBPU_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__28137\,
            DIN => \N__28136\,
            DOUT => \N__28135\,
            PACKAGEPIN => \USBPU_wire\
        );

    \USBPU_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__28137\,
            PADOUT => \N__28136\,
            PADIN => \N__28135\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \scl_output_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__28128\,
            DIN => \N__28127\,
            DOUT => \N__28126\,
            PACKAGEPIN => SCL
        );

    \scl_output_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__28128\,
            PADOUT => \N__28127\,
            PADIN => \N__28126\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \sda_output_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__28119\,
            DIN => \N__28118\,
            DOUT => \N__28117\,
            PACKAGEPIN => SDA
        );

    \sda_output_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__28119\,
            PADOUT => \N__28118\,
            PADIN => \N__28117\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__24374\
        );

    \CLK_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__28110\,
            DIN => \N__28109\,
            DOUT => \N__28108\,
            PACKAGEPIN => \CLK_wire\
        );

    \CLK_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__28110\,
            PADOUT => \N__28109\,
            PADIN => \N__28108\,
            CLOCKENABLE => 'H',
            DIN0 => \CLK_pad_gb_input\,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \I__6599\ : CascadeMux
    port map (
            O => \N__28091\,
            I => \N__28088\
        );

    \I__6598\ : InMux
    port map (
            O => \N__28088\,
            I => \N__28085\
        );

    \I__6597\ : LocalMux
    port map (
            O => \N__28085\,
            I => \N__28082\
        );

    \I__6596\ : Span4Mux_h
    port map (
            O => \N__28082\,
            I => \N__28079\
        );

    \I__6595\ : Odrv4
    port map (
            O => \N__28079\,
            I => \eeprom.n3072\
        );

    \I__6594\ : InMux
    port map (
            O => \N__28076\,
            I => \eeprom.n3662\
        );

    \I__6593\ : InMux
    port map (
            O => \N__28073\,
            I => \N__28069\
        );

    \I__6592\ : InMux
    port map (
            O => \N__28072\,
            I => \N__28066\
        );

    \I__6591\ : LocalMux
    port map (
            O => \N__28069\,
            I => \N__28063\
        );

    \I__6590\ : LocalMux
    port map (
            O => \N__28066\,
            I => \N__28057\
        );

    \I__6589\ : Span4Mux_h
    port map (
            O => \N__28063\,
            I => \N__28057\
        );

    \I__6588\ : InMux
    port map (
            O => \N__28062\,
            I => \N__28054\
        );

    \I__6587\ : Odrv4
    port map (
            O => \N__28057\,
            I => \eeprom.n3004\
        );

    \I__6586\ : LocalMux
    port map (
            O => \N__28054\,
            I => \eeprom.n3004\
        );

    \I__6585\ : CascadeMux
    port map (
            O => \N__28049\,
            I => \N__28046\
        );

    \I__6584\ : InMux
    port map (
            O => \N__28046\,
            I => \N__28043\
        );

    \I__6583\ : LocalMux
    port map (
            O => \N__28043\,
            I => \N__28040\
        );

    \I__6582\ : Odrv4
    port map (
            O => \N__28040\,
            I => \eeprom.n3071\
        );

    \I__6581\ : InMux
    port map (
            O => \N__28037\,
            I => \eeprom.n3663\
        );

    \I__6580\ : InMux
    port map (
            O => \N__28034\,
            I => \N__28031\
        );

    \I__6579\ : LocalMux
    port map (
            O => \N__28031\,
            I => \N__28027\
        );

    \I__6578\ : CascadeMux
    port map (
            O => \N__28030\,
            I => \N__28023\
        );

    \I__6577\ : Span4Mux_v
    port map (
            O => \N__28027\,
            I => \N__28020\
        );

    \I__6576\ : InMux
    port map (
            O => \N__28026\,
            I => \N__28015\
        );

    \I__6575\ : InMux
    port map (
            O => \N__28023\,
            I => \N__28015\
        );

    \I__6574\ : Odrv4
    port map (
            O => \N__28020\,
            I => \eeprom.n3003\
        );

    \I__6573\ : LocalMux
    port map (
            O => \N__28015\,
            I => \eeprom.n3003\
        );

    \I__6572\ : InMux
    port map (
            O => \N__28010\,
            I => \N__28007\
        );

    \I__6571\ : LocalMux
    port map (
            O => \N__28007\,
            I => \N__28004\
        );

    \I__6570\ : Span4Mux_h
    port map (
            O => \N__28004\,
            I => \N__28001\
        );

    \I__6569\ : Odrv4
    port map (
            O => \N__28001\,
            I => \eeprom.n3070\
        );

    \I__6568\ : InMux
    port map (
            O => \N__27998\,
            I => \bfn_16_25_0_\
        );

    \I__6567\ : InMux
    port map (
            O => \N__27995\,
            I => \N__27991\
        );

    \I__6566\ : InMux
    port map (
            O => \N__27994\,
            I => \N__27988\
        );

    \I__6565\ : LocalMux
    port map (
            O => \N__27991\,
            I => \N__27984\
        );

    \I__6564\ : LocalMux
    port map (
            O => \N__27988\,
            I => \N__27981\
        );

    \I__6563\ : InMux
    port map (
            O => \N__27987\,
            I => \N__27978\
        );

    \I__6562\ : Span12Mux_s9_v
    port map (
            O => \N__27984\,
            I => \N__27975\
        );

    \I__6561\ : Span4Mux_v
    port map (
            O => \N__27981\,
            I => \N__27970\
        );

    \I__6560\ : LocalMux
    port map (
            O => \N__27978\,
            I => \N__27970\
        );

    \I__6559\ : Odrv12
    port map (
            O => \N__27975\,
            I => \eeprom.n3002\
        );

    \I__6558\ : Odrv4
    port map (
            O => \N__27970\,
            I => \eeprom.n3002\
        );

    \I__6557\ : CascadeMux
    port map (
            O => \N__27965\,
            I => \N__27962\
        );

    \I__6556\ : InMux
    port map (
            O => \N__27962\,
            I => \N__27959\
        );

    \I__6555\ : LocalMux
    port map (
            O => \N__27959\,
            I => \N__27956\
        );

    \I__6554\ : Span4Mux_v
    port map (
            O => \N__27956\,
            I => \N__27953\
        );

    \I__6553\ : Odrv4
    port map (
            O => \N__27953\,
            I => \eeprom.n3069\
        );

    \I__6552\ : InMux
    port map (
            O => \N__27950\,
            I => \eeprom.n3665\
        );

    \I__6551\ : InMux
    port map (
            O => \N__27947\,
            I => \N__27944\
        );

    \I__6550\ : LocalMux
    port map (
            O => \N__27944\,
            I => \N__27940\
        );

    \I__6549\ : CascadeMux
    port map (
            O => \N__27943\,
            I => \N__27937\
        );

    \I__6548\ : Span4Mux_h
    port map (
            O => \N__27940\,
            I => \N__27934\
        );

    \I__6547\ : InMux
    port map (
            O => \N__27937\,
            I => \N__27931\
        );

    \I__6546\ : Span4Mux_h
    port map (
            O => \N__27934\,
            I => \N__27928\
        );

    \I__6545\ : LocalMux
    port map (
            O => \N__27931\,
            I => \N__27925\
        );

    \I__6544\ : Odrv4
    port map (
            O => \N__27928\,
            I => \eeprom.n3001\
        );

    \I__6543\ : Odrv4
    port map (
            O => \N__27925\,
            I => \eeprom.n3001\
        );

    \I__6542\ : CascadeMux
    port map (
            O => \N__27920\,
            I => \N__27916\
        );

    \I__6541\ : CascadeMux
    port map (
            O => \N__27919\,
            I => \N__27912\
        );

    \I__6540\ : InMux
    port map (
            O => \N__27916\,
            I => \N__27904\
        );

    \I__6539\ : CascadeMux
    port map (
            O => \N__27915\,
            I => \N__27899\
        );

    \I__6538\ : InMux
    port map (
            O => \N__27912\,
            I => \N__27894\
        );

    \I__6537\ : InMux
    port map (
            O => \N__27911\,
            I => \N__27894\
        );

    \I__6536\ : CascadeMux
    port map (
            O => \N__27910\,
            I => \N__27891\
        );

    \I__6535\ : CascadeMux
    port map (
            O => \N__27909\,
            I => \N__27883\
        );

    \I__6534\ : CascadeMux
    port map (
            O => \N__27908\,
            I => \N__27878\
        );

    \I__6533\ : CascadeMux
    port map (
            O => \N__27907\,
            I => \N__27875\
        );

    \I__6532\ : LocalMux
    port map (
            O => \N__27904\,
            I => \N__27871\
        );

    \I__6531\ : InMux
    port map (
            O => \N__27903\,
            I => \N__27864\
        );

    \I__6530\ : InMux
    port map (
            O => \N__27902\,
            I => \N__27864\
        );

    \I__6529\ : InMux
    port map (
            O => \N__27899\,
            I => \N__27864\
        );

    \I__6528\ : LocalMux
    port map (
            O => \N__27894\,
            I => \N__27861\
        );

    \I__6527\ : InMux
    port map (
            O => \N__27891\,
            I => \N__27856\
        );

    \I__6526\ : InMux
    port map (
            O => \N__27890\,
            I => \N__27856\
        );

    \I__6525\ : InMux
    port map (
            O => \N__27889\,
            I => \N__27851\
        );

    \I__6524\ : InMux
    port map (
            O => \N__27888\,
            I => \N__27851\
        );

    \I__6523\ : InMux
    port map (
            O => \N__27887\,
            I => \N__27848\
        );

    \I__6522\ : InMux
    port map (
            O => \N__27886\,
            I => \N__27839\
        );

    \I__6521\ : InMux
    port map (
            O => \N__27883\,
            I => \N__27839\
        );

    \I__6520\ : InMux
    port map (
            O => \N__27882\,
            I => \N__27839\
        );

    \I__6519\ : InMux
    port map (
            O => \N__27881\,
            I => \N__27839\
        );

    \I__6518\ : InMux
    port map (
            O => \N__27878\,
            I => \N__27832\
        );

    \I__6517\ : InMux
    port map (
            O => \N__27875\,
            I => \N__27832\
        );

    \I__6516\ : InMux
    port map (
            O => \N__27874\,
            I => \N__27832\
        );

    \I__6515\ : Span4Mux_h
    port map (
            O => \N__27871\,
            I => \N__27829\
        );

    \I__6514\ : LocalMux
    port map (
            O => \N__27864\,
            I => \N__27824\
        );

    \I__6513\ : Span4Mux_h
    port map (
            O => \N__27861\,
            I => \N__27824\
        );

    \I__6512\ : LocalMux
    port map (
            O => \N__27856\,
            I => \eeprom.n3034\
        );

    \I__6511\ : LocalMux
    port map (
            O => \N__27851\,
            I => \eeprom.n3034\
        );

    \I__6510\ : LocalMux
    port map (
            O => \N__27848\,
            I => \eeprom.n3034\
        );

    \I__6509\ : LocalMux
    port map (
            O => \N__27839\,
            I => \eeprom.n3034\
        );

    \I__6508\ : LocalMux
    port map (
            O => \N__27832\,
            I => \eeprom.n3034\
        );

    \I__6507\ : Odrv4
    port map (
            O => \N__27829\,
            I => \eeprom.n3034\
        );

    \I__6506\ : Odrv4
    port map (
            O => \N__27824\,
            I => \eeprom.n3034\
        );

    \I__6505\ : InMux
    port map (
            O => \N__27809\,
            I => \eeprom.n3666\
        );

    \I__6504\ : InMux
    port map (
            O => \N__27806\,
            I => \N__27802\
        );

    \I__6503\ : InMux
    port map (
            O => \N__27805\,
            I => \N__27799\
        );

    \I__6502\ : LocalMux
    port map (
            O => \N__27802\,
            I => \N__27794\
        );

    \I__6501\ : LocalMux
    port map (
            O => \N__27799\,
            I => \N__27794\
        );

    \I__6500\ : Span4Mux_v
    port map (
            O => \N__27794\,
            I => \N__27791\
        );

    \I__6499\ : Odrv4
    port map (
            O => \N__27791\,
            I => \eeprom.n3100\
        );

    \I__6498\ : CascadeMux
    port map (
            O => \N__27788\,
            I => \N__27770\
        );

    \I__6497\ : CascadeMux
    port map (
            O => \N__27787\,
            I => \N__27762\
        );

    \I__6496\ : CascadeMux
    port map (
            O => \N__27786\,
            I => \N__27757\
        );

    \I__6495\ : CascadeMux
    port map (
            O => \N__27785\,
            I => \N__27739\
        );

    \I__6494\ : CascadeMux
    port map (
            O => \N__27784\,
            I => \N__27736\
        );

    \I__6493\ : CascadeMux
    port map (
            O => \N__27783\,
            I => \N__27733\
        );

    \I__6492\ : InMux
    port map (
            O => \N__27782\,
            I => \N__27716\
        );

    \I__6491\ : InMux
    port map (
            O => \N__27781\,
            I => \N__27716\
        );

    \I__6490\ : InMux
    port map (
            O => \N__27780\,
            I => \N__27701\
        );

    \I__6489\ : InMux
    port map (
            O => \N__27779\,
            I => \N__27701\
        );

    \I__6488\ : InMux
    port map (
            O => \N__27778\,
            I => \N__27694\
        );

    \I__6487\ : InMux
    port map (
            O => \N__27777\,
            I => \N__27694\
        );

    \I__6486\ : InMux
    port map (
            O => \N__27776\,
            I => \N__27694\
        );

    \I__6485\ : InMux
    port map (
            O => \N__27775\,
            I => \N__27683\
        );

    \I__6484\ : InMux
    port map (
            O => \N__27774\,
            I => \N__27683\
        );

    \I__6483\ : InMux
    port map (
            O => \N__27773\,
            I => \N__27683\
        );

    \I__6482\ : InMux
    port map (
            O => \N__27770\,
            I => \N__27683\
        );

    \I__6481\ : InMux
    port map (
            O => \N__27769\,
            I => \N__27683\
        );

    \I__6480\ : CascadeMux
    port map (
            O => \N__27768\,
            I => \N__27680\
        );

    \I__6479\ : CascadeMux
    port map (
            O => \N__27767\,
            I => \N__27677\
        );

    \I__6478\ : CascadeMux
    port map (
            O => \N__27766\,
            I => \N__27674\
        );

    \I__6477\ : CascadeMux
    port map (
            O => \N__27765\,
            I => \N__27671\
        );

    \I__6476\ : InMux
    port map (
            O => \N__27762\,
            I => \N__27659\
        );

    \I__6475\ : InMux
    port map (
            O => \N__27761\,
            I => \N__27659\
        );

    \I__6474\ : InMux
    port map (
            O => \N__27760\,
            I => \N__27659\
        );

    \I__6473\ : InMux
    port map (
            O => \N__27757\,
            I => \N__27659\
        );

    \I__6472\ : InMux
    port map (
            O => \N__27756\,
            I => \N__27659\
        );

    \I__6471\ : InMux
    port map (
            O => \N__27755\,
            I => \N__27654\
        );

    \I__6470\ : InMux
    port map (
            O => \N__27754\,
            I => \N__27654\
        );

    \I__6469\ : CascadeMux
    port map (
            O => \N__27753\,
            I => \N__27650\
        );

    \I__6468\ : CascadeMux
    port map (
            O => \N__27752\,
            I => \N__27644\
        );

    \I__6467\ : CascadeMux
    port map (
            O => \N__27751\,
            I => \N__27638\
        );

    \I__6466\ : CascadeMux
    port map (
            O => \N__27750\,
            I => \N__27635\
        );

    \I__6465\ : InMux
    port map (
            O => \N__27749\,
            I => \N__27630\
        );

    \I__6464\ : InMux
    port map (
            O => \N__27748\,
            I => \N__27630\
        );

    \I__6463\ : CascadeMux
    port map (
            O => \N__27747\,
            I => \N__27624\
        );

    \I__6462\ : CascadeMux
    port map (
            O => \N__27746\,
            I => \N__27621\
        );

    \I__6461\ : CascadeMux
    port map (
            O => \N__27745\,
            I => \N__27617\
        );

    \I__6460\ : CascadeMux
    port map (
            O => \N__27744\,
            I => \N__27614\
        );

    \I__6459\ : CascadeMux
    port map (
            O => \N__27743\,
            I => \N__27608\
        );

    \I__6458\ : InMux
    port map (
            O => \N__27742\,
            I => \N__27599\
        );

    \I__6457\ : InMux
    port map (
            O => \N__27739\,
            I => \N__27599\
        );

    \I__6456\ : InMux
    port map (
            O => \N__27736\,
            I => \N__27596\
        );

    \I__6455\ : InMux
    port map (
            O => \N__27733\,
            I => \N__27591\
        );

    \I__6454\ : InMux
    port map (
            O => \N__27732\,
            I => \N__27591\
        );

    \I__6453\ : InMux
    port map (
            O => \N__27731\,
            I => \N__27583\
        );

    \I__6452\ : InMux
    port map (
            O => \N__27730\,
            I => \N__27578\
        );

    \I__6451\ : CascadeMux
    port map (
            O => \N__27729\,
            I => \N__27575\
        );

    \I__6450\ : InMux
    port map (
            O => \N__27728\,
            I => \N__27570\
        );

    \I__6449\ : InMux
    port map (
            O => \N__27727\,
            I => \N__27570\
        );

    \I__6448\ : CascadeMux
    port map (
            O => \N__27726\,
            I => \N__27566\
        );

    \I__6447\ : CascadeMux
    port map (
            O => \N__27725\,
            I => \N__27561\
        );

    \I__6446\ : CascadeMux
    port map (
            O => \N__27724\,
            I => \N__27557\
        );

    \I__6445\ : CascadeMux
    port map (
            O => \N__27723\,
            I => \N__27553\
        );

    \I__6444\ : CascadeMux
    port map (
            O => \N__27722\,
            I => \N__27550\
        );

    \I__6443\ : CascadeMux
    port map (
            O => \N__27721\,
            I => \N__27547\
        );

    \I__6442\ : LocalMux
    port map (
            O => \N__27716\,
            I => \N__27538\
        );

    \I__6441\ : InMux
    port map (
            O => \N__27715\,
            I => \N__27529\
        );

    \I__6440\ : InMux
    port map (
            O => \N__27714\,
            I => \N__27529\
        );

    \I__6439\ : InMux
    port map (
            O => \N__27713\,
            I => \N__27529\
        );

    \I__6438\ : InMux
    port map (
            O => \N__27712\,
            I => \N__27529\
        );

    \I__6437\ : InMux
    port map (
            O => \N__27711\,
            I => \N__27520\
        );

    \I__6436\ : InMux
    port map (
            O => \N__27710\,
            I => \N__27520\
        );

    \I__6435\ : InMux
    port map (
            O => \N__27709\,
            I => \N__27520\
        );

    \I__6434\ : InMux
    port map (
            O => \N__27708\,
            I => \N__27520\
        );

    \I__6433\ : CascadeMux
    port map (
            O => \N__27707\,
            I => \N__27515\
        );

    \I__6432\ : CascadeMux
    port map (
            O => \N__27706\,
            I => \N__27510\
        );

    \I__6431\ : LocalMux
    port map (
            O => \N__27701\,
            I => \N__27504\
        );

    \I__6430\ : LocalMux
    port map (
            O => \N__27694\,
            I => \N__27504\
        );

    \I__6429\ : LocalMux
    port map (
            O => \N__27683\,
            I => \N__27501\
        );

    \I__6428\ : InMux
    port map (
            O => \N__27680\,
            I => \N__27490\
        );

    \I__6427\ : InMux
    port map (
            O => \N__27677\,
            I => \N__27490\
        );

    \I__6426\ : InMux
    port map (
            O => \N__27674\,
            I => \N__27490\
        );

    \I__6425\ : InMux
    port map (
            O => \N__27671\,
            I => \N__27490\
        );

    \I__6424\ : InMux
    port map (
            O => \N__27670\,
            I => \N__27490\
        );

    \I__6423\ : LocalMux
    port map (
            O => \N__27659\,
            I => \N__27485\
        );

    \I__6422\ : LocalMux
    port map (
            O => \N__27654\,
            I => \N__27485\
        );

    \I__6421\ : InMux
    port map (
            O => \N__27653\,
            I => \N__27476\
        );

    \I__6420\ : InMux
    port map (
            O => \N__27650\,
            I => \N__27476\
        );

    \I__6419\ : InMux
    port map (
            O => \N__27649\,
            I => \N__27476\
        );

    \I__6418\ : InMux
    port map (
            O => \N__27648\,
            I => \N__27476\
        );

    \I__6417\ : InMux
    port map (
            O => \N__27647\,
            I => \N__27467\
        );

    \I__6416\ : InMux
    port map (
            O => \N__27644\,
            I => \N__27467\
        );

    \I__6415\ : InMux
    port map (
            O => \N__27643\,
            I => \N__27467\
        );

    \I__6414\ : InMux
    port map (
            O => \N__27642\,
            I => \N__27467\
        );

    \I__6413\ : InMux
    port map (
            O => \N__27641\,
            I => \N__27460\
        );

    \I__6412\ : InMux
    port map (
            O => \N__27638\,
            I => \N__27460\
        );

    \I__6411\ : InMux
    port map (
            O => \N__27635\,
            I => \N__27460\
        );

    \I__6410\ : LocalMux
    port map (
            O => \N__27630\,
            I => \N__27456\
        );

    \I__6409\ : InMux
    port map (
            O => \N__27629\,
            I => \N__27453\
        );

    \I__6408\ : InMux
    port map (
            O => \N__27628\,
            I => \N__27448\
        );

    \I__6407\ : InMux
    port map (
            O => \N__27627\,
            I => \N__27448\
        );

    \I__6406\ : InMux
    port map (
            O => \N__27624\,
            I => \N__27443\
        );

    \I__6405\ : InMux
    port map (
            O => \N__27621\,
            I => \N__27443\
        );

    \I__6404\ : InMux
    port map (
            O => \N__27620\,
            I => \N__27436\
        );

    \I__6403\ : InMux
    port map (
            O => \N__27617\,
            I => \N__27436\
        );

    \I__6402\ : InMux
    port map (
            O => \N__27614\,
            I => \N__27436\
        );

    \I__6401\ : InMux
    port map (
            O => \N__27613\,
            I => \N__27431\
        );

    \I__6400\ : InMux
    port map (
            O => \N__27612\,
            I => \N__27431\
        );

    \I__6399\ : InMux
    port map (
            O => \N__27611\,
            I => \N__27428\
        );

    \I__6398\ : InMux
    port map (
            O => \N__27608\,
            I => \N__27423\
        );

    \I__6397\ : InMux
    port map (
            O => \N__27607\,
            I => \N__27423\
        );

    \I__6396\ : CascadeMux
    port map (
            O => \N__27606\,
            I => \N__27418\
        );

    \I__6395\ : CascadeMux
    port map (
            O => \N__27605\,
            I => \N__27415\
        );

    \I__6394\ : CascadeMux
    port map (
            O => \N__27604\,
            I => \N__27412\
        );

    \I__6393\ : LocalMux
    port map (
            O => \N__27599\,
            I => \N__27407\
        );

    \I__6392\ : LocalMux
    port map (
            O => \N__27596\,
            I => \N__27402\
        );

    \I__6391\ : LocalMux
    port map (
            O => \N__27591\,
            I => \N__27402\
        );

    \I__6390\ : InMux
    port map (
            O => \N__27590\,
            I => \N__27397\
        );

    \I__6389\ : InMux
    port map (
            O => \N__27589\,
            I => \N__27397\
        );

    \I__6388\ : CascadeMux
    port map (
            O => \N__27588\,
            I => \N__27394\
        );

    \I__6387\ : CascadeMux
    port map (
            O => \N__27587\,
            I => \N__27390\
        );

    \I__6386\ : CascadeMux
    port map (
            O => \N__27586\,
            I => \N__27387\
        );

    \I__6385\ : LocalMux
    port map (
            O => \N__27583\,
            I => \N__27378\
        );

    \I__6384\ : InMux
    port map (
            O => \N__27582\,
            I => \N__27375\
        );

    \I__6383\ : CascadeMux
    port map (
            O => \N__27581\,
            I => \N__27372\
        );

    \I__6382\ : LocalMux
    port map (
            O => \N__27578\,
            I => \N__27368\
        );

    \I__6381\ : InMux
    port map (
            O => \N__27575\,
            I => \N__27365\
        );

    \I__6380\ : LocalMux
    port map (
            O => \N__27570\,
            I => \N__27362\
        );

    \I__6379\ : InMux
    port map (
            O => \N__27569\,
            I => \N__27357\
        );

    \I__6378\ : InMux
    port map (
            O => \N__27566\,
            I => \N__27357\
        );

    \I__6377\ : InMux
    port map (
            O => \N__27565\,
            I => \N__27348\
        );

    \I__6376\ : InMux
    port map (
            O => \N__27564\,
            I => \N__27348\
        );

    \I__6375\ : InMux
    port map (
            O => \N__27561\,
            I => \N__27348\
        );

    \I__6374\ : InMux
    port map (
            O => \N__27560\,
            I => \N__27348\
        );

    \I__6373\ : InMux
    port map (
            O => \N__27557\,
            I => \N__27345\
        );

    \I__6372\ : InMux
    port map (
            O => \N__27556\,
            I => \N__27342\
        );

    \I__6371\ : InMux
    port map (
            O => \N__27553\,
            I => \N__27335\
        );

    \I__6370\ : InMux
    port map (
            O => \N__27550\,
            I => \N__27335\
        );

    \I__6369\ : InMux
    port map (
            O => \N__27547\,
            I => \N__27335\
        );

    \I__6368\ : CascadeMux
    port map (
            O => \N__27546\,
            I => \N__27327\
        );

    \I__6367\ : CascadeMux
    port map (
            O => \N__27545\,
            I => \N__27322\
        );

    \I__6366\ : CascadeMux
    port map (
            O => \N__27544\,
            I => \N__27319\
        );

    \I__6365\ : CascadeMux
    port map (
            O => \N__27543\,
            I => \N__27315\
        );

    \I__6364\ : CascadeMux
    port map (
            O => \N__27542\,
            I => \N__27312\
        );

    \I__6363\ : CascadeMux
    port map (
            O => \N__27541\,
            I => \N__27307\
        );

    \I__6362\ : Span4Mux_v
    port map (
            O => \N__27538\,
            I => \N__27295\
        );

    \I__6361\ : LocalMux
    port map (
            O => \N__27529\,
            I => \N__27295\
        );

    \I__6360\ : LocalMux
    port map (
            O => \N__27520\,
            I => \N__27295\
        );

    \I__6359\ : InMux
    port map (
            O => \N__27519\,
            I => \N__27290\
        );

    \I__6358\ : InMux
    port map (
            O => \N__27518\,
            I => \N__27290\
        );

    \I__6357\ : InMux
    port map (
            O => \N__27515\,
            I => \N__27279\
        );

    \I__6356\ : InMux
    port map (
            O => \N__27514\,
            I => \N__27279\
        );

    \I__6355\ : InMux
    port map (
            O => \N__27513\,
            I => \N__27279\
        );

    \I__6354\ : InMux
    port map (
            O => \N__27510\,
            I => \N__27279\
        );

    \I__6353\ : InMux
    port map (
            O => \N__27509\,
            I => \N__27279\
        );

    \I__6352\ : Span4Mux_h
    port map (
            O => \N__27504\,
            I => \N__27272\
        );

    \I__6351\ : Span4Mux_h
    port map (
            O => \N__27501\,
            I => \N__27272\
        );

    \I__6350\ : LocalMux
    port map (
            O => \N__27490\,
            I => \N__27272\
        );

    \I__6349\ : Span4Mux_v
    port map (
            O => \N__27485\,
            I => \N__27263\
        );

    \I__6348\ : LocalMux
    port map (
            O => \N__27476\,
            I => \N__27263\
        );

    \I__6347\ : LocalMux
    port map (
            O => \N__27467\,
            I => \N__27263\
        );

    \I__6346\ : LocalMux
    port map (
            O => \N__27460\,
            I => \N__27263\
        );

    \I__6345\ : InMux
    port map (
            O => \N__27459\,
            I => \N__27260\
        );

    \I__6344\ : Span4Mux_v
    port map (
            O => \N__27456\,
            I => \N__27255\
        );

    \I__6343\ : LocalMux
    port map (
            O => \N__27453\,
            I => \N__27255\
        );

    \I__6342\ : LocalMux
    port map (
            O => \N__27448\,
            I => \N__27252\
        );

    \I__6341\ : LocalMux
    port map (
            O => \N__27443\,
            I => \N__27247\
        );

    \I__6340\ : LocalMux
    port map (
            O => \N__27436\,
            I => \N__27247\
        );

    \I__6339\ : LocalMux
    port map (
            O => \N__27431\,
            I => \N__27240\
        );

    \I__6338\ : LocalMux
    port map (
            O => \N__27428\,
            I => \N__27240\
        );

    \I__6337\ : LocalMux
    port map (
            O => \N__27423\,
            I => \N__27240\
        );

    \I__6336\ : InMux
    port map (
            O => \N__27422\,
            I => \N__27235\
        );

    \I__6335\ : InMux
    port map (
            O => \N__27421\,
            I => \N__27235\
        );

    \I__6334\ : InMux
    port map (
            O => \N__27418\,
            I => \N__27226\
        );

    \I__6333\ : InMux
    port map (
            O => \N__27415\,
            I => \N__27226\
        );

    \I__6332\ : InMux
    port map (
            O => \N__27412\,
            I => \N__27226\
        );

    \I__6331\ : InMux
    port map (
            O => \N__27411\,
            I => \N__27226\
        );

    \I__6330\ : InMux
    port map (
            O => \N__27410\,
            I => \N__27223\
        );

    \I__6329\ : Span4Mux_s3_h
    port map (
            O => \N__27407\,
            I => \N__27218\
        );

    \I__6328\ : Span4Mux_v
    port map (
            O => \N__27402\,
            I => \N__27218\
        );

    \I__6327\ : LocalMux
    port map (
            O => \N__27397\,
            I => \N__27215\
        );

    \I__6326\ : InMux
    port map (
            O => \N__27394\,
            I => \N__27206\
        );

    \I__6325\ : InMux
    port map (
            O => \N__27393\,
            I => \N__27206\
        );

    \I__6324\ : InMux
    port map (
            O => \N__27390\,
            I => \N__27206\
        );

    \I__6323\ : InMux
    port map (
            O => \N__27387\,
            I => \N__27206\
        );

    \I__6322\ : CascadeMux
    port map (
            O => \N__27386\,
            I => \N__27202\
        );

    \I__6321\ : CascadeMux
    port map (
            O => \N__27385\,
            I => \N__27199\
        );

    \I__6320\ : CascadeMux
    port map (
            O => \N__27384\,
            I => \N__27196\
        );

    \I__6319\ : InMux
    port map (
            O => \N__27383\,
            I => \N__27182\
        );

    \I__6318\ : CascadeMux
    port map (
            O => \N__27382\,
            I => \N__27176\
        );

    \I__6317\ : CascadeMux
    port map (
            O => \N__27381\,
            I => \N__27171\
        );

    \I__6316\ : Span4Mux_v
    port map (
            O => \N__27378\,
            I => \N__27166\
        );

    \I__6315\ : LocalMux
    port map (
            O => \N__27375\,
            I => \N__27166\
        );

    \I__6314\ : InMux
    port map (
            O => \N__27372\,
            I => \N__27163\
        );

    \I__6313\ : InMux
    port map (
            O => \N__27371\,
            I => \N__27160\
        );

    \I__6312\ : Span4Mux_v
    port map (
            O => \N__27368\,
            I => \N__27155\
        );

    \I__6311\ : LocalMux
    port map (
            O => \N__27365\,
            I => \N__27155\
        );

    \I__6310\ : Span4Mux_v
    port map (
            O => \N__27362\,
            I => \N__27142\
        );

    \I__6309\ : LocalMux
    port map (
            O => \N__27357\,
            I => \N__27142\
        );

    \I__6308\ : LocalMux
    port map (
            O => \N__27348\,
            I => \N__27142\
        );

    \I__6307\ : LocalMux
    port map (
            O => \N__27345\,
            I => \N__27142\
        );

    \I__6306\ : LocalMux
    port map (
            O => \N__27342\,
            I => \N__27142\
        );

    \I__6305\ : LocalMux
    port map (
            O => \N__27335\,
            I => \N__27142\
        );

    \I__6304\ : CascadeMux
    port map (
            O => \N__27334\,
            I => \N__27139\
        );

    \I__6303\ : CascadeMux
    port map (
            O => \N__27333\,
            I => \N__27136\
        );

    \I__6302\ : CascadeMux
    port map (
            O => \N__27332\,
            I => \N__27133\
        );

    \I__6301\ : CascadeMux
    port map (
            O => \N__27331\,
            I => \N__27130\
        );

    \I__6300\ : CascadeMux
    port map (
            O => \N__27330\,
            I => \N__27127\
        );

    \I__6299\ : InMux
    port map (
            O => \N__27327\,
            I => \N__27123\
        );

    \I__6298\ : InMux
    port map (
            O => \N__27326\,
            I => \N__27118\
        );

    \I__6297\ : InMux
    port map (
            O => \N__27325\,
            I => \N__27118\
        );

    \I__6296\ : InMux
    port map (
            O => \N__27322\,
            I => \N__27109\
        );

    \I__6295\ : InMux
    port map (
            O => \N__27319\,
            I => \N__27109\
        );

    \I__6294\ : InMux
    port map (
            O => \N__27318\,
            I => \N__27109\
        );

    \I__6293\ : InMux
    port map (
            O => \N__27315\,
            I => \N__27109\
        );

    \I__6292\ : InMux
    port map (
            O => \N__27312\,
            I => \N__27106\
        );

    \I__6291\ : InMux
    port map (
            O => \N__27311\,
            I => \N__27103\
        );

    \I__6290\ : InMux
    port map (
            O => \N__27310\,
            I => \N__27098\
        );

    \I__6289\ : InMux
    port map (
            O => \N__27307\,
            I => \N__27098\
        );

    \I__6288\ : CascadeMux
    port map (
            O => \N__27306\,
            I => \N__27095\
        );

    \I__6287\ : CascadeMux
    port map (
            O => \N__27305\,
            I => \N__27092\
        );

    \I__6286\ : CascadeMux
    port map (
            O => \N__27304\,
            I => \N__27088\
        );

    \I__6285\ : CascadeMux
    port map (
            O => \N__27303\,
            I => \N__27085\
        );

    \I__6284\ : CascadeMux
    port map (
            O => \N__27302\,
            I => \N__27081\
        );

    \I__6283\ : Span4Mux_h
    port map (
            O => \N__27295\,
            I => \N__27066\
        );

    \I__6282\ : LocalMux
    port map (
            O => \N__27290\,
            I => \N__27066\
        );

    \I__6281\ : LocalMux
    port map (
            O => \N__27279\,
            I => \N__27066\
        );

    \I__6280\ : Span4Mux_v
    port map (
            O => \N__27272\,
            I => \N__27059\
        );

    \I__6279\ : Span4Mux_h
    port map (
            O => \N__27263\,
            I => \N__27059\
        );

    \I__6278\ : LocalMux
    port map (
            O => \N__27260\,
            I => \N__27059\
        );

    \I__6277\ : Span4Mux_v
    port map (
            O => \N__27255\,
            I => \N__27048\
        );

    \I__6276\ : Span4Mux_v
    port map (
            O => \N__27252\,
            I => \N__27048\
        );

    \I__6275\ : Span4Mux_h
    port map (
            O => \N__27247\,
            I => \N__27048\
        );

    \I__6274\ : Span4Mux_v
    port map (
            O => \N__27240\,
            I => \N__27048\
        );

    \I__6273\ : LocalMux
    port map (
            O => \N__27235\,
            I => \N__27048\
        );

    \I__6272\ : LocalMux
    port map (
            O => \N__27226\,
            I => \N__27043\
        );

    \I__6271\ : LocalMux
    port map (
            O => \N__27223\,
            I => \N__27043\
        );

    \I__6270\ : Span4Mux_h
    port map (
            O => \N__27218\,
            I => \N__27036\
        );

    \I__6269\ : Span4Mux_v
    port map (
            O => \N__27215\,
            I => \N__27036\
        );

    \I__6268\ : LocalMux
    port map (
            O => \N__27206\,
            I => \N__27036\
        );

    \I__6267\ : InMux
    port map (
            O => \N__27205\,
            I => \N__27031\
        );

    \I__6266\ : InMux
    port map (
            O => \N__27202\,
            I => \N__27031\
        );

    \I__6265\ : InMux
    port map (
            O => \N__27199\,
            I => \N__27026\
        );

    \I__6264\ : InMux
    port map (
            O => \N__27196\,
            I => \N__27026\
        );

    \I__6263\ : CascadeMux
    port map (
            O => \N__27195\,
            I => \N__27021\
        );

    \I__6262\ : CascadeMux
    port map (
            O => \N__27194\,
            I => \N__27018\
        );

    \I__6261\ : CascadeMux
    port map (
            O => \N__27193\,
            I => \N__27013\
        );

    \I__6260\ : CascadeMux
    port map (
            O => \N__27192\,
            I => \N__27010\
        );

    \I__6259\ : CascadeMux
    port map (
            O => \N__27191\,
            I => \N__27005\
        );

    \I__6258\ : CascadeMux
    port map (
            O => \N__27190\,
            I => \N__27002\
        );

    \I__6257\ : CascadeMux
    port map (
            O => \N__27189\,
            I => \N__26999\
        );

    \I__6256\ : CascadeMux
    port map (
            O => \N__27188\,
            I => \N__26995\
        );

    \I__6255\ : CascadeMux
    port map (
            O => \N__27187\,
            I => \N__26992\
        );

    \I__6254\ : CascadeMux
    port map (
            O => \N__27186\,
            I => \N__26989\
        );

    \I__6253\ : CascadeMux
    port map (
            O => \N__27185\,
            I => \N__26984\
        );

    \I__6252\ : LocalMux
    port map (
            O => \N__27182\,
            I => \N__26981\
        );

    \I__6251\ : InMux
    port map (
            O => \N__27181\,
            I => \N__26978\
        );

    \I__6250\ : InMux
    port map (
            O => \N__27180\,
            I => \N__26973\
        );

    \I__6249\ : InMux
    port map (
            O => \N__27179\,
            I => \N__26973\
        );

    \I__6248\ : InMux
    port map (
            O => \N__27176\,
            I => \N__26964\
        );

    \I__6247\ : InMux
    port map (
            O => \N__27175\,
            I => \N__26964\
        );

    \I__6246\ : InMux
    port map (
            O => \N__27174\,
            I => \N__26964\
        );

    \I__6245\ : InMux
    port map (
            O => \N__27171\,
            I => \N__26964\
        );

    \I__6244\ : Sp12to4
    port map (
            O => \N__27166\,
            I => \N__26957\
        );

    \I__6243\ : LocalMux
    port map (
            O => \N__27163\,
            I => \N__26957\
        );

    \I__6242\ : LocalMux
    port map (
            O => \N__27160\,
            I => \N__26957\
        );

    \I__6241\ : Span4Mux_h
    port map (
            O => \N__27155\,
            I => \N__26952\
        );

    \I__6240\ : Span4Mux_v
    port map (
            O => \N__27142\,
            I => \N__26952\
        );

    \I__6239\ : InMux
    port map (
            O => \N__27139\,
            I => \N__26947\
        );

    \I__6238\ : InMux
    port map (
            O => \N__27136\,
            I => \N__26947\
        );

    \I__6237\ : InMux
    port map (
            O => \N__27133\,
            I => \N__26938\
        );

    \I__6236\ : InMux
    port map (
            O => \N__27130\,
            I => \N__26938\
        );

    \I__6235\ : InMux
    port map (
            O => \N__27127\,
            I => \N__26938\
        );

    \I__6234\ : InMux
    port map (
            O => \N__27126\,
            I => \N__26938\
        );

    \I__6233\ : LocalMux
    port map (
            O => \N__27123\,
            I => \N__26933\
        );

    \I__6232\ : LocalMux
    port map (
            O => \N__27118\,
            I => \N__26922\
        );

    \I__6231\ : LocalMux
    port map (
            O => \N__27109\,
            I => \N__26922\
        );

    \I__6230\ : LocalMux
    port map (
            O => \N__27106\,
            I => \N__26922\
        );

    \I__6229\ : LocalMux
    port map (
            O => \N__27103\,
            I => \N__26922\
        );

    \I__6228\ : LocalMux
    port map (
            O => \N__27098\,
            I => \N__26922\
        );

    \I__6227\ : InMux
    port map (
            O => \N__27095\,
            I => \N__26919\
        );

    \I__6226\ : InMux
    port map (
            O => \N__27092\,
            I => \N__26904\
        );

    \I__6225\ : InMux
    port map (
            O => \N__27091\,
            I => \N__26904\
        );

    \I__6224\ : InMux
    port map (
            O => \N__27088\,
            I => \N__26904\
        );

    \I__6223\ : InMux
    port map (
            O => \N__27085\,
            I => \N__26904\
        );

    \I__6222\ : InMux
    port map (
            O => \N__27084\,
            I => \N__26904\
        );

    \I__6221\ : InMux
    port map (
            O => \N__27081\,
            I => \N__26904\
        );

    \I__6220\ : InMux
    port map (
            O => \N__27080\,
            I => \N__26904\
        );

    \I__6219\ : CascadeMux
    port map (
            O => \N__27079\,
            I => \N__26901\
        );

    \I__6218\ : CascadeMux
    port map (
            O => \N__27078\,
            I => \N__26898\
        );

    \I__6217\ : CascadeMux
    port map (
            O => \N__27077\,
            I => \N__26895\
        );

    \I__6216\ : CascadeMux
    port map (
            O => \N__27076\,
            I => \N__26892\
        );

    \I__6215\ : CascadeMux
    port map (
            O => \N__27075\,
            I => \N__26889\
        );

    \I__6214\ : CascadeMux
    port map (
            O => \N__27074\,
            I => \N__26886\
        );

    \I__6213\ : CascadeMux
    port map (
            O => \N__27073\,
            I => \N__26882\
        );

    \I__6212\ : Span4Mux_v
    port map (
            O => \N__27066\,
            I => \N__26877\
        );

    \I__6211\ : Span4Mux_v
    port map (
            O => \N__27059\,
            I => \N__26870\
        );

    \I__6210\ : Span4Mux_h
    port map (
            O => \N__27048\,
            I => \N__26870\
        );

    \I__6209\ : Span4Mux_v
    port map (
            O => \N__27043\,
            I => \N__26870\
        );

    \I__6208\ : Span4Mux_h
    port map (
            O => \N__27036\,
            I => \N__26863\
        );

    \I__6207\ : LocalMux
    port map (
            O => \N__27031\,
            I => \N__26863\
        );

    \I__6206\ : LocalMux
    port map (
            O => \N__27026\,
            I => \N__26863\
        );

    \I__6205\ : InMux
    port map (
            O => \N__27025\,
            I => \N__26858\
        );

    \I__6204\ : InMux
    port map (
            O => \N__27024\,
            I => \N__26858\
        );

    \I__6203\ : InMux
    port map (
            O => \N__27021\,
            I => \N__26849\
        );

    \I__6202\ : InMux
    port map (
            O => \N__27018\,
            I => \N__26849\
        );

    \I__6201\ : InMux
    port map (
            O => \N__27017\,
            I => \N__26849\
        );

    \I__6200\ : InMux
    port map (
            O => \N__27016\,
            I => \N__26849\
        );

    \I__6199\ : InMux
    port map (
            O => \N__27013\,
            I => \N__26840\
        );

    \I__6198\ : InMux
    port map (
            O => \N__27010\,
            I => \N__26840\
        );

    \I__6197\ : InMux
    port map (
            O => \N__27009\,
            I => \N__26840\
        );

    \I__6196\ : InMux
    port map (
            O => \N__27008\,
            I => \N__26840\
        );

    \I__6195\ : InMux
    port map (
            O => \N__27005\,
            I => \N__26833\
        );

    \I__6194\ : InMux
    port map (
            O => \N__27002\,
            I => \N__26833\
        );

    \I__6193\ : InMux
    port map (
            O => \N__26999\,
            I => \N__26833\
        );

    \I__6192\ : InMux
    port map (
            O => \N__26998\,
            I => \N__26822\
        );

    \I__6191\ : InMux
    port map (
            O => \N__26995\,
            I => \N__26822\
        );

    \I__6190\ : InMux
    port map (
            O => \N__26992\,
            I => \N__26822\
        );

    \I__6189\ : InMux
    port map (
            O => \N__26989\,
            I => \N__26822\
        );

    \I__6188\ : InMux
    port map (
            O => \N__26988\,
            I => \N__26822\
        );

    \I__6187\ : InMux
    port map (
            O => \N__26987\,
            I => \N__26817\
        );

    \I__6186\ : InMux
    port map (
            O => \N__26984\,
            I => \N__26817\
        );

    \I__6185\ : Span12Mux_v
    port map (
            O => \N__26981\,
            I => \N__26800\
        );

    \I__6184\ : LocalMux
    port map (
            O => \N__26978\,
            I => \N__26800\
        );

    \I__6183\ : LocalMux
    port map (
            O => \N__26973\,
            I => \N__26800\
        );

    \I__6182\ : LocalMux
    port map (
            O => \N__26964\,
            I => \N__26800\
        );

    \I__6181\ : Span12Mux_s10_v
    port map (
            O => \N__26957\,
            I => \N__26800\
        );

    \I__6180\ : Sp12to4
    port map (
            O => \N__26952\,
            I => \N__26800\
        );

    \I__6179\ : LocalMux
    port map (
            O => \N__26947\,
            I => \N__26800\
        );

    \I__6178\ : LocalMux
    port map (
            O => \N__26938\,
            I => \N__26800\
        );

    \I__6177\ : InMux
    port map (
            O => \N__26937\,
            I => \N__26795\
        );

    \I__6176\ : InMux
    port map (
            O => \N__26936\,
            I => \N__26795\
        );

    \I__6175\ : Span4Mux_h
    port map (
            O => \N__26933\,
            I => \N__26786\
        );

    \I__6174\ : Span4Mux_v
    port map (
            O => \N__26922\,
            I => \N__26786\
        );

    \I__6173\ : LocalMux
    port map (
            O => \N__26919\,
            I => \N__26786\
        );

    \I__6172\ : LocalMux
    port map (
            O => \N__26904\,
            I => \N__26786\
        );

    \I__6171\ : InMux
    port map (
            O => \N__26901\,
            I => \N__26779\
        );

    \I__6170\ : InMux
    port map (
            O => \N__26898\,
            I => \N__26779\
        );

    \I__6169\ : InMux
    port map (
            O => \N__26895\,
            I => \N__26779\
        );

    \I__6168\ : InMux
    port map (
            O => \N__26892\,
            I => \N__26768\
        );

    \I__6167\ : InMux
    port map (
            O => \N__26889\,
            I => \N__26768\
        );

    \I__6166\ : InMux
    port map (
            O => \N__26886\,
            I => \N__26768\
        );

    \I__6165\ : InMux
    port map (
            O => \N__26885\,
            I => \N__26768\
        );

    \I__6164\ : InMux
    port map (
            O => \N__26882\,
            I => \N__26768\
        );

    \I__6163\ : CascadeMux
    port map (
            O => \N__26881\,
            I => \N__26765\
        );

    \I__6162\ : CascadeMux
    port map (
            O => \N__26880\,
            I => \N__26761\
        );

    \I__6161\ : Span4Mux_v
    port map (
            O => \N__26877\,
            I => \N__26756\
        );

    \I__6160\ : Span4Mux_h
    port map (
            O => \N__26870\,
            I => \N__26756\
        );

    \I__6159\ : Span4Mux_h
    port map (
            O => \N__26863\,
            I => \N__26753\
        );

    \I__6158\ : LocalMux
    port map (
            O => \N__26858\,
            I => \N__26740\
        );

    \I__6157\ : LocalMux
    port map (
            O => \N__26849\,
            I => \N__26740\
        );

    \I__6156\ : LocalMux
    port map (
            O => \N__26840\,
            I => \N__26740\
        );

    \I__6155\ : LocalMux
    port map (
            O => \N__26833\,
            I => \N__26740\
        );

    \I__6154\ : LocalMux
    port map (
            O => \N__26822\,
            I => \N__26740\
        );

    \I__6153\ : LocalMux
    port map (
            O => \N__26817\,
            I => \N__26740\
        );

    \I__6152\ : Span12Mux_h
    port map (
            O => \N__26800\,
            I => \N__26735\
        );

    \I__6151\ : LocalMux
    port map (
            O => \N__26795\,
            I => \N__26735\
        );

    \I__6150\ : Span4Mux_h
    port map (
            O => \N__26786\,
            I => \N__26728\
        );

    \I__6149\ : LocalMux
    port map (
            O => \N__26779\,
            I => \N__26728\
        );

    \I__6148\ : LocalMux
    port map (
            O => \N__26768\,
            I => \N__26728\
        );

    \I__6147\ : InMux
    port map (
            O => \N__26765\,
            I => \N__26725\
        );

    \I__6146\ : InMux
    port map (
            O => \N__26764\,
            I => \N__26720\
        );

    \I__6145\ : InMux
    port map (
            O => \N__26761\,
            I => \N__26720\
        );

    \I__6144\ : Odrv4
    port map (
            O => \N__26756\,
            I => \CONSTANT_ONE_NET\
        );

    \I__6143\ : Odrv4
    port map (
            O => \N__26753\,
            I => \CONSTANT_ONE_NET\
        );

    \I__6142\ : Odrv12
    port map (
            O => \N__26740\,
            I => \CONSTANT_ONE_NET\
        );

    \I__6141\ : Odrv12
    port map (
            O => \N__26735\,
            I => \CONSTANT_ONE_NET\
        );

    \I__6140\ : Odrv4
    port map (
            O => \N__26728\,
            I => \CONSTANT_ONE_NET\
        );

    \I__6139\ : LocalMux
    port map (
            O => \N__26725\,
            I => \CONSTANT_ONE_NET\
        );

    \I__6138\ : LocalMux
    port map (
            O => \N__26720\,
            I => \CONSTANT_ONE_NET\
        );

    \I__6137\ : CascadeMux
    port map (
            O => \N__26705\,
            I => \N__26700\
        );

    \I__6136\ : InMux
    port map (
            O => \N__26704\,
            I => \N__26697\
        );

    \I__6135\ : InMux
    port map (
            O => \N__26703\,
            I => \N__26694\
        );

    \I__6134\ : InMux
    port map (
            O => \N__26700\,
            I => \N__26691\
        );

    \I__6133\ : LocalMux
    port map (
            O => \N__26697\,
            I => \N__26684\
        );

    \I__6132\ : LocalMux
    port map (
            O => \N__26694\,
            I => \N__26684\
        );

    \I__6131\ : LocalMux
    port map (
            O => \N__26691\,
            I => \N__26684\
        );

    \I__6130\ : Odrv12
    port map (
            O => \N__26684\,
            I => \eeprom.n3012\
        );

    \I__6129\ : InMux
    port map (
            O => \N__26681\,
            I => \N__26678\
        );

    \I__6128\ : LocalMux
    port map (
            O => \N__26678\,
            I => \eeprom.n3079\
        );

    \I__6127\ : InMux
    port map (
            O => \N__26675\,
            I => \eeprom.n3655\
        );

    \I__6126\ : InMux
    port map (
            O => \N__26672\,
            I => \N__26668\
        );

    \I__6125\ : InMux
    port map (
            O => \N__26671\,
            I => \N__26664\
        );

    \I__6124\ : LocalMux
    port map (
            O => \N__26668\,
            I => \N__26661\
        );

    \I__6123\ : InMux
    port map (
            O => \N__26667\,
            I => \N__26658\
        );

    \I__6122\ : LocalMux
    port map (
            O => \N__26664\,
            I => \eeprom.n3011\
        );

    \I__6121\ : Odrv4
    port map (
            O => \N__26661\,
            I => \eeprom.n3011\
        );

    \I__6120\ : LocalMux
    port map (
            O => \N__26658\,
            I => \eeprom.n3011\
        );

    \I__6119\ : CascadeMux
    port map (
            O => \N__26651\,
            I => \N__26648\
        );

    \I__6118\ : InMux
    port map (
            O => \N__26648\,
            I => \N__26645\
        );

    \I__6117\ : LocalMux
    port map (
            O => \N__26645\,
            I => \eeprom.n3078\
        );

    \I__6116\ : InMux
    port map (
            O => \N__26642\,
            I => \bfn_16_24_0_\
        );

    \I__6115\ : InMux
    port map (
            O => \N__26639\,
            I => \N__26636\
        );

    \I__6114\ : LocalMux
    port map (
            O => \N__26636\,
            I => \N__26631\
        );

    \I__6113\ : InMux
    port map (
            O => \N__26635\,
            I => \N__26628\
        );

    \I__6112\ : CascadeMux
    port map (
            O => \N__26634\,
            I => \N__26625\
        );

    \I__6111\ : Span4Mux_h
    port map (
            O => \N__26631\,
            I => \N__26620\
        );

    \I__6110\ : LocalMux
    port map (
            O => \N__26628\,
            I => \N__26620\
        );

    \I__6109\ : InMux
    port map (
            O => \N__26625\,
            I => \N__26617\
        );

    \I__6108\ : Span4Mux_h
    port map (
            O => \N__26620\,
            I => \N__26614\
        );

    \I__6107\ : LocalMux
    port map (
            O => \N__26617\,
            I => \N__26611\
        );

    \I__6106\ : Odrv4
    port map (
            O => \N__26614\,
            I => \eeprom.n3010\
        );

    \I__6105\ : Odrv12
    port map (
            O => \N__26611\,
            I => \eeprom.n3010\
        );

    \I__6104\ : CascadeMux
    port map (
            O => \N__26606\,
            I => \N__26603\
        );

    \I__6103\ : InMux
    port map (
            O => \N__26603\,
            I => \N__26600\
        );

    \I__6102\ : LocalMux
    port map (
            O => \N__26600\,
            I => \eeprom.n3077\
        );

    \I__6101\ : InMux
    port map (
            O => \N__26597\,
            I => \eeprom.n3657\
        );

    \I__6100\ : InMux
    port map (
            O => \N__26594\,
            I => \N__26590\
        );

    \I__6099\ : InMux
    port map (
            O => \N__26593\,
            I => \N__26587\
        );

    \I__6098\ : LocalMux
    port map (
            O => \N__26590\,
            I => \N__26583\
        );

    \I__6097\ : LocalMux
    port map (
            O => \N__26587\,
            I => \N__26580\
        );

    \I__6096\ : InMux
    port map (
            O => \N__26586\,
            I => \N__26577\
        );

    \I__6095\ : Span4Mux_h
    port map (
            O => \N__26583\,
            I => \N__26574\
        );

    \I__6094\ : Span4Mux_h
    port map (
            O => \N__26580\,
            I => \N__26571\
        );

    \I__6093\ : LocalMux
    port map (
            O => \N__26577\,
            I => \N__26568\
        );

    \I__6092\ : Odrv4
    port map (
            O => \N__26574\,
            I => \eeprom.n3009\
        );

    \I__6091\ : Odrv4
    port map (
            O => \N__26571\,
            I => \eeprom.n3009\
        );

    \I__6090\ : Odrv12
    port map (
            O => \N__26568\,
            I => \eeprom.n3009\
        );

    \I__6089\ : CascadeMux
    port map (
            O => \N__26561\,
            I => \N__26558\
        );

    \I__6088\ : InMux
    port map (
            O => \N__26558\,
            I => \N__26555\
        );

    \I__6087\ : LocalMux
    port map (
            O => \N__26555\,
            I => \N__26552\
        );

    \I__6086\ : Span4Mux_h
    port map (
            O => \N__26552\,
            I => \N__26549\
        );

    \I__6085\ : Odrv4
    port map (
            O => \N__26549\,
            I => \eeprom.n3076\
        );

    \I__6084\ : InMux
    port map (
            O => \N__26546\,
            I => \eeprom.n3658\
        );

    \I__6083\ : CascadeMux
    port map (
            O => \N__26543\,
            I => \N__26540\
        );

    \I__6082\ : InMux
    port map (
            O => \N__26540\,
            I => \N__26535\
        );

    \I__6081\ : InMux
    port map (
            O => \N__26539\,
            I => \N__26532\
        );

    \I__6080\ : InMux
    port map (
            O => \N__26538\,
            I => \N__26529\
        );

    \I__6079\ : LocalMux
    port map (
            O => \N__26535\,
            I => \eeprom.n3008\
        );

    \I__6078\ : LocalMux
    port map (
            O => \N__26532\,
            I => \eeprom.n3008\
        );

    \I__6077\ : LocalMux
    port map (
            O => \N__26529\,
            I => \eeprom.n3008\
        );

    \I__6076\ : InMux
    port map (
            O => \N__26522\,
            I => \N__26519\
        );

    \I__6075\ : LocalMux
    port map (
            O => \N__26519\,
            I => \eeprom.n3075\
        );

    \I__6074\ : InMux
    port map (
            O => \N__26516\,
            I => \eeprom.n3659\
        );

    \I__6073\ : InMux
    port map (
            O => \N__26513\,
            I => \N__26508\
        );

    \I__6072\ : InMux
    port map (
            O => \N__26512\,
            I => \N__26505\
        );

    \I__6071\ : InMux
    port map (
            O => \N__26511\,
            I => \N__26502\
        );

    \I__6070\ : LocalMux
    port map (
            O => \N__26508\,
            I => \N__26499\
        );

    \I__6069\ : LocalMux
    port map (
            O => \N__26505\,
            I => \N__26496\
        );

    \I__6068\ : LocalMux
    port map (
            O => \N__26502\,
            I => \N__26493\
        );

    \I__6067\ : Span4Mux_h
    port map (
            O => \N__26499\,
            I => \N__26490\
        );

    \I__6066\ : Odrv4
    port map (
            O => \N__26496\,
            I => \eeprom.n3007\
        );

    \I__6065\ : Odrv12
    port map (
            O => \N__26493\,
            I => \eeprom.n3007\
        );

    \I__6064\ : Odrv4
    port map (
            O => \N__26490\,
            I => \eeprom.n3007\
        );

    \I__6063\ : CascadeMux
    port map (
            O => \N__26483\,
            I => \N__26480\
        );

    \I__6062\ : InMux
    port map (
            O => \N__26480\,
            I => \N__26477\
        );

    \I__6061\ : LocalMux
    port map (
            O => \N__26477\,
            I => \N__26474\
        );

    \I__6060\ : Odrv4
    port map (
            O => \N__26474\,
            I => \eeprom.n3074\
        );

    \I__6059\ : InMux
    port map (
            O => \N__26471\,
            I => \eeprom.n3660\
        );

    \I__6058\ : InMux
    port map (
            O => \N__26468\,
            I => \N__26464\
        );

    \I__6057\ : InMux
    port map (
            O => \N__26467\,
            I => \N__26461\
        );

    \I__6056\ : LocalMux
    port map (
            O => \N__26464\,
            I => \N__26457\
        );

    \I__6055\ : LocalMux
    port map (
            O => \N__26461\,
            I => \N__26454\
        );

    \I__6054\ : InMux
    port map (
            O => \N__26460\,
            I => \N__26451\
        );

    \I__6053\ : Odrv4
    port map (
            O => \N__26457\,
            I => \eeprom.n3006\
        );

    \I__6052\ : Odrv4
    port map (
            O => \N__26454\,
            I => \eeprom.n3006\
        );

    \I__6051\ : LocalMux
    port map (
            O => \N__26451\,
            I => \eeprom.n3006\
        );

    \I__6050\ : CascadeMux
    port map (
            O => \N__26444\,
            I => \N__26441\
        );

    \I__6049\ : InMux
    port map (
            O => \N__26441\,
            I => \N__26438\
        );

    \I__6048\ : LocalMux
    port map (
            O => \N__26438\,
            I => \N__26435\
        );

    \I__6047\ : Span4Mux_v
    port map (
            O => \N__26435\,
            I => \N__26432\
        );

    \I__6046\ : Odrv4
    port map (
            O => \N__26432\,
            I => \eeprom.n3073\
        );

    \I__6045\ : InMux
    port map (
            O => \N__26429\,
            I => \eeprom.n3661\
        );

    \I__6044\ : InMux
    port map (
            O => \N__26426\,
            I => \N__26423\
        );

    \I__6043\ : LocalMux
    port map (
            O => \N__26423\,
            I => \N__26420\
        );

    \I__6042\ : Span4Mux_h
    port map (
            O => \N__26420\,
            I => \N__26415\
        );

    \I__6041\ : InMux
    port map (
            O => \N__26419\,
            I => \N__26410\
        );

    \I__6040\ : InMux
    port map (
            O => \N__26418\,
            I => \N__26410\
        );

    \I__6039\ : Span4Mux_h
    port map (
            O => \N__26415\,
            I => \N__26407\
        );

    \I__6038\ : LocalMux
    port map (
            O => \N__26410\,
            I => \N__26404\
        );

    \I__6037\ : Odrv4
    port map (
            O => \N__26407\,
            I => \eeprom.n3005\
        );

    \I__6036\ : Odrv4
    port map (
            O => \N__26404\,
            I => \eeprom.n3005\
        );

    \I__6035\ : CascadeMux
    port map (
            O => \N__26399\,
            I => \eeprom.n4766_cascade_\
        );

    \I__6034\ : InMux
    port map (
            O => \N__26396\,
            I => \N__26393\
        );

    \I__6033\ : LocalMux
    port map (
            O => \N__26393\,
            I => \eeprom.n4903\
        );

    \I__6032\ : InMux
    port map (
            O => \N__26390\,
            I => \N__26387\
        );

    \I__6031\ : LocalMux
    port map (
            O => \N__26387\,
            I => \N__26382\
        );

    \I__6030\ : InMux
    port map (
            O => \N__26386\,
            I => \N__26379\
        );

    \I__6029\ : InMux
    port map (
            O => \N__26385\,
            I => \N__26376\
        );

    \I__6028\ : Span4Mux_v
    port map (
            O => \N__26382\,
            I => \N__26369\
        );

    \I__6027\ : LocalMux
    port map (
            O => \N__26379\,
            I => \N__26369\
        );

    \I__6026\ : LocalMux
    port map (
            O => \N__26376\,
            I => \N__26369\
        );

    \I__6025\ : Span4Mux_h
    port map (
            O => \N__26369\,
            I => \N__26366\
        );

    \I__6024\ : Span4Mux_h
    port map (
            O => \N__26366\,
            I => \N__26363\
        );

    \I__6023\ : Span4Mux_h
    port map (
            O => \N__26363\,
            I => \N__26360\
        );

    \I__6022\ : Span4Mux_h
    port map (
            O => \N__26360\,
            I => \N__26357\
        );

    \I__6021\ : Odrv4
    port map (
            O => \N__26357\,
            I => \eeprom.n3019\
        );

    \I__6020\ : InMux
    port map (
            O => \N__26354\,
            I => \N__26351\
        );

    \I__6019\ : LocalMux
    port map (
            O => \N__26351\,
            I => \N__26348\
        );

    \I__6018\ : Span4Mux_v
    port map (
            O => \N__26348\,
            I => \N__26345\
        );

    \I__6017\ : Odrv4
    port map (
            O => \N__26345\,
            I => \eeprom.n3086\
        );

    \I__6016\ : InMux
    port map (
            O => \N__26342\,
            I => \bfn_16_23_0_\
        );

    \I__6015\ : InMux
    port map (
            O => \N__26339\,
            I => \N__26336\
        );

    \I__6014\ : LocalMux
    port map (
            O => \N__26336\,
            I => \N__26332\
        );

    \I__6013\ : CascadeMux
    port map (
            O => \N__26335\,
            I => \N__26328\
        );

    \I__6012\ : Span4Mux_h
    port map (
            O => \N__26332\,
            I => \N__26325\
        );

    \I__6011\ : InMux
    port map (
            O => \N__26331\,
            I => \N__26322\
        );

    \I__6010\ : InMux
    port map (
            O => \N__26328\,
            I => \N__26319\
        );

    \I__6009\ : Odrv4
    port map (
            O => \N__26325\,
            I => \eeprom.n3018\
        );

    \I__6008\ : LocalMux
    port map (
            O => \N__26322\,
            I => \eeprom.n3018\
        );

    \I__6007\ : LocalMux
    port map (
            O => \N__26319\,
            I => \eeprom.n3018\
        );

    \I__6006\ : InMux
    port map (
            O => \N__26312\,
            I => \N__26309\
        );

    \I__6005\ : LocalMux
    port map (
            O => \N__26309\,
            I => \N__26306\
        );

    \I__6004\ : Span4Mux_h
    port map (
            O => \N__26306\,
            I => \N__26303\
        );

    \I__6003\ : Odrv4
    port map (
            O => \N__26303\,
            I => \eeprom.n3085\
        );

    \I__6002\ : InMux
    port map (
            O => \N__26300\,
            I => \eeprom.n3649\
        );

    \I__6001\ : CascadeMux
    port map (
            O => \N__26297\,
            I => \N__26294\
        );

    \I__6000\ : InMux
    port map (
            O => \N__26294\,
            I => \N__26290\
        );

    \I__5999\ : InMux
    port map (
            O => \N__26293\,
            I => \N__26287\
        );

    \I__5998\ : LocalMux
    port map (
            O => \N__26290\,
            I => \N__26284\
        );

    \I__5997\ : LocalMux
    port map (
            O => \N__26287\,
            I => \N__26278\
        );

    \I__5996\ : Span4Mux_h
    port map (
            O => \N__26284\,
            I => \N__26278\
        );

    \I__5995\ : InMux
    port map (
            O => \N__26283\,
            I => \N__26275\
        );

    \I__5994\ : Span4Mux_h
    port map (
            O => \N__26278\,
            I => \N__26272\
        );

    \I__5993\ : LocalMux
    port map (
            O => \N__26275\,
            I => \eeprom.n3017\
        );

    \I__5992\ : Odrv4
    port map (
            O => \N__26272\,
            I => \eeprom.n3017\
        );

    \I__5991\ : InMux
    port map (
            O => \N__26267\,
            I => \N__26264\
        );

    \I__5990\ : LocalMux
    port map (
            O => \N__26264\,
            I => \N__26261\
        );

    \I__5989\ : Span4Mux_h
    port map (
            O => \N__26261\,
            I => \N__26258\
        );

    \I__5988\ : Span4Mux_h
    port map (
            O => \N__26258\,
            I => \N__26255\
        );

    \I__5987\ : Odrv4
    port map (
            O => \N__26255\,
            I => \eeprom.n3084\
        );

    \I__5986\ : InMux
    port map (
            O => \N__26252\,
            I => \eeprom.n3650\
        );

    \I__5985\ : CascadeMux
    port map (
            O => \N__26249\,
            I => \N__26246\
        );

    \I__5984\ : InMux
    port map (
            O => \N__26246\,
            I => \N__26241\
        );

    \I__5983\ : InMux
    port map (
            O => \N__26245\,
            I => \N__26238\
        );

    \I__5982\ : InMux
    port map (
            O => \N__26244\,
            I => \N__26235\
        );

    \I__5981\ : LocalMux
    port map (
            O => \N__26241\,
            I => \N__26232\
        );

    \I__5980\ : LocalMux
    port map (
            O => \N__26238\,
            I => \N__26229\
        );

    \I__5979\ : LocalMux
    port map (
            O => \N__26235\,
            I => \N__26224\
        );

    \I__5978\ : Span4Mux_h
    port map (
            O => \N__26232\,
            I => \N__26224\
        );

    \I__5977\ : Span4Mux_h
    port map (
            O => \N__26229\,
            I => \N__26221\
        );

    \I__5976\ : Span4Mux_h
    port map (
            O => \N__26224\,
            I => \N__26218\
        );

    \I__5975\ : Odrv4
    port map (
            O => \N__26221\,
            I => \eeprom.n3016\
        );

    \I__5974\ : Odrv4
    port map (
            O => \N__26218\,
            I => \eeprom.n3016\
        );

    \I__5973\ : CascadeMux
    port map (
            O => \N__26213\,
            I => \N__26210\
        );

    \I__5972\ : InMux
    port map (
            O => \N__26210\,
            I => \N__26207\
        );

    \I__5971\ : LocalMux
    port map (
            O => \N__26207\,
            I => \N__26204\
        );

    \I__5970\ : Span4Mux_h
    port map (
            O => \N__26204\,
            I => \N__26201\
        );

    \I__5969\ : Odrv4
    port map (
            O => \N__26201\,
            I => \eeprom.n3083\
        );

    \I__5968\ : InMux
    port map (
            O => \N__26198\,
            I => \eeprom.n3651\
        );

    \I__5967\ : CascadeMux
    port map (
            O => \N__26195\,
            I => \N__26192\
        );

    \I__5966\ : InMux
    port map (
            O => \N__26192\,
            I => \N__26188\
        );

    \I__5965\ : InMux
    port map (
            O => \N__26191\,
            I => \N__26185\
        );

    \I__5964\ : LocalMux
    port map (
            O => \N__26188\,
            I => \N__26181\
        );

    \I__5963\ : LocalMux
    port map (
            O => \N__26185\,
            I => \N__26178\
        );

    \I__5962\ : InMux
    port map (
            O => \N__26184\,
            I => \N__26175\
        );

    \I__5961\ : Span4Mux_v
    port map (
            O => \N__26181\,
            I => \N__26172\
        );

    \I__5960\ : Odrv4
    port map (
            O => \N__26178\,
            I => \eeprom.n3015\
        );

    \I__5959\ : LocalMux
    port map (
            O => \N__26175\,
            I => \eeprom.n3015\
        );

    \I__5958\ : Odrv4
    port map (
            O => \N__26172\,
            I => \eeprom.n3015\
        );

    \I__5957\ : InMux
    port map (
            O => \N__26165\,
            I => \N__26162\
        );

    \I__5956\ : LocalMux
    port map (
            O => \N__26162\,
            I => \N__26159\
        );

    \I__5955\ : Span4Mux_h
    port map (
            O => \N__26159\,
            I => \N__26156\
        );

    \I__5954\ : Odrv4
    port map (
            O => \N__26156\,
            I => \eeprom.n3082\
        );

    \I__5953\ : InMux
    port map (
            O => \N__26153\,
            I => \eeprom.n3652\
        );

    \I__5952\ : CascadeMux
    port map (
            O => \N__26150\,
            I => \N__26147\
        );

    \I__5951\ : InMux
    port map (
            O => \N__26147\,
            I => \N__26142\
        );

    \I__5950\ : InMux
    port map (
            O => \N__26146\,
            I => \N__26139\
        );

    \I__5949\ : InMux
    port map (
            O => \N__26145\,
            I => \N__26136\
        );

    \I__5948\ : LocalMux
    port map (
            O => \N__26142\,
            I => \N__26133\
        );

    \I__5947\ : LocalMux
    port map (
            O => \N__26139\,
            I => \N__26130\
        );

    \I__5946\ : LocalMux
    port map (
            O => \N__26136\,
            I => \N__26125\
        );

    \I__5945\ : Span4Mux_h
    port map (
            O => \N__26133\,
            I => \N__26125\
        );

    \I__5944\ : Span4Mux_v
    port map (
            O => \N__26130\,
            I => \N__26120\
        );

    \I__5943\ : Span4Mux_h
    port map (
            O => \N__26125\,
            I => \N__26120\
        );

    \I__5942\ : Odrv4
    port map (
            O => \N__26120\,
            I => \eeprom.n3014\
        );

    \I__5941\ : CascadeMux
    port map (
            O => \N__26117\,
            I => \N__26114\
        );

    \I__5940\ : InMux
    port map (
            O => \N__26114\,
            I => \N__26111\
        );

    \I__5939\ : LocalMux
    port map (
            O => \N__26111\,
            I => \N__26108\
        );

    \I__5938\ : Span4Mux_v
    port map (
            O => \N__26108\,
            I => \N__26105\
        );

    \I__5937\ : Span4Mux_h
    port map (
            O => \N__26105\,
            I => \N__26102\
        );

    \I__5936\ : Odrv4
    port map (
            O => \N__26102\,
            I => \eeprom.n3081\
        );

    \I__5935\ : InMux
    port map (
            O => \N__26099\,
            I => \eeprom.n3653\
        );

    \I__5934\ : CascadeMux
    port map (
            O => \N__26096\,
            I => \N__26093\
        );

    \I__5933\ : InMux
    port map (
            O => \N__26093\,
            I => \N__26089\
        );

    \I__5932\ : CascadeMux
    port map (
            O => \N__26092\,
            I => \N__26085\
        );

    \I__5931\ : LocalMux
    port map (
            O => \N__26089\,
            I => \N__26082\
        );

    \I__5930\ : InMux
    port map (
            O => \N__26088\,
            I => \N__26077\
        );

    \I__5929\ : InMux
    port map (
            O => \N__26085\,
            I => \N__26077\
        );

    \I__5928\ : Span4Mux_h
    port map (
            O => \N__26082\,
            I => \N__26074\
        );

    \I__5927\ : LocalMux
    port map (
            O => \N__26077\,
            I => \eeprom.n3013\
        );

    \I__5926\ : Odrv4
    port map (
            O => \N__26074\,
            I => \eeprom.n3013\
        );

    \I__5925\ : InMux
    port map (
            O => \N__26069\,
            I => \N__26066\
        );

    \I__5924\ : LocalMux
    port map (
            O => \N__26066\,
            I => \N__26063\
        );

    \I__5923\ : Odrv4
    port map (
            O => \N__26063\,
            I => \eeprom.n3080\
        );

    \I__5922\ : InMux
    port map (
            O => \N__26060\,
            I => \eeprom.n3654\
        );

    \I__5921\ : InMux
    port map (
            O => \N__26057\,
            I => \N__26052\
        );

    \I__5920\ : CascadeMux
    port map (
            O => \N__26056\,
            I => \N__26049\
        );

    \I__5919\ : InMux
    port map (
            O => \N__26055\,
            I => \N__26046\
        );

    \I__5918\ : LocalMux
    port map (
            O => \N__26052\,
            I => \N__26043\
        );

    \I__5917\ : InMux
    port map (
            O => \N__26049\,
            I => \N__26040\
        );

    \I__5916\ : LocalMux
    port map (
            O => \N__26046\,
            I => \eeprom.n3613_adj_342\
        );

    \I__5915\ : Odrv4
    port map (
            O => \N__26043\,
            I => \eeprom.n3613_adj_342\
        );

    \I__5914\ : LocalMux
    port map (
            O => \N__26040\,
            I => \eeprom.n3613_adj_342\
        );

    \I__5913\ : CascadeMux
    port map (
            O => \N__26033\,
            I => \N__26030\
        );

    \I__5912\ : InMux
    port map (
            O => \N__26030\,
            I => \N__26027\
        );

    \I__5911\ : LocalMux
    port map (
            O => \N__26027\,
            I => \N__26024\
        );

    \I__5910\ : Odrv4
    port map (
            O => \N__26024\,
            I => \eeprom.n1347\
        );

    \I__5909\ : InMux
    port map (
            O => \N__26021\,
            I => \eeprom.n3515\
        );

    \I__5908\ : InMux
    port map (
            O => \N__26018\,
            I => \N__26015\
        );

    \I__5907\ : LocalMux
    port map (
            O => \N__26015\,
            I => \N__26011\
        );

    \I__5906\ : InMux
    port map (
            O => \N__26014\,
            I => \N__26008\
        );

    \I__5905\ : Odrv4
    port map (
            O => \N__26011\,
            I => \eeprom.n3612_adj_339\
        );

    \I__5904\ : LocalMux
    port map (
            O => \N__26008\,
            I => \eeprom.n3612_adj_339\
        );

    \I__5903\ : InMux
    port map (
            O => \N__26003\,
            I => \eeprom.n3516\
        );

    \I__5902\ : InMux
    port map (
            O => \N__26000\,
            I => \N__25997\
        );

    \I__5901\ : LocalMux
    port map (
            O => \N__25997\,
            I => \eeprom.n1350\
        );

    \I__5900\ : InMux
    port map (
            O => \N__25994\,
            I => \N__25990\
        );

    \I__5899\ : CascadeMux
    port map (
            O => \N__25993\,
            I => \N__25987\
        );

    \I__5898\ : LocalMux
    port map (
            O => \N__25990\,
            I => \N__25984\
        );

    \I__5897\ : InMux
    port map (
            O => \N__25987\,
            I => \N__25981\
        );

    \I__5896\ : Span4Mux_v
    port map (
            O => \N__25984\,
            I => \N__25975\
        );

    \I__5895\ : LocalMux
    port map (
            O => \N__25981\,
            I => \N__25975\
        );

    \I__5894\ : InMux
    port map (
            O => \N__25980\,
            I => \N__25972\
        );

    \I__5893\ : Odrv4
    port map (
            O => \N__25975\,
            I => \eeprom.n3616_adj_345\
        );

    \I__5892\ : LocalMux
    port map (
            O => \N__25972\,
            I => \eeprom.n3616_adj_345\
        );

    \I__5891\ : InMux
    port map (
            O => \N__25967\,
            I => \N__25964\
        );

    \I__5890\ : LocalMux
    port map (
            O => \N__25964\,
            I => \eeprom.n3715_adj_441\
        );

    \I__5889\ : CascadeMux
    port map (
            O => \N__25961\,
            I => \eeprom.n3715_adj_441_cascade_\
        );

    \I__5888\ : InMux
    port map (
            O => \N__25958\,
            I => \N__25955\
        );

    \I__5887\ : LocalMux
    port map (
            O => \N__25955\,
            I => \eeprom.n4912\
        );

    \I__5886\ : InMux
    port map (
            O => \N__25952\,
            I => \N__25949\
        );

    \I__5885\ : LocalMux
    port map (
            O => \N__25949\,
            I => \N__25945\
        );

    \I__5884\ : InMux
    port map (
            O => \N__25948\,
            I => \N__25942\
        );

    \I__5883\ : Span4Mux_h
    port map (
            O => \N__25945\,
            I => \N__25939\
        );

    \I__5882\ : LocalMux
    port map (
            O => \N__25942\,
            I => \eeprom.n1346\
        );

    \I__5881\ : Odrv4
    port map (
            O => \N__25939\,
            I => \eeprom.n1346\
        );

    \I__5880\ : CascadeMux
    port map (
            O => \N__25934\,
            I => \N__25931\
        );

    \I__5879\ : InMux
    port map (
            O => \N__25931\,
            I => \N__25928\
        );

    \I__5878\ : LocalMux
    port map (
            O => \N__25928\,
            I => \eeprom.n3711_adj_456\
        );

    \I__5877\ : InMux
    port map (
            O => \N__25925\,
            I => \N__25922\
        );

    \I__5876\ : LocalMux
    port map (
            O => \N__25922\,
            I => \eeprom.n1352\
        );

    \I__5875\ : CascadeMux
    port map (
            O => \N__25919\,
            I => \N__25916\
        );

    \I__5874\ : InMux
    port map (
            O => \N__25916\,
            I => \N__25913\
        );

    \I__5873\ : LocalMux
    port map (
            O => \N__25913\,
            I => \N__25909\
        );

    \I__5872\ : InMux
    port map (
            O => \N__25912\,
            I => \N__25906\
        );

    \I__5871\ : Odrv4
    port map (
            O => \N__25909\,
            I => \eeprom.n3618_adj_350\
        );

    \I__5870\ : LocalMux
    port map (
            O => \N__25906\,
            I => \eeprom.n3618_adj_350\
        );

    \I__5869\ : CascadeMux
    port map (
            O => \N__25901\,
            I => \N__25898\
        );

    \I__5868\ : InMux
    port map (
            O => \N__25898\,
            I => \N__25895\
        );

    \I__5867\ : LocalMux
    port map (
            O => \N__25895\,
            I => \eeprom.n3717_adj_438\
        );

    \I__5866\ : CascadeMux
    port map (
            O => \N__25892\,
            I => \eeprom.n3717_adj_438_cascade_\
        );

    \I__5865\ : InMux
    port map (
            O => \N__25889\,
            I => \N__25886\
        );

    \I__5864\ : LocalMux
    port map (
            O => \N__25886\,
            I => \eeprom.n4906\
        );

    \I__5863\ : InMux
    port map (
            O => \N__25883\,
            I => \N__25880\
        );

    \I__5862\ : LocalMux
    port map (
            O => \N__25880\,
            I => \eeprom.n1353\
        );

    \I__5861\ : InMux
    port map (
            O => \N__25877\,
            I => \N__25872\
        );

    \I__5860\ : InMux
    port map (
            O => \N__25876\,
            I => \N__25869\
        );

    \I__5859\ : InMux
    port map (
            O => \N__25875\,
            I => \N__25866\
        );

    \I__5858\ : LocalMux
    port map (
            O => \N__25872\,
            I => \N__25863\
        );

    \I__5857\ : LocalMux
    port map (
            O => \N__25869\,
            I => \N__25860\
        );

    \I__5856\ : LocalMux
    port map (
            O => \N__25866\,
            I => \N__25857\
        );

    \I__5855\ : Span4Mux_h
    port map (
            O => \N__25863\,
            I => \N__25852\
        );

    \I__5854\ : Span4Mux_v
    port map (
            O => \N__25860\,
            I => \N__25852\
        );

    \I__5853\ : Span12Mux_v
    port map (
            O => \N__25857\,
            I => \N__25849\
        );

    \I__5852\ : Span4Mux_h
    port map (
            O => \N__25852\,
            I => \N__25846\
        );

    \I__5851\ : Span12Mux_h
    port map (
            O => \N__25849\,
            I => \N__25843\
        );

    \I__5850\ : Span4Mux_h
    port map (
            O => \N__25846\,
            I => \N__25840\
        );

    \I__5849\ : Odrv12
    port map (
            O => \N__25843\,
            I => \eeprom.n3619_adj_352\
        );

    \I__5848\ : Odrv4
    port map (
            O => \N__25840\,
            I => \eeprom.n3619_adj_352\
        );

    \I__5847\ : CascadeMux
    port map (
            O => \N__25835\,
            I => \N__25829\
        );

    \I__5846\ : CascadeMux
    port map (
            O => \N__25834\,
            I => \N__25826\
        );

    \I__5845\ : InMux
    port map (
            O => \N__25833\,
            I => \N__25821\
        );

    \I__5844\ : CascadeMux
    port map (
            O => \N__25832\,
            I => \N__25818\
        );

    \I__5843\ : InMux
    port map (
            O => \N__25829\,
            I => \N__25807\
        );

    \I__5842\ : InMux
    port map (
            O => \N__25826\,
            I => \N__25807\
        );

    \I__5841\ : InMux
    port map (
            O => \N__25825\,
            I => \N__25807\
        );

    \I__5840\ : InMux
    port map (
            O => \N__25824\,
            I => \N__25807\
        );

    \I__5839\ : LocalMux
    port map (
            O => \N__25821\,
            I => \N__25804\
        );

    \I__5838\ : InMux
    port map (
            O => \N__25818\,
            I => \N__25799\
        );

    \I__5837\ : InMux
    port map (
            O => \N__25817\,
            I => \N__25799\
        );

    \I__5836\ : InMux
    port map (
            O => \N__25816\,
            I => \N__25796\
        );

    \I__5835\ : LocalMux
    port map (
            O => \N__25807\,
            I => \N__25793\
        );

    \I__5834\ : Odrv4
    port map (
            O => \N__25804\,
            I => \eeprom.n3628_adj_437\
        );

    \I__5833\ : LocalMux
    port map (
            O => \N__25799\,
            I => \eeprom.n3628_adj_437\
        );

    \I__5832\ : LocalMux
    port map (
            O => \N__25796\,
            I => \eeprom.n3628_adj_437\
        );

    \I__5831\ : Odrv4
    port map (
            O => \N__25793\,
            I => \eeprom.n3628_adj_437\
        );

    \I__5830\ : CascadeMux
    port map (
            O => \N__25784\,
            I => \N__25781\
        );

    \I__5829\ : InMux
    port map (
            O => \N__25781\,
            I => \N__25778\
        );

    \I__5828\ : LocalMux
    port map (
            O => \N__25778\,
            I => \eeprom.n4766\
        );

    \I__5827\ : InMux
    port map (
            O => \N__25775\,
            I => \N__25772\
        );

    \I__5826\ : LocalMux
    port map (
            O => \N__25772\,
            I => \eeprom.n3565_adj_338\
        );

    \I__5825\ : InMux
    port map (
            O => \N__25769\,
            I => \eeprom.n3769\
        );

    \I__5824\ : CascadeMux
    port map (
            O => \N__25766\,
            I => \N__25763\
        );

    \I__5823\ : InMux
    port map (
            O => \N__25763\,
            I => \N__25759\
        );

    \I__5822\ : InMux
    port map (
            O => \N__25762\,
            I => \N__25756\
        );

    \I__5821\ : LocalMux
    port map (
            O => \N__25759\,
            I => \N__25753\
        );

    \I__5820\ : LocalMux
    port map (
            O => \N__25756\,
            I => \N__25750\
        );

    \I__5819\ : Span4Mux_h
    port map (
            O => \N__25753\,
            I => \N__25747\
        );

    \I__5818\ : Span4Mux_h
    port map (
            O => \N__25750\,
            I => \N__25744\
        );

    \I__5817\ : Odrv4
    port map (
            O => \N__25747\,
            I => \eeprom.n3497\
        );

    \I__5816\ : Odrv4
    port map (
            O => \N__25744\,
            I => \eeprom.n3497\
        );

    \I__5815\ : InMux
    port map (
            O => \N__25739\,
            I => \N__25736\
        );

    \I__5814\ : LocalMux
    port map (
            O => \N__25736\,
            I => \N__25733\
        );

    \I__5813\ : Span4Mux_h
    port map (
            O => \N__25733\,
            I => \N__25730\
        );

    \I__5812\ : Odrv4
    port map (
            O => \N__25730\,
            I => \eeprom.n3564_adj_337\
        );

    \I__5811\ : InMux
    port map (
            O => \N__25727\,
            I => \eeprom.n3770\
        );

    \I__5810\ : InMux
    port map (
            O => \N__25724\,
            I => \N__25720\
        );

    \I__5809\ : InMux
    port map (
            O => \N__25723\,
            I => \N__25717\
        );

    \I__5808\ : LocalMux
    port map (
            O => \N__25720\,
            I => \N__25714\
        );

    \I__5807\ : LocalMux
    port map (
            O => \N__25717\,
            I => \N__25711\
        );

    \I__5806\ : Odrv4
    port map (
            O => \N__25714\,
            I => \eeprom.n3496\
        );

    \I__5805\ : Odrv4
    port map (
            O => \N__25711\,
            I => \eeprom.n3496\
        );

    \I__5804\ : CascadeMux
    port map (
            O => \N__25706\,
            I => \N__25700\
        );

    \I__5803\ : CascadeMux
    port map (
            O => \N__25705\,
            I => \N__25697\
        );

    \I__5802\ : CascadeMux
    port map (
            O => \N__25704\,
            I => \N__25693\
        );

    \I__5801\ : CascadeMux
    port map (
            O => \N__25703\,
            I => \N__25690\
        );

    \I__5800\ : InMux
    port map (
            O => \N__25700\,
            I => \N__25686\
        );

    \I__5799\ : InMux
    port map (
            O => \N__25697\,
            I => \N__25673\
        );

    \I__5798\ : InMux
    port map (
            O => \N__25696\,
            I => \N__25673\
        );

    \I__5797\ : InMux
    port map (
            O => \N__25693\,
            I => \N__25665\
        );

    \I__5796\ : InMux
    port map (
            O => \N__25690\,
            I => \N__25665\
        );

    \I__5795\ : InMux
    port map (
            O => \N__25689\,
            I => \N__25665\
        );

    \I__5794\ : LocalMux
    port map (
            O => \N__25686\,
            I => \N__25656\
        );

    \I__5793\ : InMux
    port map (
            O => \N__25685\,
            I => \N__25649\
        );

    \I__5792\ : InMux
    port map (
            O => \N__25684\,
            I => \N__25649\
        );

    \I__5791\ : InMux
    port map (
            O => \N__25683\,
            I => \N__25649\
        );

    \I__5790\ : InMux
    port map (
            O => \N__25682\,
            I => \N__25642\
        );

    \I__5789\ : InMux
    port map (
            O => \N__25681\,
            I => \N__25642\
        );

    \I__5788\ : InMux
    port map (
            O => \N__25680\,
            I => \N__25642\
        );

    \I__5787\ : InMux
    port map (
            O => \N__25679\,
            I => \N__25637\
        );

    \I__5786\ : InMux
    port map (
            O => \N__25678\,
            I => \N__25637\
        );

    \I__5785\ : LocalMux
    port map (
            O => \N__25673\,
            I => \N__25634\
        );

    \I__5784\ : CascadeMux
    port map (
            O => \N__25672\,
            I => \N__25629\
        );

    \I__5783\ : LocalMux
    port map (
            O => \N__25665\,
            I => \N__25625\
        );

    \I__5782\ : InMux
    port map (
            O => \N__25664\,
            I => \N__25616\
        );

    \I__5781\ : InMux
    port map (
            O => \N__25663\,
            I => \N__25616\
        );

    \I__5780\ : InMux
    port map (
            O => \N__25662\,
            I => \N__25616\
        );

    \I__5779\ : InMux
    port map (
            O => \N__25661\,
            I => \N__25616\
        );

    \I__5778\ : InMux
    port map (
            O => \N__25660\,
            I => \N__25613\
        );

    \I__5777\ : InMux
    port map (
            O => \N__25659\,
            I => \N__25610\
        );

    \I__5776\ : Span4Mux_h
    port map (
            O => \N__25656\,
            I => \N__25599\
        );

    \I__5775\ : LocalMux
    port map (
            O => \N__25649\,
            I => \N__25599\
        );

    \I__5774\ : LocalMux
    port map (
            O => \N__25642\,
            I => \N__25599\
        );

    \I__5773\ : LocalMux
    port map (
            O => \N__25637\,
            I => \N__25599\
        );

    \I__5772\ : Span4Mux_v
    port map (
            O => \N__25634\,
            I => \N__25599\
        );

    \I__5771\ : InMux
    port map (
            O => \N__25633\,
            I => \N__25590\
        );

    \I__5770\ : InMux
    port map (
            O => \N__25632\,
            I => \N__25590\
        );

    \I__5769\ : InMux
    port map (
            O => \N__25629\,
            I => \N__25590\
        );

    \I__5768\ : InMux
    port map (
            O => \N__25628\,
            I => \N__25590\
        );

    \I__5767\ : Span4Mux_h
    port map (
            O => \N__25625\,
            I => \N__25587\
        );

    \I__5766\ : LocalMux
    port map (
            O => \N__25616\,
            I => \eeprom.n3529_adj_336\
        );

    \I__5765\ : LocalMux
    port map (
            O => \N__25613\,
            I => \eeprom.n3529_adj_336\
        );

    \I__5764\ : LocalMux
    port map (
            O => \N__25610\,
            I => \eeprom.n3529_adj_336\
        );

    \I__5763\ : Odrv4
    port map (
            O => \N__25599\,
            I => \eeprom.n3529_adj_336\
        );

    \I__5762\ : LocalMux
    port map (
            O => \N__25590\,
            I => \eeprom.n3529_adj_336\
        );

    \I__5761\ : Odrv4
    port map (
            O => \N__25587\,
            I => \eeprom.n3529_adj_336\
        );

    \I__5760\ : InMux
    port map (
            O => \N__25574\,
            I => \eeprom.n3771\
        );

    \I__5759\ : InMux
    port map (
            O => \N__25571\,
            I => \N__25568\
        );

    \I__5758\ : LocalMux
    port map (
            O => \N__25568\,
            I => \eeprom.n4765\
        );

    \I__5757\ : InMux
    port map (
            O => \N__25565\,
            I => \bfn_16_20_0_\
        );

    \I__5756\ : InMux
    port map (
            O => \N__25562\,
            I => \eeprom.n3510\
        );

    \I__5755\ : InMux
    port map (
            O => \N__25559\,
            I => \N__25555\
        );

    \I__5754\ : InMux
    port map (
            O => \N__25558\,
            I => \N__25552\
        );

    \I__5753\ : LocalMux
    port map (
            O => \N__25555\,
            I => \N__25549\
        );

    \I__5752\ : LocalMux
    port map (
            O => \N__25552\,
            I => \eeprom.n3617_adj_346\
        );

    \I__5751\ : Odrv4
    port map (
            O => \N__25549\,
            I => \eeprom.n3617_adj_346\
        );

    \I__5750\ : InMux
    port map (
            O => \N__25544\,
            I => \N__25541\
        );

    \I__5749\ : LocalMux
    port map (
            O => \N__25541\,
            I => \eeprom.n1351\
        );

    \I__5748\ : InMux
    port map (
            O => \N__25538\,
            I => \eeprom.n3511\
        );

    \I__5747\ : InMux
    port map (
            O => \N__25535\,
            I => \eeprom.n3512\
        );

    \I__5746\ : CascadeMux
    port map (
            O => \N__25532\,
            I => \N__25529\
        );

    \I__5745\ : InMux
    port map (
            O => \N__25529\,
            I => \N__25526\
        );

    \I__5744\ : LocalMux
    port map (
            O => \N__25526\,
            I => \N__25522\
        );

    \I__5743\ : InMux
    port map (
            O => \N__25525\,
            I => \N__25519\
        );

    \I__5742\ : Odrv4
    port map (
            O => \N__25522\,
            I => \eeprom.n3615_adj_344\
        );

    \I__5741\ : LocalMux
    port map (
            O => \N__25519\,
            I => \eeprom.n3615_adj_344\
        );

    \I__5740\ : InMux
    port map (
            O => \N__25514\,
            I => \N__25511\
        );

    \I__5739\ : LocalMux
    port map (
            O => \N__25511\,
            I => \N__25508\
        );

    \I__5738\ : Odrv4
    port map (
            O => \N__25508\,
            I => \eeprom.n1349\
        );

    \I__5737\ : InMux
    port map (
            O => \N__25505\,
            I => \eeprom.n3513\
        );

    \I__5736\ : InMux
    port map (
            O => \N__25502\,
            I => \N__25498\
        );

    \I__5735\ : InMux
    port map (
            O => \N__25501\,
            I => \N__25495\
        );

    \I__5734\ : LocalMux
    port map (
            O => \N__25498\,
            I => \N__25491\
        );

    \I__5733\ : LocalMux
    port map (
            O => \N__25495\,
            I => \N__25488\
        );

    \I__5732\ : InMux
    port map (
            O => \N__25494\,
            I => \N__25485\
        );

    \I__5731\ : Odrv4
    port map (
            O => \N__25491\,
            I => \eeprom.n3614_adj_343\
        );

    \I__5730\ : Odrv4
    port map (
            O => \N__25488\,
            I => \eeprom.n3614_adj_343\
        );

    \I__5729\ : LocalMux
    port map (
            O => \N__25485\,
            I => \eeprom.n3614_adj_343\
        );

    \I__5728\ : InMux
    port map (
            O => \N__25478\,
            I => \N__25475\
        );

    \I__5727\ : LocalMux
    port map (
            O => \N__25475\,
            I => \N__25472\
        );

    \I__5726\ : Odrv4
    port map (
            O => \N__25472\,
            I => \eeprom.n1348\
        );

    \I__5725\ : InMux
    port map (
            O => \N__25469\,
            I => \eeprom.n3514\
        );

    \I__5724\ : InMux
    port map (
            O => \N__25466\,
            I => \N__25463\
        );

    \I__5723\ : LocalMux
    port map (
            O => \N__25463\,
            I => \N__25459\
        );

    \I__5722\ : InMux
    port map (
            O => \N__25462\,
            I => \N__25456\
        );

    \I__5721\ : Span4Mux_h
    port map (
            O => \N__25459\,
            I => \N__25453\
        );

    \I__5720\ : LocalMux
    port map (
            O => \N__25456\,
            I => \N__25450\
        );

    \I__5719\ : Odrv4
    port map (
            O => \N__25453\,
            I => \eeprom.n3505\
        );

    \I__5718\ : Odrv12
    port map (
            O => \N__25450\,
            I => \eeprom.n3505\
        );

    \I__5717\ : InMux
    port map (
            O => \N__25445\,
            I => \N__25442\
        );

    \I__5716\ : LocalMux
    port map (
            O => \N__25442\,
            I => \N__25439\
        );

    \I__5715\ : Span4Mux_h
    port map (
            O => \N__25439\,
            I => \N__25436\
        );

    \I__5714\ : Odrv4
    port map (
            O => \N__25436\,
            I => \eeprom.n3572_adj_354\
        );

    \I__5713\ : InMux
    port map (
            O => \N__25433\,
            I => \eeprom.n3762\
        );

    \I__5712\ : InMux
    port map (
            O => \N__25430\,
            I => \N__25426\
        );

    \I__5711\ : InMux
    port map (
            O => \N__25429\,
            I => \N__25422\
        );

    \I__5710\ : LocalMux
    port map (
            O => \N__25426\,
            I => \N__25419\
        );

    \I__5709\ : InMux
    port map (
            O => \N__25425\,
            I => \N__25416\
        );

    \I__5708\ : LocalMux
    port map (
            O => \N__25422\,
            I => \eeprom.n3504\
        );

    \I__5707\ : Odrv4
    port map (
            O => \N__25419\,
            I => \eeprom.n3504\
        );

    \I__5706\ : LocalMux
    port map (
            O => \N__25416\,
            I => \eeprom.n3504\
        );

    \I__5705\ : InMux
    port map (
            O => \N__25409\,
            I => \N__25406\
        );

    \I__5704\ : LocalMux
    port map (
            O => \N__25406\,
            I => \N__25403\
        );

    \I__5703\ : Span4Mux_h
    port map (
            O => \N__25403\,
            I => \N__25400\
        );

    \I__5702\ : Odrv4
    port map (
            O => \N__25400\,
            I => \eeprom.n3571_adj_353\
        );

    \I__5701\ : InMux
    port map (
            O => \N__25397\,
            I => \eeprom.n3763\
        );

    \I__5700\ : InMux
    port map (
            O => \N__25394\,
            I => \N__25390\
        );

    \I__5699\ : InMux
    port map (
            O => \N__25393\,
            I => \N__25386\
        );

    \I__5698\ : LocalMux
    port map (
            O => \N__25390\,
            I => \N__25383\
        );

    \I__5697\ : CascadeMux
    port map (
            O => \N__25389\,
            I => \N__25380\
        );

    \I__5696\ : LocalMux
    port map (
            O => \N__25386\,
            I => \N__25377\
        );

    \I__5695\ : Span4Mux_h
    port map (
            O => \N__25383\,
            I => \N__25374\
        );

    \I__5694\ : InMux
    port map (
            O => \N__25380\,
            I => \N__25371\
        );

    \I__5693\ : Span4Mux_h
    port map (
            O => \N__25377\,
            I => \N__25368\
        );

    \I__5692\ : Odrv4
    port map (
            O => \N__25374\,
            I => \eeprom.n3503\
        );

    \I__5691\ : LocalMux
    port map (
            O => \N__25371\,
            I => \eeprom.n3503\
        );

    \I__5690\ : Odrv4
    port map (
            O => \N__25368\,
            I => \eeprom.n3503\
        );

    \I__5689\ : InMux
    port map (
            O => \N__25361\,
            I => \N__25358\
        );

    \I__5688\ : LocalMux
    port map (
            O => \N__25358\,
            I => \N__25355\
        );

    \I__5687\ : Odrv12
    port map (
            O => \N__25355\,
            I => \eeprom.n3570_adj_349\
        );

    \I__5686\ : InMux
    port map (
            O => \N__25352\,
            I => \bfn_16_19_0_\
        );

    \I__5685\ : InMux
    port map (
            O => \N__25349\,
            I => \N__25345\
        );

    \I__5684\ : InMux
    port map (
            O => \N__25348\,
            I => \N__25342\
        );

    \I__5683\ : LocalMux
    port map (
            O => \N__25345\,
            I => \N__25336\
        );

    \I__5682\ : LocalMux
    port map (
            O => \N__25342\,
            I => \N__25336\
        );

    \I__5681\ : InMux
    port map (
            O => \N__25341\,
            I => \N__25333\
        );

    \I__5680\ : Odrv4
    port map (
            O => \N__25336\,
            I => \eeprom.n3502\
        );

    \I__5679\ : LocalMux
    port map (
            O => \N__25333\,
            I => \eeprom.n3502\
        );

    \I__5678\ : CascadeMux
    port map (
            O => \N__25328\,
            I => \N__25325\
        );

    \I__5677\ : InMux
    port map (
            O => \N__25325\,
            I => \N__25322\
        );

    \I__5676\ : LocalMux
    port map (
            O => \N__25322\,
            I => \eeprom.n3569_adj_348\
        );

    \I__5675\ : InMux
    port map (
            O => \N__25319\,
            I => \eeprom.n3765\
        );

    \I__5674\ : InMux
    port map (
            O => \N__25316\,
            I => \N__25313\
        );

    \I__5673\ : LocalMux
    port map (
            O => \N__25313\,
            I => \N__25309\
        );

    \I__5672\ : InMux
    port map (
            O => \N__25312\,
            I => \N__25305\
        );

    \I__5671\ : Span4Mux_h
    port map (
            O => \N__25309\,
            I => \N__25302\
        );

    \I__5670\ : InMux
    port map (
            O => \N__25308\,
            I => \N__25299\
        );

    \I__5669\ : LocalMux
    port map (
            O => \N__25305\,
            I => \eeprom.n3501\
        );

    \I__5668\ : Odrv4
    port map (
            O => \N__25302\,
            I => \eeprom.n3501\
        );

    \I__5667\ : LocalMux
    port map (
            O => \N__25299\,
            I => \eeprom.n3501\
        );

    \I__5666\ : InMux
    port map (
            O => \N__25292\,
            I => \N__25289\
        );

    \I__5665\ : LocalMux
    port map (
            O => \N__25289\,
            I => \N__25286\
        );

    \I__5664\ : Span4Mux_h
    port map (
            O => \N__25286\,
            I => \N__25283\
        );

    \I__5663\ : Odrv4
    port map (
            O => \N__25283\,
            I => \eeprom.n3568_adj_347\
        );

    \I__5662\ : InMux
    port map (
            O => \N__25280\,
            I => \eeprom.n3766\
        );

    \I__5661\ : InMux
    port map (
            O => \N__25277\,
            I => \N__25273\
        );

    \I__5660\ : CascadeMux
    port map (
            O => \N__25276\,
            I => \N__25270\
        );

    \I__5659\ : LocalMux
    port map (
            O => \N__25273\,
            I => \N__25267\
        );

    \I__5658\ : InMux
    port map (
            O => \N__25270\,
            I => \N__25264\
        );

    \I__5657\ : Span4Mux_v
    port map (
            O => \N__25267\,
            I => \N__25261\
        );

    \I__5656\ : LocalMux
    port map (
            O => \N__25264\,
            I => \eeprom.n3500\
        );

    \I__5655\ : Odrv4
    port map (
            O => \N__25261\,
            I => \eeprom.n3500\
        );

    \I__5654\ : InMux
    port map (
            O => \N__25256\,
            I => \N__25253\
        );

    \I__5653\ : LocalMux
    port map (
            O => \N__25253\,
            I => \N__25250\
        );

    \I__5652\ : Span4Mux_h
    port map (
            O => \N__25250\,
            I => \N__25247\
        );

    \I__5651\ : Odrv4
    port map (
            O => \N__25247\,
            I => \eeprom.n3567_adj_341\
        );

    \I__5650\ : InMux
    port map (
            O => \N__25244\,
            I => \eeprom.n3767\
        );

    \I__5649\ : InMux
    port map (
            O => \N__25241\,
            I => \N__25236\
        );

    \I__5648\ : InMux
    port map (
            O => \N__25240\,
            I => \N__25233\
        );

    \I__5647\ : InMux
    port map (
            O => \N__25239\,
            I => \N__25230\
        );

    \I__5646\ : LocalMux
    port map (
            O => \N__25236\,
            I => \N__25227\
        );

    \I__5645\ : LocalMux
    port map (
            O => \N__25233\,
            I => \N__25224\
        );

    \I__5644\ : LocalMux
    port map (
            O => \N__25230\,
            I => \eeprom.n3499\
        );

    \I__5643\ : Odrv12
    port map (
            O => \N__25227\,
            I => \eeprom.n3499\
        );

    \I__5642\ : Odrv4
    port map (
            O => \N__25224\,
            I => \eeprom.n3499\
        );

    \I__5641\ : CascadeMux
    port map (
            O => \N__25217\,
            I => \N__25214\
        );

    \I__5640\ : InMux
    port map (
            O => \N__25214\,
            I => \N__25211\
        );

    \I__5639\ : LocalMux
    port map (
            O => \N__25211\,
            I => \N__25208\
        );

    \I__5638\ : Span4Mux_v
    port map (
            O => \N__25208\,
            I => \N__25205\
        );

    \I__5637\ : Odrv4
    port map (
            O => \N__25205\,
            I => \eeprom.n3566_adj_340\
        );

    \I__5636\ : InMux
    port map (
            O => \N__25202\,
            I => \eeprom.n3768\
        );

    \I__5635\ : InMux
    port map (
            O => \N__25199\,
            I => \N__25195\
        );

    \I__5634\ : InMux
    port map (
            O => \N__25198\,
            I => \N__25192\
        );

    \I__5633\ : LocalMux
    port map (
            O => \N__25195\,
            I => \N__25187\
        );

    \I__5632\ : LocalMux
    port map (
            O => \N__25192\,
            I => \N__25187\
        );

    \I__5631\ : Span4Mux_h
    port map (
            O => \N__25187\,
            I => \N__25183\
        );

    \I__5630\ : InMux
    port map (
            O => \N__25186\,
            I => \N__25180\
        );

    \I__5629\ : Odrv4
    port map (
            O => \N__25183\,
            I => \eeprom.n3498\
        );

    \I__5628\ : LocalMux
    port map (
            O => \N__25180\,
            I => \eeprom.n3498\
        );

    \I__5627\ : CascadeMux
    port map (
            O => \N__25175\,
            I => \N__25171\
        );

    \I__5626\ : CascadeMux
    port map (
            O => \N__25174\,
            I => \N__25168\
        );

    \I__5625\ : InMux
    port map (
            O => \N__25171\,
            I => \N__25165\
        );

    \I__5624\ : InMux
    port map (
            O => \N__25168\,
            I => \N__25162\
        );

    \I__5623\ : LocalMux
    port map (
            O => \N__25165\,
            I => \N__25158\
        );

    \I__5622\ : LocalMux
    port map (
            O => \N__25162\,
            I => \N__25155\
        );

    \I__5621\ : InMux
    port map (
            O => \N__25161\,
            I => \N__25152\
        );

    \I__5620\ : Span4Mux_v
    port map (
            O => \N__25158\,
            I => \N__25149\
        );

    \I__5619\ : Span4Mux_h
    port map (
            O => \N__25155\,
            I => \N__25144\
        );

    \I__5618\ : LocalMux
    port map (
            O => \N__25152\,
            I => \N__25144\
        );

    \I__5617\ : Odrv4
    port map (
            O => \N__25149\,
            I => \eeprom.n3513_adj_366\
        );

    \I__5616\ : Odrv4
    port map (
            O => \N__25144\,
            I => \eeprom.n3513_adj_366\
        );

    \I__5615\ : InMux
    port map (
            O => \N__25139\,
            I => \N__25136\
        );

    \I__5614\ : LocalMux
    port map (
            O => \N__25136\,
            I => \N__25133\
        );

    \I__5613\ : Span4Mux_v
    port map (
            O => \N__25133\,
            I => \N__25130\
        );

    \I__5612\ : Odrv4
    port map (
            O => \N__25130\,
            I => \eeprom.n3580_adj_365\
        );

    \I__5611\ : InMux
    port map (
            O => \N__25127\,
            I => \eeprom.n3754\
        );

    \I__5610\ : CascadeMux
    port map (
            O => \N__25124\,
            I => \N__25120\
        );

    \I__5609\ : InMux
    port map (
            O => \N__25123\,
            I => \N__25117\
        );

    \I__5608\ : InMux
    port map (
            O => \N__25120\,
            I => \N__25114\
        );

    \I__5607\ : LocalMux
    port map (
            O => \N__25117\,
            I => \N__25110\
        );

    \I__5606\ : LocalMux
    port map (
            O => \N__25114\,
            I => \N__25107\
        );

    \I__5605\ : InMux
    port map (
            O => \N__25113\,
            I => \N__25104\
        );

    \I__5604\ : Odrv4
    port map (
            O => \N__25110\,
            I => \eeprom.n3512_adj_364\
        );

    \I__5603\ : Odrv4
    port map (
            O => \N__25107\,
            I => \eeprom.n3512_adj_364\
        );

    \I__5602\ : LocalMux
    port map (
            O => \N__25104\,
            I => \eeprom.n3512_adj_364\
        );

    \I__5601\ : CascadeMux
    port map (
            O => \N__25097\,
            I => \N__25094\
        );

    \I__5600\ : InMux
    port map (
            O => \N__25094\,
            I => \N__25091\
        );

    \I__5599\ : LocalMux
    port map (
            O => \N__25091\,
            I => \N__25088\
        );

    \I__5598\ : Span4Mux_h
    port map (
            O => \N__25088\,
            I => \N__25085\
        );

    \I__5597\ : Odrv4
    port map (
            O => \N__25085\,
            I => \eeprom.n3579_adj_363\
        );

    \I__5596\ : InMux
    port map (
            O => \N__25082\,
            I => \eeprom.n3755\
        );

    \I__5595\ : CascadeMux
    port map (
            O => \N__25079\,
            I => \N__25076\
        );

    \I__5594\ : InMux
    port map (
            O => \N__25076\,
            I => \N__25073\
        );

    \I__5593\ : LocalMux
    port map (
            O => \N__25073\,
            I => \N__25068\
        );

    \I__5592\ : InMux
    port map (
            O => \N__25072\,
            I => \N__25065\
        );

    \I__5591\ : InMux
    port map (
            O => \N__25071\,
            I => \N__25062\
        );

    \I__5590\ : Span4Mux_h
    port map (
            O => \N__25068\,
            I => \N__25059\
        );

    \I__5589\ : LocalMux
    port map (
            O => \N__25065\,
            I => \eeprom.n3511_adj_362\
        );

    \I__5588\ : LocalMux
    port map (
            O => \N__25062\,
            I => \eeprom.n3511_adj_362\
        );

    \I__5587\ : Odrv4
    port map (
            O => \N__25059\,
            I => \eeprom.n3511_adj_362\
        );

    \I__5586\ : InMux
    port map (
            O => \N__25052\,
            I => \N__25049\
        );

    \I__5585\ : LocalMux
    port map (
            O => \N__25049\,
            I => \N__25046\
        );

    \I__5584\ : Span4Mux_h
    port map (
            O => \N__25046\,
            I => \N__25043\
        );

    \I__5583\ : Odrv4
    port map (
            O => \N__25043\,
            I => \eeprom.n3578_adj_361\
        );

    \I__5582\ : InMux
    port map (
            O => \N__25040\,
            I => \bfn_16_18_0_\
        );

    \I__5581\ : CascadeMux
    port map (
            O => \N__25037\,
            I => \N__25034\
        );

    \I__5580\ : InMux
    port map (
            O => \N__25034\,
            I => \N__25030\
        );

    \I__5579\ : CascadeMux
    port map (
            O => \N__25033\,
            I => \N__25027\
        );

    \I__5578\ : LocalMux
    port map (
            O => \N__25030\,
            I => \N__25023\
        );

    \I__5577\ : InMux
    port map (
            O => \N__25027\,
            I => \N__25018\
        );

    \I__5576\ : InMux
    port map (
            O => \N__25026\,
            I => \N__25018\
        );

    \I__5575\ : Odrv4
    port map (
            O => \N__25023\,
            I => \eeprom.n3510_adj_360\
        );

    \I__5574\ : LocalMux
    port map (
            O => \N__25018\,
            I => \eeprom.n3510_adj_360\
        );

    \I__5573\ : InMux
    port map (
            O => \N__25013\,
            I => \N__25010\
        );

    \I__5572\ : LocalMux
    port map (
            O => \N__25010\,
            I => \N__25007\
        );

    \I__5571\ : Span4Mux_h
    port map (
            O => \N__25007\,
            I => \N__25004\
        );

    \I__5570\ : Odrv4
    port map (
            O => \N__25004\,
            I => \eeprom.n3577_adj_359\
        );

    \I__5569\ : InMux
    port map (
            O => \N__25001\,
            I => \eeprom.n3757\
        );

    \I__5568\ : CascadeMux
    port map (
            O => \N__24998\,
            I => \N__24995\
        );

    \I__5567\ : InMux
    port map (
            O => \N__24995\,
            I => \N__24991\
        );

    \I__5566\ : CascadeMux
    port map (
            O => \N__24994\,
            I => \N__24988\
        );

    \I__5565\ : LocalMux
    port map (
            O => \N__24991\,
            I => \N__24985\
        );

    \I__5564\ : InMux
    port map (
            O => \N__24988\,
            I => \N__24981\
        );

    \I__5563\ : Span4Mux_h
    port map (
            O => \N__24985\,
            I => \N__24978\
        );

    \I__5562\ : InMux
    port map (
            O => \N__24984\,
            I => \N__24975\
        );

    \I__5561\ : LocalMux
    port map (
            O => \N__24981\,
            I => \eeprom.n3509\
        );

    \I__5560\ : Odrv4
    port map (
            O => \N__24978\,
            I => \eeprom.n3509\
        );

    \I__5559\ : LocalMux
    port map (
            O => \N__24975\,
            I => \eeprom.n3509\
        );

    \I__5558\ : InMux
    port map (
            O => \N__24968\,
            I => \N__24965\
        );

    \I__5557\ : LocalMux
    port map (
            O => \N__24965\,
            I => \N__24962\
        );

    \I__5556\ : Span4Mux_h
    port map (
            O => \N__24962\,
            I => \N__24959\
        );

    \I__5555\ : Odrv4
    port map (
            O => \N__24959\,
            I => \eeprom.n3576_adj_358\
        );

    \I__5554\ : InMux
    port map (
            O => \N__24956\,
            I => \eeprom.n3758\
        );

    \I__5553\ : CascadeMux
    port map (
            O => \N__24953\,
            I => \N__24950\
        );

    \I__5552\ : InMux
    port map (
            O => \N__24950\,
            I => \N__24947\
        );

    \I__5551\ : LocalMux
    port map (
            O => \N__24947\,
            I => \N__24943\
        );

    \I__5550\ : InMux
    port map (
            O => \N__24946\,
            I => \N__24940\
        );

    \I__5549\ : Odrv12
    port map (
            O => \N__24943\,
            I => \eeprom.n3508\
        );

    \I__5548\ : LocalMux
    port map (
            O => \N__24940\,
            I => \eeprom.n3508\
        );

    \I__5547\ : InMux
    port map (
            O => \N__24935\,
            I => \N__24932\
        );

    \I__5546\ : LocalMux
    port map (
            O => \N__24932\,
            I => \N__24929\
        );

    \I__5545\ : Odrv4
    port map (
            O => \N__24929\,
            I => \eeprom.n3575_adj_357\
        );

    \I__5544\ : InMux
    port map (
            O => \N__24926\,
            I => \eeprom.n3759\
        );

    \I__5543\ : InMux
    port map (
            O => \N__24923\,
            I => \N__24919\
        );

    \I__5542\ : CascadeMux
    port map (
            O => \N__24922\,
            I => \N__24915\
        );

    \I__5541\ : LocalMux
    port map (
            O => \N__24919\,
            I => \N__24912\
        );

    \I__5540\ : InMux
    port map (
            O => \N__24918\,
            I => \N__24907\
        );

    \I__5539\ : InMux
    port map (
            O => \N__24915\,
            I => \N__24907\
        );

    \I__5538\ : Odrv4
    port map (
            O => \N__24912\,
            I => \eeprom.n3507\
        );

    \I__5537\ : LocalMux
    port map (
            O => \N__24907\,
            I => \eeprom.n3507\
        );

    \I__5536\ : CascadeMux
    port map (
            O => \N__24902\,
            I => \N__24899\
        );

    \I__5535\ : InMux
    port map (
            O => \N__24899\,
            I => \N__24896\
        );

    \I__5534\ : LocalMux
    port map (
            O => \N__24896\,
            I => \N__24893\
        );

    \I__5533\ : Span4Mux_v
    port map (
            O => \N__24893\,
            I => \N__24890\
        );

    \I__5532\ : Odrv4
    port map (
            O => \N__24890\,
            I => \eeprom.n3574_adj_356\
        );

    \I__5531\ : InMux
    port map (
            O => \N__24887\,
            I => \eeprom.n3760\
        );

    \I__5530\ : InMux
    port map (
            O => \N__24884\,
            I => \N__24880\
        );

    \I__5529\ : InMux
    port map (
            O => \N__24883\,
            I => \N__24877\
        );

    \I__5528\ : LocalMux
    port map (
            O => \N__24880\,
            I => \N__24874\
        );

    \I__5527\ : LocalMux
    port map (
            O => \N__24877\,
            I => \N__24871\
        );

    \I__5526\ : Span4Mux_h
    port map (
            O => \N__24874\,
            I => \N__24865\
        );

    \I__5525\ : Span4Mux_h
    port map (
            O => \N__24871\,
            I => \N__24865\
        );

    \I__5524\ : InMux
    port map (
            O => \N__24870\,
            I => \N__24862\
        );

    \I__5523\ : Odrv4
    port map (
            O => \N__24865\,
            I => \eeprom.n3506\
        );

    \I__5522\ : LocalMux
    port map (
            O => \N__24862\,
            I => \eeprom.n3506\
        );

    \I__5521\ : InMux
    port map (
            O => \N__24857\,
            I => \N__24854\
        );

    \I__5520\ : LocalMux
    port map (
            O => \N__24854\,
            I => \eeprom.n3573_adj_355\
        );

    \I__5519\ : InMux
    port map (
            O => \N__24851\,
            I => \eeprom.n3761\
        );

    \I__5518\ : InMux
    port map (
            O => \N__24848\,
            I => \N__24845\
        );

    \I__5517\ : LocalMux
    port map (
            O => \N__24845\,
            I => \N__24842\
        );

    \I__5516\ : Span4Mux_v
    port map (
            O => \N__24842\,
            I => \N__24839\
        );

    \I__5515\ : Odrv4
    port map (
            O => \N__24839\,
            I => \eeprom.n2986\
        );

    \I__5514\ : InMux
    port map (
            O => \N__24836\,
            I => \N__24833\
        );

    \I__5513\ : LocalMux
    port map (
            O => \N__24833\,
            I => \N__24829\
        );

    \I__5512\ : InMux
    port map (
            O => \N__24832\,
            I => \N__24826\
        );

    \I__5511\ : Span4Mux_h
    port map (
            O => \N__24829\,
            I => \N__24822\
        );

    \I__5510\ : LocalMux
    port map (
            O => \N__24826\,
            I => \N__24819\
        );

    \I__5509\ : InMux
    port map (
            O => \N__24825\,
            I => \N__24816\
        );

    \I__5508\ : Span4Mux_h
    port map (
            O => \N__24822\,
            I => \N__24811\
        );

    \I__5507\ : Span4Mux_v
    port map (
            O => \N__24819\,
            I => \N__24811\
        );

    \I__5506\ : LocalMux
    port map (
            O => \N__24816\,
            I => \N__24808\
        );

    \I__5505\ : Span4Mux_h
    port map (
            O => \N__24811\,
            I => \N__24803\
        );

    \I__5504\ : Span4Mux_h
    port map (
            O => \N__24808\,
            I => \N__24803\
        );

    \I__5503\ : Span4Mux_h
    port map (
            O => \N__24803\,
            I => \N__24800\
        );

    \I__5502\ : Odrv4
    port map (
            O => \N__24800\,
            I => \eeprom.n2919\
        );

    \I__5501\ : CascadeMux
    port map (
            O => \N__24797\,
            I => \N__24793\
        );

    \I__5500\ : InMux
    port map (
            O => \N__24796\,
            I => \N__24790\
        );

    \I__5499\ : InMux
    port map (
            O => \N__24793\,
            I => \N__24787\
        );

    \I__5498\ : LocalMux
    port map (
            O => \N__24790\,
            I => \N__24784\
        );

    \I__5497\ : LocalMux
    port map (
            O => \N__24787\,
            I => \N__24781\
        );

    \I__5496\ : Odrv12
    port map (
            O => \N__24784\,
            I => \eeprom.n2909\
        );

    \I__5495\ : Odrv4
    port map (
            O => \N__24781\,
            I => \eeprom.n2909\
        );

    \I__5494\ : InMux
    port map (
            O => \N__24776\,
            I => \N__24773\
        );

    \I__5493\ : LocalMux
    port map (
            O => \N__24773\,
            I => \N__24770\
        );

    \I__5492\ : Span4Mux_v
    port map (
            O => \N__24770\,
            I => \N__24767\
        );

    \I__5491\ : Odrv4
    port map (
            O => \N__24767\,
            I => \eeprom.n2976\
        );

    \I__5490\ : CascadeMux
    port map (
            O => \N__24764\,
            I => \N__24754\
        );

    \I__5489\ : InMux
    port map (
            O => \N__24763\,
            I => \N__24750\
        );

    \I__5488\ : InMux
    port map (
            O => \N__24762\,
            I => \N__24747\
        );

    \I__5487\ : InMux
    port map (
            O => \N__24761\,
            I => \N__24742\
        );

    \I__5486\ : InMux
    port map (
            O => \N__24760\,
            I => \N__24742\
        );

    \I__5485\ : CascadeMux
    port map (
            O => \N__24759\,
            I => \N__24738\
        );

    \I__5484\ : CascadeMux
    port map (
            O => \N__24758\,
            I => \N__24732\
        );

    \I__5483\ : CascadeMux
    port map (
            O => \N__24757\,
            I => \N__24729\
        );

    \I__5482\ : InMux
    port map (
            O => \N__24754\,
            I => \N__24722\
        );

    \I__5481\ : InMux
    port map (
            O => \N__24753\,
            I => \N__24722\
        );

    \I__5480\ : LocalMux
    port map (
            O => \N__24750\,
            I => \N__24719\
        );

    \I__5479\ : LocalMux
    port map (
            O => \N__24747\,
            I => \N__24714\
        );

    \I__5478\ : LocalMux
    port map (
            O => \N__24742\,
            I => \N__24714\
        );

    \I__5477\ : InMux
    port map (
            O => \N__24741\,
            I => \N__24707\
        );

    \I__5476\ : InMux
    port map (
            O => \N__24738\,
            I => \N__24707\
        );

    \I__5475\ : InMux
    port map (
            O => \N__24737\,
            I => \N__24707\
        );

    \I__5474\ : CascadeMux
    port map (
            O => \N__24736\,
            I => \N__24702\
        );

    \I__5473\ : InMux
    port map (
            O => \N__24735\,
            I => \N__24698\
        );

    \I__5472\ : InMux
    port map (
            O => \N__24732\,
            I => \N__24689\
        );

    \I__5471\ : InMux
    port map (
            O => \N__24729\,
            I => \N__24689\
        );

    \I__5470\ : InMux
    port map (
            O => \N__24728\,
            I => \N__24689\
        );

    \I__5469\ : InMux
    port map (
            O => \N__24727\,
            I => \N__24689\
        );

    \I__5468\ : LocalMux
    port map (
            O => \N__24722\,
            I => \N__24680\
        );

    \I__5467\ : Span4Mux_v
    port map (
            O => \N__24719\,
            I => \N__24680\
        );

    \I__5466\ : Span4Mux_h
    port map (
            O => \N__24714\,
            I => \N__24680\
        );

    \I__5465\ : LocalMux
    port map (
            O => \N__24707\,
            I => \N__24680\
        );

    \I__5464\ : InMux
    port map (
            O => \N__24706\,
            I => \N__24671\
        );

    \I__5463\ : InMux
    port map (
            O => \N__24705\,
            I => \N__24671\
        );

    \I__5462\ : InMux
    port map (
            O => \N__24702\,
            I => \N__24671\
        );

    \I__5461\ : InMux
    port map (
            O => \N__24701\,
            I => \N__24671\
        );

    \I__5460\ : LocalMux
    port map (
            O => \N__24698\,
            I => \N__24668\
        );

    \I__5459\ : LocalMux
    port map (
            O => \N__24689\,
            I => \eeprom.n2935\
        );

    \I__5458\ : Odrv4
    port map (
            O => \N__24680\,
            I => \eeprom.n2935\
        );

    \I__5457\ : LocalMux
    port map (
            O => \N__24671\,
            I => \eeprom.n2935\
        );

    \I__5456\ : Odrv4
    port map (
            O => \N__24668\,
            I => \eeprom.n2935\
        );

    \I__5455\ : InMux
    port map (
            O => \N__24659\,
            I => \N__24655\
        );

    \I__5454\ : InMux
    port map (
            O => \N__24658\,
            I => \N__24651\
        );

    \I__5453\ : LocalMux
    port map (
            O => \N__24655\,
            I => \N__24648\
        );

    \I__5452\ : InMux
    port map (
            O => \N__24654\,
            I => \N__24645\
        );

    \I__5451\ : LocalMux
    port map (
            O => \N__24651\,
            I => \N__24642\
        );

    \I__5450\ : Span12Mux_v
    port map (
            O => \N__24648\,
            I => \N__24639\
        );

    \I__5449\ : LocalMux
    port map (
            O => \N__24645\,
            I => \N__24636\
        );

    \I__5448\ : Span4Mux_v
    port map (
            O => \N__24642\,
            I => \N__24633\
        );

    \I__5447\ : Span12Mux_h
    port map (
            O => \N__24639\,
            I => \N__24630\
        );

    \I__5446\ : Span12Mux_v
    port map (
            O => \N__24636\,
            I => \N__24625\
        );

    \I__5445\ : Sp12to4
    port map (
            O => \N__24633\,
            I => \N__24625\
        );

    \I__5444\ : Odrv12
    port map (
            O => \N__24630\,
            I => \eeprom.n3519_adj_379\
        );

    \I__5443\ : Odrv12
    port map (
            O => \N__24625\,
            I => \eeprom.n3519_adj_379\
        );

    \I__5442\ : InMux
    port map (
            O => \N__24620\,
            I => \N__24617\
        );

    \I__5441\ : LocalMux
    port map (
            O => \N__24617\,
            I => \N__24614\
        );

    \I__5440\ : Span4Mux_h
    port map (
            O => \N__24614\,
            I => \N__24611\
        );

    \I__5439\ : Odrv4
    port map (
            O => \N__24611\,
            I => \eeprom.n3586_adj_378\
        );

    \I__5438\ : InMux
    port map (
            O => \N__24608\,
            I => \bfn_16_17_0_\
        );

    \I__5437\ : CascadeMux
    port map (
            O => \N__24605\,
            I => \N__24601\
        );

    \I__5436\ : InMux
    port map (
            O => \N__24604\,
            I => \N__24597\
        );

    \I__5435\ : InMux
    port map (
            O => \N__24601\,
            I => \N__24594\
        );

    \I__5434\ : InMux
    port map (
            O => \N__24600\,
            I => \N__24591\
        );

    \I__5433\ : LocalMux
    port map (
            O => \N__24597\,
            I => \eeprom.n3518_adj_376\
        );

    \I__5432\ : LocalMux
    port map (
            O => \N__24594\,
            I => \eeprom.n3518_adj_376\
        );

    \I__5431\ : LocalMux
    port map (
            O => \N__24591\,
            I => \eeprom.n3518_adj_376\
        );

    \I__5430\ : InMux
    port map (
            O => \N__24584\,
            I => \N__24581\
        );

    \I__5429\ : LocalMux
    port map (
            O => \N__24581\,
            I => \eeprom.n3585_adj_375\
        );

    \I__5428\ : InMux
    port map (
            O => \N__24578\,
            I => \eeprom.n3749\
        );

    \I__5427\ : CascadeMux
    port map (
            O => \N__24575\,
            I => \N__24571\
        );

    \I__5426\ : InMux
    port map (
            O => \N__24574\,
            I => \N__24568\
        );

    \I__5425\ : InMux
    port map (
            O => \N__24571\,
            I => \N__24565\
        );

    \I__5424\ : LocalMux
    port map (
            O => \N__24568\,
            I => \eeprom.n3517_adj_374\
        );

    \I__5423\ : LocalMux
    port map (
            O => \N__24565\,
            I => \eeprom.n3517_adj_374\
        );

    \I__5422\ : InMux
    port map (
            O => \N__24560\,
            I => \N__24557\
        );

    \I__5421\ : LocalMux
    port map (
            O => \N__24557\,
            I => \eeprom.n3584_adj_373\
        );

    \I__5420\ : InMux
    port map (
            O => \N__24554\,
            I => \eeprom.n3750\
        );

    \I__5419\ : CascadeMux
    port map (
            O => \N__24551\,
            I => \N__24547\
        );

    \I__5418\ : CascadeMux
    port map (
            O => \N__24550\,
            I => \N__24544\
        );

    \I__5417\ : InMux
    port map (
            O => \N__24547\,
            I => \N__24540\
        );

    \I__5416\ : InMux
    port map (
            O => \N__24544\,
            I => \N__24537\
        );

    \I__5415\ : InMux
    port map (
            O => \N__24543\,
            I => \N__24534\
        );

    \I__5414\ : LocalMux
    port map (
            O => \N__24540\,
            I => \eeprom.n3516_adj_372\
        );

    \I__5413\ : LocalMux
    port map (
            O => \N__24537\,
            I => \eeprom.n3516_adj_372\
        );

    \I__5412\ : LocalMux
    port map (
            O => \N__24534\,
            I => \eeprom.n3516_adj_372\
        );

    \I__5411\ : InMux
    port map (
            O => \N__24527\,
            I => \N__24524\
        );

    \I__5410\ : LocalMux
    port map (
            O => \N__24524\,
            I => \eeprom.n3583_adj_371\
        );

    \I__5409\ : InMux
    port map (
            O => \N__24521\,
            I => \eeprom.n3751\
        );

    \I__5408\ : CascadeMux
    port map (
            O => \N__24518\,
            I => \N__24514\
        );

    \I__5407\ : InMux
    port map (
            O => \N__24517\,
            I => \N__24511\
        );

    \I__5406\ : InMux
    port map (
            O => \N__24514\,
            I => \N__24508\
        );

    \I__5405\ : LocalMux
    port map (
            O => \N__24511\,
            I => \eeprom.n3515_adj_370\
        );

    \I__5404\ : LocalMux
    port map (
            O => \N__24508\,
            I => \eeprom.n3515_adj_370\
        );

    \I__5403\ : CascadeMux
    port map (
            O => \N__24503\,
            I => \N__24500\
        );

    \I__5402\ : InMux
    port map (
            O => \N__24500\,
            I => \N__24497\
        );

    \I__5401\ : LocalMux
    port map (
            O => \N__24497\,
            I => \eeprom.n3582_adj_369\
        );

    \I__5400\ : InMux
    port map (
            O => \N__24494\,
            I => \eeprom.n3752\
        );

    \I__5399\ : CascadeMux
    port map (
            O => \N__24491\,
            I => \N__24488\
        );

    \I__5398\ : InMux
    port map (
            O => \N__24488\,
            I => \N__24484\
        );

    \I__5397\ : InMux
    port map (
            O => \N__24487\,
            I => \N__24480\
        );

    \I__5396\ : LocalMux
    port map (
            O => \N__24484\,
            I => \N__24477\
        );

    \I__5395\ : InMux
    port map (
            O => \N__24483\,
            I => \N__24474\
        );

    \I__5394\ : LocalMux
    port map (
            O => \N__24480\,
            I => \N__24471\
        );

    \I__5393\ : Span4Mux_h
    port map (
            O => \N__24477\,
            I => \N__24466\
        );

    \I__5392\ : LocalMux
    port map (
            O => \N__24474\,
            I => \N__24466\
        );

    \I__5391\ : Odrv12
    port map (
            O => \N__24471\,
            I => \eeprom.n3514_adj_368\
        );

    \I__5390\ : Odrv4
    port map (
            O => \N__24466\,
            I => \eeprom.n3514_adj_368\
        );

    \I__5389\ : CascadeMux
    port map (
            O => \N__24461\,
            I => \N__24458\
        );

    \I__5388\ : InMux
    port map (
            O => \N__24458\,
            I => \N__24455\
        );

    \I__5387\ : LocalMux
    port map (
            O => \N__24455\,
            I => \N__24452\
        );

    \I__5386\ : Span4Mux_h
    port map (
            O => \N__24452\,
            I => \N__24449\
        );

    \I__5385\ : Odrv4
    port map (
            O => \N__24449\,
            I => \eeprom.n3581_adj_367\
        );

    \I__5384\ : InMux
    port map (
            O => \N__24446\,
            I => \eeprom.n3753\
        );

    \I__5383\ : InMux
    port map (
            O => \N__24443\,
            I => \N__24440\
        );

    \I__5382\ : LocalMux
    port map (
            O => \N__24440\,
            I => \N__24437\
        );

    \I__5381\ : Odrv12
    port map (
            O => \N__24437\,
            I => \eeprom.number_of_bytes_7_N_68_6\
        );

    \I__5380\ : InMux
    port map (
            O => \N__24434\,
            I => \N__24431\
        );

    \I__5379\ : LocalMux
    port map (
            O => \N__24431\,
            I => \eeprom.number_of_bytes_7_N_68_8\
        );

    \I__5378\ : CascadeMux
    port map (
            O => \N__24428\,
            I => \eeprom.n4301_cascade_\
        );

    \I__5377\ : InMux
    port map (
            O => \N__24425\,
            I => \N__24422\
        );

    \I__5376\ : LocalMux
    port map (
            O => \N__24422\,
            I => \N__24419\
        );

    \I__5375\ : Odrv4
    port map (
            O => \N__24419\,
            I => \eeprom.number_of_bytes_7_N_68_7\
        );

    \I__5374\ : InMux
    port map (
            O => \N__24416\,
            I => \N__24413\
        );

    \I__5373\ : LocalMux
    port map (
            O => \N__24413\,
            I => \eeprom.number_of_bytes_7_N_68_9\
        );

    \I__5372\ : InMux
    port map (
            O => \N__24410\,
            I => \N__24407\
        );

    \I__5371\ : LocalMux
    port map (
            O => \N__24407\,
            I => \eeprom.number_of_bytes_7_N_68_10\
        );

    \I__5370\ : CascadeMux
    port map (
            O => \N__24404\,
            I => \eeprom.n4307_cascade_\
        );

    \I__5369\ : InMux
    port map (
            O => \N__24401\,
            I => \N__24398\
        );

    \I__5368\ : LocalMux
    port map (
            O => \N__24398\,
            I => \eeprom.number_of_bytes_7_N_68_11\
        );

    \I__5367\ : InMux
    port map (
            O => \N__24395\,
            I => \N__24392\
        );

    \I__5366\ : LocalMux
    port map (
            O => \N__24392\,
            I => \eeprom.number_of_bytes_7_N_68_12\
        );

    \I__5365\ : InMux
    port map (
            O => \N__24389\,
            I => \N__24386\
        );

    \I__5364\ : LocalMux
    port map (
            O => \N__24386\,
            I => \eeprom.number_of_bytes_7_N_68_13\
        );

    \I__5363\ : CascadeMux
    port map (
            O => \N__24383\,
            I => \eeprom.n4313_cascade_\
        );

    \I__5362\ : InMux
    port map (
            O => \N__24380\,
            I => \N__24377\
        );

    \I__5361\ : LocalMux
    port map (
            O => \N__24377\,
            I => \eeprom.number_of_bytes_7_N_68_14\
        );

    \I__5360\ : IoInMux
    port map (
            O => \N__24374\,
            I => \N__24371\
        );

    \I__5359\ : LocalMux
    port map (
            O => \N__24371\,
            I => \N__24368\
        );

    \I__5358\ : IoSpan4Mux
    port map (
            O => \N__24368\,
            I => \N__24365\
        );

    \I__5357\ : Span4Mux_s3_h
    port map (
            O => \N__24365\,
            I => \N__24362\
        );

    \I__5356\ : Sp12to4
    port map (
            O => \N__24362\,
            I => \N__24359\
        );

    \I__5355\ : Span12Mux_h
    port map (
            O => \N__24359\,
            I => \N__24356\
        );

    \I__5354\ : Span12Mux_v
    port map (
            O => \N__24356\,
            I => \N__24353\
        );

    \I__5353\ : Odrv12
    port map (
            O => \N__24353\,
            I => sda_enable
        );

    \I__5352\ : ClkMux
    port map (
            O => \N__24350\,
            I => \N__24323\
        );

    \I__5351\ : ClkMux
    port map (
            O => \N__24349\,
            I => \N__24323\
        );

    \I__5350\ : ClkMux
    port map (
            O => \N__24348\,
            I => \N__24323\
        );

    \I__5349\ : ClkMux
    port map (
            O => \N__24347\,
            I => \N__24323\
        );

    \I__5348\ : ClkMux
    port map (
            O => \N__24346\,
            I => \N__24323\
        );

    \I__5347\ : ClkMux
    port map (
            O => \N__24345\,
            I => \N__24323\
        );

    \I__5346\ : ClkMux
    port map (
            O => \N__24344\,
            I => \N__24323\
        );

    \I__5345\ : ClkMux
    port map (
            O => \N__24343\,
            I => \N__24323\
        );

    \I__5344\ : ClkMux
    port map (
            O => \N__24342\,
            I => \N__24323\
        );

    \I__5343\ : GlobalMux
    port map (
            O => \N__24323\,
            I => \N__24320\
        );

    \I__5342\ : gio2CtrlBuf
    port map (
            O => \N__24320\,
            I => \CLK_N\
        );

    \I__5341\ : InMux
    port map (
            O => \N__24317\,
            I => \N__24314\
        );

    \I__5340\ : LocalMux
    port map (
            O => \N__24314\,
            I => \N__24311\
        );

    \I__5339\ : Odrv4
    port map (
            O => \N__24311\,
            I => \eeprom.number_of_bytes_7_N_68_2\
        );

    \I__5338\ : InMux
    port map (
            O => \N__24308\,
            I => \N__24305\
        );

    \I__5337\ : LocalMux
    port map (
            O => \N__24305\,
            I => \N__24302\
        );

    \I__5336\ : Odrv12
    port map (
            O => \N__24302\,
            I => \eeprom.number_of_bytes_7_N_68_0\
        );

    \I__5335\ : InMux
    port map (
            O => \N__24299\,
            I => \N__24296\
        );

    \I__5334\ : LocalMux
    port map (
            O => \N__24296\,
            I => \N__24293\
        );

    \I__5333\ : Odrv12
    port map (
            O => \N__24293\,
            I => \eeprom.number_of_bytes_7_N_68_1\
        );

    \I__5332\ : InMux
    port map (
            O => \N__24290\,
            I => \N__24287\
        );

    \I__5331\ : LocalMux
    port map (
            O => \N__24287\,
            I => \eeprom.n4295\
        );

    \I__5330\ : CascadeMux
    port map (
            O => \N__24284\,
            I => \N__24280\
        );

    \I__5329\ : InMux
    port map (
            O => \N__24283\,
            I => \N__24277\
        );

    \I__5328\ : InMux
    port map (
            O => \N__24280\,
            I => \N__24274\
        );

    \I__5327\ : LocalMux
    port map (
            O => \N__24277\,
            I => \N__24270\
        );

    \I__5326\ : LocalMux
    port map (
            O => \N__24274\,
            I => \N__24267\
        );

    \I__5325\ : CascadeMux
    port map (
            O => \N__24273\,
            I => \N__24264\
        );

    \I__5324\ : Span4Mux_h
    port map (
            O => \N__24270\,
            I => \N__24261\
        );

    \I__5323\ : Span4Mux_h
    port map (
            O => \N__24267\,
            I => \N__24258\
        );

    \I__5322\ : InMux
    port map (
            O => \N__24264\,
            I => \N__24255\
        );

    \I__5321\ : Odrv4
    port map (
            O => \N__24261\,
            I => \eeprom.n3111\
        );

    \I__5320\ : Odrv4
    port map (
            O => \N__24258\,
            I => \eeprom.n3111\
        );

    \I__5319\ : LocalMux
    port map (
            O => \N__24255\,
            I => \eeprom.n3111\
        );

    \I__5318\ : InMux
    port map (
            O => \N__24248\,
            I => \N__24245\
        );

    \I__5317\ : LocalMux
    port map (
            O => \N__24245\,
            I => \N__24241\
        );

    \I__5316\ : CascadeMux
    port map (
            O => \N__24244\,
            I => \N__24238\
        );

    \I__5315\ : Span4Mux_v
    port map (
            O => \N__24241\,
            I => \N__24235\
        );

    \I__5314\ : InMux
    port map (
            O => \N__24238\,
            I => \N__24232\
        );

    \I__5313\ : Span4Mux_h
    port map (
            O => \N__24235\,
            I => \N__24228\
        );

    \I__5312\ : LocalMux
    port map (
            O => \N__24232\,
            I => \N__24225\
        );

    \I__5311\ : InMux
    port map (
            O => \N__24231\,
            I => \N__24222\
        );

    \I__5310\ : Odrv4
    port map (
            O => \N__24228\,
            I => \eeprom.n3109\
        );

    \I__5309\ : Odrv4
    port map (
            O => \N__24225\,
            I => \eeprom.n3109\
        );

    \I__5308\ : LocalMux
    port map (
            O => \N__24222\,
            I => \eeprom.n3109\
        );

    \I__5307\ : InMux
    port map (
            O => \N__24215\,
            I => \N__24212\
        );

    \I__5306\ : LocalMux
    port map (
            O => \N__24212\,
            I => \N__24209\
        );

    \I__5305\ : Span4Mux_v
    port map (
            O => \N__24209\,
            I => \N__24205\
        );

    \I__5304\ : InMux
    port map (
            O => \N__24208\,
            I => \N__24202\
        );

    \I__5303\ : Span4Mux_h
    port map (
            O => \N__24205\,
            I => \N__24198\
        );

    \I__5302\ : LocalMux
    port map (
            O => \N__24202\,
            I => \N__24195\
        );

    \I__5301\ : InMux
    port map (
            O => \N__24201\,
            I => \N__24192\
        );

    \I__5300\ : Odrv4
    port map (
            O => \N__24198\,
            I => \eeprom.n3110\
        );

    \I__5299\ : Odrv4
    port map (
            O => \N__24195\,
            I => \eeprom.n3110\
        );

    \I__5298\ : LocalMux
    port map (
            O => \N__24192\,
            I => \eeprom.n3110\
        );

    \I__5297\ : CascadeMux
    port map (
            O => \N__24185\,
            I => \N__24182\
        );

    \I__5296\ : InMux
    port map (
            O => \N__24182\,
            I => \N__24179\
        );

    \I__5295\ : LocalMux
    port map (
            O => \N__24179\,
            I => \N__24175\
        );

    \I__5294\ : InMux
    port map (
            O => \N__24178\,
            I => \N__24172\
        );

    \I__5293\ : Span4Mux_h
    port map (
            O => \N__24175\,
            I => \N__24168\
        );

    \I__5292\ : LocalMux
    port map (
            O => \N__24172\,
            I => \N__24165\
        );

    \I__5291\ : InMux
    port map (
            O => \N__24171\,
            I => \N__24162\
        );

    \I__5290\ : Odrv4
    port map (
            O => \N__24168\,
            I => \eeprom.n3107\
        );

    \I__5289\ : Odrv4
    port map (
            O => \N__24165\,
            I => \eeprom.n3107\
        );

    \I__5288\ : LocalMux
    port map (
            O => \N__24162\,
            I => \eeprom.n3107\
        );

    \I__5287\ : InMux
    port map (
            O => \N__24155\,
            I => \N__24152\
        );

    \I__5286\ : LocalMux
    port map (
            O => \N__24152\,
            I => \N__24149\
        );

    \I__5285\ : Odrv4
    port map (
            O => \N__24149\,
            I => \eeprom.n4909\
        );

    \I__5284\ : CascadeMux
    port map (
            O => \N__24146\,
            I => \N__24143\
        );

    \I__5283\ : InMux
    port map (
            O => \N__24143\,
            I => \N__24140\
        );

    \I__5282\ : LocalMux
    port map (
            O => \N__24140\,
            I => \N__24137\
        );

    \I__5281\ : Odrv4
    port map (
            O => \N__24137\,
            I => \eeprom.n3716_adj_439\
        );

    \I__5280\ : InMux
    port map (
            O => \N__24134\,
            I => \eeprom.n3780\
        );

    \I__5279\ : InMux
    port map (
            O => \N__24131\,
            I => \eeprom.n3781\
        );

    \I__5278\ : InMux
    port map (
            O => \N__24128\,
            I => \N__24125\
        );

    \I__5277\ : LocalMux
    port map (
            O => \N__24125\,
            I => \N__24122\
        );

    \I__5276\ : Odrv4
    port map (
            O => \N__24122\,
            I => \eeprom.n4915\
        );

    \I__5275\ : CascadeMux
    port map (
            O => \N__24119\,
            I => \N__24116\
        );

    \I__5274\ : InMux
    port map (
            O => \N__24116\,
            I => \N__24113\
        );

    \I__5273\ : LocalMux
    port map (
            O => \N__24113\,
            I => \N__24110\
        );

    \I__5272\ : Odrv4
    port map (
            O => \N__24110\,
            I => \eeprom.n3714_adj_442\
        );

    \I__5271\ : InMux
    port map (
            O => \N__24107\,
            I => \eeprom.n3782\
        );

    \I__5270\ : InMux
    port map (
            O => \N__24104\,
            I => \eeprom.n3783\
        );

    \I__5269\ : InMux
    port map (
            O => \N__24101\,
            I => \N__24098\
        );

    \I__5268\ : LocalMux
    port map (
            O => \N__24098\,
            I => \eeprom.n4921\
        );

    \I__5267\ : CascadeMux
    port map (
            O => \N__24095\,
            I => \N__24092\
        );

    \I__5266\ : InMux
    port map (
            O => \N__24092\,
            I => \N__24088\
        );

    \I__5265\ : InMux
    port map (
            O => \N__24091\,
            I => \N__24085\
        );

    \I__5264\ : LocalMux
    port map (
            O => \N__24088\,
            I => \eeprom.n3712_adj_444\
        );

    \I__5263\ : LocalMux
    port map (
            O => \N__24085\,
            I => \eeprom.n3712_adj_444\
        );

    \I__5262\ : InMux
    port map (
            O => \N__24080\,
            I => \eeprom.n3784\
        );

    \I__5261\ : CascadeMux
    port map (
            O => \N__24077\,
            I => \N__24071\
        );

    \I__5260\ : CascadeMux
    port map (
            O => \N__24076\,
            I => \N__24067\
        );

    \I__5259\ : CascadeMux
    port map (
            O => \N__24075\,
            I => \N__24063\
        );

    \I__5258\ : InMux
    port map (
            O => \N__24074\,
            I => \N__24044\
        );

    \I__5257\ : InMux
    port map (
            O => \N__24071\,
            I => \N__24044\
        );

    \I__5256\ : InMux
    port map (
            O => \N__24070\,
            I => \N__24044\
        );

    \I__5255\ : InMux
    port map (
            O => \N__24067\,
            I => \N__24044\
        );

    \I__5254\ : InMux
    port map (
            O => \N__24066\,
            I => \N__24044\
        );

    \I__5253\ : InMux
    port map (
            O => \N__24063\,
            I => \N__24044\
        );

    \I__5252\ : InMux
    port map (
            O => \N__24062\,
            I => \N__24044\
        );

    \I__5251\ : CascadeMux
    port map (
            O => \N__24061\,
            I => \N__24038\
        );

    \I__5250\ : CascadeMux
    port map (
            O => \N__24060\,
            I => \N__24034\
        );

    \I__5249\ : InMux
    port map (
            O => \N__24059\,
            I => \N__24030\
        );

    \I__5248\ : LocalMux
    port map (
            O => \N__24044\,
            I => \N__24027\
        );

    \I__5247\ : InMux
    port map (
            O => \N__24043\,
            I => \N__24024\
        );

    \I__5246\ : InMux
    port map (
            O => \N__24042\,
            I => \N__24011\
        );

    \I__5245\ : InMux
    port map (
            O => \N__24041\,
            I => \N__24011\
        );

    \I__5244\ : InMux
    port map (
            O => \N__24038\,
            I => \N__24011\
        );

    \I__5243\ : InMux
    port map (
            O => \N__24037\,
            I => \N__24011\
        );

    \I__5242\ : InMux
    port map (
            O => \N__24034\,
            I => \N__24011\
        );

    \I__5241\ : InMux
    port map (
            O => \N__24033\,
            I => \N__24011\
        );

    \I__5240\ : LocalMux
    port map (
            O => \N__24030\,
            I => \N__24008\
        );

    \I__5239\ : Span4Mux_h
    port map (
            O => \N__24027\,
            I => \N__24005\
        );

    \I__5238\ : LocalMux
    port map (
            O => \N__24024\,
            I => \N__23999\
        );

    \I__5237\ : LocalMux
    port map (
            O => \N__24011\,
            I => \N__23999\
        );

    \I__5236\ : Span12Mux_v
    port map (
            O => \N__24008\,
            I => \N__23996\
        );

    \I__5235\ : Span4Mux_h
    port map (
            O => \N__24005\,
            I => \N__23993\
        );

    \I__5234\ : InMux
    port map (
            O => \N__24004\,
            I => \N__23990\
        );

    \I__5233\ : Span12Mux_h
    port map (
            O => \N__23999\,
            I => \N__23987\
        );

    \I__5232\ : Span12Mux_h
    port map (
            O => \N__23996\,
            I => \N__23984\
        );

    \I__5231\ : Span4Mux_h
    port map (
            O => \N__23993\,
            I => \N__23981\
        );

    \I__5230\ : LocalMux
    port map (
            O => \N__23990\,
            I => \N__23978\
        );

    \I__5229\ : Odrv12
    port map (
            O => \N__23987\,
            I => \eeprom.n2\
        );

    \I__5228\ : Odrv12
    port map (
            O => \N__23984\,
            I => \eeprom.n2\
        );

    \I__5227\ : Odrv4
    port map (
            O => \N__23981\,
            I => \eeprom.n2\
        );

    \I__5226\ : Odrv4
    port map (
            O => \N__23978\,
            I => \eeprom.n2\
        );

    \I__5225\ : InMux
    port map (
            O => \N__23969\,
            I => \N__23966\
        );

    \I__5224\ : LocalMux
    port map (
            O => \N__23966\,
            I => \eeprom.n4924\
        );

    \I__5223\ : InMux
    port map (
            O => \N__23963\,
            I => \eeprom.n3785\
        );

    \I__5222\ : CascadeMux
    port map (
            O => \N__23960\,
            I => \N__23956\
        );

    \I__5221\ : InMux
    port map (
            O => \N__23959\,
            I => \N__23951\
        );

    \I__5220\ : InMux
    port map (
            O => \N__23956\,
            I => \N__23951\
        );

    \I__5219\ : LocalMux
    port map (
            O => \N__23951\,
            I => \eeprom.n3713_adj_443\
        );

    \I__5218\ : InMux
    port map (
            O => \N__23948\,
            I => \N__23945\
        );

    \I__5217\ : LocalMux
    port map (
            O => \N__23945\,
            I => \eeprom.n4918\
        );

    \I__5216\ : InMux
    port map (
            O => \N__23942\,
            I => \N__23939\
        );

    \I__5215\ : LocalMux
    port map (
            O => \N__23939\,
            I => \N__23936\
        );

    \I__5214\ : Odrv4
    port map (
            O => \N__23936\,
            I => \eeprom.number_of_bytes_7_N_68_5\
        );

    \I__5213\ : InMux
    port map (
            O => \N__23933\,
            I => \N__23930\
        );

    \I__5212\ : LocalMux
    port map (
            O => \N__23930\,
            I => \N__23927\
        );

    \I__5211\ : Odrv12
    port map (
            O => \N__23927\,
            I => \eeprom.number_of_bytes_7_N_68_4\
        );

    \I__5210\ : CascadeMux
    port map (
            O => \N__23924\,
            I => \N__23921\
        );

    \I__5209\ : InMux
    port map (
            O => \N__23921\,
            I => \N__23918\
        );

    \I__5208\ : LocalMux
    port map (
            O => \N__23918\,
            I => \N__23915\
        );

    \I__5207\ : Odrv12
    port map (
            O => \N__23915\,
            I => \eeprom.number_of_bytes_7_N_68_3\
        );

    \I__5206\ : InMux
    port map (
            O => \N__23912\,
            I => \N__23909\
        );

    \I__5205\ : LocalMux
    port map (
            O => \N__23909\,
            I => \N__23905\
        );

    \I__5204\ : InMux
    port map (
            O => \N__23908\,
            I => \N__23902\
        );

    \I__5203\ : Span4Mux_v
    port map (
            O => \N__23905\,
            I => \N__23898\
        );

    \I__5202\ : LocalMux
    port map (
            O => \N__23902\,
            I => \N__23895\
        );

    \I__5201\ : InMux
    port map (
            O => \N__23901\,
            I => \N__23892\
        );

    \I__5200\ : Span4Mux_h
    port map (
            O => \N__23898\,
            I => \N__23886\
        );

    \I__5199\ : Span4Mux_v
    port map (
            O => \N__23895\,
            I => \N__23886\
        );

    \I__5198\ : LocalMux
    port map (
            O => \N__23892\,
            I => \N__23883\
        );

    \I__5197\ : InMux
    port map (
            O => \N__23891\,
            I => \N__23880\
        );

    \I__5196\ : Sp12to4
    port map (
            O => \N__23886\,
            I => \N__23877\
        );

    \I__5195\ : Span4Mux_v
    port map (
            O => \N__23883\,
            I => \N__23874\
        );

    \I__5194\ : LocalMux
    port map (
            O => \N__23880\,
            I => \eeprom.delay_counter_1\
        );

    \I__5193\ : Odrv12
    port map (
            O => \N__23877\,
            I => \eeprom.delay_counter_1\
        );

    \I__5192\ : Odrv4
    port map (
            O => \N__23874\,
            I => \eeprom.delay_counter_1\
        );

    \I__5191\ : InMux
    port map (
            O => \N__23867\,
            I => \N__23864\
        );

    \I__5190\ : LocalMux
    port map (
            O => \N__23864\,
            I => \N__23861\
        );

    \I__5189\ : Span12Mux_h
    port map (
            O => \N__23861\,
            I => \N__23858\
        );

    \I__5188\ : Odrv12
    port map (
            O => \N__23858\,
            I => \eeprom.n3724_adj_335\
        );

    \I__5187\ : InMux
    port map (
            O => \N__23855\,
            I => \eeprom.n3772\
        );

    \I__5186\ : InMux
    port map (
            O => \N__23852\,
            I => \N__23849\
        );

    \I__5185\ : LocalMux
    port map (
            O => \N__23849\,
            I => \N__23846\
        );

    \I__5184\ : Span4Mux_v
    port map (
            O => \N__23846\,
            I => \N__23842\
        );

    \I__5183\ : InMux
    port map (
            O => \N__23845\,
            I => \N__23839\
        );

    \I__5182\ : Span4Mux_v
    port map (
            O => \N__23842\,
            I => \N__23835\
        );

    \I__5181\ : LocalMux
    port map (
            O => \N__23839\,
            I => \N__23832\
        );

    \I__5180\ : CascadeMux
    port map (
            O => \N__23838\,
            I => \N__23829\
        );

    \I__5179\ : Sp12to4
    port map (
            O => \N__23835\,
            I => \N__23823\
        );

    \I__5178\ : Span12Mux_v
    port map (
            O => \N__23832\,
            I => \N__23823\
        );

    \I__5177\ : InMux
    port map (
            O => \N__23829\,
            I => \N__23820\
        );

    \I__5176\ : InMux
    port map (
            O => \N__23828\,
            I => \N__23817\
        );

    \I__5175\ : Span12Mux_h
    port map (
            O => \N__23823\,
            I => \N__23814\
        );

    \I__5174\ : LocalMux
    port map (
            O => \N__23820\,
            I => \N__23811\
        );

    \I__5173\ : LocalMux
    port map (
            O => \N__23817\,
            I => \eeprom.delay_counter_2\
        );

    \I__5172\ : Odrv12
    port map (
            O => \N__23814\,
            I => \eeprom.delay_counter_2\
        );

    \I__5171\ : Odrv4
    port map (
            O => \N__23811\,
            I => \eeprom.delay_counter_2\
        );

    \I__5170\ : CascadeMux
    port map (
            O => \N__23804\,
            I => \N__23801\
        );

    \I__5169\ : InMux
    port map (
            O => \N__23801\,
            I => \N__23798\
        );

    \I__5168\ : LocalMux
    port map (
            O => \N__23798\,
            I => \N__23795\
        );

    \I__5167\ : Odrv4
    port map (
            O => \N__23795\,
            I => \eeprom.n3723_adj_334\
        );

    \I__5166\ : InMux
    port map (
            O => \N__23792\,
            I => \eeprom.n3773\
        );

    \I__5165\ : InMux
    port map (
            O => \N__23789\,
            I => \N__23785\
        );

    \I__5164\ : CascadeMux
    port map (
            O => \N__23788\,
            I => \N__23782\
        );

    \I__5163\ : LocalMux
    port map (
            O => \N__23785\,
            I => \N__23779\
        );

    \I__5162\ : InMux
    port map (
            O => \N__23782\,
            I => \N__23776\
        );

    \I__5161\ : Span12Mux_h
    port map (
            O => \N__23779\,
            I => \N__23773\
        );

    \I__5160\ : LocalMux
    port map (
            O => \N__23776\,
            I => \N__23769\
        );

    \I__5159\ : Span12Mux_h
    port map (
            O => \N__23773\,
            I => \N__23765\
        );

    \I__5158\ : InMux
    port map (
            O => \N__23772\,
            I => \N__23762\
        );

    \I__5157\ : Span4Mux_v
    port map (
            O => \N__23769\,
            I => \N__23759\
        );

    \I__5156\ : InMux
    port map (
            O => \N__23768\,
            I => \N__23756\
        );

    \I__5155\ : Odrv12
    port map (
            O => \N__23765\,
            I => \eeprom.delay_counter_3\
        );

    \I__5154\ : LocalMux
    port map (
            O => \N__23762\,
            I => \eeprom.delay_counter_3\
        );

    \I__5153\ : Odrv4
    port map (
            O => \N__23759\,
            I => \eeprom.delay_counter_3\
        );

    \I__5152\ : LocalMux
    port map (
            O => \N__23756\,
            I => \eeprom.delay_counter_3\
        );

    \I__5151\ : InMux
    port map (
            O => \N__23747\,
            I => \N__23744\
        );

    \I__5150\ : LocalMux
    port map (
            O => \N__23744\,
            I => \N__23741\
        );

    \I__5149\ : Span4Mux_v
    port map (
            O => \N__23741\,
            I => \N__23738\
        );

    \I__5148\ : Span4Mux_h
    port map (
            O => \N__23738\,
            I => \N__23735\
        );

    \I__5147\ : Span4Mux_h
    port map (
            O => \N__23735\,
            I => \N__23732\
        );

    \I__5146\ : Odrv4
    port map (
            O => \N__23732\,
            I => \eeprom.n3722_adj_433\
        );

    \I__5145\ : InMux
    port map (
            O => \N__23729\,
            I => \eeprom.n3774\
        );

    \I__5144\ : InMux
    port map (
            O => \N__23726\,
            I => \N__23723\
        );

    \I__5143\ : LocalMux
    port map (
            O => \N__23723\,
            I => \N__23719\
        );

    \I__5142\ : InMux
    port map (
            O => \N__23722\,
            I => \N__23716\
        );

    \I__5141\ : Span4Mux_v
    port map (
            O => \N__23719\,
            I => \N__23711\
        );

    \I__5140\ : LocalMux
    port map (
            O => \N__23716\,
            I => \N__23711\
        );

    \I__5139\ : Span4Mux_h
    port map (
            O => \N__23711\,
            I => \N__23707\
        );

    \I__5138\ : InMux
    port map (
            O => \N__23710\,
            I => \N__23704\
        );

    \I__5137\ : Span4Mux_h
    port map (
            O => \N__23707\,
            I => \N__23698\
        );

    \I__5136\ : LocalMux
    port map (
            O => \N__23704\,
            I => \N__23698\
        );

    \I__5135\ : InMux
    port map (
            O => \N__23703\,
            I => \N__23695\
        );

    \I__5134\ : Span4Mux_h
    port map (
            O => \N__23698\,
            I => \N__23692\
        );

    \I__5133\ : LocalMux
    port map (
            O => \N__23695\,
            I => \eeprom.delay_counter_4\
        );

    \I__5132\ : Odrv4
    port map (
            O => \N__23692\,
            I => \eeprom.delay_counter_4\
        );

    \I__5131\ : CascadeMux
    port map (
            O => \N__23687\,
            I => \N__23684\
        );

    \I__5130\ : InMux
    port map (
            O => \N__23684\,
            I => \N__23681\
        );

    \I__5129\ : LocalMux
    port map (
            O => \N__23681\,
            I => \N__23678\
        );

    \I__5128\ : Odrv4
    port map (
            O => \N__23678\,
            I => \eeprom.n3721_adj_434\
        );

    \I__5127\ : InMux
    port map (
            O => \N__23675\,
            I => \eeprom.n3775\
        );

    \I__5126\ : InMux
    port map (
            O => \N__23672\,
            I => \N__23669\
        );

    \I__5125\ : LocalMux
    port map (
            O => \N__23669\,
            I => \N__23666\
        );

    \I__5124\ : Span4Mux_h
    port map (
            O => \N__23666\,
            I => \N__23662\
        );

    \I__5123\ : InMux
    port map (
            O => \N__23665\,
            I => \N__23659\
        );

    \I__5122\ : Span4Mux_h
    port map (
            O => \N__23662\,
            I => \N__23653\
        );

    \I__5121\ : LocalMux
    port map (
            O => \N__23659\,
            I => \N__23653\
        );

    \I__5120\ : CascadeMux
    port map (
            O => \N__23658\,
            I => \N__23650\
        );

    \I__5119\ : Span4Mux_h
    port map (
            O => \N__23653\,
            I => \N__23646\
        );

    \I__5118\ : InMux
    port map (
            O => \N__23650\,
            I => \N__23643\
        );

    \I__5117\ : InMux
    port map (
            O => \N__23649\,
            I => \N__23640\
        );

    \I__5116\ : Span4Mux_h
    port map (
            O => \N__23646\,
            I => \N__23635\
        );

    \I__5115\ : LocalMux
    port map (
            O => \N__23643\,
            I => \N__23635\
        );

    \I__5114\ : LocalMux
    port map (
            O => \N__23640\,
            I => \eeprom.delay_counter_5\
        );

    \I__5113\ : Odrv4
    port map (
            O => \N__23635\,
            I => \eeprom.delay_counter_5\
        );

    \I__5112\ : InMux
    port map (
            O => \N__23630\,
            I => \N__23627\
        );

    \I__5111\ : LocalMux
    port map (
            O => \N__23627\,
            I => \N__23624\
        );

    \I__5110\ : Odrv12
    port map (
            O => \N__23624\,
            I => \eeprom.n3720_adj_435\
        );

    \I__5109\ : InMux
    port map (
            O => \N__23621\,
            I => \eeprom.n3776\
        );

    \I__5108\ : InMux
    port map (
            O => \N__23618\,
            I => \N__23615\
        );

    \I__5107\ : LocalMux
    port map (
            O => \N__23615\,
            I => \N__23612\
        );

    \I__5106\ : Span4Mux_h
    port map (
            O => \N__23612\,
            I => \N__23608\
        );

    \I__5105\ : InMux
    port map (
            O => \N__23611\,
            I => \N__23605\
        );

    \I__5104\ : Span4Mux_h
    port map (
            O => \N__23608\,
            I => \N__23600\
        );

    \I__5103\ : LocalMux
    port map (
            O => \N__23605\,
            I => \N__23600\
        );

    \I__5102\ : Span4Mux_h
    port map (
            O => \N__23600\,
            I => \N__23596\
        );

    \I__5101\ : InMux
    port map (
            O => \N__23599\,
            I => \N__23592\
        );

    \I__5100\ : Span4Mux_h
    port map (
            O => \N__23596\,
            I => \N__23589\
        );

    \I__5099\ : InMux
    port map (
            O => \N__23595\,
            I => \N__23586\
        );

    \I__5098\ : LocalMux
    port map (
            O => \N__23592\,
            I => \eeprom.delay_counter_6\
        );

    \I__5097\ : Odrv4
    port map (
            O => \N__23589\,
            I => \eeprom.delay_counter_6\
        );

    \I__5096\ : LocalMux
    port map (
            O => \N__23586\,
            I => \eeprom.delay_counter_6\
        );

    \I__5095\ : CascadeMux
    port map (
            O => \N__23579\,
            I => \N__23576\
        );

    \I__5094\ : InMux
    port map (
            O => \N__23576\,
            I => \N__23573\
        );

    \I__5093\ : LocalMux
    port map (
            O => \N__23573\,
            I => \N__23570\
        );

    \I__5092\ : Span12Mux_h
    port map (
            O => \N__23570\,
            I => \N__23567\
        );

    \I__5091\ : Odrv12
    port map (
            O => \N__23567\,
            I => \eeprom.n3719_adj_436\
        );

    \I__5090\ : InMux
    port map (
            O => \N__23564\,
            I => \eeprom.n3777\
        );

    \I__5089\ : InMux
    port map (
            O => \N__23561\,
            I => \eeprom.n3778\
        );

    \I__5088\ : InMux
    port map (
            O => \N__23558\,
            I => \bfn_15_21_0_\
        );

    \I__5087\ : CascadeMux
    port map (
            O => \N__23555\,
            I => \eeprom.n3617_adj_346_cascade_\
        );

    \I__5086\ : InMux
    port map (
            O => \N__23552\,
            I => \N__23549\
        );

    \I__5085\ : LocalMux
    port map (
            O => \N__23549\,
            I => \eeprom.n4619\
        );

    \I__5084\ : CascadeMux
    port map (
            O => \N__23546\,
            I => \eeprom.n4427_cascade_\
        );

    \I__5083\ : InMux
    port map (
            O => \N__23543\,
            I => \N__23540\
        );

    \I__5082\ : LocalMux
    port map (
            O => \N__23540\,
            I => \eeprom.n3596_adj_454\
        );

    \I__5081\ : CascadeMux
    port map (
            O => \N__23537\,
            I => \eeprom.n28_adj_455_cascade_\
        );

    \I__5080\ : InMux
    port map (
            O => \N__23534\,
            I => \N__23531\
        );

    \I__5079\ : LocalMux
    port map (
            O => \N__23531\,
            I => \eeprom.n4567\
        );

    \I__5078\ : CascadeMux
    port map (
            O => \N__23528\,
            I => \eeprom.n3628_adj_437_cascade_\
        );

    \I__5077\ : CascadeMux
    port map (
            O => \N__23525\,
            I => \eeprom.n3716_adj_439_cascade_\
        );

    \I__5076\ : InMux
    port map (
            O => \N__23522\,
            I => \N__23519\
        );

    \I__5075\ : LocalMux
    port map (
            O => \N__23519\,
            I => \eeprom.n3605_adj_453\
        );

    \I__5074\ : CascadeMux
    port map (
            O => \N__23516\,
            I => \eeprom.n3618_adj_350_cascade_\
        );

    \I__5073\ : InMux
    port map (
            O => \N__23513\,
            I => \N__23510\
        );

    \I__5072\ : LocalMux
    port map (
            O => \N__23510\,
            I => \eeprom.n4623\
        );

    \I__5071\ : InMux
    port map (
            O => \N__23507\,
            I => \N__23504\
        );

    \I__5070\ : LocalMux
    port map (
            O => \N__23504\,
            I => \eeprom.n4425\
        );

    \I__5069\ : InMux
    port map (
            O => \N__23501\,
            I => \N__23498\
        );

    \I__5068\ : LocalMux
    port map (
            O => \N__23498\,
            I => \N__23495\
        );

    \I__5067\ : Span4Mux_v
    port map (
            O => \N__23495\,
            I => \N__23492\
        );

    \I__5066\ : Span4Mux_h
    port map (
            O => \N__23492\,
            I => \N__23489\
        );

    \I__5065\ : Span4Mux_h
    port map (
            O => \N__23489\,
            I => \N__23485\
        );

    \I__5064\ : InMux
    port map (
            O => \N__23488\,
            I => \N__23482\
        );

    \I__5063\ : Span4Mux_h
    port map (
            O => \N__23485\,
            I => \N__23476\
        );

    \I__5062\ : LocalMux
    port map (
            O => \N__23482\,
            I => \N__23476\
        );

    \I__5061\ : InMux
    port map (
            O => \N__23481\,
            I => \N__23472\
        );

    \I__5060\ : Span4Mux_v
    port map (
            O => \N__23476\,
            I => \N__23469\
        );

    \I__5059\ : InMux
    port map (
            O => \N__23475\,
            I => \N__23466\
        );

    \I__5058\ : LocalMux
    port map (
            O => \N__23472\,
            I => \eeprom.delay_counter_0\
        );

    \I__5057\ : Odrv4
    port map (
            O => \N__23469\,
            I => \eeprom.delay_counter_0\
        );

    \I__5056\ : LocalMux
    port map (
            O => \N__23466\,
            I => \eeprom.delay_counter_0\
        );

    \I__5055\ : CascadeMux
    port map (
            O => \N__23459\,
            I => \N__23456\
        );

    \I__5054\ : InMux
    port map (
            O => \N__23456\,
            I => \N__23453\
        );

    \I__5053\ : LocalMux
    port map (
            O => \N__23453\,
            I => \N__23450\
        );

    \I__5052\ : Span12Mux_v
    port map (
            O => \N__23450\,
            I => \N__23447\
        );

    \I__5051\ : Span12Mux_h
    port map (
            O => \N__23447\,
            I => \N__23444\
        );

    \I__5050\ : Odrv12
    port map (
            O => \N__23444\,
            I => \eeprom.n1166\
        );

    \I__5049\ : InMux
    port map (
            O => \N__23441\,
            I => \bfn_15_20_0_\
        );

    \I__5048\ : CascadeMux
    port map (
            O => \N__23438\,
            I => \eeprom.n3515_adj_370_cascade_\
        );

    \I__5047\ : CascadeMux
    port map (
            O => \N__23435\,
            I => \N__23432\
        );

    \I__5046\ : InMux
    port map (
            O => \N__23432\,
            I => \N__23429\
        );

    \I__5045\ : LocalMux
    port map (
            O => \N__23429\,
            I => \eeprom.n4727\
        );

    \I__5044\ : InMux
    port map (
            O => \N__23426\,
            I => \N__23422\
        );

    \I__5043\ : InMux
    port map (
            O => \N__23425\,
            I => \N__23418\
        );

    \I__5042\ : LocalMux
    port map (
            O => \N__23422\,
            I => \N__23415\
        );

    \I__5041\ : InMux
    port map (
            O => \N__23421\,
            I => \N__23412\
        );

    \I__5040\ : LocalMux
    port map (
            O => \N__23418\,
            I => \N__23409\
        );

    \I__5039\ : Span12Mux_v
    port map (
            O => \N__23415\,
            I => \N__23406\
        );

    \I__5038\ : LocalMux
    port map (
            O => \N__23412\,
            I => \N__23403\
        );

    \I__5037\ : Span4Mux_v
    port map (
            O => \N__23409\,
            I => \N__23400\
        );

    \I__5036\ : Span12Mux_h
    port map (
            O => \N__23406\,
            I => \N__23397\
        );

    \I__5035\ : Span12Mux_v
    port map (
            O => \N__23403\,
            I => \N__23392\
        );

    \I__5034\ : Sp12to4
    port map (
            O => \N__23400\,
            I => \N__23392\
        );

    \I__5033\ : Odrv12
    port map (
            O => \N__23397\,
            I => \eeprom.n3419\
        );

    \I__5032\ : Odrv12
    port map (
            O => \N__23392\,
            I => \eeprom.n3419\
        );

    \I__5031\ : InMux
    port map (
            O => \N__23387\,
            I => \N__23384\
        );

    \I__5030\ : LocalMux
    port map (
            O => \N__23384\,
            I => \eeprom.n3486\
        );

    \I__5029\ : InMux
    port map (
            O => \N__23381\,
            I => \N__23378\
        );

    \I__5028\ : LocalMux
    port map (
            O => \N__23378\,
            I => \eeprom.n3471_adj_386\
        );

    \I__5027\ : CascadeMux
    port map (
            O => \N__23375\,
            I => \N__23366\
        );

    \I__5026\ : InMux
    port map (
            O => \N__23374\,
            I => \N__23354\
        );

    \I__5025\ : InMux
    port map (
            O => \N__23373\,
            I => \N__23354\
        );

    \I__5024\ : InMux
    port map (
            O => \N__23372\,
            I => \N__23354\
        );

    \I__5023\ : CascadeMux
    port map (
            O => \N__23371\,
            I => \N__23349\
        );

    \I__5022\ : CascadeMux
    port map (
            O => \N__23370\,
            I => \N__23342\
        );

    \I__5021\ : CascadeMux
    port map (
            O => \N__23369\,
            I => \N__23338\
        );

    \I__5020\ : InMux
    port map (
            O => \N__23366\,
            I => \N__23333\
        );

    \I__5019\ : InMux
    port map (
            O => \N__23365\,
            I => \N__23333\
        );

    \I__5018\ : CascadeMux
    port map (
            O => \N__23364\,
            I => \N__23328\
        );

    \I__5017\ : CascadeMux
    port map (
            O => \N__23363\,
            I => \N__23325\
        );

    \I__5016\ : InMux
    port map (
            O => \N__23362\,
            I => \N__23319\
        );

    \I__5015\ : InMux
    port map (
            O => \N__23361\,
            I => \N__23319\
        );

    \I__5014\ : LocalMux
    port map (
            O => \N__23354\,
            I => \N__23316\
        );

    \I__5013\ : InMux
    port map (
            O => \N__23353\,
            I => \N__23313\
        );

    \I__5012\ : InMux
    port map (
            O => \N__23352\,
            I => \N__23306\
        );

    \I__5011\ : InMux
    port map (
            O => \N__23349\,
            I => \N__23306\
        );

    \I__5010\ : InMux
    port map (
            O => \N__23348\,
            I => \N__23306\
        );

    \I__5009\ : InMux
    port map (
            O => \N__23347\,
            I => \N__23299\
        );

    \I__5008\ : InMux
    port map (
            O => \N__23346\,
            I => \N__23299\
        );

    \I__5007\ : InMux
    port map (
            O => \N__23345\,
            I => \N__23299\
        );

    \I__5006\ : InMux
    port map (
            O => \N__23342\,
            I => \N__23294\
        );

    \I__5005\ : InMux
    port map (
            O => \N__23341\,
            I => \N__23294\
        );

    \I__5004\ : InMux
    port map (
            O => \N__23338\,
            I => \N__23291\
        );

    \I__5003\ : LocalMux
    port map (
            O => \N__23333\,
            I => \N__23288\
        );

    \I__5002\ : InMux
    port map (
            O => \N__23332\,
            I => \N__23277\
        );

    \I__5001\ : InMux
    port map (
            O => \N__23331\,
            I => \N__23277\
        );

    \I__5000\ : InMux
    port map (
            O => \N__23328\,
            I => \N__23277\
        );

    \I__4999\ : InMux
    port map (
            O => \N__23325\,
            I => \N__23277\
        );

    \I__4998\ : InMux
    port map (
            O => \N__23324\,
            I => \N__23277\
        );

    \I__4997\ : LocalMux
    port map (
            O => \N__23319\,
            I => \N__23272\
        );

    \I__4996\ : Span4Mux_h
    port map (
            O => \N__23316\,
            I => \N__23272\
        );

    \I__4995\ : LocalMux
    port map (
            O => \N__23313\,
            I => \eeprom.n3430\
        );

    \I__4994\ : LocalMux
    port map (
            O => \N__23306\,
            I => \eeprom.n3430\
        );

    \I__4993\ : LocalMux
    port map (
            O => \N__23299\,
            I => \eeprom.n3430\
        );

    \I__4992\ : LocalMux
    port map (
            O => \N__23294\,
            I => \eeprom.n3430\
        );

    \I__4991\ : LocalMux
    port map (
            O => \N__23291\,
            I => \eeprom.n3430\
        );

    \I__4990\ : Odrv4
    port map (
            O => \N__23288\,
            I => \eeprom.n3430\
        );

    \I__4989\ : LocalMux
    port map (
            O => \N__23277\,
            I => \eeprom.n3430\
        );

    \I__4988\ : Odrv4
    port map (
            O => \N__23272\,
            I => \eeprom.n3430\
        );

    \I__4987\ : CascadeMux
    port map (
            O => \N__23255\,
            I => \N__23251\
        );

    \I__4986\ : InMux
    port map (
            O => \N__23254\,
            I => \N__23248\
        );

    \I__4985\ : InMux
    port map (
            O => \N__23251\,
            I => \N__23245\
        );

    \I__4984\ : LocalMux
    port map (
            O => \N__23248\,
            I => \N__23239\
        );

    \I__4983\ : LocalMux
    port map (
            O => \N__23245\,
            I => \N__23239\
        );

    \I__4982\ : InMux
    port map (
            O => \N__23244\,
            I => \N__23236\
        );

    \I__4981\ : Odrv12
    port map (
            O => \N__23239\,
            I => \eeprom.n3404\
        );

    \I__4980\ : LocalMux
    port map (
            O => \N__23236\,
            I => \eeprom.n3404\
        );

    \I__4979\ : CascadeMux
    port map (
            O => \N__23231\,
            I => \eeprom.n3615_adj_344_cascade_\
        );

    \I__4978\ : CascadeMux
    port map (
            O => \N__23228\,
            I => \eeprom.n3714_adj_442_cascade_\
        );

    \I__4977\ : CascadeMux
    port map (
            O => \N__23225\,
            I => \eeprom.n3034_cascade_\
        );

    \I__4976\ : InMux
    port map (
            O => \N__23222\,
            I => \N__23217\
        );

    \I__4975\ : InMux
    port map (
            O => \N__23221\,
            I => \N__23214\
        );

    \I__4974\ : InMux
    port map (
            O => \N__23220\,
            I => \N__23211\
        );

    \I__4973\ : LocalMux
    port map (
            O => \N__23217\,
            I => \N__23208\
        );

    \I__4972\ : LocalMux
    port map (
            O => \N__23214\,
            I => \N__23205\
        );

    \I__4971\ : LocalMux
    port map (
            O => \N__23211\,
            I => \N__23202\
        );

    \I__4970\ : Span4Mux_h
    port map (
            O => \N__23208\,
            I => \N__23199\
        );

    \I__4969\ : Span4Mux_v
    port map (
            O => \N__23205\,
            I => \N__23194\
        );

    \I__4968\ : Span4Mux_h
    port map (
            O => \N__23202\,
            I => \N__23194\
        );

    \I__4967\ : Odrv4
    port map (
            O => \N__23199\,
            I => \eeprom.n3112\
        );

    \I__4966\ : Odrv4
    port map (
            O => \N__23194\,
            I => \eeprom.n3112\
        );

    \I__4965\ : InMux
    port map (
            O => \N__23189\,
            I => \N__23185\
        );

    \I__4964\ : CascadeMux
    port map (
            O => \N__23188\,
            I => \N__23182\
        );

    \I__4963\ : LocalMux
    port map (
            O => \N__23185\,
            I => \N__23179\
        );

    \I__4962\ : InMux
    port map (
            O => \N__23182\,
            I => \N__23175\
        );

    \I__4961\ : Span4Mux_v
    port map (
            O => \N__23179\,
            I => \N__23172\
        );

    \I__4960\ : InMux
    port map (
            O => \N__23178\,
            I => \N__23169\
        );

    \I__4959\ : LocalMux
    port map (
            O => \N__23175\,
            I => \N__23166\
        );

    \I__4958\ : Odrv4
    port map (
            O => \N__23172\,
            I => \eeprom.n2912\
        );

    \I__4957\ : LocalMux
    port map (
            O => \N__23169\,
            I => \eeprom.n2912\
        );

    \I__4956\ : Odrv4
    port map (
            O => \N__23166\,
            I => \eeprom.n2912\
        );

    \I__4955\ : CascadeMux
    port map (
            O => \N__23159\,
            I => \N__23156\
        );

    \I__4954\ : InMux
    port map (
            O => \N__23156\,
            I => \N__23153\
        );

    \I__4953\ : LocalMux
    port map (
            O => \N__23153\,
            I => \N__23150\
        );

    \I__4952\ : Span4Mux_h
    port map (
            O => \N__23150\,
            I => \N__23147\
        );

    \I__4951\ : Odrv4
    port map (
            O => \N__23147\,
            I => \eeprom.n2979\
        );

    \I__4950\ : InMux
    port map (
            O => \N__23144\,
            I => \N__23141\
        );

    \I__4949\ : LocalMux
    port map (
            O => \N__23141\,
            I => \N__23136\
        );

    \I__4948\ : InMux
    port map (
            O => \N__23140\,
            I => \N__23131\
        );

    \I__4947\ : InMux
    port map (
            O => \N__23139\,
            I => \N__23131\
        );

    \I__4946\ : Odrv4
    port map (
            O => \N__23136\,
            I => \eeprom.n3103\
        );

    \I__4945\ : LocalMux
    port map (
            O => \N__23131\,
            I => \eeprom.n3103\
        );

    \I__4944\ : InMux
    port map (
            O => \N__23126\,
            I => \N__23123\
        );

    \I__4943\ : LocalMux
    port map (
            O => \N__23123\,
            I => \N__23120\
        );

    \I__4942\ : Span4Mux_h
    port map (
            O => \N__23120\,
            I => \N__23117\
        );

    \I__4941\ : Odrv4
    port map (
            O => \N__23117\,
            I => \eeprom.n4137\
        );

    \I__4940\ : InMux
    port map (
            O => \N__23114\,
            I => \N__23110\
        );

    \I__4939\ : CascadeMux
    port map (
            O => \N__23113\,
            I => \N__23107\
        );

    \I__4938\ : LocalMux
    port map (
            O => \N__23110\,
            I => \N__23103\
        );

    \I__4937\ : InMux
    port map (
            O => \N__23107\,
            I => \N__23100\
        );

    \I__4936\ : InMux
    port map (
            O => \N__23106\,
            I => \N__23097\
        );

    \I__4935\ : Span4Mux_h
    port map (
            O => \N__23103\,
            I => \N__23092\
        );

    \I__4934\ : LocalMux
    port map (
            O => \N__23100\,
            I => \N__23092\
        );

    \I__4933\ : LocalMux
    port map (
            O => \N__23097\,
            I => \eeprom.n3417\
        );

    \I__4932\ : Odrv4
    port map (
            O => \N__23092\,
            I => \eeprom.n3417\
        );

    \I__4931\ : CascadeMux
    port map (
            O => \N__23087\,
            I => \N__23084\
        );

    \I__4930\ : InMux
    port map (
            O => \N__23084\,
            I => \N__23081\
        );

    \I__4929\ : LocalMux
    port map (
            O => \N__23081\,
            I => \eeprom.n3484_adj_406\
        );

    \I__4928\ : CascadeMux
    port map (
            O => \N__23078\,
            I => \N__23074\
        );

    \I__4927\ : InMux
    port map (
            O => \N__23077\,
            I => \N__23070\
        );

    \I__4926\ : InMux
    port map (
            O => \N__23074\,
            I => \N__23067\
        );

    \I__4925\ : InMux
    port map (
            O => \N__23073\,
            I => \N__23064\
        );

    \I__4924\ : LocalMux
    port map (
            O => \N__23070\,
            I => \N__23059\
        );

    \I__4923\ : LocalMux
    port map (
            O => \N__23067\,
            I => \N__23059\
        );

    \I__4922\ : LocalMux
    port map (
            O => \N__23064\,
            I => \eeprom.n3418\
        );

    \I__4921\ : Odrv4
    port map (
            O => \N__23059\,
            I => \eeprom.n3418\
        );

    \I__4920\ : CascadeMux
    port map (
            O => \N__23054\,
            I => \N__23051\
        );

    \I__4919\ : InMux
    port map (
            O => \N__23051\,
            I => \N__23048\
        );

    \I__4918\ : LocalMux
    port map (
            O => \N__23048\,
            I => \eeprom.n3485\
        );

    \I__4917\ : CascadeMux
    port map (
            O => \N__23045\,
            I => \eeprom.n3517_adj_374_cascade_\
        );

    \I__4916\ : InMux
    port map (
            O => \N__23042\,
            I => \N__23039\
        );

    \I__4915\ : LocalMux
    port map (
            O => \N__23039\,
            I => \eeprom.n4729\
        );

    \I__4914\ : CascadeMux
    port map (
            O => \N__23036\,
            I => \N__23032\
        );

    \I__4913\ : InMux
    port map (
            O => \N__23035\,
            I => \N__23028\
        );

    \I__4912\ : InMux
    port map (
            O => \N__23032\,
            I => \N__23025\
        );

    \I__4911\ : InMux
    port map (
            O => \N__23031\,
            I => \N__23022\
        );

    \I__4910\ : LocalMux
    port map (
            O => \N__23028\,
            I => \N__23017\
        );

    \I__4909\ : LocalMux
    port map (
            O => \N__23025\,
            I => \N__23017\
        );

    \I__4908\ : LocalMux
    port map (
            O => \N__23022\,
            I => \eeprom.n3416\
        );

    \I__4907\ : Odrv12
    port map (
            O => \N__23017\,
            I => \eeprom.n3416\
        );

    \I__4906\ : CascadeMux
    port map (
            O => \N__23012\,
            I => \N__23009\
        );

    \I__4905\ : InMux
    port map (
            O => \N__23009\,
            I => \N__23006\
        );

    \I__4904\ : LocalMux
    port map (
            O => \N__23006\,
            I => \eeprom.n3483_adj_404\
        );

    \I__4903\ : InMux
    port map (
            O => \N__23003\,
            I => \N__23000\
        );

    \I__4902\ : LocalMux
    port map (
            O => \N__23000\,
            I => \N__22997\
        );

    \I__4901\ : Span12Mux_h
    port map (
            O => \N__22997\,
            I => \N__22994\
        );

    \I__4900\ : Odrv12
    port map (
            O => \N__22994\,
            I => \eeprom.n31_adj_476\
        );

    \I__4899\ : InMux
    port map (
            O => \N__22991\,
            I => \N__22987\
        );

    \I__4898\ : InMux
    port map (
            O => \N__22990\,
            I => \N__22984\
        );

    \I__4897\ : LocalMux
    port map (
            O => \N__22987\,
            I => \N__22980\
        );

    \I__4896\ : LocalMux
    port map (
            O => \N__22984\,
            I => \N__22974\
        );

    \I__4895\ : InMux
    port map (
            O => \N__22983\,
            I => \N__22971\
        );

    \I__4894\ : Span4Mux_v
    port map (
            O => \N__22980\,
            I => \N__22966\
        );

    \I__4893\ : InMux
    port map (
            O => \N__22979\,
            I => \N__22963\
        );

    \I__4892\ : InMux
    port map (
            O => \N__22978\,
            I => \N__22960\
        );

    \I__4891\ : InMux
    port map (
            O => \N__22977\,
            I => \N__22951\
        );

    \I__4890\ : Span4Mux_h
    port map (
            O => \N__22974\,
            I => \N__22944\
        );

    \I__4889\ : LocalMux
    port map (
            O => \N__22971\,
            I => \N__22944\
        );

    \I__4888\ : InMux
    port map (
            O => \N__22970\,
            I => \N__22939\
        );

    \I__4887\ : InMux
    port map (
            O => \N__22969\,
            I => \N__22935\
        );

    \I__4886\ : Span4Mux_h
    port map (
            O => \N__22966\,
            I => \N__22930\
        );

    \I__4885\ : LocalMux
    port map (
            O => \N__22963\,
            I => \N__22930\
        );

    \I__4884\ : LocalMux
    port map (
            O => \N__22960\,
            I => \N__22927\
        );

    \I__4883\ : InMux
    port map (
            O => \N__22959\,
            I => \N__22924\
        );

    \I__4882\ : InMux
    port map (
            O => \N__22958\,
            I => \N__22917\
        );

    \I__4881\ : InMux
    port map (
            O => \N__22957\,
            I => \N__22912\
        );

    \I__4880\ : InMux
    port map (
            O => \N__22956\,
            I => \N__22912\
        );

    \I__4879\ : InMux
    port map (
            O => \N__22955\,
            I => \N__22907\
        );

    \I__4878\ : InMux
    port map (
            O => \N__22954\,
            I => \N__22907\
        );

    \I__4877\ : LocalMux
    port map (
            O => \N__22951\,
            I => \N__22903\
        );

    \I__4876\ : InMux
    port map (
            O => \N__22950\,
            I => \N__22898\
        );

    \I__4875\ : InMux
    port map (
            O => \N__22949\,
            I => \N__22898\
        );

    \I__4874\ : Span4Mux_v
    port map (
            O => \N__22944\,
            I => \N__22895\
        );

    \I__4873\ : InMux
    port map (
            O => \N__22943\,
            I => \N__22892\
        );

    \I__4872\ : InMux
    port map (
            O => \N__22942\,
            I => \N__22889\
        );

    \I__4871\ : LocalMux
    port map (
            O => \N__22939\,
            I => \N__22885\
        );

    \I__4870\ : InMux
    port map (
            O => \N__22938\,
            I => \N__22882\
        );

    \I__4869\ : LocalMux
    port map (
            O => \N__22935\,
            I => \N__22879\
        );

    \I__4868\ : Span4Mux_h
    port map (
            O => \N__22930\,
            I => \N__22874\
        );

    \I__4867\ : Span4Mux_v
    port map (
            O => \N__22927\,
            I => \N__22874\
        );

    \I__4866\ : LocalMux
    port map (
            O => \N__22924\,
            I => \N__22871\
        );

    \I__4865\ : InMux
    port map (
            O => \N__22923\,
            I => \N__22862\
        );

    \I__4864\ : InMux
    port map (
            O => \N__22922\,
            I => \N__22862\
        );

    \I__4863\ : InMux
    port map (
            O => \N__22921\,
            I => \N__22862\
        );

    \I__4862\ : InMux
    port map (
            O => \N__22920\,
            I => \N__22862\
        );

    \I__4861\ : LocalMux
    port map (
            O => \N__22917\,
            I => \N__22855\
        );

    \I__4860\ : LocalMux
    port map (
            O => \N__22912\,
            I => \N__22855\
        );

    \I__4859\ : LocalMux
    port map (
            O => \N__22907\,
            I => \N__22855\
        );

    \I__4858\ : InMux
    port map (
            O => \N__22906\,
            I => \N__22842\
        );

    \I__4857\ : Span12Mux_h
    port map (
            O => \N__22903\,
            I => \N__22831\
        );

    \I__4856\ : LocalMux
    port map (
            O => \N__22898\,
            I => \N__22831\
        );

    \I__4855\ : Sp12to4
    port map (
            O => \N__22895\,
            I => \N__22831\
        );

    \I__4854\ : LocalMux
    port map (
            O => \N__22892\,
            I => \N__22831\
        );

    \I__4853\ : LocalMux
    port map (
            O => \N__22889\,
            I => \N__22831\
        );

    \I__4852\ : InMux
    port map (
            O => \N__22888\,
            I => \N__22828\
        );

    \I__4851\ : Span4Mux_v
    port map (
            O => \N__22885\,
            I => \N__22819\
        );

    \I__4850\ : LocalMux
    port map (
            O => \N__22882\,
            I => \N__22819\
        );

    \I__4849\ : Span4Mux_v
    port map (
            O => \N__22879\,
            I => \N__22819\
        );

    \I__4848\ : Span4Mux_h
    port map (
            O => \N__22874\,
            I => \N__22819\
        );

    \I__4847\ : Span4Mux_h
    port map (
            O => \N__22871\,
            I => \N__22812\
        );

    \I__4846\ : LocalMux
    port map (
            O => \N__22862\,
            I => \N__22812\
        );

    \I__4845\ : Span4Mux_h
    port map (
            O => \N__22855\,
            I => \N__22812\
        );

    \I__4844\ : InMux
    port map (
            O => \N__22854\,
            I => \N__22803\
        );

    \I__4843\ : InMux
    port map (
            O => \N__22853\,
            I => \N__22803\
        );

    \I__4842\ : InMux
    port map (
            O => \N__22852\,
            I => \N__22803\
        );

    \I__4841\ : InMux
    port map (
            O => \N__22851\,
            I => \N__22803\
        );

    \I__4840\ : InMux
    port map (
            O => \N__22850\,
            I => \N__22794\
        );

    \I__4839\ : InMux
    port map (
            O => \N__22849\,
            I => \N__22794\
        );

    \I__4838\ : InMux
    port map (
            O => \N__22848\,
            I => \N__22794\
        );

    \I__4837\ : InMux
    port map (
            O => \N__22847\,
            I => \N__22794\
        );

    \I__4836\ : InMux
    port map (
            O => \N__22846\,
            I => \N__22789\
        );

    \I__4835\ : InMux
    port map (
            O => \N__22845\,
            I => \N__22789\
        );

    \I__4834\ : LocalMux
    port map (
            O => \N__22842\,
            I => \eeprom.delay_counter_31\
        );

    \I__4833\ : Odrv12
    port map (
            O => \N__22831\,
            I => \eeprom.delay_counter_31\
        );

    \I__4832\ : LocalMux
    port map (
            O => \N__22828\,
            I => \eeprom.delay_counter_31\
        );

    \I__4831\ : Odrv4
    port map (
            O => \N__22819\,
            I => \eeprom.delay_counter_31\
        );

    \I__4830\ : Odrv4
    port map (
            O => \N__22812\,
            I => \eeprom.delay_counter_31\
        );

    \I__4829\ : LocalMux
    port map (
            O => \N__22803\,
            I => \eeprom.delay_counter_31\
        );

    \I__4828\ : LocalMux
    port map (
            O => \N__22794\,
            I => \eeprom.delay_counter_31\
        );

    \I__4827\ : LocalMux
    port map (
            O => \N__22789\,
            I => \eeprom.delay_counter_31\
        );

    \I__4826\ : InMux
    port map (
            O => \N__22772\,
            I => \N__22769\
        );

    \I__4825\ : LocalMux
    port map (
            O => \N__22769\,
            I => \N__22766\
        );

    \I__4824\ : Span4Mux_h
    port map (
            O => \N__22766\,
            I => \N__22763\
        );

    \I__4823\ : Odrv4
    port map (
            O => \N__22763\,
            I => \eeprom.n24_adj_459\
        );

    \I__4822\ : CascadeMux
    port map (
            O => \N__22760\,
            I => \eeprom.n4559_cascade_\
        );

    \I__4821\ : CascadeMux
    port map (
            O => \N__22757\,
            I => \eeprom.n4563_cascade_\
        );

    \I__4820\ : InMux
    port map (
            O => \N__22754\,
            I => \N__22751\
        );

    \I__4819\ : LocalMux
    port map (
            O => \N__22751\,
            I => \eeprom.n21_adj_422\
        );

    \I__4818\ : CascadeMux
    port map (
            O => \N__22748\,
            I => \eeprom.n17_adj_421_cascade_\
        );

    \I__4817\ : CascadeMux
    port map (
            O => \N__22745\,
            I => \eeprom.n24_cascade_\
        );

    \I__4816\ : InMux
    port map (
            O => \N__22742\,
            I => \N__22739\
        );

    \I__4815\ : LocalMux
    port map (
            O => \N__22739\,
            I => \eeprom.n20_adj_423\
        );

    \I__4814\ : InMux
    port map (
            O => \N__22736\,
            I => \eeprom.n3747\
        );

    \I__4813\ : InMux
    port map (
            O => \N__22733\,
            I => \N__22729\
        );

    \I__4812\ : InMux
    port map (
            O => \N__22732\,
            I => \N__22726\
        );

    \I__4811\ : LocalMux
    port map (
            O => \N__22729\,
            I => \N__22723\
        );

    \I__4810\ : LocalMux
    port map (
            O => \N__22726\,
            I => \N__22720\
        );

    \I__4809\ : Span4Mux_h
    port map (
            O => \N__22723\,
            I => \N__22715\
        );

    \I__4808\ : Span4Mux_v
    port map (
            O => \N__22720\,
            I => \N__22715\
        );

    \I__4807\ : Odrv4
    port map (
            O => \N__22715\,
            I => \eeprom.n3397\
        );

    \I__4806\ : InMux
    port map (
            O => \N__22712\,
            I => \eeprom.n3748\
        );

    \I__4805\ : CascadeMux
    port map (
            O => \N__22709\,
            I => \N__22706\
        );

    \I__4804\ : InMux
    port map (
            O => \N__22706\,
            I => \N__22703\
        );

    \I__4803\ : LocalMux
    port map (
            O => \N__22703\,
            I => \eeprom.n4583\
        );

    \I__4802\ : CascadeMux
    port map (
            O => \N__22700\,
            I => \eeprom.n31_cascade_\
        );

    \I__4801\ : InMux
    port map (
            O => \N__22697\,
            I => \N__22694\
        );

    \I__4800\ : LocalMux
    port map (
            O => \N__22694\,
            I => \eeprom.n4433\
        );

    \I__4799\ : InMux
    port map (
            O => \N__22691\,
            I => \N__22688\
        );

    \I__4798\ : LocalMux
    port map (
            O => \N__22688\,
            I => \eeprom.n3598_adj_452\
        );

    \I__4797\ : CascadeMux
    port map (
            O => \N__22685\,
            I => \N__22681\
        );

    \I__4796\ : InMux
    port map (
            O => \N__22684\,
            I => \N__22678\
        );

    \I__4795\ : InMux
    port map (
            O => \N__22681\,
            I => \N__22675\
        );

    \I__4794\ : LocalMux
    port map (
            O => \N__22678\,
            I => \N__22669\
        );

    \I__4793\ : LocalMux
    port map (
            O => \N__22675\,
            I => \N__22669\
        );

    \I__4792\ : InMux
    port map (
            O => \N__22674\,
            I => \N__22666\
        );

    \I__4791\ : Odrv4
    port map (
            O => \N__22669\,
            I => \eeprom.n3405\
        );

    \I__4790\ : LocalMux
    port map (
            O => \N__22666\,
            I => \eeprom.n3405\
        );

    \I__4789\ : InMux
    port map (
            O => \N__22661\,
            I => \N__22658\
        );

    \I__4788\ : LocalMux
    port map (
            O => \N__22658\,
            I => \N__22655\
        );

    \I__4787\ : Odrv4
    port map (
            O => \N__22655\,
            I => \eeprom.n3472_adj_387\
        );

    \I__4786\ : InMux
    port map (
            O => \N__22652\,
            I => \eeprom.n3740\
        );

    \I__4785\ : InMux
    port map (
            O => \N__22649\,
            I => \eeprom.n3741\
        );

    \I__4784\ : CascadeMux
    port map (
            O => \N__22646\,
            I => \N__22642\
        );

    \I__4783\ : InMux
    port map (
            O => \N__22645\,
            I => \N__22639\
        );

    \I__4782\ : InMux
    port map (
            O => \N__22642\,
            I => \N__22636\
        );

    \I__4781\ : LocalMux
    port map (
            O => \N__22639\,
            I => \N__22630\
        );

    \I__4780\ : LocalMux
    port map (
            O => \N__22636\,
            I => \N__22630\
        );

    \I__4779\ : InMux
    port map (
            O => \N__22635\,
            I => \N__22627\
        );

    \I__4778\ : Span4Mux_v
    port map (
            O => \N__22630\,
            I => \N__22622\
        );

    \I__4777\ : LocalMux
    port map (
            O => \N__22627\,
            I => \N__22622\
        );

    \I__4776\ : Odrv4
    port map (
            O => \N__22622\,
            I => \eeprom.n3403\
        );

    \I__4775\ : InMux
    port map (
            O => \N__22619\,
            I => \N__22616\
        );

    \I__4774\ : LocalMux
    port map (
            O => \N__22616\,
            I => \eeprom.n3470_adj_385\
        );

    \I__4773\ : InMux
    port map (
            O => \N__22613\,
            I => \bfn_14_19_0_\
        );

    \I__4772\ : InMux
    port map (
            O => \N__22610\,
            I => \N__22607\
        );

    \I__4771\ : LocalMux
    port map (
            O => \N__22607\,
            I => \N__22602\
        );

    \I__4770\ : InMux
    port map (
            O => \N__22606\,
            I => \N__22597\
        );

    \I__4769\ : InMux
    port map (
            O => \N__22605\,
            I => \N__22597\
        );

    \I__4768\ : Odrv4
    port map (
            O => \N__22602\,
            I => \eeprom.n3402\
        );

    \I__4767\ : LocalMux
    port map (
            O => \N__22597\,
            I => \eeprom.n3402\
        );

    \I__4766\ : CascadeMux
    port map (
            O => \N__22592\,
            I => \N__22589\
        );

    \I__4765\ : InMux
    port map (
            O => \N__22589\,
            I => \N__22586\
        );

    \I__4764\ : LocalMux
    port map (
            O => \N__22586\,
            I => \N__22583\
        );

    \I__4763\ : Span4Mux_h
    port map (
            O => \N__22583\,
            I => \N__22580\
        );

    \I__4762\ : Odrv4
    port map (
            O => \N__22580\,
            I => \eeprom.n3469_adj_384\
        );

    \I__4761\ : InMux
    port map (
            O => \N__22577\,
            I => \eeprom.n3743\
        );

    \I__4760\ : CascadeMux
    port map (
            O => \N__22574\,
            I => \N__22571\
        );

    \I__4759\ : InMux
    port map (
            O => \N__22571\,
            I => \N__22567\
        );

    \I__4758\ : CascadeMux
    port map (
            O => \N__22570\,
            I => \N__22564\
        );

    \I__4757\ : LocalMux
    port map (
            O => \N__22567\,
            I => \N__22560\
        );

    \I__4756\ : InMux
    port map (
            O => \N__22564\,
            I => \N__22555\
        );

    \I__4755\ : InMux
    port map (
            O => \N__22563\,
            I => \N__22555\
        );

    \I__4754\ : Span4Mux_v
    port map (
            O => \N__22560\,
            I => \N__22552\
        );

    \I__4753\ : LocalMux
    port map (
            O => \N__22555\,
            I => \N__22549\
        );

    \I__4752\ : Odrv4
    port map (
            O => \N__22552\,
            I => \eeprom.n3401\
        );

    \I__4751\ : Odrv4
    port map (
            O => \N__22549\,
            I => \eeprom.n3401\
        );

    \I__4750\ : InMux
    port map (
            O => \N__22544\,
            I => \N__22541\
        );

    \I__4749\ : LocalMux
    port map (
            O => \N__22541\,
            I => \N__22538\
        );

    \I__4748\ : Span4Mux_h
    port map (
            O => \N__22538\,
            I => \N__22535\
        );

    \I__4747\ : Odrv4
    port map (
            O => \N__22535\,
            I => \eeprom.n3468_adj_383\
        );

    \I__4746\ : InMux
    port map (
            O => \N__22532\,
            I => \eeprom.n3744\
        );

    \I__4745\ : CascadeMux
    port map (
            O => \N__22529\,
            I => \N__22525\
        );

    \I__4744\ : InMux
    port map (
            O => \N__22528\,
            I => \N__22521\
        );

    \I__4743\ : InMux
    port map (
            O => \N__22525\,
            I => \N__22518\
        );

    \I__4742\ : CascadeMux
    port map (
            O => \N__22524\,
            I => \N__22515\
        );

    \I__4741\ : LocalMux
    port map (
            O => \N__22521\,
            I => \N__22510\
        );

    \I__4740\ : LocalMux
    port map (
            O => \N__22518\,
            I => \N__22510\
        );

    \I__4739\ : InMux
    port map (
            O => \N__22515\,
            I => \N__22507\
        );

    \I__4738\ : Odrv12
    port map (
            O => \N__22510\,
            I => \eeprom.n3400\
        );

    \I__4737\ : LocalMux
    port map (
            O => \N__22507\,
            I => \eeprom.n3400\
        );

    \I__4736\ : CascadeMux
    port map (
            O => \N__22502\,
            I => \N__22499\
        );

    \I__4735\ : InMux
    port map (
            O => \N__22499\,
            I => \N__22496\
        );

    \I__4734\ : LocalMux
    port map (
            O => \N__22496\,
            I => \eeprom.n3467_adj_382\
        );

    \I__4733\ : InMux
    port map (
            O => \N__22493\,
            I => \eeprom.n3745\
        );

    \I__4732\ : CascadeMux
    port map (
            O => \N__22490\,
            I => \N__22486\
        );

    \I__4731\ : InMux
    port map (
            O => \N__22489\,
            I => \N__22483\
        );

    \I__4730\ : InMux
    port map (
            O => \N__22486\,
            I => \N__22480\
        );

    \I__4729\ : LocalMux
    port map (
            O => \N__22483\,
            I => \N__22476\
        );

    \I__4728\ : LocalMux
    port map (
            O => \N__22480\,
            I => \N__22473\
        );

    \I__4727\ : InMux
    port map (
            O => \N__22479\,
            I => \N__22470\
        );

    \I__4726\ : Span4Mux_v
    port map (
            O => \N__22476\,
            I => \N__22463\
        );

    \I__4725\ : Span4Mux_v
    port map (
            O => \N__22473\,
            I => \N__22463\
        );

    \I__4724\ : LocalMux
    port map (
            O => \N__22470\,
            I => \N__22463\
        );

    \I__4723\ : Span4Mux_h
    port map (
            O => \N__22463\,
            I => \N__22460\
        );

    \I__4722\ : Odrv4
    port map (
            O => \N__22460\,
            I => \eeprom.n3399\
        );

    \I__4721\ : InMux
    port map (
            O => \N__22457\,
            I => \N__22454\
        );

    \I__4720\ : LocalMux
    port map (
            O => \N__22454\,
            I => \N__22451\
        );

    \I__4719\ : Odrv4
    port map (
            O => \N__22451\,
            I => \eeprom.n3466_adj_381\
        );

    \I__4718\ : InMux
    port map (
            O => \N__22448\,
            I => \eeprom.n3746\
        );

    \I__4717\ : InMux
    port map (
            O => \N__22445\,
            I => \N__22440\
        );

    \I__4716\ : InMux
    port map (
            O => \N__22444\,
            I => \N__22437\
        );

    \I__4715\ : CascadeMux
    port map (
            O => \N__22443\,
            I => \N__22434\
        );

    \I__4714\ : LocalMux
    port map (
            O => \N__22440\,
            I => \N__22431\
        );

    \I__4713\ : LocalMux
    port map (
            O => \N__22437\,
            I => \N__22428\
        );

    \I__4712\ : InMux
    port map (
            O => \N__22434\,
            I => \N__22425\
        );

    \I__4711\ : Odrv4
    port map (
            O => \N__22431\,
            I => \eeprom.n3398\
        );

    \I__4710\ : Odrv4
    port map (
            O => \N__22428\,
            I => \eeprom.n3398\
        );

    \I__4709\ : LocalMux
    port map (
            O => \N__22425\,
            I => \eeprom.n3398\
        );

    \I__4708\ : CascadeMux
    port map (
            O => \N__22418\,
            I => \N__22415\
        );

    \I__4707\ : InMux
    port map (
            O => \N__22415\,
            I => \N__22412\
        );

    \I__4706\ : LocalMux
    port map (
            O => \N__22412\,
            I => \N__22409\
        );

    \I__4705\ : Odrv4
    port map (
            O => \N__22409\,
            I => \eeprom.n3465_adj_380\
        );

    \I__4704\ : CascadeMux
    port map (
            O => \N__22406\,
            I => \N__22402\
        );

    \I__4703\ : CascadeMux
    port map (
            O => \N__22405\,
            I => \N__22399\
        );

    \I__4702\ : InMux
    port map (
            O => \N__22402\,
            I => \N__22396\
        );

    \I__4701\ : InMux
    port map (
            O => \N__22399\,
            I => \N__22393\
        );

    \I__4700\ : LocalMux
    port map (
            O => \N__22396\,
            I => \N__22388\
        );

    \I__4699\ : LocalMux
    port map (
            O => \N__22393\,
            I => \N__22388\
        );

    \I__4698\ : Odrv4
    port map (
            O => \N__22388\,
            I => \eeprom.n3413\
        );

    \I__4697\ : InMux
    port map (
            O => \N__22385\,
            I => \N__22382\
        );

    \I__4696\ : LocalMux
    port map (
            O => \N__22382\,
            I => \eeprom.n3480_adj_398\
        );

    \I__4695\ : InMux
    port map (
            O => \N__22379\,
            I => \eeprom.n3732\
        );

    \I__4694\ : CascadeMux
    port map (
            O => \N__22376\,
            I => \N__22373\
        );

    \I__4693\ : InMux
    port map (
            O => \N__22373\,
            I => \N__22370\
        );

    \I__4692\ : LocalMux
    port map (
            O => \N__22370\,
            I => \N__22366\
        );

    \I__4691\ : InMux
    port map (
            O => \N__22369\,
            I => \N__22363\
        );

    \I__4690\ : Span4Mux_v
    port map (
            O => \N__22366\,
            I => \N__22360\
        );

    \I__4689\ : LocalMux
    port map (
            O => \N__22363\,
            I => \eeprom.n3412\
        );

    \I__4688\ : Odrv4
    port map (
            O => \N__22360\,
            I => \eeprom.n3412\
        );

    \I__4687\ : InMux
    port map (
            O => \N__22355\,
            I => \N__22352\
        );

    \I__4686\ : LocalMux
    port map (
            O => \N__22352\,
            I => \N__22349\
        );

    \I__4685\ : Span4Mux_h
    port map (
            O => \N__22349\,
            I => \N__22346\
        );

    \I__4684\ : Odrv4
    port map (
            O => \N__22346\,
            I => \eeprom.n3479_adj_394\
        );

    \I__4683\ : InMux
    port map (
            O => \N__22343\,
            I => \eeprom.n3733\
        );

    \I__4682\ : CascadeMux
    port map (
            O => \N__22340\,
            I => \N__22335\
        );

    \I__4681\ : InMux
    port map (
            O => \N__22339\,
            I => \N__22332\
        );

    \I__4680\ : InMux
    port map (
            O => \N__22338\,
            I => \N__22329\
        );

    \I__4679\ : InMux
    port map (
            O => \N__22335\,
            I => \N__22326\
        );

    \I__4678\ : LocalMux
    port map (
            O => \N__22332\,
            I => \N__22319\
        );

    \I__4677\ : LocalMux
    port map (
            O => \N__22329\,
            I => \N__22319\
        );

    \I__4676\ : LocalMux
    port map (
            O => \N__22326\,
            I => \N__22319\
        );

    \I__4675\ : Odrv12
    port map (
            O => \N__22319\,
            I => \eeprom.n3411\
        );

    \I__4674\ : CascadeMux
    port map (
            O => \N__22316\,
            I => \N__22313\
        );

    \I__4673\ : InMux
    port map (
            O => \N__22313\,
            I => \N__22310\
        );

    \I__4672\ : LocalMux
    port map (
            O => \N__22310\,
            I => \eeprom.n3478_adj_393\
        );

    \I__4671\ : InMux
    port map (
            O => \N__22307\,
            I => \bfn_14_18_0_\
        );

    \I__4670\ : CascadeMux
    port map (
            O => \N__22304\,
            I => \N__22301\
        );

    \I__4669\ : InMux
    port map (
            O => \N__22301\,
            I => \N__22298\
        );

    \I__4668\ : LocalMux
    port map (
            O => \N__22298\,
            I => \N__22294\
        );

    \I__4667\ : InMux
    port map (
            O => \N__22297\,
            I => \N__22291\
        );

    \I__4666\ : Odrv4
    port map (
            O => \N__22294\,
            I => \eeprom.n3410\
        );

    \I__4665\ : LocalMux
    port map (
            O => \N__22291\,
            I => \eeprom.n3410\
        );

    \I__4664\ : InMux
    port map (
            O => \N__22286\,
            I => \N__22283\
        );

    \I__4663\ : LocalMux
    port map (
            O => \N__22283\,
            I => \N__22280\
        );

    \I__4662\ : Odrv4
    port map (
            O => \N__22280\,
            I => \eeprom.n3477_adj_392\
        );

    \I__4661\ : InMux
    port map (
            O => \N__22277\,
            I => \eeprom.n3735\
        );

    \I__4660\ : CascadeMux
    port map (
            O => \N__22274\,
            I => \N__22271\
        );

    \I__4659\ : InMux
    port map (
            O => \N__22271\,
            I => \N__22266\
        );

    \I__4658\ : InMux
    port map (
            O => \N__22270\,
            I => \N__22261\
        );

    \I__4657\ : InMux
    port map (
            O => \N__22269\,
            I => \N__22261\
        );

    \I__4656\ : LocalMux
    port map (
            O => \N__22266\,
            I => \N__22258\
        );

    \I__4655\ : LocalMux
    port map (
            O => \N__22261\,
            I => \eeprom.n3409\
        );

    \I__4654\ : Odrv4
    port map (
            O => \N__22258\,
            I => \eeprom.n3409\
        );

    \I__4653\ : InMux
    port map (
            O => \N__22253\,
            I => \N__22250\
        );

    \I__4652\ : LocalMux
    port map (
            O => \N__22250\,
            I => \N__22247\
        );

    \I__4651\ : Odrv4
    port map (
            O => \N__22247\,
            I => \eeprom.n3476_adj_391\
        );

    \I__4650\ : InMux
    port map (
            O => \N__22244\,
            I => \eeprom.n3736\
        );

    \I__4649\ : CascadeMux
    port map (
            O => \N__22241\,
            I => \N__22237\
        );

    \I__4648\ : InMux
    port map (
            O => \N__22240\,
            I => \N__22234\
        );

    \I__4647\ : InMux
    port map (
            O => \N__22237\,
            I => \N__22231\
        );

    \I__4646\ : LocalMux
    port map (
            O => \N__22234\,
            I => \N__22227\
        );

    \I__4645\ : LocalMux
    port map (
            O => \N__22231\,
            I => \N__22224\
        );

    \I__4644\ : InMux
    port map (
            O => \N__22230\,
            I => \N__22221\
        );

    \I__4643\ : Odrv4
    port map (
            O => \N__22227\,
            I => \eeprom.n3408\
        );

    \I__4642\ : Odrv12
    port map (
            O => \N__22224\,
            I => \eeprom.n3408\
        );

    \I__4641\ : LocalMux
    port map (
            O => \N__22221\,
            I => \eeprom.n3408\
        );

    \I__4640\ : CascadeMux
    port map (
            O => \N__22214\,
            I => \N__22211\
        );

    \I__4639\ : InMux
    port map (
            O => \N__22211\,
            I => \N__22208\
        );

    \I__4638\ : LocalMux
    port map (
            O => \N__22208\,
            I => \N__22205\
        );

    \I__4637\ : Odrv4
    port map (
            O => \N__22205\,
            I => \eeprom.n3475_adj_390\
        );

    \I__4636\ : InMux
    port map (
            O => \N__22202\,
            I => \eeprom.n3737\
        );

    \I__4635\ : CascadeMux
    port map (
            O => \N__22199\,
            I => \N__22195\
        );

    \I__4634\ : CascadeMux
    port map (
            O => \N__22198\,
            I => \N__22192\
        );

    \I__4633\ : InMux
    port map (
            O => \N__22195\,
            I => \N__22189\
        );

    \I__4632\ : InMux
    port map (
            O => \N__22192\,
            I => \N__22186\
        );

    \I__4631\ : LocalMux
    port map (
            O => \N__22189\,
            I => \N__22183\
        );

    \I__4630\ : LocalMux
    port map (
            O => \N__22186\,
            I => \eeprom.n3407\
        );

    \I__4629\ : Odrv4
    port map (
            O => \N__22183\,
            I => \eeprom.n3407\
        );

    \I__4628\ : InMux
    port map (
            O => \N__22178\,
            I => \N__22175\
        );

    \I__4627\ : LocalMux
    port map (
            O => \N__22175\,
            I => \N__22172\
        );

    \I__4626\ : Odrv4
    port map (
            O => \N__22172\,
            I => \eeprom.n3474_adj_389\
        );

    \I__4625\ : InMux
    port map (
            O => \N__22169\,
            I => \eeprom.n3738\
        );

    \I__4624\ : CascadeMux
    port map (
            O => \N__22166\,
            I => \N__22162\
        );

    \I__4623\ : InMux
    port map (
            O => \N__22165\,
            I => \N__22159\
        );

    \I__4622\ : InMux
    port map (
            O => \N__22162\,
            I => \N__22156\
        );

    \I__4621\ : LocalMux
    port map (
            O => \N__22159\,
            I => \N__22150\
        );

    \I__4620\ : LocalMux
    port map (
            O => \N__22156\,
            I => \N__22150\
        );

    \I__4619\ : InMux
    port map (
            O => \N__22155\,
            I => \N__22147\
        );

    \I__4618\ : Odrv12
    port map (
            O => \N__22150\,
            I => \eeprom.n3406\
        );

    \I__4617\ : LocalMux
    port map (
            O => \N__22147\,
            I => \eeprom.n3406\
        );

    \I__4616\ : CascadeMux
    port map (
            O => \N__22142\,
            I => \N__22139\
        );

    \I__4615\ : InMux
    port map (
            O => \N__22139\,
            I => \N__22136\
        );

    \I__4614\ : LocalMux
    port map (
            O => \N__22136\,
            I => \N__22133\
        );

    \I__4613\ : Odrv12
    port map (
            O => \N__22133\,
            I => \eeprom.n3473_adj_388\
        );

    \I__4612\ : InMux
    port map (
            O => \N__22130\,
            I => \eeprom.n3739\
        );

    \I__4611\ : InMux
    port map (
            O => \N__22127\,
            I => \N__22122\
        );

    \I__4610\ : InMux
    port map (
            O => \N__22126\,
            I => \N__22119\
        );

    \I__4609\ : CascadeMux
    port map (
            O => \N__22125\,
            I => \N__22116\
        );

    \I__4608\ : LocalMux
    port map (
            O => \N__22122\,
            I => \N__22113\
        );

    \I__4607\ : LocalMux
    port map (
            O => \N__22119\,
            I => \N__22110\
        );

    \I__4606\ : InMux
    port map (
            O => \N__22116\,
            I => \N__22107\
        );

    \I__4605\ : Odrv12
    port map (
            O => \N__22113\,
            I => \eeprom.n2907\
        );

    \I__4604\ : Odrv4
    port map (
            O => \N__22110\,
            I => \eeprom.n2907\
        );

    \I__4603\ : LocalMux
    port map (
            O => \N__22107\,
            I => \eeprom.n2907\
        );

    \I__4602\ : CascadeMux
    port map (
            O => \N__22100\,
            I => \N__22097\
        );

    \I__4601\ : InMux
    port map (
            O => \N__22097\,
            I => \N__22094\
        );

    \I__4600\ : LocalMux
    port map (
            O => \N__22094\,
            I => \N__22091\
        );

    \I__4599\ : Span4Mux_v
    port map (
            O => \N__22091\,
            I => \N__22088\
        );

    \I__4598\ : Odrv4
    port map (
            O => \N__22088\,
            I => \eeprom.n2974\
        );

    \I__4597\ : InMux
    port map (
            O => \N__22085\,
            I => \N__22082\
        );

    \I__4596\ : LocalMux
    port map (
            O => \N__22082\,
            I => \N__22077\
        );

    \I__4595\ : CascadeMux
    port map (
            O => \N__22081\,
            I => \N__22074\
        );

    \I__4594\ : InMux
    port map (
            O => \N__22080\,
            I => \N__22071\
        );

    \I__4593\ : Span4Mux_v
    port map (
            O => \N__22077\,
            I => \N__22068\
        );

    \I__4592\ : InMux
    port map (
            O => \N__22074\,
            I => \N__22065\
        );

    \I__4591\ : LocalMux
    port map (
            O => \N__22071\,
            I => \N__22062\
        );

    \I__4590\ : Odrv4
    port map (
            O => \N__22068\,
            I => \eeprom.n2914\
        );

    \I__4589\ : LocalMux
    port map (
            O => \N__22065\,
            I => \eeprom.n2914\
        );

    \I__4588\ : Odrv12
    port map (
            O => \N__22062\,
            I => \eeprom.n2914\
        );

    \I__4587\ : InMux
    port map (
            O => \N__22055\,
            I => \N__22052\
        );

    \I__4586\ : LocalMux
    port map (
            O => \N__22052\,
            I => \N__22049\
        );

    \I__4585\ : Span4Mux_h
    port map (
            O => \N__22049\,
            I => \N__22046\
        );

    \I__4584\ : Odrv4
    port map (
            O => \N__22046\,
            I => \eeprom.n2981\
        );

    \I__4583\ : CascadeMux
    port map (
            O => \N__22043\,
            I => \N__22039\
        );

    \I__4582\ : InMux
    port map (
            O => \N__22042\,
            I => \N__22035\
        );

    \I__4581\ : InMux
    port map (
            O => \N__22039\,
            I => \N__22030\
        );

    \I__4580\ : InMux
    port map (
            O => \N__22038\,
            I => \N__22030\
        );

    \I__4579\ : LocalMux
    port map (
            O => \N__22035\,
            I => \eeprom.n3101\
        );

    \I__4578\ : LocalMux
    port map (
            O => \N__22030\,
            I => \eeprom.n3101\
        );

    \I__4577\ : InMux
    port map (
            O => \N__22025\,
            I => \bfn_14_17_0_\
        );

    \I__4576\ : InMux
    port map (
            O => \N__22022\,
            I => \eeprom.n3727\
        );

    \I__4575\ : InMux
    port map (
            O => \N__22019\,
            I => \eeprom.n3728\
        );

    \I__4574\ : InMux
    port map (
            O => \N__22016\,
            I => \eeprom.n3729\
        );

    \I__4573\ : CascadeMux
    port map (
            O => \N__22013\,
            I => \N__22009\
        );

    \I__4572\ : CascadeMux
    port map (
            O => \N__22012\,
            I => \N__22006\
        );

    \I__4571\ : InMux
    port map (
            O => \N__22009\,
            I => \N__22003\
        );

    \I__4570\ : InMux
    port map (
            O => \N__22006\,
            I => \N__21999\
        );

    \I__4569\ : LocalMux
    port map (
            O => \N__22003\,
            I => \N__21996\
        );

    \I__4568\ : InMux
    port map (
            O => \N__22002\,
            I => \N__21993\
        );

    \I__4567\ : LocalMux
    port map (
            O => \N__21999\,
            I => \eeprom.n3415\
        );

    \I__4566\ : Odrv4
    port map (
            O => \N__21996\,
            I => \eeprom.n3415\
        );

    \I__4565\ : LocalMux
    port map (
            O => \N__21993\,
            I => \eeprom.n3415\
        );

    \I__4564\ : InMux
    port map (
            O => \N__21986\,
            I => \N__21983\
        );

    \I__4563\ : LocalMux
    port map (
            O => \N__21983\,
            I => \eeprom.n3482_adj_401\
        );

    \I__4562\ : InMux
    port map (
            O => \N__21980\,
            I => \eeprom.n3730\
        );

    \I__4561\ : InMux
    port map (
            O => \N__21977\,
            I => \N__21973\
        );

    \I__4560\ : InMux
    port map (
            O => \N__21976\,
            I => \N__21970\
        );

    \I__4559\ : LocalMux
    port map (
            O => \N__21973\,
            I => \N__21967\
        );

    \I__4558\ : LocalMux
    port map (
            O => \N__21970\,
            I => \eeprom.n3414\
        );

    \I__4557\ : Odrv4
    port map (
            O => \N__21967\,
            I => \eeprom.n3414\
        );

    \I__4556\ : InMux
    port map (
            O => \N__21962\,
            I => \N__21959\
        );

    \I__4555\ : LocalMux
    port map (
            O => \N__21959\,
            I => \eeprom.n3481_adj_399\
        );

    \I__4554\ : InMux
    port map (
            O => \N__21956\,
            I => \eeprom.n3731\
        );

    \I__4553\ : InMux
    port map (
            O => \N__21953\,
            I => \N__21948\
        );

    \I__4552\ : InMux
    port map (
            O => \N__21952\,
            I => \N__21945\
        );

    \I__4551\ : InMux
    port map (
            O => \N__21951\,
            I => \N__21942\
        );

    \I__4550\ : LocalMux
    port map (
            O => \N__21948\,
            I => \N__21937\
        );

    \I__4549\ : LocalMux
    port map (
            O => \N__21945\,
            I => \N__21937\
        );

    \I__4548\ : LocalMux
    port map (
            O => \N__21942\,
            I => \eeprom.n3104\
        );

    \I__4547\ : Odrv4
    port map (
            O => \N__21937\,
            I => \eeprom.n3104\
        );

    \I__4546\ : InMux
    port map (
            O => \N__21932\,
            I => \N__21929\
        );

    \I__4545\ : LocalMux
    port map (
            O => \N__21929\,
            I => \eeprom.n3170\
        );

    \I__4544\ : InMux
    port map (
            O => \N__21926\,
            I => \N__21922\
        );

    \I__4543\ : InMux
    port map (
            O => \N__21925\,
            I => \N__21919\
        );

    \I__4542\ : LocalMux
    port map (
            O => \N__21922\,
            I => \N__21916\
        );

    \I__4541\ : LocalMux
    port map (
            O => \N__21919\,
            I => \N__21913\
        );

    \I__4540\ : Span4Mux_h
    port map (
            O => \N__21916\,
            I => \N__21909\
        );

    \I__4539\ : Span4Mux_h
    port map (
            O => \N__21913\,
            I => \N__21906\
        );

    \I__4538\ : InMux
    port map (
            O => \N__21912\,
            I => \N__21903\
        );

    \I__4537\ : Odrv4
    port map (
            O => \N__21909\,
            I => \eeprom.n3202\
        );

    \I__4536\ : Odrv4
    port map (
            O => \N__21906\,
            I => \eeprom.n3202\
        );

    \I__4535\ : LocalMux
    port map (
            O => \N__21903\,
            I => \eeprom.n3202\
        );

    \I__4534\ : InMux
    port map (
            O => \N__21896\,
            I => \N__21893\
        );

    \I__4533\ : LocalMux
    port map (
            O => \N__21893\,
            I => \eeprom.n3168\
        );

    \I__4532\ : InMux
    port map (
            O => \N__21890\,
            I => \N__21886\
        );

    \I__4531\ : InMux
    port map (
            O => \N__21889\,
            I => \N__21883\
        );

    \I__4530\ : LocalMux
    port map (
            O => \N__21886\,
            I => \N__21880\
        );

    \I__4529\ : LocalMux
    port map (
            O => \N__21883\,
            I => \N__21877\
        );

    \I__4528\ : Span4Mux_h
    port map (
            O => \N__21880\,
            I => \N__21873\
        );

    \I__4527\ : Span4Mux_h
    port map (
            O => \N__21877\,
            I => \N__21870\
        );

    \I__4526\ : InMux
    port map (
            O => \N__21876\,
            I => \N__21867\
        );

    \I__4525\ : Odrv4
    port map (
            O => \N__21873\,
            I => \eeprom.n3200\
        );

    \I__4524\ : Odrv4
    port map (
            O => \N__21870\,
            I => \eeprom.n3200\
        );

    \I__4523\ : LocalMux
    port map (
            O => \N__21867\,
            I => \eeprom.n3200\
        );

    \I__4522\ : InMux
    port map (
            O => \N__21860\,
            I => \N__21857\
        );

    \I__4521\ : LocalMux
    port map (
            O => \N__21857\,
            I => \N__21854\
        );

    \I__4520\ : Span4Mux_h
    port map (
            O => \N__21854\,
            I => \N__21851\
        );

    \I__4519\ : Odrv4
    port map (
            O => \N__21851\,
            I => \eeprom.n2983\
        );

    \I__4518\ : CascadeMux
    port map (
            O => \N__21848\,
            I => \N__21845\
        );

    \I__4517\ : InMux
    port map (
            O => \N__21845\,
            I => \N__21841\
        );

    \I__4516\ : CascadeMux
    port map (
            O => \N__21844\,
            I => \N__21838\
        );

    \I__4515\ : LocalMux
    port map (
            O => \N__21841\,
            I => \N__21835\
        );

    \I__4514\ : InMux
    port map (
            O => \N__21838\,
            I => \N__21832\
        );

    \I__4513\ : Span4Mux_h
    port map (
            O => \N__21835\,
            I => \N__21826\
        );

    \I__4512\ : LocalMux
    port map (
            O => \N__21832\,
            I => \N__21826\
        );

    \I__4511\ : InMux
    port map (
            O => \N__21831\,
            I => \N__21823\
        );

    \I__4510\ : Odrv4
    port map (
            O => \N__21826\,
            I => \eeprom.n2916\
        );

    \I__4509\ : LocalMux
    port map (
            O => \N__21823\,
            I => \eeprom.n2916\
        );

    \I__4508\ : InMux
    port map (
            O => \N__21818\,
            I => \N__21814\
        );

    \I__4507\ : InMux
    port map (
            O => \N__21817\,
            I => \N__21811\
        );

    \I__4506\ : LocalMux
    port map (
            O => \N__21814\,
            I => \N__21808\
        );

    \I__4505\ : LocalMux
    port map (
            O => \N__21811\,
            I => \eeprom.n3106\
        );

    \I__4504\ : Odrv4
    port map (
            O => \N__21808\,
            I => \eeprom.n3106\
        );

    \I__4503\ : InMux
    port map (
            O => \N__21803\,
            I => \N__21800\
        );

    \I__4502\ : LocalMux
    port map (
            O => \N__21800\,
            I => \eeprom.n3173\
        );

    \I__4501\ : CascadeMux
    port map (
            O => \N__21797\,
            I => \eeprom.n3106_cascade_\
        );

    \I__4500\ : CascadeMux
    port map (
            O => \N__21794\,
            I => \N__21785\
        );

    \I__4499\ : InMux
    port map (
            O => \N__21793\,
            I => \N__21781\
        );

    \I__4498\ : CascadeMux
    port map (
            O => \N__21792\,
            I => \N__21778\
        );

    \I__4497\ : CascadeMux
    port map (
            O => \N__21791\,
            I => \N__21773\
        );

    \I__4496\ : InMux
    port map (
            O => \N__21790\,
            I => \N__21766\
        );

    \I__4495\ : InMux
    port map (
            O => \N__21789\,
            I => \N__21766\
        );

    \I__4494\ : InMux
    port map (
            O => \N__21788\,
            I => \N__21758\
        );

    \I__4493\ : InMux
    port map (
            O => \N__21785\,
            I => \N__21753\
        );

    \I__4492\ : InMux
    port map (
            O => \N__21784\,
            I => \N__21753\
        );

    \I__4491\ : LocalMux
    port map (
            O => \N__21781\,
            I => \N__21750\
        );

    \I__4490\ : InMux
    port map (
            O => \N__21778\,
            I => \N__21747\
        );

    \I__4489\ : CascadeMux
    port map (
            O => \N__21777\,
            I => \N__21743\
        );

    \I__4488\ : InMux
    port map (
            O => \N__21776\,
            I => \N__21738\
        );

    \I__4487\ : InMux
    port map (
            O => \N__21773\,
            I => \N__21731\
        );

    \I__4486\ : InMux
    port map (
            O => \N__21772\,
            I => \N__21731\
        );

    \I__4485\ : InMux
    port map (
            O => \N__21771\,
            I => \N__21731\
        );

    \I__4484\ : LocalMux
    port map (
            O => \N__21766\,
            I => \N__21728\
        );

    \I__4483\ : InMux
    port map (
            O => \N__21765\,
            I => \N__21721\
        );

    \I__4482\ : InMux
    port map (
            O => \N__21764\,
            I => \N__21721\
        );

    \I__4481\ : InMux
    port map (
            O => \N__21763\,
            I => \N__21721\
        );

    \I__4480\ : InMux
    port map (
            O => \N__21762\,
            I => \N__21716\
        );

    \I__4479\ : InMux
    port map (
            O => \N__21761\,
            I => \N__21716\
        );

    \I__4478\ : LocalMux
    port map (
            O => \N__21758\,
            I => \N__21711\
        );

    \I__4477\ : LocalMux
    port map (
            O => \N__21753\,
            I => \N__21711\
        );

    \I__4476\ : Span4Mux_h
    port map (
            O => \N__21750\,
            I => \N__21706\
        );

    \I__4475\ : LocalMux
    port map (
            O => \N__21747\,
            I => \N__21706\
        );

    \I__4474\ : InMux
    port map (
            O => \N__21746\,
            I => \N__21697\
        );

    \I__4473\ : InMux
    port map (
            O => \N__21743\,
            I => \N__21697\
        );

    \I__4472\ : InMux
    port map (
            O => \N__21742\,
            I => \N__21697\
        );

    \I__4471\ : InMux
    port map (
            O => \N__21741\,
            I => \N__21697\
        );

    \I__4470\ : LocalMux
    port map (
            O => \N__21738\,
            I => \eeprom.n3133\
        );

    \I__4469\ : LocalMux
    port map (
            O => \N__21731\,
            I => \eeprom.n3133\
        );

    \I__4468\ : Odrv4
    port map (
            O => \N__21728\,
            I => \eeprom.n3133\
        );

    \I__4467\ : LocalMux
    port map (
            O => \N__21721\,
            I => \eeprom.n3133\
        );

    \I__4466\ : LocalMux
    port map (
            O => \N__21716\,
            I => \eeprom.n3133\
        );

    \I__4465\ : Odrv4
    port map (
            O => \N__21711\,
            I => \eeprom.n3133\
        );

    \I__4464\ : Odrv4
    port map (
            O => \N__21706\,
            I => \eeprom.n3133\
        );

    \I__4463\ : LocalMux
    port map (
            O => \N__21697\,
            I => \eeprom.n3133\
        );

    \I__4462\ : InMux
    port map (
            O => \N__21680\,
            I => \N__21677\
        );

    \I__4461\ : LocalMux
    port map (
            O => \N__21677\,
            I => \N__21673\
        );

    \I__4460\ : InMux
    port map (
            O => \N__21676\,
            I => \N__21670\
        );

    \I__4459\ : Span4Mux_v
    port map (
            O => \N__21673\,
            I => \N__21667\
        );

    \I__4458\ : LocalMux
    port map (
            O => \N__21670\,
            I => \N__21664\
        );

    \I__4457\ : Span4Mux_h
    port map (
            O => \N__21667\,
            I => \N__21661\
        );

    \I__4456\ : Span4Mux_h
    port map (
            O => \N__21664\,
            I => \N__21658\
        );

    \I__4455\ : Odrv4
    port map (
            O => \N__21661\,
            I => \eeprom.n3205\
        );

    \I__4454\ : Odrv4
    port map (
            O => \N__21658\,
            I => \eeprom.n3205\
        );

    \I__4453\ : CascadeMux
    port map (
            O => \N__21653\,
            I => \eeprom.n3205_cascade_\
        );

    \I__4452\ : InMux
    port map (
            O => \N__21650\,
            I => \N__21647\
        );

    \I__4451\ : LocalMux
    port map (
            O => \N__21647\,
            I => \N__21644\
        );

    \I__4450\ : Span4Mux_v
    port map (
            O => \N__21644\,
            I => \N__21640\
        );

    \I__4449\ : InMux
    port map (
            O => \N__21643\,
            I => \N__21637\
        );

    \I__4448\ : Odrv4
    port map (
            O => \N__21640\,
            I => \eeprom.n3199\
        );

    \I__4447\ : LocalMux
    port map (
            O => \N__21637\,
            I => \eeprom.n3199\
        );

    \I__4446\ : InMux
    port map (
            O => \N__21632\,
            I => \N__21629\
        );

    \I__4445\ : LocalMux
    port map (
            O => \N__21629\,
            I => \N__21626\
        );

    \I__4444\ : Span4Mux_h
    port map (
            O => \N__21626\,
            I => \N__21623\
        );

    \I__4443\ : Span4Mux_v
    port map (
            O => \N__21623\,
            I => \N__21620\
        );

    \I__4442\ : Odrv4
    port map (
            O => \N__21620\,
            I => \eeprom.n16_adj_479\
        );

    \I__4441\ : CascadeMux
    port map (
            O => \N__21617\,
            I => \N__21612\
        );

    \I__4440\ : CascadeMux
    port map (
            O => \N__21616\,
            I => \N__21609\
        );

    \I__4439\ : CascadeMux
    port map (
            O => \N__21615\,
            I => \N__21606\
        );

    \I__4438\ : InMux
    port map (
            O => \N__21612\,
            I => \N__21603\
        );

    \I__4437\ : InMux
    port map (
            O => \N__21609\,
            I => \N__21598\
        );

    \I__4436\ : InMux
    port map (
            O => \N__21606\,
            I => \N__21598\
        );

    \I__4435\ : LocalMux
    port map (
            O => \N__21603\,
            I => \eeprom.n3115\
        );

    \I__4434\ : LocalMux
    port map (
            O => \N__21598\,
            I => \eeprom.n3115\
        );

    \I__4433\ : InMux
    port map (
            O => \N__21593\,
            I => \N__21590\
        );

    \I__4432\ : LocalMux
    port map (
            O => \N__21590\,
            I => \N__21587\
        );

    \I__4431\ : Odrv4
    port map (
            O => \N__21587\,
            I => \eeprom.n3169\
        );

    \I__4430\ : InMux
    port map (
            O => \N__21584\,
            I => \N__21581\
        );

    \I__4429\ : LocalMux
    port map (
            O => \N__21581\,
            I => \N__21577\
        );

    \I__4428\ : InMux
    port map (
            O => \N__21580\,
            I => \N__21574\
        );

    \I__4427\ : Span4Mux_h
    port map (
            O => \N__21577\,
            I => \N__21571\
        );

    \I__4426\ : LocalMux
    port map (
            O => \N__21574\,
            I => \N__21568\
        );

    \I__4425\ : Odrv4
    port map (
            O => \N__21571\,
            I => \eeprom.n3201\
        );

    \I__4424\ : Odrv12
    port map (
            O => \N__21568\,
            I => \eeprom.n3201\
        );

    \I__4423\ : InMux
    port map (
            O => \N__21563\,
            I => \N__21560\
        );

    \I__4422\ : LocalMux
    port map (
            O => \N__21560\,
            I => \N__21556\
        );

    \I__4421\ : InMux
    port map (
            O => \N__21559\,
            I => \N__21553\
        );

    \I__4420\ : Span4Mux_h
    port map (
            O => \N__21556\,
            I => \N__21549\
        );

    \I__4419\ : LocalMux
    port map (
            O => \N__21553\,
            I => \N__21546\
        );

    \I__4418\ : InMux
    port map (
            O => \N__21552\,
            I => \N__21543\
        );

    \I__4417\ : Odrv4
    port map (
            O => \N__21549\,
            I => \eeprom.n3207\
        );

    \I__4416\ : Odrv12
    port map (
            O => \N__21546\,
            I => \eeprom.n3207\
        );

    \I__4415\ : LocalMux
    port map (
            O => \N__21543\,
            I => \eeprom.n3207\
        );

    \I__4414\ : CascadeMux
    port map (
            O => \N__21536\,
            I => \eeprom.n3201_cascade_\
        );

    \I__4413\ : InMux
    port map (
            O => \N__21533\,
            I => \N__21530\
        );

    \I__4412\ : LocalMux
    port map (
            O => \N__21530\,
            I => \N__21527\
        );

    \I__4411\ : Span4Mux_h
    port map (
            O => \N__21527\,
            I => \N__21524\
        );

    \I__4410\ : Odrv4
    port map (
            O => \N__21524\,
            I => \eeprom.n24_adj_481\
        );

    \I__4409\ : InMux
    port map (
            O => \N__21521\,
            I => \N__21518\
        );

    \I__4408\ : LocalMux
    port map (
            O => \N__21518\,
            I => \N__21514\
        );

    \I__4407\ : CascadeMux
    port map (
            O => \N__21517\,
            I => \N__21511\
        );

    \I__4406\ : Span4Mux_v
    port map (
            O => \N__21514\,
            I => \N__21507\
        );

    \I__4405\ : InMux
    port map (
            O => \N__21511\,
            I => \N__21504\
        );

    \I__4404\ : InMux
    port map (
            O => \N__21510\,
            I => \N__21501\
        );

    \I__4403\ : Odrv4
    port map (
            O => \N__21507\,
            I => \eeprom.n3114\
        );

    \I__4402\ : LocalMux
    port map (
            O => \N__21504\,
            I => \eeprom.n3114\
        );

    \I__4401\ : LocalMux
    port map (
            O => \N__21501\,
            I => \eeprom.n3114\
        );

    \I__4400\ : InMux
    port map (
            O => \N__21494\,
            I => \N__21490\
        );

    \I__4399\ : InMux
    port map (
            O => \N__21493\,
            I => \N__21487\
        );

    \I__4398\ : LocalMux
    port map (
            O => \N__21490\,
            I => \N__21482\
        );

    \I__4397\ : LocalMux
    port map (
            O => \N__21487\,
            I => \N__21482\
        );

    \I__4396\ : Span4Mux_h
    port map (
            O => \N__21482\,
            I => \N__21478\
        );

    \I__4395\ : InMux
    port map (
            O => \N__21481\,
            I => \N__21475\
        );

    \I__4394\ : Odrv4
    port map (
            O => \N__21478\,
            I => \eeprom.n2905\
        );

    \I__4393\ : LocalMux
    port map (
            O => \N__21475\,
            I => \eeprom.n2905\
        );

    \I__4392\ : CascadeMux
    port map (
            O => \N__21470\,
            I => \N__21467\
        );

    \I__4391\ : InMux
    port map (
            O => \N__21467\,
            I => \N__21464\
        );

    \I__4390\ : LocalMux
    port map (
            O => \N__21464\,
            I => \N__21461\
        );

    \I__4389\ : Odrv4
    port map (
            O => \N__21461\,
            I => \eeprom.n2972\
        );

    \I__4388\ : InMux
    port map (
            O => \N__21458\,
            I => \N__21455\
        );

    \I__4387\ : LocalMux
    port map (
            O => \N__21455\,
            I => \N__21450\
        );

    \I__4386\ : CascadeMux
    port map (
            O => \N__21454\,
            I => \N__21447\
        );

    \I__4385\ : CascadeMux
    port map (
            O => \N__21453\,
            I => \N__21444\
        );

    \I__4384\ : Span4Mux_v
    port map (
            O => \N__21450\,
            I => \N__21441\
        );

    \I__4383\ : InMux
    port map (
            O => \N__21447\,
            I => \N__21438\
        );

    \I__4382\ : InMux
    port map (
            O => \N__21444\,
            I => \N__21435\
        );

    \I__4381\ : Odrv4
    port map (
            O => \N__21441\,
            I => \eeprom.n3118\
        );

    \I__4380\ : LocalMux
    port map (
            O => \N__21438\,
            I => \eeprom.n3118\
        );

    \I__4379\ : LocalMux
    port map (
            O => \N__21435\,
            I => \eeprom.n3118\
        );

    \I__4378\ : InMux
    port map (
            O => \N__21428\,
            I => \N__21424\
        );

    \I__4377\ : InMux
    port map (
            O => \N__21427\,
            I => \N__21421\
        );

    \I__4376\ : LocalMux
    port map (
            O => \N__21424\,
            I => \eeprom.n3102\
        );

    \I__4375\ : LocalMux
    port map (
            O => \N__21421\,
            I => \eeprom.n3102\
        );

    \I__4374\ : CascadeMux
    port map (
            O => \N__21416\,
            I => \eeprom.n3102_cascade_\
        );

    \I__4373\ : InMux
    port map (
            O => \N__21413\,
            I => \N__21410\
        );

    \I__4372\ : LocalMux
    port map (
            O => \N__21410\,
            I => \N__21407\
        );

    \I__4371\ : Odrv4
    port map (
            O => \N__21407\,
            I => \eeprom.n22_adj_465\
        );

    \I__4370\ : InMux
    port map (
            O => \N__21404\,
            I => \N__21401\
        );

    \I__4369\ : LocalMux
    port map (
            O => \N__21401\,
            I => \eeprom.n3600_adj_449\
        );

    \I__4368\ : InMux
    port map (
            O => \N__21398\,
            I => \N__21395\
        );

    \I__4367\ : LocalMux
    port map (
            O => \N__21395\,
            I => \eeprom.n4581\
        );

    \I__4366\ : CascadeMux
    port map (
            O => \N__21392\,
            I => \N__21387\
        );

    \I__4365\ : InMux
    port map (
            O => \N__21391\,
            I => \N__21384\
        );

    \I__4364\ : InMux
    port map (
            O => \N__21390\,
            I => \N__21381\
        );

    \I__4363\ : InMux
    port map (
            O => \N__21387\,
            I => \N__21378\
        );

    \I__4362\ : LocalMux
    port map (
            O => \N__21384\,
            I => \eeprom.n3117\
        );

    \I__4361\ : LocalMux
    port map (
            O => \N__21381\,
            I => \eeprom.n3117\
        );

    \I__4360\ : LocalMux
    port map (
            O => \N__21378\,
            I => \eeprom.n3117\
        );

    \I__4359\ : InMux
    port map (
            O => \N__21371\,
            I => \N__21367\
        );

    \I__4358\ : InMux
    port map (
            O => \N__21370\,
            I => \N__21364\
        );

    \I__4357\ : LocalMux
    port map (
            O => \N__21367\,
            I => \N__21361\
        );

    \I__4356\ : LocalMux
    port map (
            O => \N__21364\,
            I => \eeprom.n3108\
        );

    \I__4355\ : Odrv4
    port map (
            O => \N__21361\,
            I => \eeprom.n3108\
        );

    \I__4354\ : InMux
    port map (
            O => \N__21356\,
            I => \N__21353\
        );

    \I__4353\ : LocalMux
    port map (
            O => \N__21353\,
            I => \N__21350\
        );

    \I__4352\ : Odrv4
    port map (
            O => \N__21350\,
            I => \eeprom.n3175\
        );

    \I__4351\ : CascadeMux
    port map (
            O => \N__21347\,
            I => \eeprom.n3108_cascade_\
        );

    \I__4350\ : CascadeMux
    port map (
            O => \N__21344\,
            I => \N__21341\
        );

    \I__4349\ : InMux
    port map (
            O => \N__21341\,
            I => \N__21337\
        );

    \I__4348\ : InMux
    port map (
            O => \N__21340\,
            I => \N__21334\
        );

    \I__4347\ : LocalMux
    port map (
            O => \N__21337\,
            I => \N__21331\
        );

    \I__4346\ : LocalMux
    port map (
            O => \N__21334\,
            I => \eeprom.n3105\
        );

    \I__4345\ : Odrv4
    port map (
            O => \N__21331\,
            I => \eeprom.n3105\
        );

    \I__4344\ : InMux
    port map (
            O => \N__21326\,
            I => \N__21323\
        );

    \I__4343\ : LocalMux
    port map (
            O => \N__21323\,
            I => \N__21320\
        );

    \I__4342\ : Span4Mux_h
    port map (
            O => \N__21320\,
            I => \N__21317\
        );

    \I__4341\ : Odrv4
    port map (
            O => \N__21317\,
            I => \eeprom.n3172\
        );

    \I__4340\ : CascadeMux
    port map (
            O => \N__21314\,
            I => \eeprom.n3105_cascade_\
        );

    \I__4339\ : InMux
    port map (
            O => \N__21311\,
            I => \N__21307\
        );

    \I__4338\ : InMux
    port map (
            O => \N__21310\,
            I => \N__21303\
        );

    \I__4337\ : LocalMux
    port map (
            O => \N__21307\,
            I => \N__21300\
        );

    \I__4336\ : InMux
    port map (
            O => \N__21306\,
            I => \N__21297\
        );

    \I__4335\ : LocalMux
    port map (
            O => \N__21303\,
            I => \N__21294\
        );

    \I__4334\ : Span4Mux_h
    port map (
            O => \N__21300\,
            I => \N__21291\
        );

    \I__4333\ : LocalMux
    port map (
            O => \N__21297\,
            I => \N__21288\
        );

    \I__4332\ : Span4Mux_h
    port map (
            O => \N__21294\,
            I => \N__21285\
        );

    \I__4331\ : Odrv4
    port map (
            O => \N__21291\,
            I => \eeprom.n3204\
        );

    \I__4330\ : Odrv12
    port map (
            O => \N__21288\,
            I => \eeprom.n3204\
        );

    \I__4329\ : Odrv4
    port map (
            O => \N__21285\,
            I => \eeprom.n3204\
        );

    \I__4328\ : CascadeMux
    port map (
            O => \N__21278\,
            I => \N__21275\
        );

    \I__4327\ : InMux
    port map (
            O => \N__21275\,
            I => \N__21272\
        );

    \I__4326\ : LocalMux
    port map (
            O => \N__21272\,
            I => \eeprom.n3179\
        );

    \I__4325\ : InMux
    port map (
            O => \N__21269\,
            I => \N__21266\
        );

    \I__4324\ : LocalMux
    port map (
            O => \N__21266\,
            I => \N__21261\
        );

    \I__4323\ : InMux
    port map (
            O => \N__21265\,
            I => \N__21258\
        );

    \I__4322\ : CascadeMux
    port map (
            O => \N__21264\,
            I => \N__21255\
        );

    \I__4321\ : Span4Mux_v
    port map (
            O => \N__21261\,
            I => \N__21252\
        );

    \I__4320\ : LocalMux
    port map (
            O => \N__21258\,
            I => \N__21249\
        );

    \I__4319\ : InMux
    port map (
            O => \N__21255\,
            I => \N__21246\
        );

    \I__4318\ : Span4Mux_h
    port map (
            O => \N__21252\,
            I => \N__21241\
        );

    \I__4317\ : Span4Mux_v
    port map (
            O => \N__21249\,
            I => \N__21241\
        );

    \I__4316\ : LocalMux
    port map (
            O => \N__21246\,
            I => \N__21238\
        );

    \I__4315\ : Odrv4
    port map (
            O => \N__21241\,
            I => \eeprom.n3211\
        );

    \I__4314\ : Odrv12
    port map (
            O => \N__21238\,
            I => \eeprom.n3211\
        );

    \I__4313\ : InMux
    port map (
            O => \N__21233\,
            I => \N__21230\
        );

    \I__4312\ : LocalMux
    port map (
            O => \N__21230\,
            I => \eeprom.n31_adj_496\
        );

    \I__4311\ : InMux
    port map (
            O => \N__21227\,
            I => \N__21224\
        );

    \I__4310\ : LocalMux
    port map (
            O => \N__21224\,
            I => \eeprom.n29_adj_497\
        );

    \I__4309\ : CascadeMux
    port map (
            O => \N__21221\,
            I => \eeprom.n30_adj_495_cascade_\
        );

    \I__4308\ : InMux
    port map (
            O => \N__21218\,
            I => \N__21215\
        );

    \I__4307\ : LocalMux
    port map (
            O => \N__21215\,
            I => \N__21212\
        );

    \I__4306\ : Odrv4
    port map (
            O => \N__21212\,
            I => \eeprom.n32_adj_494\
        );

    \I__4305\ : CascadeMux
    port map (
            O => \N__21209\,
            I => \eeprom.n3606_adj_446_cascade_\
        );

    \I__4304\ : CascadeMux
    port map (
            O => \N__21206\,
            I => \eeprom.n4451_cascade_\
        );

    \I__4303\ : InMux
    port map (
            O => \N__21203\,
            I => \N__21200\
        );

    \I__4302\ : LocalMux
    port map (
            O => \N__21200\,
            I => \eeprom.n4453\
        );

    \I__4301\ : CascadeMux
    port map (
            O => \N__21197\,
            I => \eeprom.n3599_adj_450_cascade_\
        );

    \I__4300\ : InMux
    port map (
            O => \N__21194\,
            I => \N__21191\
        );

    \I__4299\ : LocalMux
    port map (
            O => \N__21191\,
            I => \N__21188\
        );

    \I__4298\ : Odrv4
    port map (
            O => \N__21188\,
            I => \eeprom.n4429\
        );

    \I__4297\ : InMux
    port map (
            O => \N__21185\,
            I => \N__21182\
        );

    \I__4296\ : LocalMux
    port map (
            O => \N__21182\,
            I => \N__21179\
        );

    \I__4295\ : Span4Mux_v
    port map (
            O => \N__21179\,
            I => \N__21176\
        );

    \I__4294\ : Sp12to4
    port map (
            O => \N__21176\,
            I => \N__21173\
        );

    \I__4293\ : Odrv12
    port map (
            O => \N__21173\,
            I => \eeprom.n29\
        );

    \I__4292\ : CascadeMux
    port map (
            O => \N__21170\,
            I => \eeprom.n28_adj_493_cascade_\
        );

    \I__4291\ : CascadeMux
    port map (
            O => \N__21167\,
            I => \eeprom.n18_adj_488_cascade_\
        );

    \I__4290\ : InMux
    port map (
            O => \N__21164\,
            I => \N__21161\
        );

    \I__4289\ : LocalMux
    port map (
            O => \N__21161\,
            I => \N__21158\
        );

    \I__4288\ : Odrv4
    port map (
            O => \N__21158\,
            I => \eeprom.n29_adj_491\
        );

    \I__4287\ : InMux
    port map (
            O => \N__21155\,
            I => \N__21152\
        );

    \I__4286\ : LocalMux
    port map (
            O => \N__21152\,
            I => \eeprom.n28_adj_490\
        );

    \I__4285\ : CascadeMux
    port map (
            O => \N__21149\,
            I => \eeprom.n30_adj_489_cascade_\
        );

    \I__4284\ : InMux
    port map (
            O => \N__21146\,
            I => \N__21143\
        );

    \I__4283\ : LocalMux
    port map (
            O => \N__21143\,
            I => \N__21140\
        );

    \I__4282\ : Odrv4
    port map (
            O => \N__21140\,
            I => \eeprom.n27_adj_492\
        );

    \I__4281\ : CascadeMux
    port map (
            O => \N__21137\,
            I => \eeprom.n3430_cascade_\
        );

    \I__4280\ : InMux
    port map (
            O => \N__21134\,
            I => \N__21131\
        );

    \I__4279\ : LocalMux
    port map (
            O => \N__21131\,
            I => \eeprom.n3609_adj_445\
        );

    \I__4278\ : CascadeMux
    port map (
            O => \N__21128\,
            I => \eeprom.n3508_cascade_\
        );

    \I__4277\ : InMux
    port map (
            O => \N__21125\,
            I => \eeprom.n3685\
        );

    \I__4276\ : InMux
    port map (
            O => \N__21122\,
            I => \N__21119\
        );

    \I__4275\ : LocalMux
    port map (
            O => \N__21119\,
            I => \N__21116\
        );

    \I__4274\ : Odrv4
    port map (
            O => \N__21116\,
            I => \eeprom.n2971\
        );

    \I__4273\ : CascadeMux
    port map (
            O => \N__21113\,
            I => \N__21110\
        );

    \I__4272\ : InMux
    port map (
            O => \N__21110\,
            I => \N__21107\
        );

    \I__4271\ : LocalMux
    port map (
            O => \N__21107\,
            I => \N__21103\
        );

    \I__4270\ : InMux
    port map (
            O => \N__21106\,
            I => \N__21100\
        );

    \I__4269\ : Span4Mux_v
    port map (
            O => \N__21103\,
            I => \N__21095\
        );

    \I__4268\ : LocalMux
    port map (
            O => \N__21100\,
            I => \N__21095\
        );

    \I__4267\ : Span4Mux_h
    port map (
            O => \N__21095\,
            I => \N__21092\
        );

    \I__4266\ : Odrv4
    port map (
            O => \N__21092\,
            I => \eeprom.n2904\
        );

    \I__4265\ : InMux
    port map (
            O => \N__21089\,
            I => \N__21086\
        );

    \I__4264\ : LocalMux
    port map (
            O => \N__21086\,
            I => \N__21083\
        );

    \I__4263\ : Odrv4
    port map (
            O => \N__21083\,
            I => \eeprom.n2977\
        );

    \I__4262\ : CascadeMux
    port map (
            O => \N__21080\,
            I => \N__21077\
        );

    \I__4261\ : InMux
    port map (
            O => \N__21077\,
            I => \N__21073\
        );

    \I__4260\ : InMux
    port map (
            O => \N__21076\,
            I => \N__21069\
        );

    \I__4259\ : LocalMux
    port map (
            O => \N__21073\,
            I => \N__21066\
        );

    \I__4258\ : InMux
    port map (
            O => \N__21072\,
            I => \N__21063\
        );

    \I__4257\ : LocalMux
    port map (
            O => \N__21069\,
            I => \eeprom.n2910\
        );

    \I__4256\ : Odrv4
    port map (
            O => \N__21066\,
            I => \eeprom.n2910\
        );

    \I__4255\ : LocalMux
    port map (
            O => \N__21063\,
            I => \eeprom.n2910\
        );

    \I__4254\ : CascadeMux
    port map (
            O => \N__21056\,
            I => \eeprom.n3497_cascade_\
        );

    \I__4253\ : CascadeMux
    port map (
            O => \N__21053\,
            I => \N__21050\
        );

    \I__4252\ : InMux
    port map (
            O => \N__21050\,
            I => \N__21047\
        );

    \I__4251\ : LocalMux
    port map (
            O => \N__21047\,
            I => \N__21044\
        );

    \I__4250\ : Span4Mux_v
    port map (
            O => \N__21044\,
            I => \N__21041\
        );

    \I__4249\ : Odrv4
    port map (
            O => \N__21041\,
            I => \eeprom.n3176\
        );

    \I__4248\ : InMux
    port map (
            O => \N__21038\,
            I => \eeprom.n3676\
        );

    \I__4247\ : InMux
    port map (
            O => \N__21035\,
            I => \eeprom.n3677\
        );

    \I__4246\ : InMux
    port map (
            O => \N__21032\,
            I => \N__21029\
        );

    \I__4245\ : LocalMux
    port map (
            O => \N__21029\,
            I => \N__21026\
        );

    \I__4244\ : Odrv12
    port map (
            O => \N__21026\,
            I => \eeprom.n3174\
        );

    \I__4243\ : InMux
    port map (
            O => \N__21023\,
            I => \eeprom.n3678\
        );

    \I__4242\ : InMux
    port map (
            O => \N__21020\,
            I => \eeprom.n3679\
        );

    \I__4241\ : InMux
    port map (
            O => \N__21017\,
            I => \eeprom.n3680\
        );

    \I__4240\ : InMux
    port map (
            O => \N__21014\,
            I => \N__21011\
        );

    \I__4239\ : LocalMux
    port map (
            O => \N__21011\,
            I => \N__21008\
        );

    \I__4238\ : Odrv12
    port map (
            O => \N__21008\,
            I => \eeprom.n3171\
        );

    \I__4237\ : InMux
    port map (
            O => \N__21005\,
            I => \eeprom.n3681\
        );

    \I__4236\ : InMux
    port map (
            O => \N__21002\,
            I => \bfn_12_24_0_\
        );

    \I__4235\ : InMux
    port map (
            O => \N__20999\,
            I => \eeprom.n3683\
        );

    \I__4234\ : InMux
    port map (
            O => \N__20996\,
            I => \eeprom.n3684\
        );

    \I__4233\ : CascadeMux
    port map (
            O => \N__20993\,
            I => \N__20990\
        );

    \I__4232\ : InMux
    port map (
            O => \N__20990\,
            I => \N__20987\
        );

    \I__4231\ : LocalMux
    port map (
            O => \N__20987\,
            I => \N__20984\
        );

    \I__4230\ : Odrv4
    port map (
            O => \N__20984\,
            I => \eeprom.n3184\
        );

    \I__4229\ : InMux
    port map (
            O => \N__20981\,
            I => \eeprom.n3668\
        );

    \I__4228\ : CascadeMux
    port map (
            O => \N__20978\,
            I => \N__20975\
        );

    \I__4227\ : InMux
    port map (
            O => \N__20975\,
            I => \N__20971\
        );

    \I__4226\ : InMux
    port map (
            O => \N__20974\,
            I => \N__20968\
        );

    \I__4225\ : LocalMux
    port map (
            O => \N__20971\,
            I => \N__20965\
        );

    \I__4224\ : LocalMux
    port map (
            O => \N__20968\,
            I => \eeprom.n3116\
        );

    \I__4223\ : Odrv4
    port map (
            O => \N__20965\,
            I => \eeprom.n3116\
        );

    \I__4222\ : InMux
    port map (
            O => \N__20960\,
            I => \N__20957\
        );

    \I__4221\ : LocalMux
    port map (
            O => \N__20957\,
            I => \N__20954\
        );

    \I__4220\ : Odrv4
    port map (
            O => \N__20954\,
            I => \eeprom.n3183\
        );

    \I__4219\ : InMux
    port map (
            O => \N__20951\,
            I => \eeprom.n3669\
        );

    \I__4218\ : InMux
    port map (
            O => \N__20948\,
            I => \N__20945\
        );

    \I__4217\ : LocalMux
    port map (
            O => \N__20945\,
            I => \eeprom.n3182\
        );

    \I__4216\ : InMux
    port map (
            O => \N__20942\,
            I => \eeprom.n3670\
        );

    \I__4215\ : CascadeMux
    port map (
            O => \N__20939\,
            I => \N__20936\
        );

    \I__4214\ : InMux
    port map (
            O => \N__20936\,
            I => \N__20933\
        );

    \I__4213\ : LocalMux
    port map (
            O => \N__20933\,
            I => \N__20930\
        );

    \I__4212\ : Odrv4
    port map (
            O => \N__20930\,
            I => \eeprom.n3181\
        );

    \I__4211\ : InMux
    port map (
            O => \N__20927\,
            I => \eeprom.n3671\
        );

    \I__4210\ : CascadeMux
    port map (
            O => \N__20924\,
            I => \N__20921\
        );

    \I__4209\ : InMux
    port map (
            O => \N__20921\,
            I => \N__20918\
        );

    \I__4208\ : LocalMux
    port map (
            O => \N__20918\,
            I => \N__20914\
        );

    \I__4207\ : InMux
    port map (
            O => \N__20917\,
            I => \N__20911\
        );

    \I__4206\ : Odrv4
    port map (
            O => \N__20914\,
            I => \eeprom.n3113\
        );

    \I__4205\ : LocalMux
    port map (
            O => \N__20911\,
            I => \eeprom.n3113\
        );

    \I__4204\ : InMux
    port map (
            O => \N__20906\,
            I => \N__20903\
        );

    \I__4203\ : LocalMux
    port map (
            O => \N__20903\,
            I => \N__20900\
        );

    \I__4202\ : Span4Mux_h
    port map (
            O => \N__20900\,
            I => \N__20897\
        );

    \I__4201\ : Odrv4
    port map (
            O => \N__20897\,
            I => \eeprom.n3180\
        );

    \I__4200\ : InMux
    port map (
            O => \N__20894\,
            I => \eeprom.n3672\
        );

    \I__4199\ : InMux
    port map (
            O => \N__20891\,
            I => \eeprom.n3673\
        );

    \I__4198\ : InMux
    port map (
            O => \N__20888\,
            I => \N__20885\
        );

    \I__4197\ : LocalMux
    port map (
            O => \N__20885\,
            I => \N__20882\
        );

    \I__4196\ : Span4Mux_h
    port map (
            O => \N__20882\,
            I => \N__20879\
        );

    \I__4195\ : Odrv4
    port map (
            O => \N__20879\,
            I => \eeprom.n3178\
        );

    \I__4194\ : InMux
    port map (
            O => \N__20876\,
            I => \bfn_12_23_0_\
        );

    \I__4193\ : CascadeMux
    port map (
            O => \N__20873\,
            I => \N__20870\
        );

    \I__4192\ : InMux
    port map (
            O => \N__20870\,
            I => \N__20867\
        );

    \I__4191\ : LocalMux
    port map (
            O => \N__20867\,
            I => \N__20864\
        );

    \I__4190\ : Span4Mux_h
    port map (
            O => \N__20864\,
            I => \N__20861\
        );

    \I__4189\ : Odrv4
    port map (
            O => \N__20861\,
            I => \eeprom.n3177\
        );

    \I__4188\ : InMux
    port map (
            O => \N__20858\,
            I => \eeprom.n3675\
        );

    \I__4187\ : CascadeMux
    port map (
            O => \N__20855\,
            I => \eeprom.n18_adj_432_cascade_\
        );

    \I__4186\ : CascadeMux
    port map (
            O => \N__20852\,
            I => \eeprom.n26_adj_466_cascade_\
        );

    \I__4185\ : CascadeMux
    port map (
            O => \N__20849\,
            I => \eeprom.n4711_cascade_\
        );

    \I__4184\ : InMux
    port map (
            O => \N__20846\,
            I => \N__20843\
        );

    \I__4183\ : LocalMux
    port map (
            O => \N__20843\,
            I => \eeprom.n4715\
        );

    \I__4182\ : CascadeMux
    port map (
            O => \N__20840\,
            I => \N__20837\
        );

    \I__4181\ : InMux
    port map (
            O => \N__20837\,
            I => \N__20834\
        );

    \I__4180\ : LocalMux
    port map (
            O => \N__20834\,
            I => \N__20831\
        );

    \I__4179\ : Span4Mux_v
    port map (
            O => \N__20831\,
            I => \N__20826\
        );

    \I__4178\ : InMux
    port map (
            O => \N__20830\,
            I => \N__20823\
        );

    \I__4177\ : CascadeMux
    port map (
            O => \N__20829\,
            I => \N__20820\
        );

    \I__4176\ : Span4Mux_h
    port map (
            O => \N__20826\,
            I => \N__20817\
        );

    \I__4175\ : LocalMux
    port map (
            O => \N__20823\,
            I => \N__20814\
        );

    \I__4174\ : InMux
    port map (
            O => \N__20820\,
            I => \N__20811\
        );

    \I__4173\ : Odrv4
    port map (
            O => \N__20817\,
            I => \eeprom.n3206\
        );

    \I__4172\ : Odrv4
    port map (
            O => \N__20814\,
            I => \eeprom.n3206\
        );

    \I__4171\ : LocalMux
    port map (
            O => \N__20811\,
            I => \eeprom.n3206\
        );

    \I__4170\ : InMux
    port map (
            O => \N__20804\,
            I => \N__20800\
        );

    \I__4169\ : CascadeMux
    port map (
            O => \N__20803\,
            I => \N__20797\
        );

    \I__4168\ : LocalMux
    port map (
            O => \N__20800\,
            I => \N__20793\
        );

    \I__4167\ : InMux
    port map (
            O => \N__20797\,
            I => \N__20790\
        );

    \I__4166\ : CascadeMux
    port map (
            O => \N__20796\,
            I => \N__20787\
        );

    \I__4165\ : Span4Mux_v
    port map (
            O => \N__20793\,
            I => \N__20782\
        );

    \I__4164\ : LocalMux
    port map (
            O => \N__20790\,
            I => \N__20782\
        );

    \I__4163\ : InMux
    port map (
            O => \N__20787\,
            I => \N__20779\
        );

    \I__4162\ : Span4Mux_h
    port map (
            O => \N__20782\,
            I => \N__20776\
        );

    \I__4161\ : LocalMux
    port map (
            O => \N__20779\,
            I => \N__20773\
        );

    \I__4160\ : Odrv4
    port map (
            O => \N__20776\,
            I => \eeprom.n3214\
        );

    \I__4159\ : Odrv4
    port map (
            O => \N__20773\,
            I => \eeprom.n3214\
        );

    \I__4158\ : InMux
    port map (
            O => \N__20768\,
            I => \N__20764\
        );

    \I__4157\ : InMux
    port map (
            O => \N__20767\,
            I => \N__20760\
        );

    \I__4156\ : LocalMux
    port map (
            O => \N__20764\,
            I => \N__20757\
        );

    \I__4155\ : InMux
    port map (
            O => \N__20763\,
            I => \N__20754\
        );

    \I__4154\ : LocalMux
    port map (
            O => \N__20760\,
            I => \N__20751\
        );

    \I__4153\ : Span4Mux_v
    port map (
            O => \N__20757\,
            I => \N__20748\
        );

    \I__4152\ : LocalMux
    port map (
            O => \N__20754\,
            I => \N__20745\
        );

    \I__4151\ : Span4Mux_h
    port map (
            O => \N__20751\,
            I => \N__20742\
        );

    \I__4150\ : Span4Mux_v
    port map (
            O => \N__20748\,
            I => \N__20737\
        );

    \I__4149\ : Span4Mux_v
    port map (
            O => \N__20745\,
            I => \N__20737\
        );

    \I__4148\ : Span4Mux_h
    port map (
            O => \N__20742\,
            I => \N__20734\
        );

    \I__4147\ : Span4Mux_h
    port map (
            O => \N__20737\,
            I => \N__20731\
        );

    \I__4146\ : Odrv4
    port map (
            O => \N__20734\,
            I => \eeprom.n3119\
        );

    \I__4145\ : Odrv4
    port map (
            O => \N__20731\,
            I => \eeprom.n3119\
        );

    \I__4144\ : InMux
    port map (
            O => \N__20726\,
            I => \N__20723\
        );

    \I__4143\ : LocalMux
    port map (
            O => \N__20723\,
            I => \N__20720\
        );

    \I__4142\ : Span4Mux_v
    port map (
            O => \N__20720\,
            I => \N__20717\
        );

    \I__4141\ : Span4Mux_h
    port map (
            O => \N__20717\,
            I => \N__20714\
        );

    \I__4140\ : Odrv4
    port map (
            O => \N__20714\,
            I => \eeprom.n3186\
        );

    \I__4139\ : InMux
    port map (
            O => \N__20711\,
            I => \bfn_12_22_0_\
        );

    \I__4138\ : CascadeMux
    port map (
            O => \N__20708\,
            I => \N__20705\
        );

    \I__4137\ : InMux
    port map (
            O => \N__20705\,
            I => \N__20702\
        );

    \I__4136\ : LocalMux
    port map (
            O => \N__20702\,
            I => \N__20699\
        );

    \I__4135\ : Odrv4
    port map (
            O => \N__20699\,
            I => \eeprom.n3185\
        );

    \I__4134\ : InMux
    port map (
            O => \N__20696\,
            I => \eeprom.n3667\
        );

    \I__4133\ : CascadeMux
    port map (
            O => \N__20693\,
            I => \N__20689\
        );

    \I__4132\ : InMux
    port map (
            O => \N__20692\,
            I => \N__20685\
        );

    \I__4131\ : InMux
    port map (
            O => \N__20689\,
            I => \N__20682\
        );

    \I__4130\ : InMux
    port map (
            O => \N__20688\,
            I => \N__20679\
        );

    \I__4129\ : LocalMux
    port map (
            O => \N__20685\,
            I => \N__20674\
        );

    \I__4128\ : LocalMux
    port map (
            O => \N__20682\,
            I => \N__20674\
        );

    \I__4127\ : LocalMux
    port map (
            O => \N__20679\,
            I => \N__20671\
        );

    \I__4126\ : Odrv4
    port map (
            O => \N__20674\,
            I => \eeprom.n3303\
        );

    \I__4125\ : Odrv4
    port map (
            O => \N__20671\,
            I => \eeprom.n3303\
        );

    \I__4124\ : InMux
    port map (
            O => \N__20666\,
            I => \N__20663\
        );

    \I__4123\ : LocalMux
    port map (
            O => \N__20663\,
            I => \N__20660\
        );

    \I__4122\ : Odrv4
    port map (
            O => \N__20660\,
            I => \eeprom.n3370\
        );

    \I__4121\ : InMux
    port map (
            O => \N__20657\,
            I => \N__20654\
        );

    \I__4120\ : LocalMux
    port map (
            O => \N__20654\,
            I => \N__20651\
        );

    \I__4119\ : Odrv4
    port map (
            O => \N__20651\,
            I => \eeprom.n3366\
        );

    \I__4118\ : CascadeMux
    port map (
            O => \N__20648\,
            I => \N__20644\
        );

    \I__4117\ : CascadeMux
    port map (
            O => \N__20647\,
            I => \N__20640\
        );

    \I__4116\ : InMux
    port map (
            O => \N__20644\,
            I => \N__20637\
        );

    \I__4115\ : InMux
    port map (
            O => \N__20643\,
            I => \N__20634\
        );

    \I__4114\ : InMux
    port map (
            O => \N__20640\,
            I => \N__20631\
        );

    \I__4113\ : LocalMux
    port map (
            O => \N__20637\,
            I => \N__20626\
        );

    \I__4112\ : LocalMux
    port map (
            O => \N__20634\,
            I => \N__20626\
        );

    \I__4111\ : LocalMux
    port map (
            O => \N__20631\,
            I => \N__20623\
        );

    \I__4110\ : Span4Mux_v
    port map (
            O => \N__20626\,
            I => \N__20620\
        );

    \I__4109\ : Odrv4
    port map (
            O => \N__20623\,
            I => \eeprom.n3299\
        );

    \I__4108\ : Odrv4
    port map (
            O => \N__20620\,
            I => \eeprom.n3299\
        );

    \I__4107\ : CascadeMux
    port map (
            O => \N__20615\,
            I => \N__20612\
        );

    \I__4106\ : InMux
    port map (
            O => \N__20612\,
            I => \N__20603\
        );

    \I__4105\ : CascadeMux
    port map (
            O => \N__20611\,
            I => \N__20600\
        );

    \I__4104\ : CascadeMux
    port map (
            O => \N__20610\,
            I => \N__20592\
        );

    \I__4103\ : CascadeMux
    port map (
            O => \N__20609\,
            I => \N__20589\
        );

    \I__4102\ : CascadeMux
    port map (
            O => \N__20608\,
            I => \N__20582\
        );

    \I__4101\ : InMux
    port map (
            O => \N__20607\,
            I => \N__20573\
        );

    \I__4100\ : InMux
    port map (
            O => \N__20606\,
            I => \N__20573\
        );

    \I__4099\ : LocalMux
    port map (
            O => \N__20603\,
            I => \N__20570\
        );

    \I__4098\ : InMux
    port map (
            O => \N__20600\,
            I => \N__20567\
        );

    \I__4097\ : CascadeMux
    port map (
            O => \N__20599\,
            I => \N__20564\
        );

    \I__4096\ : CascadeMux
    port map (
            O => \N__20598\,
            I => \N__20561\
        );

    \I__4095\ : CascadeMux
    port map (
            O => \N__20597\,
            I => \N__20558\
        );

    \I__4094\ : InMux
    port map (
            O => \N__20596\,
            I => \N__20554\
        );

    \I__4093\ : InMux
    port map (
            O => \N__20595\,
            I => \N__20551\
        );

    \I__4092\ : InMux
    port map (
            O => \N__20592\,
            I => \N__20544\
        );

    \I__4091\ : InMux
    port map (
            O => \N__20589\,
            I => \N__20544\
        );

    \I__4090\ : InMux
    port map (
            O => \N__20588\,
            I => \N__20544\
        );

    \I__4089\ : InMux
    port map (
            O => \N__20587\,
            I => \N__20539\
        );

    \I__4088\ : InMux
    port map (
            O => \N__20586\,
            I => \N__20539\
        );

    \I__4087\ : InMux
    port map (
            O => \N__20585\,
            I => \N__20532\
        );

    \I__4086\ : InMux
    port map (
            O => \N__20582\,
            I => \N__20532\
        );

    \I__4085\ : InMux
    port map (
            O => \N__20581\,
            I => \N__20532\
        );

    \I__4084\ : InMux
    port map (
            O => \N__20580\,
            I => \N__20527\
        );

    \I__4083\ : InMux
    port map (
            O => \N__20579\,
            I => \N__20527\
        );

    \I__4082\ : InMux
    port map (
            O => \N__20578\,
            I => \N__20524\
        );

    \I__4081\ : LocalMux
    port map (
            O => \N__20573\,
            I => \N__20519\
        );

    \I__4080\ : Span4Mux_v
    port map (
            O => \N__20570\,
            I => \N__20519\
        );

    \I__4079\ : LocalMux
    port map (
            O => \N__20567\,
            I => \N__20516\
        );

    \I__4078\ : InMux
    port map (
            O => \N__20564\,
            I => \N__20507\
        );

    \I__4077\ : InMux
    port map (
            O => \N__20561\,
            I => \N__20507\
        );

    \I__4076\ : InMux
    port map (
            O => \N__20558\,
            I => \N__20507\
        );

    \I__4075\ : InMux
    port map (
            O => \N__20557\,
            I => \N__20507\
        );

    \I__4074\ : LocalMux
    port map (
            O => \N__20554\,
            I => \eeprom.n3331\
        );

    \I__4073\ : LocalMux
    port map (
            O => \N__20551\,
            I => \eeprom.n3331\
        );

    \I__4072\ : LocalMux
    port map (
            O => \N__20544\,
            I => \eeprom.n3331\
        );

    \I__4071\ : LocalMux
    port map (
            O => \N__20539\,
            I => \eeprom.n3331\
        );

    \I__4070\ : LocalMux
    port map (
            O => \N__20532\,
            I => \eeprom.n3331\
        );

    \I__4069\ : LocalMux
    port map (
            O => \N__20527\,
            I => \eeprom.n3331\
        );

    \I__4068\ : LocalMux
    port map (
            O => \N__20524\,
            I => \eeprom.n3331\
        );

    \I__4067\ : Odrv4
    port map (
            O => \N__20519\,
            I => \eeprom.n3331\
        );

    \I__4066\ : Odrv4
    port map (
            O => \N__20516\,
            I => \eeprom.n3331\
        );

    \I__4065\ : LocalMux
    port map (
            O => \N__20507\,
            I => \eeprom.n3331\
        );

    \I__4064\ : CascadeMux
    port map (
            O => \N__20486\,
            I => \eeprom.n3500_cascade_\
        );

    \I__4063\ : InMux
    port map (
            O => \N__20483\,
            I => \N__20479\
        );

    \I__4062\ : CascadeMux
    port map (
            O => \N__20482\,
            I => \N__20476\
        );

    \I__4061\ : LocalMux
    port map (
            O => \N__20479\,
            I => \N__20473\
        );

    \I__4060\ : InMux
    port map (
            O => \N__20476\,
            I => \N__20470\
        );

    \I__4059\ : Span4Mux_h
    port map (
            O => \N__20473\,
            I => \N__20466\
        );

    \I__4058\ : LocalMux
    port map (
            O => \N__20470\,
            I => \N__20463\
        );

    \I__4057\ : InMux
    port map (
            O => \N__20469\,
            I => \N__20460\
        );

    \I__4056\ : Odrv4
    port map (
            O => \N__20466\,
            I => \eeprom.n3216\
        );

    \I__4055\ : Odrv4
    port map (
            O => \N__20463\,
            I => \eeprom.n3216\
        );

    \I__4054\ : LocalMux
    port map (
            O => \N__20460\,
            I => \eeprom.n3216\
        );

    \I__4053\ : CascadeMux
    port map (
            O => \N__20453\,
            I => \N__20450\
        );

    \I__4052\ : InMux
    port map (
            O => \N__20450\,
            I => \N__20446\
        );

    \I__4051\ : InMux
    port map (
            O => \N__20449\,
            I => \N__20443\
        );

    \I__4050\ : LocalMux
    port map (
            O => \N__20446\,
            I => \N__20438\
        );

    \I__4049\ : LocalMux
    port map (
            O => \N__20443\,
            I => \N__20438\
        );

    \I__4048\ : Span4Mux_h
    port map (
            O => \N__20438\,
            I => \N__20434\
        );

    \I__4047\ : InMux
    port map (
            O => \N__20437\,
            I => \N__20431\
        );

    \I__4046\ : Odrv4
    port map (
            O => \N__20434\,
            I => \eeprom.n3203\
        );

    \I__4045\ : LocalMux
    port map (
            O => \N__20431\,
            I => \eeprom.n3203\
        );

    \I__4044\ : CascadeMux
    port map (
            O => \N__20426\,
            I => \N__20422\
        );

    \I__4043\ : CascadeMux
    port map (
            O => \N__20425\,
            I => \N__20419\
        );

    \I__4042\ : InMux
    port map (
            O => \N__20422\,
            I => \N__20416\
        );

    \I__4041\ : InMux
    port map (
            O => \N__20419\,
            I => \N__20412\
        );

    \I__4040\ : LocalMux
    port map (
            O => \N__20416\,
            I => \N__20409\
        );

    \I__4039\ : InMux
    port map (
            O => \N__20415\,
            I => \N__20406\
        );

    \I__4038\ : LocalMux
    port map (
            O => \N__20412\,
            I => \eeprom.n3217\
        );

    \I__4037\ : Odrv12
    port map (
            O => \N__20409\,
            I => \eeprom.n3217\
        );

    \I__4036\ : LocalMux
    port map (
            O => \N__20406\,
            I => \eeprom.n3217\
        );

    \I__4035\ : CascadeMux
    port map (
            O => \N__20399\,
            I => \eeprom.n3410_cascade_\
        );

    \I__4034\ : CascadeMux
    port map (
            O => \N__20396\,
            I => \eeprom.n3505_cascade_\
        );

    \I__4033\ : InMux
    port map (
            O => \N__20393\,
            I => \N__20390\
        );

    \I__4032\ : LocalMux
    port map (
            O => \N__20390\,
            I => \N__20387\
        );

    \I__4031\ : Span4Mux_h
    port map (
            O => \N__20387\,
            I => \N__20382\
        );

    \I__4030\ : InMux
    port map (
            O => \N__20386\,
            I => \N__20379\
        );

    \I__4029\ : InMux
    port map (
            O => \N__20385\,
            I => \N__20376\
        );

    \I__4028\ : Odrv4
    port map (
            O => \N__20382\,
            I => \eeprom.n3310\
        );

    \I__4027\ : LocalMux
    port map (
            O => \N__20379\,
            I => \eeprom.n3310\
        );

    \I__4026\ : LocalMux
    port map (
            O => \N__20376\,
            I => \eeprom.n3310\
        );

    \I__4025\ : CascadeMux
    port map (
            O => \N__20369\,
            I => \N__20366\
        );

    \I__4024\ : InMux
    port map (
            O => \N__20366\,
            I => \N__20363\
        );

    \I__4023\ : LocalMux
    port map (
            O => \N__20363\,
            I => \N__20360\
        );

    \I__4022\ : Odrv4
    port map (
            O => \N__20360\,
            I => \eeprom.n3377\
        );

    \I__4021\ : CascadeMux
    port map (
            O => \N__20357\,
            I => \eeprom.n3608_adj_451_cascade_\
        );

    \I__4020\ : InMux
    port map (
            O => \N__20354\,
            I => \N__20349\
        );

    \I__4019\ : CascadeMux
    port map (
            O => \N__20353\,
            I => \N__20346\
        );

    \I__4018\ : InMux
    port map (
            O => \N__20352\,
            I => \N__20343\
        );

    \I__4017\ : LocalMux
    port map (
            O => \N__20349\,
            I => \N__20340\
        );

    \I__4016\ : InMux
    port map (
            O => \N__20346\,
            I => \N__20337\
        );

    \I__4015\ : LocalMux
    port map (
            O => \N__20343\,
            I => \N__20334\
        );

    \I__4014\ : Span4Mux_h
    port map (
            O => \N__20340\,
            I => \N__20331\
        );

    \I__4013\ : LocalMux
    port map (
            O => \N__20337\,
            I => \N__20328\
        );

    \I__4012\ : Odrv12
    port map (
            O => \N__20334\,
            I => \eeprom.n3313\
        );

    \I__4011\ : Odrv4
    port map (
            O => \N__20331\,
            I => \eeprom.n3313\
        );

    \I__4010\ : Odrv4
    port map (
            O => \N__20328\,
            I => \eeprom.n3313\
        );

    \I__4009\ : CascadeMux
    port map (
            O => \N__20321\,
            I => \N__20318\
        );

    \I__4008\ : InMux
    port map (
            O => \N__20318\,
            I => \N__20315\
        );

    \I__4007\ : LocalMux
    port map (
            O => \N__20315\,
            I => \N__20312\
        );

    \I__4006\ : Span4Mux_h
    port map (
            O => \N__20312\,
            I => \N__20309\
        );

    \I__4005\ : Odrv4
    port map (
            O => \N__20309\,
            I => \eeprom.n3380\
        );

    \I__4004\ : CascadeMux
    port map (
            O => \N__20306\,
            I => \eeprom.n3412_cascade_\
        );

    \I__4003\ : CascadeMux
    port map (
            O => \N__20303\,
            I => \eeprom.n3414_cascade_\
        );

    \I__4002\ : CascadeMux
    port map (
            O => \N__20300\,
            I => \eeprom.n4689_cascade_\
        );

    \I__4001\ : CascadeMux
    port map (
            O => \N__20297\,
            I => \eeprom.n4144_cascade_\
        );

    \I__4000\ : InMux
    port map (
            O => \N__20294\,
            I => \N__20291\
        );

    \I__3999\ : LocalMux
    port map (
            O => \N__20291\,
            I => \N__20288\
        );

    \I__3998\ : Span4Mux_h
    port map (
            O => \N__20288\,
            I => \N__20285\
        );

    \I__3997\ : Odrv4
    port map (
            O => \N__20285\,
            I => \eeprom.n3386\
        );

    \I__3996\ : InMux
    port map (
            O => \N__20282\,
            I => \N__20278\
        );

    \I__3995\ : InMux
    port map (
            O => \N__20281\,
            I => \N__20275\
        );

    \I__3994\ : LocalMux
    port map (
            O => \N__20278\,
            I => \N__20269\
        );

    \I__3993\ : LocalMux
    port map (
            O => \N__20275\,
            I => \N__20269\
        );

    \I__3992\ : InMux
    port map (
            O => \N__20274\,
            I => \N__20266\
        );

    \I__3991\ : Span4Mux_h
    port map (
            O => \N__20269\,
            I => \N__20263\
        );

    \I__3990\ : LocalMux
    port map (
            O => \N__20266\,
            I => \N__20260\
        );

    \I__3989\ : Span4Mux_h
    port map (
            O => \N__20263\,
            I => \N__20257\
        );

    \I__3988\ : Span4Mux_v
    port map (
            O => \N__20260\,
            I => \N__20254\
        );

    \I__3987\ : Odrv4
    port map (
            O => \N__20257\,
            I => \eeprom.n3319\
        );

    \I__3986\ : Odrv4
    port map (
            O => \N__20254\,
            I => \eeprom.n3319\
        );

    \I__3985\ : CascadeMux
    port map (
            O => \N__20249\,
            I => \N__20245\
        );

    \I__3984\ : InMux
    port map (
            O => \N__20248\,
            I => \N__20241\
        );

    \I__3983\ : InMux
    port map (
            O => \N__20245\,
            I => \N__20238\
        );

    \I__3982\ : InMux
    port map (
            O => \N__20244\,
            I => \N__20235\
        );

    \I__3981\ : LocalMux
    port map (
            O => \N__20241\,
            I => \N__20230\
        );

    \I__3980\ : LocalMux
    port map (
            O => \N__20238\,
            I => \N__20230\
        );

    \I__3979\ : LocalMux
    port map (
            O => \N__20235\,
            I => \N__20227\
        );

    \I__3978\ : Span4Mux_h
    port map (
            O => \N__20230\,
            I => \N__20224\
        );

    \I__3977\ : Odrv4
    port map (
            O => \N__20227\,
            I => \eeprom.n3316\
        );

    \I__3976\ : Odrv4
    port map (
            O => \N__20224\,
            I => \eeprom.n3316\
        );

    \I__3975\ : CascadeMux
    port map (
            O => \N__20219\,
            I => \N__20216\
        );

    \I__3974\ : InMux
    port map (
            O => \N__20216\,
            I => \N__20213\
        );

    \I__3973\ : LocalMux
    port map (
            O => \N__20213\,
            I => \N__20210\
        );

    \I__3972\ : Odrv4
    port map (
            O => \N__20210\,
            I => \eeprom.n3383\
        );

    \I__3971\ : InMux
    port map (
            O => \N__20207\,
            I => \N__20203\
        );

    \I__3970\ : CascadeMux
    port map (
            O => \N__20206\,
            I => \N__20200\
        );

    \I__3969\ : LocalMux
    port map (
            O => \N__20203\,
            I => \N__20197\
        );

    \I__3968\ : InMux
    port map (
            O => \N__20200\,
            I => \N__20194\
        );

    \I__3967\ : Odrv12
    port map (
            O => \N__20197\,
            I => \eeprom.n3314\
        );

    \I__3966\ : LocalMux
    port map (
            O => \N__20194\,
            I => \eeprom.n3314\
        );

    \I__3965\ : InMux
    port map (
            O => \N__20189\,
            I => \N__20186\
        );

    \I__3964\ : LocalMux
    port map (
            O => \N__20186\,
            I => \N__20183\
        );

    \I__3963\ : Odrv4
    port map (
            O => \N__20183\,
            I => \eeprom.n3381\
        );

    \I__3962\ : CascadeMux
    port map (
            O => \N__20180\,
            I => \eeprom.n3413_cascade_\
        );

    \I__3961\ : InMux
    port map (
            O => \N__20177\,
            I => \N__20174\
        );

    \I__3960\ : LocalMux
    port map (
            O => \N__20174\,
            I => \eeprom.n4687\
        );

    \I__3959\ : InMux
    port map (
            O => \N__20171\,
            I => \N__20168\
        );

    \I__3958\ : LocalMux
    port map (
            O => \N__20168\,
            I => \N__20165\
        );

    \I__3957\ : Odrv12
    port map (
            O => \N__20165\,
            I => \eeprom.n3378\
        );

    \I__3956\ : CascadeMux
    port map (
            O => \N__20162\,
            I => \N__20159\
        );

    \I__3955\ : InMux
    port map (
            O => \N__20159\,
            I => \N__20156\
        );

    \I__3954\ : LocalMux
    port map (
            O => \N__20156\,
            I => \N__20152\
        );

    \I__3953\ : CascadeMux
    port map (
            O => \N__20155\,
            I => \N__20148\
        );

    \I__3952\ : Span4Mux_h
    port map (
            O => \N__20152\,
            I => \N__20145\
        );

    \I__3951\ : InMux
    port map (
            O => \N__20151\,
            I => \N__20142\
        );

    \I__3950\ : InMux
    port map (
            O => \N__20148\,
            I => \N__20139\
        );

    \I__3949\ : Odrv4
    port map (
            O => \N__20145\,
            I => \eeprom.n3311\
        );

    \I__3948\ : LocalMux
    port map (
            O => \N__20142\,
            I => \eeprom.n3311\
        );

    \I__3947\ : LocalMux
    port map (
            O => \N__20139\,
            I => \eeprom.n3311\
        );

    \I__3946\ : CascadeMux
    port map (
            O => \N__20132\,
            I => \N__20127\
        );

    \I__3945\ : CascadeMux
    port map (
            O => \N__20131\,
            I => \N__20124\
        );

    \I__3944\ : InMux
    port map (
            O => \N__20130\,
            I => \N__20121\
        );

    \I__3943\ : InMux
    port map (
            O => \N__20127\,
            I => \N__20118\
        );

    \I__3942\ : InMux
    port map (
            O => \N__20124\,
            I => \N__20115\
        );

    \I__3941\ : LocalMux
    port map (
            O => \N__20121\,
            I => \N__20112\
        );

    \I__3940\ : LocalMux
    port map (
            O => \N__20118\,
            I => \N__20107\
        );

    \I__3939\ : LocalMux
    port map (
            O => \N__20115\,
            I => \N__20107\
        );

    \I__3938\ : Span4Mux_v
    port map (
            O => \N__20112\,
            I => \N__20104\
        );

    \I__3937\ : Span4Mux_v
    port map (
            O => \N__20107\,
            I => \N__20101\
        );

    \I__3936\ : Odrv4
    port map (
            O => \N__20104\,
            I => \eeprom.n2817\
        );

    \I__3935\ : Odrv4
    port map (
            O => \N__20101\,
            I => \eeprom.n2817\
        );

    \I__3934\ : CascadeMux
    port map (
            O => \N__20096\,
            I => \N__20093\
        );

    \I__3933\ : InMux
    port map (
            O => \N__20093\,
            I => \N__20090\
        );

    \I__3932\ : LocalMux
    port map (
            O => \N__20090\,
            I => \N__20087\
        );

    \I__3931\ : Odrv4
    port map (
            O => \N__20087\,
            I => \eeprom.n2884\
        );

    \I__3930\ : CascadeMux
    port map (
            O => \N__20084\,
            I => \N__20081\
        );

    \I__3929\ : InMux
    port map (
            O => \N__20081\,
            I => \N__20078\
        );

    \I__3928\ : LocalMux
    port map (
            O => \N__20078\,
            I => \N__20075\
        );

    \I__3927\ : Odrv4
    port map (
            O => \N__20075\,
            I => \eeprom.n2877\
        );

    \I__3926\ : InMux
    port map (
            O => \N__20072\,
            I => \N__20067\
        );

    \I__3925\ : InMux
    port map (
            O => \N__20071\,
            I => \N__20064\
        );

    \I__3924\ : InMux
    port map (
            O => \N__20070\,
            I => \N__20061\
        );

    \I__3923\ : LocalMux
    port map (
            O => \N__20067\,
            I => \N__20056\
        );

    \I__3922\ : LocalMux
    port map (
            O => \N__20064\,
            I => \N__20056\
        );

    \I__3921\ : LocalMux
    port map (
            O => \N__20061\,
            I => \N__20053\
        );

    \I__3920\ : Span4Mux_h
    port map (
            O => \N__20056\,
            I => \N__20050\
        );

    \I__3919\ : Odrv4
    port map (
            O => \N__20053\,
            I => \eeprom.n2810\
        );

    \I__3918\ : Odrv4
    port map (
            O => \N__20050\,
            I => \eeprom.n2810\
        );

    \I__3917\ : CascadeMux
    port map (
            O => \N__20045\,
            I => \eeprom.n2909_cascade_\
        );

    \I__3916\ : InMux
    port map (
            O => \N__20042\,
            I => \N__20039\
        );

    \I__3915\ : LocalMux
    port map (
            O => \N__20039\,
            I => \eeprom.n18_adj_420\
        );

    \I__3914\ : CascadeMux
    port map (
            O => \N__20036\,
            I => \N__20033\
        );

    \I__3913\ : InMux
    port map (
            O => \N__20033\,
            I => \N__20030\
        );

    \I__3912\ : LocalMux
    port map (
            O => \N__20030\,
            I => \N__20027\
        );

    \I__3911\ : Odrv4
    port map (
            O => \N__20027\,
            I => \eeprom.n2975\
        );

    \I__3910\ : InMux
    port map (
            O => \N__20024\,
            I => \N__20019\
        );

    \I__3909\ : InMux
    port map (
            O => \N__20023\,
            I => \N__20016\
        );

    \I__3908\ : InMux
    port map (
            O => \N__20022\,
            I => \N__20013\
        );

    \I__3907\ : LocalMux
    port map (
            O => \N__20019\,
            I => \eeprom.n2908\
        );

    \I__3906\ : LocalMux
    port map (
            O => \N__20016\,
            I => \eeprom.n2908\
        );

    \I__3905\ : LocalMux
    port map (
            O => \N__20013\,
            I => \eeprom.n2908\
        );

    \I__3904\ : InMux
    port map (
            O => \N__20006\,
            I => \N__20003\
        );

    \I__3903\ : LocalMux
    port map (
            O => \N__20003\,
            I => \N__20000\
        );

    \I__3902\ : Odrv4
    port map (
            O => \N__20000\,
            I => \eeprom.n2878\
        );

    \I__3901\ : CascadeMux
    port map (
            O => \N__19997\,
            I => \N__19993\
        );

    \I__3900\ : CascadeMux
    port map (
            O => \N__19996\,
            I => \N__19990\
        );

    \I__3899\ : InMux
    port map (
            O => \N__19993\,
            I => \N__19987\
        );

    \I__3898\ : InMux
    port map (
            O => \N__19990\,
            I => \N__19984\
        );

    \I__3897\ : LocalMux
    port map (
            O => \N__19987\,
            I => \N__19980\
        );

    \I__3896\ : LocalMux
    port map (
            O => \N__19984\,
            I => \N__19977\
        );

    \I__3895\ : InMux
    port map (
            O => \N__19983\,
            I => \N__19974\
        );

    \I__3894\ : Odrv4
    port map (
            O => \N__19980\,
            I => \eeprom.n2811\
        );

    \I__3893\ : Odrv4
    port map (
            O => \N__19977\,
            I => \eeprom.n2811\
        );

    \I__3892\ : LocalMux
    port map (
            O => \N__19974\,
            I => \eeprom.n2811\
        );

    \I__3891\ : CascadeMux
    port map (
            O => \N__19967\,
            I => \N__19960\
        );

    \I__3890\ : CascadeMux
    port map (
            O => \N__19966\,
            I => \N__19955\
        );

    \I__3889\ : CascadeMux
    port map (
            O => \N__19965\,
            I => \N__19949\
        );

    \I__3888\ : CascadeMux
    port map (
            O => \N__19964\,
            I => \N__19945\
        );

    \I__3887\ : InMux
    port map (
            O => \N__19963\,
            I => \N__19936\
        );

    \I__3886\ : InMux
    port map (
            O => \N__19960\,
            I => \N__19936\
        );

    \I__3885\ : InMux
    port map (
            O => \N__19959\,
            I => \N__19936\
        );

    \I__3884\ : CascadeMux
    port map (
            O => \N__19958\,
            I => \N__19931\
        );

    \I__3883\ : InMux
    port map (
            O => \N__19955\,
            I => \N__19925\
        );

    \I__3882\ : InMux
    port map (
            O => \N__19954\,
            I => \N__19925\
        );

    \I__3881\ : InMux
    port map (
            O => \N__19953\,
            I => \N__19920\
        );

    \I__3880\ : InMux
    port map (
            O => \N__19952\,
            I => \N__19920\
        );

    \I__3879\ : InMux
    port map (
            O => \N__19949\,
            I => \N__19915\
        );

    \I__3878\ : InMux
    port map (
            O => \N__19948\,
            I => \N__19915\
        );

    \I__3877\ : InMux
    port map (
            O => \N__19945\,
            I => \N__19908\
        );

    \I__3876\ : InMux
    port map (
            O => \N__19944\,
            I => \N__19908\
        );

    \I__3875\ : InMux
    port map (
            O => \N__19943\,
            I => \N__19908\
        );

    \I__3874\ : LocalMux
    port map (
            O => \N__19936\,
            I => \N__19905\
        );

    \I__3873\ : InMux
    port map (
            O => \N__19935\,
            I => \N__19902\
        );

    \I__3872\ : InMux
    port map (
            O => \N__19934\,
            I => \N__19895\
        );

    \I__3871\ : InMux
    port map (
            O => \N__19931\,
            I => \N__19895\
        );

    \I__3870\ : InMux
    port map (
            O => \N__19930\,
            I => \N__19895\
        );

    \I__3869\ : LocalMux
    port map (
            O => \N__19925\,
            I => \N__19892\
        );

    \I__3868\ : LocalMux
    port map (
            O => \N__19920\,
            I => \eeprom.n2836\
        );

    \I__3867\ : LocalMux
    port map (
            O => \N__19915\,
            I => \eeprom.n2836\
        );

    \I__3866\ : LocalMux
    port map (
            O => \N__19908\,
            I => \eeprom.n2836\
        );

    \I__3865\ : Odrv4
    port map (
            O => \N__19905\,
            I => \eeprom.n2836\
        );

    \I__3864\ : LocalMux
    port map (
            O => \N__19902\,
            I => \eeprom.n2836\
        );

    \I__3863\ : LocalMux
    port map (
            O => \N__19895\,
            I => \eeprom.n2836\
        );

    \I__3862\ : Odrv4
    port map (
            O => \N__19892\,
            I => \eeprom.n2836\
        );

    \I__3861\ : CascadeMux
    port map (
            O => \N__19877\,
            I => \N__19874\
        );

    \I__3860\ : InMux
    port map (
            O => \N__19874\,
            I => \N__19870\
        );

    \I__3859\ : InMux
    port map (
            O => \N__19873\,
            I => \N__19866\
        );

    \I__3858\ : LocalMux
    port map (
            O => \N__19870\,
            I => \N__19863\
        );

    \I__3857\ : InMux
    port map (
            O => \N__19869\,
            I => \N__19860\
        );

    \I__3856\ : LocalMux
    port map (
            O => \N__19866\,
            I => \eeprom.n2915\
        );

    \I__3855\ : Odrv4
    port map (
            O => \N__19863\,
            I => \eeprom.n2915\
        );

    \I__3854\ : LocalMux
    port map (
            O => \N__19860\,
            I => \eeprom.n2915\
        );

    \I__3853\ : InMux
    port map (
            O => \N__19853\,
            I => \N__19850\
        );

    \I__3852\ : LocalMux
    port map (
            O => \N__19850\,
            I => \N__19847\
        );

    \I__3851\ : Odrv12
    port map (
            O => \N__19847\,
            I => \eeprom.n2982\
        );

    \I__3850\ : InMux
    port map (
            O => \N__19844\,
            I => \N__19839\
        );

    \I__3849\ : InMux
    port map (
            O => \N__19843\,
            I => \N__19836\
        );

    \I__3848\ : InMux
    port map (
            O => \N__19842\,
            I => \N__19833\
        );

    \I__3847\ : LocalMux
    port map (
            O => \N__19839\,
            I => \eeprom.n2911\
        );

    \I__3846\ : LocalMux
    port map (
            O => \N__19836\,
            I => \eeprom.n2911\
        );

    \I__3845\ : LocalMux
    port map (
            O => \N__19833\,
            I => \eeprom.n2911\
        );

    \I__3844\ : CascadeMux
    port map (
            O => \N__19826\,
            I => \N__19823\
        );

    \I__3843\ : InMux
    port map (
            O => \N__19823\,
            I => \N__19820\
        );

    \I__3842\ : LocalMux
    port map (
            O => \N__19820\,
            I => \N__19817\
        );

    \I__3841\ : Odrv4
    port map (
            O => \N__19817\,
            I => \eeprom.n2978\
        );

    \I__3840\ : InMux
    port map (
            O => \N__19814\,
            I => \N__19811\
        );

    \I__3839\ : LocalMux
    port map (
            O => \N__19811\,
            I => \N__19808\
        );

    \I__3838\ : Odrv4
    port map (
            O => \N__19808\,
            I => \eeprom.n2984\
        );

    \I__3837\ : CascadeMux
    port map (
            O => \N__19805\,
            I => \N__19802\
        );

    \I__3836\ : InMux
    port map (
            O => \N__19802\,
            I => \N__19798\
        );

    \I__3835\ : InMux
    port map (
            O => \N__19801\,
            I => \N__19795\
        );

    \I__3834\ : LocalMux
    port map (
            O => \N__19798\,
            I => \N__19792\
        );

    \I__3833\ : LocalMux
    port map (
            O => \N__19795\,
            I => \eeprom.n2917\
        );

    \I__3832\ : Odrv4
    port map (
            O => \N__19792\,
            I => \eeprom.n2917\
        );

    \I__3831\ : CascadeMux
    port map (
            O => \N__19787\,
            I => \N__19784\
        );

    \I__3830\ : InMux
    port map (
            O => \N__19784\,
            I => \N__19780\
        );

    \I__3829\ : InMux
    port map (
            O => \N__19783\,
            I => \N__19777\
        );

    \I__3828\ : LocalMux
    port map (
            O => \N__19780\,
            I => \N__19774\
        );

    \I__3827\ : LocalMux
    port map (
            O => \N__19777\,
            I => \eeprom.n3315\
        );

    \I__3826\ : Odrv4
    port map (
            O => \N__19774\,
            I => \eeprom.n3315\
        );

    \I__3825\ : InMux
    port map (
            O => \N__19769\,
            I => \N__19766\
        );

    \I__3824\ : LocalMux
    port map (
            O => \N__19766\,
            I => \N__19763\
        );

    \I__3823\ : Odrv4
    port map (
            O => \N__19763\,
            I => \eeprom.n3382\
        );

    \I__3822\ : InMux
    port map (
            O => \N__19760\,
            I => \eeprom.n3646\
        );

    \I__3821\ : InMux
    port map (
            O => \N__19757\,
            I => \bfn_11_23_0_\
        );

    \I__3820\ : InMux
    port map (
            O => \N__19754\,
            I => \N__19751\
        );

    \I__3819\ : LocalMux
    port map (
            O => \N__19751\,
            I => \N__19748\
        );

    \I__3818\ : Span4Mux_h
    port map (
            O => \N__19748\,
            I => \N__19744\
        );

    \I__3817\ : InMux
    port map (
            O => \N__19747\,
            I => \N__19741\
        );

    \I__3816\ : Odrv4
    port map (
            O => \N__19744\,
            I => \eeprom.n2902\
        );

    \I__3815\ : LocalMux
    port map (
            O => \N__19741\,
            I => \eeprom.n2902\
        );

    \I__3814\ : InMux
    port map (
            O => \N__19736\,
            I => \eeprom.n3648\
        );

    \I__3813\ : InMux
    port map (
            O => \N__19733\,
            I => \N__19728\
        );

    \I__3812\ : InMux
    port map (
            O => \N__19732\,
            I => \N__19725\
        );

    \I__3811\ : InMux
    port map (
            O => \N__19731\,
            I => \N__19722\
        );

    \I__3810\ : LocalMux
    port map (
            O => \N__19728\,
            I => \N__19719\
        );

    \I__3809\ : LocalMux
    port map (
            O => \N__19725\,
            I => \eeprom.n2906\
        );

    \I__3808\ : LocalMux
    port map (
            O => \N__19722\,
            I => \eeprom.n2906\
        );

    \I__3807\ : Odrv4
    port map (
            O => \N__19719\,
            I => \eeprom.n2906\
        );

    \I__3806\ : CascadeMux
    port map (
            O => \N__19712\,
            I => \N__19709\
        );

    \I__3805\ : InMux
    port map (
            O => \N__19709\,
            I => \N__19706\
        );

    \I__3804\ : LocalMux
    port map (
            O => \N__19706\,
            I => \eeprom.n2973\
        );

    \I__3803\ : InMux
    port map (
            O => \N__19703\,
            I => \N__19698\
        );

    \I__3802\ : InMux
    port map (
            O => \N__19702\,
            I => \N__19693\
        );

    \I__3801\ : InMux
    port map (
            O => \N__19701\,
            I => \N__19693\
        );

    \I__3800\ : LocalMux
    port map (
            O => \N__19698\,
            I => \N__19690\
        );

    \I__3799\ : LocalMux
    port map (
            O => \N__19693\,
            I => \eeprom.n2903\
        );

    \I__3798\ : Odrv4
    port map (
            O => \N__19690\,
            I => \eeprom.n2903\
        );

    \I__3797\ : InMux
    port map (
            O => \N__19685\,
            I => \N__19682\
        );

    \I__3796\ : LocalMux
    port map (
            O => \N__19682\,
            I => \eeprom.n2970\
        );

    \I__3795\ : InMux
    port map (
            O => \N__19679\,
            I => \N__19676\
        );

    \I__3794\ : LocalMux
    port map (
            O => \N__19676\,
            I => \N__19673\
        );

    \I__3793\ : Odrv4
    port map (
            O => \N__19673\,
            I => \eeprom.n2879\
        );

    \I__3792\ : InMux
    port map (
            O => \N__19670\,
            I => \N__19665\
        );

    \I__3791\ : InMux
    port map (
            O => \N__19669\,
            I => \N__19662\
        );

    \I__3790\ : InMux
    port map (
            O => \N__19668\,
            I => \N__19659\
        );

    \I__3789\ : LocalMux
    port map (
            O => \N__19665\,
            I => \N__19656\
        );

    \I__3788\ : LocalMux
    port map (
            O => \N__19662\,
            I => \N__19651\
        );

    \I__3787\ : LocalMux
    port map (
            O => \N__19659\,
            I => \N__19651\
        );

    \I__3786\ : Odrv12
    port map (
            O => \N__19656\,
            I => \eeprom.n2812\
        );

    \I__3785\ : Odrv4
    port map (
            O => \N__19651\,
            I => \eeprom.n2812\
        );

    \I__3784\ : InMux
    port map (
            O => \N__19646\,
            I => \N__19643\
        );

    \I__3783\ : LocalMux
    port map (
            O => \N__19643\,
            I => \N__19640\
        );

    \I__3782\ : Odrv4
    port map (
            O => \N__19640\,
            I => \eeprom.n2880\
        );

    \I__3781\ : CascadeMux
    port map (
            O => \N__19637\,
            I => \N__19634\
        );

    \I__3780\ : InMux
    port map (
            O => \N__19634\,
            I => \N__19630\
        );

    \I__3779\ : CascadeMux
    port map (
            O => \N__19633\,
            I => \N__19627\
        );

    \I__3778\ : LocalMux
    port map (
            O => \N__19630\,
            I => \N__19624\
        );

    \I__3777\ : InMux
    port map (
            O => \N__19627\,
            I => \N__19621\
        );

    \I__3776\ : Span4Mux_h
    port map (
            O => \N__19624\,
            I => \N__19616\
        );

    \I__3775\ : LocalMux
    port map (
            O => \N__19621\,
            I => \N__19616\
        );

    \I__3774\ : Span4Mux_h
    port map (
            O => \N__19616\,
            I => \N__19612\
        );

    \I__3773\ : InMux
    port map (
            O => \N__19615\,
            I => \N__19609\
        );

    \I__3772\ : Odrv4
    port map (
            O => \N__19612\,
            I => \eeprom.n2813\
        );

    \I__3771\ : LocalMux
    port map (
            O => \N__19609\,
            I => \eeprom.n2813\
        );

    \I__3770\ : InMux
    port map (
            O => \N__19604\,
            I => \N__19600\
        );

    \I__3769\ : InMux
    port map (
            O => \N__19603\,
            I => \N__19597\
        );

    \I__3768\ : LocalMux
    port map (
            O => \N__19600\,
            I => \N__19594\
        );

    \I__3767\ : LocalMux
    port map (
            O => \N__19597\,
            I => \eeprom.n2913\
        );

    \I__3766\ : Odrv4
    port map (
            O => \N__19594\,
            I => \eeprom.n2913\
        );

    \I__3765\ : CascadeMux
    port map (
            O => \N__19589\,
            I => \N__19586\
        );

    \I__3764\ : InMux
    port map (
            O => \N__19586\,
            I => \N__19583\
        );

    \I__3763\ : LocalMux
    port map (
            O => \N__19583\,
            I => \N__19580\
        );

    \I__3762\ : Odrv4
    port map (
            O => \N__19580\,
            I => \eeprom.n2980\
        );

    \I__3761\ : InMux
    port map (
            O => \N__19577\,
            I => \eeprom.n3637\
        );

    \I__3760\ : InMux
    port map (
            O => \N__19574\,
            I => \eeprom.n3638\
        );

    \I__3759\ : InMux
    port map (
            O => \N__19571\,
            I => \bfn_11_22_0_\
        );

    \I__3758\ : InMux
    port map (
            O => \N__19568\,
            I => \eeprom.n3640\
        );

    \I__3757\ : InMux
    port map (
            O => \N__19565\,
            I => \eeprom.n3641\
        );

    \I__3756\ : InMux
    port map (
            O => \N__19562\,
            I => \eeprom.n3642\
        );

    \I__3755\ : InMux
    port map (
            O => \N__19559\,
            I => \eeprom.n3643\
        );

    \I__3754\ : InMux
    port map (
            O => \N__19556\,
            I => \eeprom.n3644\
        );

    \I__3753\ : InMux
    port map (
            O => \N__19553\,
            I => \eeprom.n3645\
        );

    \I__3752\ : CascadeMux
    port map (
            O => \N__19550\,
            I => \N__19546\
        );

    \I__3751\ : InMux
    port map (
            O => \N__19549\,
            I => \N__19543\
        );

    \I__3750\ : InMux
    port map (
            O => \N__19546\,
            I => \N__19540\
        );

    \I__3749\ : LocalMux
    port map (
            O => \N__19543\,
            I => \N__19536\
        );

    \I__3748\ : LocalMux
    port map (
            O => \N__19540\,
            I => \N__19533\
        );

    \I__3747\ : InMux
    port map (
            O => \N__19539\,
            I => \N__19530\
        );

    \I__3746\ : Odrv4
    port map (
            O => \N__19536\,
            I => \eeprom.n3213\
        );

    \I__3745\ : Odrv4
    port map (
            O => \N__19533\,
            I => \eeprom.n3213\
        );

    \I__3744\ : LocalMux
    port map (
            O => \N__19530\,
            I => \eeprom.n3213\
        );

    \I__3743\ : CascadeMux
    port map (
            O => \N__19523\,
            I => \eeprom.n3116_cascade_\
        );

    \I__3742\ : InMux
    port map (
            O => \N__19520\,
            I => \N__19516\
        );

    \I__3741\ : CascadeMux
    port map (
            O => \N__19519\,
            I => \N__19513\
        );

    \I__3740\ : LocalMux
    port map (
            O => \N__19516\,
            I => \N__19509\
        );

    \I__3739\ : InMux
    port map (
            O => \N__19513\,
            I => \N__19506\
        );

    \I__3738\ : CascadeMux
    port map (
            O => \N__19512\,
            I => \N__19503\
        );

    \I__3737\ : Span4Mux_h
    port map (
            O => \N__19509\,
            I => \N__19500\
        );

    \I__3736\ : LocalMux
    port map (
            O => \N__19506\,
            I => \N__19497\
        );

    \I__3735\ : InMux
    port map (
            O => \N__19503\,
            I => \N__19494\
        );

    \I__3734\ : Odrv4
    port map (
            O => \N__19500\,
            I => \eeprom.n3215\
        );

    \I__3733\ : Odrv4
    port map (
            O => \N__19497\,
            I => \eeprom.n3215\
        );

    \I__3732\ : LocalMux
    port map (
            O => \N__19494\,
            I => \eeprom.n3215\
        );

    \I__3731\ : InMux
    port map (
            O => \N__19487\,
            I => \bfn_11_21_0_\
        );

    \I__3730\ : CascadeMux
    port map (
            O => \N__19484\,
            I => \N__19480\
        );

    \I__3729\ : InMux
    port map (
            O => \N__19483\,
            I => \N__19477\
        );

    \I__3728\ : InMux
    port map (
            O => \N__19480\,
            I => \N__19474\
        );

    \I__3727\ : LocalMux
    port map (
            O => \N__19477\,
            I => \N__19471\
        );

    \I__3726\ : LocalMux
    port map (
            O => \N__19474\,
            I => \eeprom.n2918\
        );

    \I__3725\ : Odrv4
    port map (
            O => \N__19471\,
            I => \eeprom.n2918\
        );

    \I__3724\ : InMux
    port map (
            O => \N__19466\,
            I => \N__19463\
        );

    \I__3723\ : LocalMux
    port map (
            O => \N__19463\,
            I => \eeprom.n2985\
        );

    \I__3722\ : InMux
    port map (
            O => \N__19460\,
            I => \eeprom.n3632\
        );

    \I__3721\ : InMux
    port map (
            O => \N__19457\,
            I => \eeprom.n3633\
        );

    \I__3720\ : InMux
    port map (
            O => \N__19454\,
            I => \eeprom.n3634\
        );

    \I__3719\ : InMux
    port map (
            O => \N__19451\,
            I => \eeprom.n3635\
        );

    \I__3718\ : InMux
    port map (
            O => \N__19448\,
            I => \eeprom.n3636\
        );

    \I__3717\ : CascadeMux
    port map (
            O => \N__19445\,
            I => \N__19442\
        );

    \I__3716\ : InMux
    port map (
            O => \N__19442\,
            I => \N__19439\
        );

    \I__3715\ : LocalMux
    port map (
            O => \N__19439\,
            I => \N__19435\
        );

    \I__3714\ : InMux
    port map (
            O => \N__19438\,
            I => \N__19432\
        );

    \I__3713\ : Span4Mux_v
    port map (
            O => \N__19435\,
            I => \N__19428\
        );

    \I__3712\ : LocalMux
    port map (
            O => \N__19432\,
            I => \N__19425\
        );

    \I__3711\ : InMux
    port map (
            O => \N__19431\,
            I => \N__19422\
        );

    \I__3710\ : Span4Mux_h
    port map (
            O => \N__19428\,
            I => \N__19419\
        );

    \I__3709\ : Sp12to4
    port map (
            O => \N__19425\,
            I => \N__19416\
        );

    \I__3708\ : LocalMux
    port map (
            O => \N__19422\,
            I => \N__19409\
        );

    \I__3707\ : Sp12to4
    port map (
            O => \N__19419\,
            I => \N__19409\
        );

    \I__3706\ : Span12Mux_v
    port map (
            O => \N__19416\,
            I => \N__19409\
        );

    \I__3705\ : Odrv12
    port map (
            O => \N__19409\,
            I => \eeprom.n3219\
        );

    \I__3704\ : CascadeMux
    port map (
            O => \N__19406\,
            I => \eeprom.n4615_cascade_\
        );

    \I__3703\ : CascadeMux
    port map (
            O => \N__19403\,
            I => \N__19400\
        );

    \I__3702\ : InMux
    port map (
            O => \N__19400\,
            I => \N__19396\
        );

    \I__3701\ : CascadeMux
    port map (
            O => \N__19399\,
            I => \N__19392\
        );

    \I__3700\ : LocalMux
    port map (
            O => \N__19396\,
            I => \N__19389\
        );

    \I__3699\ : InMux
    port map (
            O => \N__19395\,
            I => \N__19386\
        );

    \I__3698\ : InMux
    port map (
            O => \N__19392\,
            I => \N__19383\
        );

    \I__3697\ : Span4Mux_h
    port map (
            O => \N__19389\,
            I => \N__19378\
        );

    \I__3696\ : LocalMux
    port map (
            O => \N__19386\,
            I => \N__19378\
        );

    \I__3695\ : LocalMux
    port map (
            O => \N__19383\,
            I => \eeprom.n3218\
        );

    \I__3694\ : Odrv4
    port map (
            O => \N__19378\,
            I => \eeprom.n3218\
        );

    \I__3693\ : InMux
    port map (
            O => \N__19373\,
            I => \N__19370\
        );

    \I__3692\ : LocalMux
    port map (
            O => \N__19370\,
            I => \eeprom.n21_adj_477\
        );

    \I__3691\ : InMux
    port map (
            O => \N__19367\,
            I => \N__19364\
        );

    \I__3690\ : LocalMux
    port map (
            O => \N__19364\,
            I => \eeprom.n4611\
        );

    \I__3689\ : CascadeMux
    port map (
            O => \N__19361\,
            I => \N__19357\
        );

    \I__3688\ : CascadeMux
    port map (
            O => \N__19360\,
            I => \N__19354\
        );

    \I__3687\ : InMux
    port map (
            O => \N__19357\,
            I => \N__19350\
        );

    \I__3686\ : InMux
    port map (
            O => \N__19354\,
            I => \N__19347\
        );

    \I__3685\ : InMux
    port map (
            O => \N__19353\,
            I => \N__19344\
        );

    \I__3684\ : LocalMux
    port map (
            O => \N__19350\,
            I => \eeprom.n3300\
        );

    \I__3683\ : LocalMux
    port map (
            O => \N__19347\,
            I => \eeprom.n3300\
        );

    \I__3682\ : LocalMux
    port map (
            O => \N__19344\,
            I => \eeprom.n3300\
        );

    \I__3681\ : InMux
    port map (
            O => \N__19337\,
            I => \N__19333\
        );

    \I__3680\ : InMux
    port map (
            O => \N__19336\,
            I => \N__19330\
        );

    \I__3679\ : LocalMux
    port map (
            O => \N__19333\,
            I => \N__19327\
        );

    \I__3678\ : LocalMux
    port map (
            O => \N__19330\,
            I => \N__19324\
        );

    \I__3677\ : Span4Mux_v
    port map (
            O => \N__19327\,
            I => \N__19321\
        );

    \I__3676\ : Odrv4
    port map (
            O => \N__19324\,
            I => \eeprom.n3298\
        );

    \I__3675\ : Odrv4
    port map (
            O => \N__19321\,
            I => \eeprom.n3298\
        );

    \I__3674\ : InMux
    port map (
            O => \N__19316\,
            I => \N__19313\
        );

    \I__3673\ : LocalMux
    port map (
            O => \N__19313\,
            I => \eeprom.n25_adj_487\
        );

    \I__3672\ : CascadeMux
    port map (
            O => \N__19310\,
            I => \N__19305\
        );

    \I__3671\ : InMux
    port map (
            O => \N__19309\,
            I => \N__19302\
        );

    \I__3670\ : InMux
    port map (
            O => \N__19308\,
            I => \N__19297\
        );

    \I__3669\ : InMux
    port map (
            O => \N__19305\,
            I => \N__19297\
        );

    \I__3668\ : LocalMux
    port map (
            O => \N__19302\,
            I => \eeprom.n3301\
        );

    \I__3667\ : LocalMux
    port map (
            O => \N__19297\,
            I => \eeprom.n3301\
        );

    \I__3666\ : CascadeMux
    port map (
            O => \N__19292\,
            I => \N__19289\
        );

    \I__3665\ : InMux
    port map (
            O => \N__19289\,
            I => \N__19286\
        );

    \I__3664\ : LocalMux
    port map (
            O => \N__19286\,
            I => \N__19283\
        );

    \I__3663\ : Odrv4
    port map (
            O => \N__19283\,
            I => \eeprom.n3368\
        );

    \I__3662\ : InMux
    port map (
            O => \N__19280\,
            I => \N__19277\
        );

    \I__3661\ : LocalMux
    port map (
            O => \N__19277\,
            I => \N__19274\
        );

    \I__3660\ : Span4Mux_h
    port map (
            O => \N__19274\,
            I => \N__19271\
        );

    \I__3659\ : Odrv4
    port map (
            O => \N__19271\,
            I => \eeprom.n3284\
        );

    \I__3658\ : CascadeMux
    port map (
            O => \N__19268\,
            I => \N__19263\
        );

    \I__3657\ : InMux
    port map (
            O => \N__19267\,
            I => \N__19250\
        );

    \I__3656\ : InMux
    port map (
            O => \N__19266\,
            I => \N__19247\
        );

    \I__3655\ : InMux
    port map (
            O => \N__19263\,
            I => \N__19244\
        );

    \I__3654\ : CascadeMux
    port map (
            O => \N__19262\,
            I => \N__19241\
        );

    \I__3653\ : CascadeMux
    port map (
            O => \N__19261\,
            I => \N__19236\
        );

    \I__3652\ : CascadeMux
    port map (
            O => \N__19260\,
            I => \N__19233\
        );

    \I__3651\ : CascadeMux
    port map (
            O => \N__19259\,
            I => \N__19230\
        );

    \I__3650\ : CascadeMux
    port map (
            O => \N__19258\,
            I => \N__19227\
        );

    \I__3649\ : CascadeMux
    port map (
            O => \N__19257\,
            I => \N__19221\
        );

    \I__3648\ : CascadeMux
    port map (
            O => \N__19256\,
            I => \N__19218\
        );

    \I__3647\ : CascadeMux
    port map (
            O => \N__19255\,
            I => \N__19215\
        );

    \I__3646\ : CascadeMux
    port map (
            O => \N__19254\,
            I => \N__19212\
        );

    \I__3645\ : InMux
    port map (
            O => \N__19253\,
            I => \N__19208\
        );

    \I__3644\ : LocalMux
    port map (
            O => \N__19250\,
            I => \N__19201\
        );

    \I__3643\ : LocalMux
    port map (
            O => \N__19247\,
            I => \N__19201\
        );

    \I__3642\ : LocalMux
    port map (
            O => \N__19244\,
            I => \N__19201\
        );

    \I__3641\ : InMux
    port map (
            O => \N__19241\,
            I => \N__19194\
        );

    \I__3640\ : InMux
    port map (
            O => \N__19240\,
            I => \N__19194\
        );

    \I__3639\ : InMux
    port map (
            O => \N__19239\,
            I => \N__19194\
        );

    \I__3638\ : InMux
    port map (
            O => \N__19236\,
            I => \N__19188\
        );

    \I__3637\ : InMux
    port map (
            O => \N__19233\,
            I => \N__19188\
        );

    \I__3636\ : InMux
    port map (
            O => \N__19230\,
            I => \N__19179\
        );

    \I__3635\ : InMux
    port map (
            O => \N__19227\,
            I => \N__19179\
        );

    \I__3634\ : InMux
    port map (
            O => \N__19226\,
            I => \N__19179\
        );

    \I__3633\ : InMux
    port map (
            O => \N__19225\,
            I => \N__19179\
        );

    \I__3632\ : InMux
    port map (
            O => \N__19224\,
            I => \N__19168\
        );

    \I__3631\ : InMux
    port map (
            O => \N__19221\,
            I => \N__19168\
        );

    \I__3630\ : InMux
    port map (
            O => \N__19218\,
            I => \N__19168\
        );

    \I__3629\ : InMux
    port map (
            O => \N__19215\,
            I => \N__19168\
        );

    \I__3628\ : InMux
    port map (
            O => \N__19212\,
            I => \N__19168\
        );

    \I__3627\ : InMux
    port map (
            O => \N__19211\,
            I => \N__19165\
        );

    \I__3626\ : LocalMux
    port map (
            O => \N__19208\,
            I => \N__19162\
        );

    \I__3625\ : Span4Mux_v
    port map (
            O => \N__19201\,
            I => \N__19157\
        );

    \I__3624\ : LocalMux
    port map (
            O => \N__19194\,
            I => \N__19157\
        );

    \I__3623\ : InMux
    port map (
            O => \N__19193\,
            I => \N__19154\
        );

    \I__3622\ : LocalMux
    port map (
            O => \N__19188\,
            I => \eeprom.n3232\
        );

    \I__3621\ : LocalMux
    port map (
            O => \N__19179\,
            I => \eeprom.n3232\
        );

    \I__3620\ : LocalMux
    port map (
            O => \N__19168\,
            I => \eeprom.n3232\
        );

    \I__3619\ : LocalMux
    port map (
            O => \N__19165\,
            I => \eeprom.n3232\
        );

    \I__3618\ : Odrv4
    port map (
            O => \N__19162\,
            I => \eeprom.n3232\
        );

    \I__3617\ : Odrv4
    port map (
            O => \N__19157\,
            I => \eeprom.n3232\
        );

    \I__3616\ : LocalMux
    port map (
            O => \N__19154\,
            I => \eeprom.n3232\
        );

    \I__3615\ : InMux
    port map (
            O => \N__19139\,
            I => \N__19136\
        );

    \I__3614\ : LocalMux
    port map (
            O => \N__19136\,
            I => \N__19132\
        );

    \I__3613\ : InMux
    port map (
            O => \N__19135\,
            I => \N__19128\
        );

    \I__3612\ : Span4Mux_h
    port map (
            O => \N__19132\,
            I => \N__19125\
        );

    \I__3611\ : InMux
    port map (
            O => \N__19131\,
            I => \N__19122\
        );

    \I__3610\ : LocalMux
    port map (
            O => \N__19128\,
            I => \eeprom.n3210\
        );

    \I__3609\ : Odrv4
    port map (
            O => \N__19125\,
            I => \eeprom.n3210\
        );

    \I__3608\ : LocalMux
    port map (
            O => \N__19122\,
            I => \eeprom.n3210\
        );

    \I__3607\ : CascadeMux
    port map (
            O => \N__19115\,
            I => \eeprom.n3113_cascade_\
        );

    \I__3606\ : InMux
    port map (
            O => \N__19112\,
            I => \N__19107\
        );

    \I__3605\ : InMux
    port map (
            O => \N__19111\,
            I => \N__19102\
        );

    \I__3604\ : InMux
    port map (
            O => \N__19110\,
            I => \N__19102\
        );

    \I__3603\ : LocalMux
    port map (
            O => \N__19107\,
            I => \N__19099\
        );

    \I__3602\ : LocalMux
    port map (
            O => \N__19102\,
            I => \eeprom.n3212\
        );

    \I__3601\ : Odrv4
    port map (
            O => \N__19099\,
            I => \eeprom.n3212\
        );

    \I__3600\ : InMux
    port map (
            O => \N__19094\,
            I => \N__19091\
        );

    \I__3599\ : LocalMux
    port map (
            O => \N__19091\,
            I => \N__19086\
        );

    \I__3598\ : InMux
    port map (
            O => \N__19090\,
            I => \N__19083\
        );

    \I__3597\ : InMux
    port map (
            O => \N__19089\,
            I => \N__19080\
        );

    \I__3596\ : Odrv4
    port map (
            O => \N__19086\,
            I => \eeprom.n3208\
        );

    \I__3595\ : LocalMux
    port map (
            O => \N__19083\,
            I => \eeprom.n3208\
        );

    \I__3594\ : LocalMux
    port map (
            O => \N__19080\,
            I => \eeprom.n3208\
        );

    \I__3593\ : CascadeMux
    port map (
            O => \N__19073\,
            I => \N__19070\
        );

    \I__3592\ : InMux
    port map (
            O => \N__19070\,
            I => \N__19067\
        );

    \I__3591\ : LocalMux
    port map (
            O => \N__19067\,
            I => \eeprom.n25_adj_478\
        );

    \I__3590\ : CascadeMux
    port map (
            O => \N__19064\,
            I => \N__19059\
        );

    \I__3589\ : InMux
    port map (
            O => \N__19063\,
            I => \N__19056\
        );

    \I__3588\ : InMux
    port map (
            O => \N__19062\,
            I => \N__19053\
        );

    \I__3587\ : InMux
    port map (
            O => \N__19059\,
            I => \N__19050\
        );

    \I__3586\ : LocalMux
    port map (
            O => \N__19056\,
            I => \eeprom.n3317\
        );

    \I__3585\ : LocalMux
    port map (
            O => \N__19053\,
            I => \eeprom.n3317\
        );

    \I__3584\ : LocalMux
    port map (
            O => \N__19050\,
            I => \eeprom.n3317\
        );

    \I__3583\ : CascadeMux
    port map (
            O => \N__19043\,
            I => \N__19040\
        );

    \I__3582\ : InMux
    port map (
            O => \N__19040\,
            I => \N__19037\
        );

    \I__3581\ : LocalMux
    port map (
            O => \N__19037\,
            I => \N__19034\
        );

    \I__3580\ : Odrv4
    port map (
            O => \N__19034\,
            I => \eeprom.n3384\
        );

    \I__3579\ : InMux
    port map (
            O => \N__19031\,
            I => \N__19028\
        );

    \I__3578\ : LocalMux
    port map (
            O => \N__19028\,
            I => \N__19025\
        );

    \I__3577\ : Odrv4
    port map (
            O => \N__19025\,
            I => \eeprom.n3375\
        );

    \I__3576\ : InMux
    port map (
            O => \N__19022\,
            I => \N__19018\
        );

    \I__3575\ : CascadeMux
    port map (
            O => \N__19021\,
            I => \N__19014\
        );

    \I__3574\ : LocalMux
    port map (
            O => \N__19018\,
            I => \N__19011\
        );

    \I__3573\ : InMux
    port map (
            O => \N__19017\,
            I => \N__19008\
        );

    \I__3572\ : InMux
    port map (
            O => \N__19014\,
            I => \N__19005\
        );

    \I__3571\ : Odrv4
    port map (
            O => \N__19011\,
            I => \eeprom.n3308\
        );

    \I__3570\ : LocalMux
    port map (
            O => \N__19008\,
            I => \eeprom.n3308\
        );

    \I__3569\ : LocalMux
    port map (
            O => \N__19005\,
            I => \eeprom.n3308\
        );

    \I__3568\ : CascadeMux
    port map (
            O => \N__18998\,
            I => \eeprom.n3407_cascade_\
        );

    \I__3567\ : InMux
    port map (
            O => \N__18995\,
            I => \N__18992\
        );

    \I__3566\ : LocalMux
    port map (
            O => \N__18992\,
            I => \eeprom.n28_adj_484\
        );

    \I__3565\ : CascadeMux
    port map (
            O => \N__18989\,
            I => \eeprom.n27_adj_486_cascade_\
        );

    \I__3564\ : InMux
    port map (
            O => \N__18986\,
            I => \N__18983\
        );

    \I__3563\ : LocalMux
    port map (
            O => \N__18983\,
            I => \eeprom.n26_adj_485\
        );

    \I__3562\ : CascadeMux
    port map (
            O => \N__18980\,
            I => \N__18976\
        );

    \I__3561\ : CascadeMux
    port map (
            O => \N__18979\,
            I => \N__18972\
        );

    \I__3560\ : InMux
    port map (
            O => \N__18976\,
            I => \N__18969\
        );

    \I__3559\ : InMux
    port map (
            O => \N__18975\,
            I => \N__18964\
        );

    \I__3558\ : InMux
    port map (
            O => \N__18972\,
            I => \N__18964\
        );

    \I__3557\ : LocalMux
    port map (
            O => \N__18969\,
            I => \eeprom.n3306\
        );

    \I__3556\ : LocalMux
    port map (
            O => \N__18964\,
            I => \eeprom.n3306\
        );

    \I__3555\ : CascadeMux
    port map (
            O => \N__18959\,
            I => \eeprom.n3331_cascade_\
        );

    \I__3554\ : InMux
    port map (
            O => \N__18956\,
            I => \N__18953\
        );

    \I__3553\ : LocalMux
    port map (
            O => \N__18953\,
            I => \N__18950\
        );

    \I__3552\ : Odrv4
    port map (
            O => \N__18950\,
            I => \eeprom.n3373\
        );

    \I__3551\ : CascadeMux
    port map (
            O => \N__18947\,
            I => \N__18942\
        );

    \I__3550\ : InMux
    port map (
            O => \N__18946\,
            I => \N__18937\
        );

    \I__3549\ : InMux
    port map (
            O => \N__18945\,
            I => \N__18937\
        );

    \I__3548\ : InMux
    port map (
            O => \N__18942\,
            I => \N__18934\
        );

    \I__3547\ : LocalMux
    port map (
            O => \N__18937\,
            I => \eeprom.n3305\
        );

    \I__3546\ : LocalMux
    port map (
            O => \N__18934\,
            I => \eeprom.n3305\
        );

    \I__3545\ : InMux
    port map (
            O => \N__18929\,
            I => \N__18926\
        );

    \I__3544\ : LocalMux
    port map (
            O => \N__18926\,
            I => \N__18923\
        );

    \I__3543\ : Odrv4
    port map (
            O => \N__18923\,
            I => \eeprom.n3372\
        );

    \I__3542\ : InMux
    port map (
            O => \N__18920\,
            I => \N__18917\
        );

    \I__3541\ : LocalMux
    port map (
            O => \N__18917\,
            I => \N__18914\
        );

    \I__3540\ : Odrv4
    port map (
            O => \N__18914\,
            I => \eeprom.n3376\
        );

    \I__3539\ : CascadeMux
    port map (
            O => \N__18911\,
            I => \N__18907\
        );

    \I__3538\ : CascadeMux
    port map (
            O => \N__18910\,
            I => \N__18903\
        );

    \I__3537\ : InMux
    port map (
            O => \N__18907\,
            I => \N__18900\
        );

    \I__3536\ : InMux
    port map (
            O => \N__18906\,
            I => \N__18897\
        );

    \I__3535\ : InMux
    port map (
            O => \N__18903\,
            I => \N__18894\
        );

    \I__3534\ : LocalMux
    port map (
            O => \N__18900\,
            I => \eeprom.n3309\
        );

    \I__3533\ : LocalMux
    port map (
            O => \N__18897\,
            I => \eeprom.n3309\
        );

    \I__3532\ : LocalMux
    port map (
            O => \N__18894\,
            I => \eeprom.n3309\
        );

    \I__3531\ : InMux
    port map (
            O => \N__18887\,
            I => \N__18884\
        );

    \I__3530\ : LocalMux
    port map (
            O => \N__18884\,
            I => \eeprom.n4703\
        );

    \I__3529\ : CascadeMux
    port map (
            O => \N__18881\,
            I => \eeprom.n2917_cascade_\
        );

    \I__3528\ : CascadeMux
    port map (
            O => \N__18878\,
            I => \eeprom.n4707_cascade_\
        );

    \I__3527\ : InMux
    port map (
            O => \N__18875\,
            I => \N__18872\
        );

    \I__3526\ : LocalMux
    port map (
            O => \N__18872\,
            I => \eeprom.n15_adj_419\
        );

    \I__3525\ : InMux
    port map (
            O => \N__18869\,
            I => \N__18866\
        );

    \I__3524\ : LocalMux
    port map (
            O => \N__18866\,
            I => \eeprom.n2875\
        );

    \I__3523\ : InMux
    port map (
            O => \N__18863\,
            I => \N__18859\
        );

    \I__3522\ : InMux
    port map (
            O => \N__18862\,
            I => \N__18856\
        );

    \I__3521\ : LocalMux
    port map (
            O => \N__18859\,
            I => \N__18852\
        );

    \I__3520\ : LocalMux
    port map (
            O => \N__18856\,
            I => \N__18849\
        );

    \I__3519\ : InMux
    port map (
            O => \N__18855\,
            I => \N__18846\
        );

    \I__3518\ : Odrv4
    port map (
            O => \N__18852\,
            I => \eeprom.n2808\
        );

    \I__3517\ : Odrv4
    port map (
            O => \N__18849\,
            I => \eeprom.n2808\
        );

    \I__3516\ : LocalMux
    port map (
            O => \N__18846\,
            I => \eeprom.n2808\
        );

    \I__3515\ : CascadeMux
    port map (
            O => \N__18839\,
            I => \N__18836\
        );

    \I__3514\ : InMux
    port map (
            O => \N__18836\,
            I => \N__18833\
        );

    \I__3513\ : LocalMux
    port map (
            O => \N__18833\,
            I => \N__18830\
        );

    \I__3512\ : Odrv4
    port map (
            O => \N__18830\,
            I => \eeprom.n3385\
        );

    \I__3511\ : CascadeMux
    port map (
            O => \N__18827\,
            I => \N__18824\
        );

    \I__3510\ : InMux
    port map (
            O => \N__18824\,
            I => \N__18821\
        );

    \I__3509\ : LocalMux
    port map (
            O => \N__18821\,
            I => \N__18818\
        );

    \I__3508\ : Span4Mux_h
    port map (
            O => \N__18818\,
            I => \N__18815\
        );

    \I__3507\ : Odrv4
    port map (
            O => \N__18815\,
            I => \eeprom.n3283\
        );

    \I__3506\ : CascadeMux
    port map (
            O => \N__18812\,
            I => \eeprom.n3315_cascade_\
        );

    \I__3505\ : CascadeMux
    port map (
            O => \N__18809\,
            I => \N__18806\
        );

    \I__3504\ : InMux
    port map (
            O => \N__18806\,
            I => \N__18801\
        );

    \I__3503\ : InMux
    port map (
            O => \N__18805\,
            I => \N__18796\
        );

    \I__3502\ : InMux
    port map (
            O => \N__18804\,
            I => \N__18796\
        );

    \I__3501\ : LocalMux
    port map (
            O => \N__18801\,
            I => \eeprom.n3318\
        );

    \I__3500\ : LocalMux
    port map (
            O => \N__18796\,
            I => \eeprom.n3318\
        );

    \I__3499\ : CascadeMux
    port map (
            O => \N__18791\,
            I => \eeprom.n4719_cascade_\
        );

    \I__3498\ : InMux
    port map (
            O => \N__18788\,
            I => \N__18785\
        );

    \I__3497\ : LocalMux
    port map (
            O => \N__18785\,
            I => \eeprom.n4721\
        );

    \I__3496\ : CascadeMux
    port map (
            O => \N__18782\,
            I => \N__18778\
        );

    \I__3495\ : InMux
    port map (
            O => \N__18781\,
            I => \N__18774\
        );

    \I__3494\ : InMux
    port map (
            O => \N__18778\,
            I => \N__18771\
        );

    \I__3493\ : InMux
    port map (
            O => \N__18777\,
            I => \N__18768\
        );

    \I__3492\ : LocalMux
    port map (
            O => \N__18774\,
            I => \eeprom.n3304\
        );

    \I__3491\ : LocalMux
    port map (
            O => \N__18771\,
            I => \eeprom.n3304\
        );

    \I__3490\ : LocalMux
    port map (
            O => \N__18768\,
            I => \eeprom.n3304\
        );

    \I__3489\ : CascadeMux
    port map (
            O => \N__18761\,
            I => \eeprom.n4151_cascade_\
        );

    \I__3488\ : InMux
    port map (
            O => \N__18758\,
            I => \N__18753\
        );

    \I__3487\ : InMux
    port map (
            O => \N__18757\,
            I => \N__18750\
        );

    \I__3486\ : InMux
    port map (
            O => \N__18756\,
            I => \N__18747\
        );

    \I__3485\ : LocalMux
    port map (
            O => \N__18753\,
            I => \N__18744\
        );

    \I__3484\ : LocalMux
    port map (
            O => \N__18750\,
            I => \N__18739\
        );

    \I__3483\ : LocalMux
    port map (
            O => \N__18747\,
            I => \N__18739\
        );

    \I__3482\ : Span4Mux_v
    port map (
            O => \N__18744\,
            I => \N__18736\
        );

    \I__3481\ : Odrv4
    port map (
            O => \N__18739\,
            I => \eeprom.n3302\
        );

    \I__3480\ : Odrv4
    port map (
            O => \N__18736\,
            I => \eeprom.n3302\
        );

    \I__3479\ : InMux
    port map (
            O => \N__18731\,
            I => \N__18728\
        );

    \I__3478\ : LocalMux
    port map (
            O => \N__18728\,
            I => \N__18725\
        );

    \I__3477\ : Span4Mux_h
    port map (
            O => \N__18725\,
            I => \N__18722\
        );

    \I__3476\ : Odrv4
    port map (
            O => \N__18722\,
            I => \eeprom.n4529\
        );

    \I__3475\ : CascadeMux
    port map (
            O => \N__18719\,
            I => \N__18714\
        );

    \I__3474\ : InMux
    port map (
            O => \N__18718\,
            I => \N__18709\
        );

    \I__3473\ : InMux
    port map (
            O => \N__18717\,
            I => \N__18709\
        );

    \I__3472\ : InMux
    port map (
            O => \N__18714\,
            I => \N__18706\
        );

    \I__3471\ : LocalMux
    port map (
            O => \N__18709\,
            I => \N__18701\
        );

    \I__3470\ : LocalMux
    port map (
            O => \N__18706\,
            I => \N__18701\
        );

    \I__3469\ : Odrv4
    port map (
            O => \N__18701\,
            I => \eeprom.n2814\
        );

    \I__3468\ : InMux
    port map (
            O => \N__18698\,
            I => \N__18695\
        );

    \I__3467\ : LocalMux
    port map (
            O => \N__18695\,
            I => \N__18690\
        );

    \I__3466\ : InMux
    port map (
            O => \N__18694\,
            I => \N__18687\
        );

    \I__3465\ : InMux
    port map (
            O => \N__18693\,
            I => \N__18684\
        );

    \I__3464\ : Span4Mux_v
    port map (
            O => \N__18690\,
            I => \N__18677\
        );

    \I__3463\ : LocalMux
    port map (
            O => \N__18687\,
            I => \N__18677\
        );

    \I__3462\ : LocalMux
    port map (
            O => \N__18684\,
            I => \N__18677\
        );

    \I__3461\ : Span4Mux_h
    port map (
            O => \N__18677\,
            I => \N__18674\
        );

    \I__3460\ : Span4Mux_h
    port map (
            O => \N__18674\,
            I => \N__18671\
        );

    \I__3459\ : Odrv4
    port map (
            O => \N__18671\,
            I => \eeprom.n2819\
        );

    \I__3458\ : CascadeMux
    port map (
            O => \N__18668\,
            I => \eeprom.n4533_cascade_\
        );

    \I__3457\ : InMux
    port map (
            O => \N__18665\,
            I => \N__18662\
        );

    \I__3456\ : LocalMux
    port map (
            O => \N__18662\,
            I => \eeprom.n20\
        );

    \I__3455\ : CascadeMux
    port map (
            O => \N__18659\,
            I => \eeprom.n15_cascade_\
        );

    \I__3454\ : InMux
    port map (
            O => \N__18656\,
            I => \N__18649\
        );

    \I__3453\ : InMux
    port map (
            O => \N__18655\,
            I => \N__18649\
        );

    \I__3452\ : CascadeMux
    port map (
            O => \N__18654\,
            I => \N__18646\
        );

    \I__3451\ : LocalMux
    port map (
            O => \N__18649\,
            I => \N__18643\
        );

    \I__3450\ : InMux
    port map (
            O => \N__18646\,
            I => \N__18640\
        );

    \I__3449\ : Span4Mux_h
    port map (
            O => \N__18643\,
            I => \N__18635\
        );

    \I__3448\ : LocalMux
    port map (
            O => \N__18640\,
            I => \N__18635\
        );

    \I__3447\ : Odrv4
    port map (
            O => \N__18635\,
            I => \eeprom.n2816\
        );

    \I__3446\ : CascadeMux
    port map (
            O => \N__18632\,
            I => \eeprom.n2836_cascade_\
        );

    \I__3445\ : InMux
    port map (
            O => \N__18629\,
            I => \N__18626\
        );

    \I__3444\ : LocalMux
    port map (
            O => \N__18626\,
            I => \eeprom.n2883\
        );

    \I__3443\ : InMux
    port map (
            O => \N__18623\,
            I => \N__18616\
        );

    \I__3442\ : InMux
    port map (
            O => \N__18622\,
            I => \N__18616\
        );

    \I__3441\ : InMux
    port map (
            O => \N__18621\,
            I => \N__18613\
        );

    \I__3440\ : LocalMux
    port map (
            O => \N__18616\,
            I => \N__18610\
        );

    \I__3439\ : LocalMux
    port map (
            O => \N__18613\,
            I => \N__18607\
        );

    \I__3438\ : Span4Mux_h
    port map (
            O => \N__18610\,
            I => \N__18604\
        );

    \I__3437\ : Span4Mux_h
    port map (
            O => \N__18607\,
            I => \N__18601\
        );

    \I__3436\ : Odrv4
    port map (
            O => \N__18604\,
            I => \eeprom.n2809\
        );

    \I__3435\ : Odrv4
    port map (
            O => \N__18601\,
            I => \eeprom.n2809\
        );

    \I__3434\ : CascadeMux
    port map (
            O => \N__18596\,
            I => \N__18593\
        );

    \I__3433\ : InMux
    port map (
            O => \N__18593\,
            I => \N__18590\
        );

    \I__3432\ : LocalMux
    port map (
            O => \N__18590\,
            I => \eeprom.n2876\
        );

    \I__3431\ : InMux
    port map (
            O => \N__18587\,
            I => \N__18583\
        );

    \I__3430\ : InMux
    port map (
            O => \N__18586\,
            I => \N__18580\
        );

    \I__3429\ : LocalMux
    port map (
            O => \N__18583\,
            I => \N__18577\
        );

    \I__3428\ : LocalMux
    port map (
            O => \N__18580\,
            I => \eeprom.n2804\
        );

    \I__3427\ : Odrv4
    port map (
            O => \N__18577\,
            I => \eeprom.n2804\
        );

    \I__3426\ : InMux
    port map (
            O => \N__18572\,
            I => \N__18569\
        );

    \I__3425\ : LocalMux
    port map (
            O => \N__18569\,
            I => \eeprom.n2871\
        );

    \I__3424\ : InMux
    port map (
            O => \N__18566\,
            I => \N__18563\
        );

    \I__3423\ : LocalMux
    port map (
            O => \N__18563\,
            I => \eeprom.n19\
        );

    \I__3422\ : CascadeMux
    port map (
            O => \N__18560\,
            I => \eeprom.n22_cascade_\
        );

    \I__3421\ : InMux
    port map (
            O => \N__18557\,
            I => \N__18554\
        );

    \I__3420\ : LocalMux
    port map (
            O => \N__18554\,
            I => \eeprom.n2885\
        );

    \I__3419\ : CascadeMux
    port map (
            O => \N__18551\,
            I => \N__18547\
        );

    \I__3418\ : CascadeMux
    port map (
            O => \N__18550\,
            I => \N__18543\
        );

    \I__3417\ : InMux
    port map (
            O => \N__18547\,
            I => \N__18540\
        );

    \I__3416\ : InMux
    port map (
            O => \N__18546\,
            I => \N__18537\
        );

    \I__3415\ : InMux
    port map (
            O => \N__18543\,
            I => \N__18534\
        );

    \I__3414\ : LocalMux
    port map (
            O => \N__18540\,
            I => \N__18527\
        );

    \I__3413\ : LocalMux
    port map (
            O => \N__18537\,
            I => \N__18527\
        );

    \I__3412\ : LocalMux
    port map (
            O => \N__18534\,
            I => \N__18527\
        );

    \I__3411\ : Span4Mux_v
    port map (
            O => \N__18527\,
            I => \N__18524\
        );

    \I__3410\ : Odrv4
    port map (
            O => \N__18524\,
            I => \eeprom.n2818\
        );

    \I__3409\ : InMux
    port map (
            O => \N__18521\,
            I => \N__18518\
        );

    \I__3408\ : LocalMux
    port map (
            O => \N__18518\,
            I => \eeprom.n3270\
        );

    \I__3407\ : InMux
    port map (
            O => \N__18515\,
            I => \N__18512\
        );

    \I__3406\ : LocalMux
    port map (
            O => \N__18512\,
            I => \N__18508\
        );

    \I__3405\ : CascadeMux
    port map (
            O => \N__18511\,
            I => \N__18505\
        );

    \I__3404\ : Span4Mux_h
    port map (
            O => \N__18508\,
            I => \N__18501\
        );

    \I__3403\ : InMux
    port map (
            O => \N__18505\,
            I => \N__18498\
        );

    \I__3402\ : InMux
    port map (
            O => \N__18504\,
            I => \N__18495\
        );

    \I__3401\ : Sp12to4
    port map (
            O => \N__18501\,
            I => \N__18490\
        );

    \I__3400\ : LocalMux
    port map (
            O => \N__18498\,
            I => \N__18490\
        );

    \I__3399\ : LocalMux
    port map (
            O => \N__18495\,
            I => \eeprom.n2712\
        );

    \I__3398\ : Odrv12
    port map (
            O => \N__18490\,
            I => \eeprom.n2712\
        );

    \I__3397\ : InMux
    port map (
            O => \N__18485\,
            I => \N__18482\
        );

    \I__3396\ : LocalMux
    port map (
            O => \N__18482\,
            I => \N__18479\
        );

    \I__3395\ : Span4Mux_h
    port map (
            O => \N__18479\,
            I => \N__18476\
        );

    \I__3394\ : Odrv4
    port map (
            O => \N__18476\,
            I => \eeprom.n2779\
        );

    \I__3393\ : InMux
    port map (
            O => \N__18473\,
            I => \N__18469\
        );

    \I__3392\ : CascadeMux
    port map (
            O => \N__18472\,
            I => \N__18466\
        );

    \I__3391\ : LocalMux
    port map (
            O => \N__18469\,
            I => \N__18463\
        );

    \I__3390\ : InMux
    port map (
            O => \N__18466\,
            I => \N__18460\
        );

    \I__3389\ : Span4Mux_h
    port map (
            O => \N__18463\,
            I => \N__18454\
        );

    \I__3388\ : LocalMux
    port map (
            O => \N__18460\,
            I => \N__18454\
        );

    \I__3387\ : InMux
    port map (
            O => \N__18459\,
            I => \N__18451\
        );

    \I__3386\ : Odrv4
    port map (
            O => \N__18454\,
            I => \eeprom.n2707\
        );

    \I__3385\ : LocalMux
    port map (
            O => \N__18451\,
            I => \eeprom.n2707\
        );

    \I__3384\ : CascadeMux
    port map (
            O => \N__18446\,
            I => \N__18443\
        );

    \I__3383\ : InMux
    port map (
            O => \N__18443\,
            I => \N__18440\
        );

    \I__3382\ : LocalMux
    port map (
            O => \N__18440\,
            I => \N__18437\
        );

    \I__3381\ : Odrv4
    port map (
            O => \N__18437\,
            I => \eeprom.n2774\
        );

    \I__3380\ : InMux
    port map (
            O => \N__18434\,
            I => \N__18430\
        );

    \I__3379\ : CascadeMux
    port map (
            O => \N__18433\,
            I => \N__18427\
        );

    \I__3378\ : LocalMux
    port map (
            O => \N__18430\,
            I => \N__18424\
        );

    \I__3377\ : InMux
    port map (
            O => \N__18427\,
            I => \N__18421\
        );

    \I__3376\ : Span4Mux_h
    port map (
            O => \N__18424\,
            I => \N__18416\
        );

    \I__3375\ : LocalMux
    port map (
            O => \N__18421\,
            I => \N__18416\
        );

    \I__3374\ : Odrv4
    port map (
            O => \N__18416\,
            I => \eeprom.n2806\
        );

    \I__3373\ : CascadeMux
    port map (
            O => \N__18413\,
            I => \eeprom.n2806_cascade_\
        );

    \I__3372\ : InMux
    port map (
            O => \N__18410\,
            I => \N__18406\
        );

    \I__3371\ : InMux
    port map (
            O => \N__18409\,
            I => \N__18403\
        );

    \I__3370\ : LocalMux
    port map (
            O => \N__18406\,
            I => \N__18397\
        );

    \I__3369\ : LocalMux
    port map (
            O => \N__18403\,
            I => \N__18397\
        );

    \I__3368\ : InMux
    port map (
            O => \N__18402\,
            I => \N__18394\
        );

    \I__3367\ : Odrv4
    port map (
            O => \N__18397\,
            I => \eeprom.n2805\
        );

    \I__3366\ : LocalMux
    port map (
            O => \N__18394\,
            I => \eeprom.n2805\
        );

    \I__3365\ : InMux
    port map (
            O => \N__18389\,
            I => \N__18386\
        );

    \I__3364\ : LocalMux
    port map (
            O => \N__18386\,
            I => \eeprom.n18_adj_418\
        );

    \I__3363\ : InMux
    port map (
            O => \N__18383\,
            I => \N__18379\
        );

    \I__3362\ : CascadeMux
    port map (
            O => \N__18382\,
            I => \N__18376\
        );

    \I__3361\ : LocalMux
    port map (
            O => \N__18379\,
            I => \N__18373\
        );

    \I__3360\ : InMux
    port map (
            O => \N__18376\,
            I => \N__18370\
        );

    \I__3359\ : Span4Mux_v
    port map (
            O => \N__18373\,
            I => \N__18366\
        );

    \I__3358\ : LocalMux
    port map (
            O => \N__18370\,
            I => \N__18363\
        );

    \I__3357\ : InMux
    port map (
            O => \N__18369\,
            I => \N__18360\
        );

    \I__3356\ : Odrv4
    port map (
            O => \N__18366\,
            I => \eeprom.n2708\
        );

    \I__3355\ : Odrv4
    port map (
            O => \N__18363\,
            I => \eeprom.n2708\
        );

    \I__3354\ : LocalMux
    port map (
            O => \N__18360\,
            I => \eeprom.n2708\
        );

    \I__3353\ : CascadeMux
    port map (
            O => \N__18353\,
            I => \N__18350\
        );

    \I__3352\ : InMux
    port map (
            O => \N__18350\,
            I => \N__18347\
        );

    \I__3351\ : LocalMux
    port map (
            O => \N__18347\,
            I => \N__18344\
        );

    \I__3350\ : Odrv4
    port map (
            O => \N__18344\,
            I => \eeprom.n2775\
        );

    \I__3349\ : CascadeMux
    port map (
            O => \N__18341\,
            I => \N__18333\
        );

    \I__3348\ : CascadeMux
    port map (
            O => \N__18340\,
            I => \N__18328\
        );

    \I__3347\ : CascadeMux
    port map (
            O => \N__18339\,
            I => \N__18323\
        );

    \I__3346\ : CascadeMux
    port map (
            O => \N__18338\,
            I => \N__18320\
        );

    \I__3345\ : CascadeMux
    port map (
            O => \N__18337\,
            I => \N__18316\
        );

    \I__3344\ : InMux
    port map (
            O => \N__18336\,
            I => \N__18304\
        );

    \I__3343\ : InMux
    port map (
            O => \N__18333\,
            I => \N__18304\
        );

    \I__3342\ : InMux
    port map (
            O => \N__18332\,
            I => \N__18304\
        );

    \I__3341\ : InMux
    port map (
            O => \N__18331\,
            I => \N__18304\
        );

    \I__3340\ : InMux
    port map (
            O => \N__18328\,
            I => \N__18299\
        );

    \I__3339\ : InMux
    port map (
            O => \N__18327\,
            I => \N__18299\
        );

    \I__3338\ : InMux
    port map (
            O => \N__18326\,
            I => \N__18296\
        );

    \I__3337\ : InMux
    port map (
            O => \N__18323\,
            I => \N__18285\
        );

    \I__3336\ : InMux
    port map (
            O => \N__18320\,
            I => \N__18285\
        );

    \I__3335\ : InMux
    port map (
            O => \N__18319\,
            I => \N__18285\
        );

    \I__3334\ : InMux
    port map (
            O => \N__18316\,
            I => \N__18285\
        );

    \I__3333\ : InMux
    port map (
            O => \N__18315\,
            I => \N__18285\
        );

    \I__3332\ : CascadeMux
    port map (
            O => \N__18314\,
            I => \N__18282\
        );

    \I__3331\ : CascadeMux
    port map (
            O => \N__18313\,
            I => \N__18279\
        );

    \I__3330\ : LocalMux
    port map (
            O => \N__18304\,
            I => \N__18273\
        );

    \I__3329\ : LocalMux
    port map (
            O => \N__18299\,
            I => \N__18273\
        );

    \I__3328\ : LocalMux
    port map (
            O => \N__18296\,
            I => \N__18268\
        );

    \I__3327\ : LocalMux
    port map (
            O => \N__18285\,
            I => \N__18268\
        );

    \I__3326\ : InMux
    port map (
            O => \N__18282\,
            I => \N__18261\
        );

    \I__3325\ : InMux
    port map (
            O => \N__18279\,
            I => \N__18261\
        );

    \I__3324\ : InMux
    port map (
            O => \N__18278\,
            I => \N__18261\
        );

    \I__3323\ : Span4Mux_h
    port map (
            O => \N__18273\,
            I => \N__18258\
        );

    \I__3322\ : Odrv4
    port map (
            O => \N__18268\,
            I => \eeprom.n2737\
        );

    \I__3321\ : LocalMux
    port map (
            O => \N__18261\,
            I => \eeprom.n2737\
        );

    \I__3320\ : Odrv4
    port map (
            O => \N__18258\,
            I => \eeprom.n2737\
        );

    \I__3319\ : InMux
    port map (
            O => \N__18251\,
            I => \N__18248\
        );

    \I__3318\ : LocalMux
    port map (
            O => \N__18248\,
            I => \N__18244\
        );

    \I__3317\ : InMux
    port map (
            O => \N__18247\,
            I => \N__18241\
        );

    \I__3316\ : Odrv4
    port map (
            O => \N__18244\,
            I => \eeprom.n2807\
        );

    \I__3315\ : LocalMux
    port map (
            O => \N__18241\,
            I => \eeprom.n2807\
        );

    \I__3314\ : InMux
    port map (
            O => \N__18236\,
            I => \N__18233\
        );

    \I__3313\ : LocalMux
    port map (
            O => \N__18233\,
            I => \N__18230\
        );

    \I__3312\ : Odrv4
    port map (
            O => \N__18230\,
            I => \eeprom.n2874\
        );

    \I__3311\ : CascadeMux
    port map (
            O => \N__18227\,
            I => \eeprom.n2807_cascade_\
        );

    \I__3310\ : CascadeMux
    port map (
            O => \N__18224\,
            I => \N__18221\
        );

    \I__3309\ : InMux
    port map (
            O => \N__18221\,
            I => \N__18218\
        );

    \I__3308\ : LocalMux
    port map (
            O => \N__18218\,
            I => \eeprom.n2881\
        );

    \I__3307\ : CascadeMux
    port map (
            O => \N__18215\,
            I => \eeprom.n2913_cascade_\
        );

    \I__3306\ : InMux
    port map (
            O => \N__18212\,
            I => \N__18209\
        );

    \I__3305\ : LocalMux
    port map (
            O => \N__18209\,
            I => \N__18206\
        );

    \I__3304\ : Odrv4
    port map (
            O => \N__18206\,
            I => \eeprom.n3269\
        );

    \I__3303\ : InMux
    port map (
            O => \N__18203\,
            I => \N__18199\
        );

    \I__3302\ : CascadeMux
    port map (
            O => \N__18202\,
            I => \N__18196\
        );

    \I__3301\ : LocalMux
    port map (
            O => \N__18199\,
            I => \N__18193\
        );

    \I__3300\ : InMux
    port map (
            O => \N__18196\,
            I => \N__18190\
        );

    \I__3299\ : Span4Mux_v
    port map (
            O => \N__18193\,
            I => \N__18185\
        );

    \I__3298\ : LocalMux
    port map (
            O => \N__18190\,
            I => \N__18185\
        );

    \I__3297\ : Span4Mux_h
    port map (
            O => \N__18185\,
            I => \N__18182\
        );

    \I__3296\ : Odrv4
    port map (
            O => \N__18182\,
            I => \eeprom.n2815\
        );

    \I__3295\ : CascadeMux
    port map (
            O => \N__18179\,
            I => \N__18176\
        );

    \I__3294\ : InMux
    port map (
            O => \N__18176\,
            I => \N__18173\
        );

    \I__3293\ : LocalMux
    port map (
            O => \N__18173\,
            I => \N__18170\
        );

    \I__3292\ : Odrv4
    port map (
            O => \N__18170\,
            I => \eeprom.n2882\
        );

    \I__3291\ : InMux
    port map (
            O => \N__18167\,
            I => \N__18164\
        );

    \I__3290\ : LocalMux
    port map (
            O => \N__18164\,
            I => \N__18161\
        );

    \I__3289\ : Span4Mux_h
    port map (
            O => \N__18161\,
            I => \N__18158\
        );

    \I__3288\ : Odrv4
    port map (
            O => \N__18158\,
            I => \eeprom.n2886\
        );

    \I__3287\ : CascadeMux
    port map (
            O => \N__18155\,
            I => \eeprom.n2918_cascade_\
        );

    \I__3286\ : CascadeMux
    port map (
            O => \N__18152\,
            I => \N__18149\
        );

    \I__3285\ : InMux
    port map (
            O => \N__18149\,
            I => \N__18146\
        );

    \I__3284\ : LocalMux
    port map (
            O => \N__18146\,
            I => \eeprom.n3267\
        );

    \I__3283\ : InMux
    port map (
            O => \N__18143\,
            I => \N__18140\
        );

    \I__3282\ : LocalMux
    port map (
            O => \N__18140\,
            I => \N__18136\
        );

    \I__3281\ : InMux
    port map (
            O => \N__18139\,
            I => \N__18133\
        );

    \I__3280\ : Span4Mux_v
    port map (
            O => \N__18136\,
            I => \N__18129\
        );

    \I__3279\ : LocalMux
    port map (
            O => \N__18133\,
            I => \N__18126\
        );

    \I__3278\ : InMux
    port map (
            O => \N__18132\,
            I => \N__18123\
        );

    \I__3277\ : Odrv4
    port map (
            O => \N__18129\,
            I => \eeprom.n2705\
        );

    \I__3276\ : Odrv12
    port map (
            O => \N__18126\,
            I => \eeprom.n2705\
        );

    \I__3275\ : LocalMux
    port map (
            O => \N__18123\,
            I => \eeprom.n2705\
        );

    \I__3274\ : CascadeMux
    port map (
            O => \N__18116\,
            I => \N__18113\
        );

    \I__3273\ : InMux
    port map (
            O => \N__18113\,
            I => \N__18110\
        );

    \I__3272\ : LocalMux
    port map (
            O => \N__18110\,
            I => \N__18107\
        );

    \I__3271\ : Span4Mux_h
    port map (
            O => \N__18107\,
            I => \N__18104\
        );

    \I__3270\ : Odrv4
    port map (
            O => \N__18104\,
            I => \eeprom.n2772\
        );

    \I__3269\ : CascadeMux
    port map (
            O => \N__18101\,
            I => \N__18098\
        );

    \I__3268\ : InMux
    port map (
            O => \N__18098\,
            I => \N__18095\
        );

    \I__3267\ : LocalMux
    port map (
            O => \N__18095\,
            I => \N__18091\
        );

    \I__3266\ : InMux
    port map (
            O => \N__18094\,
            I => \N__18088\
        );

    \I__3265\ : Span4Mux_h
    port map (
            O => \N__18091\,
            I => \N__18085\
        );

    \I__3264\ : LocalMux
    port map (
            O => \N__18088\,
            I => \N__18082\
        );

    \I__3263\ : Odrv4
    port map (
            O => \N__18085\,
            I => \eeprom.n2803\
        );

    \I__3262\ : Odrv12
    port map (
            O => \N__18082\,
            I => \eeprom.n2803\
        );

    \I__3261\ : CascadeMux
    port map (
            O => \N__18077\,
            I => \eeprom.n2804_cascade_\
        );

    \I__3260\ : InMux
    port map (
            O => \N__18074\,
            I => \N__18071\
        );

    \I__3259\ : LocalMux
    port map (
            O => \N__18071\,
            I => \N__18068\
        );

    \I__3258\ : Odrv4
    port map (
            O => \N__18068\,
            I => \eeprom.n3276\
        );

    \I__3257\ : CascadeMux
    port map (
            O => \N__18065\,
            I => \N__18062\
        );

    \I__3256\ : InMux
    port map (
            O => \N__18062\,
            I => \N__18059\
        );

    \I__3255\ : LocalMux
    port map (
            O => \N__18059\,
            I => \eeprom.n3279\
        );

    \I__3254\ : InMux
    port map (
            O => \N__18056\,
            I => \N__18053\
        );

    \I__3253\ : LocalMux
    port map (
            O => \N__18053\,
            I => \N__18050\
        );

    \I__3252\ : Odrv4
    port map (
            O => \N__18050\,
            I => \eeprom.n3271\
        );

    \I__3251\ : CascadeMux
    port map (
            O => \N__18047\,
            I => \N__18044\
        );

    \I__3250\ : InMux
    port map (
            O => \N__18044\,
            I => \N__18041\
        );

    \I__3249\ : LocalMux
    port map (
            O => \N__18041\,
            I => \N__18038\
        );

    \I__3248\ : Odrv4
    port map (
            O => \N__18038\,
            I => \eeprom.n3277\
        );

    \I__3247\ : InMux
    port map (
            O => \N__18035\,
            I => \N__18030\
        );

    \I__3246\ : InMux
    port map (
            O => \N__18034\,
            I => \N__18025\
        );

    \I__3245\ : InMux
    port map (
            O => \N__18033\,
            I => \N__18025\
        );

    \I__3244\ : LocalMux
    port map (
            O => \N__18030\,
            I => \eeprom.n3209\
        );

    \I__3243\ : LocalMux
    port map (
            O => \N__18025\,
            I => \eeprom.n3209\
        );

    \I__3242\ : InMux
    port map (
            O => \N__18020\,
            I => \N__18017\
        );

    \I__3241\ : LocalMux
    port map (
            O => \N__18017\,
            I => \eeprom.n3369\
        );

    \I__3240\ : InMux
    port map (
            O => \N__18014\,
            I => \N__18011\
        );

    \I__3239\ : LocalMux
    port map (
            O => \N__18011\,
            I => \N__18008\
        );

    \I__3238\ : Span4Mux_h
    port map (
            O => \N__18008\,
            I => \N__18005\
        );

    \I__3237\ : Span4Mux_h
    port map (
            O => \N__18005\,
            I => \N__18002\
        );

    \I__3236\ : Span4Mux_h
    port map (
            O => \N__18002\,
            I => \N__17999\
        );

    \I__3235\ : Odrv4
    port map (
            O => \N__17999\,
            I => \eeprom.n27\
        );

    \I__3234\ : InMux
    port map (
            O => \N__17996\,
            I => \N__17993\
        );

    \I__3233\ : LocalMux
    port map (
            O => \N__17993\,
            I => \N__17990\
        );

    \I__3232\ : Odrv4
    port map (
            O => \N__17990\,
            I => \eeprom.n3268\
        );

    \I__3231\ : InMux
    port map (
            O => \N__17987\,
            I => \N__17984\
        );

    \I__3230\ : LocalMux
    port map (
            O => \N__17984\,
            I => \N__17981\
        );

    \I__3229\ : Span4Mux_v
    port map (
            O => \N__17981\,
            I => \N__17978\
        );

    \I__3228\ : Span4Mux_h
    port map (
            O => \N__17978\,
            I => \N__17975\
        );

    \I__3227\ : Span4Mux_h
    port map (
            O => \N__17975\,
            I => \N__17972\
        );

    \I__3226\ : Odrv4
    port map (
            O => \N__17972\,
            I => \eeprom.n32_adj_480\
        );

    \I__3225\ : InMux
    port map (
            O => \N__17969\,
            I => \N__17966\
        );

    \I__3224\ : LocalMux
    port map (
            O => \N__17966\,
            I => \N__17963\
        );

    \I__3223\ : Odrv4
    port map (
            O => \N__17963\,
            I => \eeprom.n3273\
        );

    \I__3222\ : InMux
    port map (
            O => \N__17960\,
            I => \N__17957\
        );

    \I__3221\ : LocalMux
    port map (
            O => \N__17957\,
            I => \N__17954\
        );

    \I__3220\ : Odrv4
    port map (
            O => \N__17954\,
            I => \eeprom.n3280\
        );

    \I__3219\ : CascadeMux
    port map (
            O => \N__17951\,
            I => \N__17947\
        );

    \I__3218\ : CascadeMux
    port map (
            O => \N__17950\,
            I => \N__17944\
        );

    \I__3217\ : InMux
    port map (
            O => \N__17947\,
            I => \N__17941\
        );

    \I__3216\ : InMux
    port map (
            O => \N__17944\,
            I => \N__17938\
        );

    \I__3215\ : LocalMux
    port map (
            O => \N__17941\,
            I => \eeprom.n3312\
        );

    \I__3214\ : LocalMux
    port map (
            O => \N__17938\,
            I => \eeprom.n3312\
        );

    \I__3213\ : InMux
    port map (
            O => \N__17933\,
            I => \N__17930\
        );

    \I__3212\ : LocalMux
    port map (
            O => \N__17930\,
            I => \eeprom.n3379\
        );

    \I__3211\ : CascadeMux
    port map (
            O => \N__17927\,
            I => \eeprom.n3312_cascade_\
        );

    \I__3210\ : InMux
    port map (
            O => \N__17924\,
            I => \N__17921\
        );

    \I__3209\ : LocalMux
    port map (
            O => \N__17921\,
            I => \N__17918\
        );

    \I__3208\ : Odrv4
    port map (
            O => \N__17918\,
            I => \eeprom.n3275\
        );

    \I__3207\ : CascadeMux
    port map (
            O => \N__17915\,
            I => \N__17911\
        );

    \I__3206\ : InMux
    port map (
            O => \N__17914\,
            I => \N__17908\
        );

    \I__3205\ : InMux
    port map (
            O => \N__17911\,
            I => \N__17905\
        );

    \I__3204\ : LocalMux
    port map (
            O => \N__17908\,
            I => \eeprom.n3307\
        );

    \I__3203\ : LocalMux
    port map (
            O => \N__17905\,
            I => \eeprom.n3307\
        );

    \I__3202\ : InMux
    port map (
            O => \N__17900\,
            I => \N__17897\
        );

    \I__3201\ : LocalMux
    port map (
            O => \N__17897\,
            I => \eeprom.n3374\
        );

    \I__3200\ : CascadeMux
    port map (
            O => \N__17894\,
            I => \eeprom.n3307_cascade_\
        );

    \I__3199\ : CascadeMux
    port map (
            O => \N__17891\,
            I => \eeprom.n28_adj_482_cascade_\
        );

    \I__3198\ : InMux
    port map (
            O => \N__17888\,
            I => \N__17885\
        );

    \I__3197\ : LocalMux
    port map (
            O => \N__17885\,
            I => \N__17882\
        );

    \I__3196\ : Odrv4
    port map (
            O => \N__17882\,
            I => \eeprom.n3278\
        );

    \I__3195\ : CascadeMux
    port map (
            O => \N__17879\,
            I => \eeprom.n3232_cascade_\
        );

    \I__3194\ : InMux
    port map (
            O => \N__17876\,
            I => \N__17873\
        );

    \I__3193\ : LocalMux
    port map (
            O => \N__17873\,
            I => \eeprom.n3367\
        );

    \I__3192\ : CascadeMux
    port map (
            O => \N__17870\,
            I => \eeprom.n2904_cascade_\
        );

    \I__3191\ : CascadeMux
    port map (
            O => \N__17867\,
            I => \N__17864\
        );

    \I__3190\ : InMux
    port map (
            O => \N__17864\,
            I => \N__17861\
        );

    \I__3189\ : LocalMux
    port map (
            O => \N__17861\,
            I => \N__17858\
        );

    \I__3188\ : Span4Mux_h
    port map (
            O => \N__17858\,
            I => \N__17855\
        );

    \I__3187\ : Odrv4
    port map (
            O => \N__17855\,
            I => \eeprom.n3286\
        );

    \I__3186\ : InMux
    port map (
            O => \N__17852\,
            I => \N__17849\
        );

    \I__3185\ : LocalMux
    port map (
            O => \N__17849\,
            I => \N__17846\
        );

    \I__3184\ : Odrv4
    port map (
            O => \N__17846\,
            I => \eeprom.n3285\
        );

    \I__3183\ : CascadeMux
    port map (
            O => \N__17843\,
            I => \N__17840\
        );

    \I__3182\ : InMux
    port map (
            O => \N__17840\,
            I => \N__17837\
        );

    \I__3181\ : LocalMux
    port map (
            O => \N__17837\,
            I => \eeprom.n3371\
        );

    \I__3180\ : InMux
    port map (
            O => \N__17834\,
            I => \N__17831\
        );

    \I__3179\ : LocalMux
    port map (
            O => \N__17831\,
            I => \N__17828\
        );

    \I__3178\ : Odrv4
    port map (
            O => \N__17828\,
            I => \eeprom.n3282\
        );

    \I__3177\ : CascadeMux
    port map (
            O => \N__17825\,
            I => \eeprom.n3314_cascade_\
        );

    \I__3176\ : InMux
    port map (
            O => \N__17822\,
            I => \N__17819\
        );

    \I__3175\ : LocalMux
    port map (
            O => \N__17819\,
            I => \N__17816\
        );

    \I__3174\ : Span4Mux_h
    port map (
            O => \N__17816\,
            I => \N__17813\
        );

    \I__3173\ : Odrv4
    port map (
            O => \N__17813\,
            I => \eeprom.n3272\
        );

    \I__3172\ : InMux
    port map (
            O => \N__17810\,
            I => \N__17807\
        );

    \I__3171\ : LocalMux
    port map (
            O => \N__17807\,
            I => \N__17804\
        );

    \I__3170\ : Odrv4
    port map (
            O => \N__17804\,
            I => \eeprom.n3274\
        );

    \I__3169\ : InMux
    port map (
            O => \N__17801\,
            I => \eeprom.n3625\
        );

    \I__3168\ : InMux
    port map (
            O => \N__17798\,
            I => \eeprom.n3626\
        );

    \I__3167\ : InMux
    port map (
            O => \N__17795\,
            I => \eeprom.n3627\
        );

    \I__3166\ : InMux
    port map (
            O => \N__17792\,
            I => \eeprom.n3628\
        );

    \I__3165\ : InMux
    port map (
            O => \N__17789\,
            I => \eeprom.n3629\
        );

    \I__3164\ : InMux
    port map (
            O => \N__17786\,
            I => \eeprom.n3630\
        );

    \I__3163\ : InMux
    port map (
            O => \N__17783\,
            I => \bfn_9_25_0_\
        );

    \I__3162\ : InMux
    port map (
            O => \N__17780\,
            I => \N__17777\
        );

    \I__3161\ : LocalMux
    port map (
            O => \N__17777\,
            I => \eeprom.n2873\
        );

    \I__3160\ : CascadeMux
    port map (
            O => \N__17774\,
            I => \N__17771\
        );

    \I__3159\ : InMux
    port map (
            O => \N__17771\,
            I => \N__17768\
        );

    \I__3158\ : LocalMux
    port map (
            O => \N__17768\,
            I => \eeprom.n2872\
        );

    \I__3157\ : InMux
    port map (
            O => \N__17765\,
            I => \bfn_9_23_0_\
        );

    \I__3156\ : InMux
    port map (
            O => \N__17762\,
            I => \eeprom.n3616\
        );

    \I__3155\ : InMux
    port map (
            O => \N__17759\,
            I => \eeprom.n3617\
        );

    \I__3154\ : InMux
    port map (
            O => \N__17756\,
            I => \eeprom.n3618\
        );

    \I__3153\ : InMux
    port map (
            O => \N__17753\,
            I => \eeprom.n3619\
        );

    \I__3152\ : InMux
    port map (
            O => \N__17750\,
            I => \eeprom.n3620\
        );

    \I__3151\ : InMux
    port map (
            O => \N__17747\,
            I => \eeprom.n3621\
        );

    \I__3150\ : InMux
    port map (
            O => \N__17744\,
            I => \eeprom.n3622\
        );

    \I__3149\ : InMux
    port map (
            O => \N__17741\,
            I => \bfn_9_24_0_\
        );

    \I__3148\ : InMux
    port map (
            O => \N__17738\,
            I => \eeprom.n3624\
        );

    \I__3147\ : InMux
    port map (
            O => \N__17735\,
            I => \eeprom.n3700\
        );

    \I__3146\ : InMux
    port map (
            O => \N__17732\,
            I => \bfn_9_22_0_\
        );

    \I__3145\ : InMux
    port map (
            O => \N__17729\,
            I => \eeprom.n3702\
        );

    \I__3144\ : InMux
    port map (
            O => \N__17726\,
            I => \eeprom.n3703\
        );

    \I__3143\ : InMux
    port map (
            O => \N__17723\,
            I => \eeprom.n3704\
        );

    \I__3142\ : InMux
    port map (
            O => \N__17720\,
            I => \eeprom.n3705\
        );

    \I__3141\ : InMux
    port map (
            O => \N__17717\,
            I => \N__17714\
        );

    \I__3140\ : LocalMux
    port map (
            O => \N__17714\,
            I => \N__17710\
        );

    \I__3139\ : InMux
    port map (
            O => \N__17713\,
            I => \N__17707\
        );

    \I__3138\ : Span4Mux_v
    port map (
            O => \N__17710\,
            I => \N__17703\
        );

    \I__3137\ : LocalMux
    port map (
            O => \N__17707\,
            I => \N__17700\
        );

    \I__3136\ : InMux
    port map (
            O => \N__17706\,
            I => \N__17697\
        );

    \I__3135\ : Odrv4
    port map (
            O => \N__17703\,
            I => \eeprom.n2706\
        );

    \I__3134\ : Odrv12
    port map (
            O => \N__17700\,
            I => \eeprom.n2706\
        );

    \I__3133\ : LocalMux
    port map (
            O => \N__17697\,
            I => \eeprom.n2706\
        );

    \I__3132\ : InMux
    port map (
            O => \N__17690\,
            I => \N__17687\
        );

    \I__3131\ : LocalMux
    port map (
            O => \N__17687\,
            I => \N__17684\
        );

    \I__3130\ : Odrv4
    port map (
            O => \N__17684\,
            I => \eeprom.n2773\
        );

    \I__3129\ : InMux
    port map (
            O => \N__17681\,
            I => \N__17677\
        );

    \I__3128\ : CascadeMux
    port map (
            O => \N__17680\,
            I => \N__17674\
        );

    \I__3127\ : LocalMux
    port map (
            O => \N__17677\,
            I => \N__17671\
        );

    \I__3126\ : InMux
    port map (
            O => \N__17674\,
            I => \N__17668\
        );

    \I__3125\ : Span4Mux_h
    port map (
            O => \N__17671\,
            I => \N__17665\
        );

    \I__3124\ : LocalMux
    port map (
            O => \N__17668\,
            I => \N__17662\
        );

    \I__3123\ : Odrv4
    port map (
            O => \N__17665\,
            I => \eeprom.n2709\
        );

    \I__3122\ : Odrv4
    port map (
            O => \N__17662\,
            I => \eeprom.n2709\
        );

    \I__3121\ : CascadeMux
    port map (
            O => \N__17657\,
            I => \N__17654\
        );

    \I__3120\ : InMux
    port map (
            O => \N__17654\,
            I => \N__17651\
        );

    \I__3119\ : LocalMux
    port map (
            O => \N__17651\,
            I => \N__17648\
        );

    \I__3118\ : Odrv4
    port map (
            O => \N__17648\,
            I => \eeprom.n2776\
        );

    \I__3117\ : InMux
    port map (
            O => \N__17645\,
            I => \eeprom.n3690\
        );

    \I__3116\ : InMux
    port map (
            O => \N__17642\,
            I => \eeprom.n3691\
        );

    \I__3115\ : InMux
    port map (
            O => \N__17639\,
            I => \eeprom.n3692\
        );

    \I__3114\ : InMux
    port map (
            O => \N__17636\,
            I => \bfn_9_21_0_\
        );

    \I__3113\ : InMux
    port map (
            O => \N__17633\,
            I => \eeprom.n3694\
        );

    \I__3112\ : InMux
    port map (
            O => \N__17630\,
            I => \eeprom.n3695\
        );

    \I__3111\ : InMux
    port map (
            O => \N__17627\,
            I => \eeprom.n3696\
        );

    \I__3110\ : InMux
    port map (
            O => \N__17624\,
            I => \eeprom.n3697\
        );

    \I__3109\ : InMux
    port map (
            O => \N__17621\,
            I => \eeprom.n3698\
        );

    \I__3108\ : InMux
    port map (
            O => \N__17618\,
            I => \eeprom.n3699\
        );

    \I__3107\ : InMux
    port map (
            O => \N__17615\,
            I => \eeprom.n3724\
        );

    \I__3106\ : InMux
    port map (
            O => \N__17612\,
            I => \eeprom.n3725\
        );

    \I__3105\ : InMux
    port map (
            O => \N__17609\,
            I => \eeprom.n3726\
        );

    \I__3104\ : InMux
    port map (
            O => \N__17606\,
            I => \bfn_9_20_0_\
        );

    \I__3103\ : InMux
    port map (
            O => \N__17603\,
            I => \eeprom.n3686\
        );

    \I__3102\ : InMux
    port map (
            O => \N__17600\,
            I => \eeprom.n3687\
        );

    \I__3101\ : InMux
    port map (
            O => \N__17597\,
            I => \eeprom.n3688\
        );

    \I__3100\ : InMux
    port map (
            O => \N__17594\,
            I => \eeprom.n3689\
        );

    \I__3099\ : CascadeMux
    port map (
            O => \N__17591\,
            I => \N__17588\
        );

    \I__3098\ : InMux
    port map (
            O => \N__17588\,
            I => \N__17585\
        );

    \I__3097\ : LocalMux
    port map (
            O => \N__17585\,
            I => \eeprom.n3281\
        );

    \I__3096\ : InMux
    port map (
            O => \N__17582\,
            I => \eeprom.n3715\
        );

    \I__3095\ : InMux
    port map (
            O => \N__17579\,
            I => \eeprom.n3716\
        );

    \I__3094\ : InMux
    port map (
            O => \N__17576\,
            I => \eeprom.n3717\
        );

    \I__3093\ : InMux
    port map (
            O => \N__17573\,
            I => \eeprom.n3718\
        );

    \I__3092\ : InMux
    port map (
            O => \N__17570\,
            I => \eeprom.n3719\
        );

    \I__3091\ : InMux
    port map (
            O => \N__17567\,
            I => \eeprom.n3720\
        );

    \I__3090\ : InMux
    port map (
            O => \N__17564\,
            I => \bfn_9_19_0_\
        );

    \I__3089\ : InMux
    port map (
            O => \N__17561\,
            I => \eeprom.n3722\
        );

    \I__3088\ : InMux
    port map (
            O => \N__17558\,
            I => \eeprom.n3723\
        );

    \I__3087\ : InMux
    port map (
            O => \N__17555\,
            I => \eeprom.n3706\
        );

    \I__3086\ : InMux
    port map (
            O => \N__17552\,
            I => \eeprom.n3707\
        );

    \I__3085\ : InMux
    port map (
            O => \N__17549\,
            I => \eeprom.n3708\
        );

    \I__3084\ : InMux
    port map (
            O => \N__17546\,
            I => \eeprom.n3709\
        );

    \I__3083\ : InMux
    port map (
            O => \N__17543\,
            I => \eeprom.n3710\
        );

    \I__3082\ : InMux
    port map (
            O => \N__17540\,
            I => \eeprom.n3711\
        );

    \I__3081\ : InMux
    port map (
            O => \N__17537\,
            I => \eeprom.n3712\
        );

    \I__3080\ : InMux
    port map (
            O => \N__17534\,
            I => \bfn_9_18_0_\
        );

    \I__3079\ : InMux
    port map (
            O => \N__17531\,
            I => \eeprom.n3714\
        );

    \I__3078\ : InMux
    port map (
            O => \N__17528\,
            I => \eeprom.n3613\
        );

    \I__3077\ : InMux
    port map (
            O => \N__17525\,
            I => \eeprom.n3614\
        );

    \I__3076\ : CascadeMux
    port map (
            O => \N__17522\,
            I => \N__17519\
        );

    \I__3075\ : InMux
    port map (
            O => \N__17519\,
            I => \N__17515\
        );

    \I__3074\ : CascadeMux
    port map (
            O => \N__17518\,
            I => \N__17512\
        );

    \I__3073\ : LocalMux
    port map (
            O => \N__17515\,
            I => \N__17509\
        );

    \I__3072\ : InMux
    port map (
            O => \N__17512\,
            I => \N__17506\
        );

    \I__3071\ : Odrv4
    port map (
            O => \N__17509\,
            I => \eeprom.n2704\
        );

    \I__3070\ : LocalMux
    port map (
            O => \N__17506\,
            I => \eeprom.n2704\
        );

    \I__3069\ : InMux
    port map (
            O => \N__17501\,
            I => \eeprom.n3615\
        );

    \I__3068\ : InMux
    port map (
            O => \N__17498\,
            I => \N__17495\
        );

    \I__3067\ : LocalMux
    port map (
            O => \N__17495\,
            I => \eeprom.n2777\
        );

    \I__3066\ : CascadeMux
    port map (
            O => \N__17492\,
            I => \N__17488\
        );

    \I__3065\ : InMux
    port map (
            O => \N__17491\,
            I => \N__17484\
        );

    \I__3064\ : InMux
    port map (
            O => \N__17488\,
            I => \N__17481\
        );

    \I__3063\ : InMux
    port map (
            O => \N__17487\,
            I => \N__17478\
        );

    \I__3062\ : LocalMux
    port map (
            O => \N__17484\,
            I => \N__17473\
        );

    \I__3061\ : LocalMux
    port map (
            O => \N__17481\,
            I => \N__17473\
        );

    \I__3060\ : LocalMux
    port map (
            O => \N__17478\,
            I => \N__17470\
        );

    \I__3059\ : Odrv4
    port map (
            O => \N__17473\,
            I => \eeprom.n2710\
        );

    \I__3058\ : Odrv4
    port map (
            O => \N__17470\,
            I => \eeprom.n2710\
        );

    \I__3057\ : InMux
    port map (
            O => \N__17465\,
            I => \N__17462\
        );

    \I__3056\ : LocalMux
    port map (
            O => \N__17462\,
            I => \eeprom.n2778\
        );

    \I__3055\ : InMux
    port map (
            O => \N__17459\,
            I => \N__17454\
        );

    \I__3054\ : InMux
    port map (
            O => \N__17458\,
            I => \N__17451\
        );

    \I__3053\ : InMux
    port map (
            O => \N__17457\,
            I => \N__17448\
        );

    \I__3052\ : LocalMux
    port map (
            O => \N__17454\,
            I => \N__17441\
        );

    \I__3051\ : LocalMux
    port map (
            O => \N__17451\,
            I => \N__17441\
        );

    \I__3050\ : LocalMux
    port map (
            O => \N__17448\,
            I => \N__17441\
        );

    \I__3049\ : Odrv12
    port map (
            O => \N__17441\,
            I => \eeprom.n2711\
        );

    \I__3048\ : InMux
    port map (
            O => \N__17438\,
            I => \N__17434\
        );

    \I__3047\ : CascadeMux
    port map (
            O => \N__17437\,
            I => \N__17431\
        );

    \I__3046\ : LocalMux
    port map (
            O => \N__17434\,
            I => \N__17427\
        );

    \I__3045\ : InMux
    port map (
            O => \N__17431\,
            I => \N__17424\
        );

    \I__3044\ : InMux
    port map (
            O => \N__17430\,
            I => \N__17421\
        );

    \I__3043\ : Span4Mux_v
    port map (
            O => \N__17427\,
            I => \N__17416\
        );

    \I__3042\ : LocalMux
    port map (
            O => \N__17424\,
            I => \N__17416\
        );

    \I__3041\ : LocalMux
    port map (
            O => \N__17421\,
            I => \eeprom.n2717\
        );

    \I__3040\ : Odrv4
    port map (
            O => \N__17416\,
            I => \eeprom.n2717\
        );

    \I__3039\ : CascadeMux
    port map (
            O => \N__17411\,
            I => \N__17408\
        );

    \I__3038\ : InMux
    port map (
            O => \N__17408\,
            I => \N__17405\
        );

    \I__3037\ : LocalMux
    port map (
            O => \N__17405\,
            I => \N__17402\
        );

    \I__3036\ : Odrv4
    port map (
            O => \N__17402\,
            I => \eeprom.n2784\
        );

    \I__3035\ : InMux
    port map (
            O => \N__17399\,
            I => \N__17396\
        );

    \I__3034\ : LocalMux
    port map (
            O => \N__17396\,
            I => \N__17393\
        );

    \I__3033\ : Odrv4
    port map (
            O => \N__17393\,
            I => \eeprom.n2782\
        );

    \I__3032\ : InMux
    port map (
            O => \N__17390\,
            I => \N__17386\
        );

    \I__3031\ : CascadeMux
    port map (
            O => \N__17389\,
            I => \N__17383\
        );

    \I__3030\ : LocalMux
    port map (
            O => \N__17386\,
            I => \N__17380\
        );

    \I__3029\ : InMux
    port map (
            O => \N__17383\,
            I => \N__17377\
        );

    \I__3028\ : Span4Mux_v
    port map (
            O => \N__17380\,
            I => \N__17371\
        );

    \I__3027\ : LocalMux
    port map (
            O => \N__17377\,
            I => \N__17371\
        );

    \I__3026\ : InMux
    port map (
            O => \N__17376\,
            I => \N__17368\
        );

    \I__3025\ : Odrv4
    port map (
            O => \N__17371\,
            I => \eeprom.n2715\
        );

    \I__3024\ : LocalMux
    port map (
            O => \N__17368\,
            I => \eeprom.n2715\
        );

    \I__3023\ : InMux
    port map (
            O => \N__17363\,
            I => \N__17359\
        );

    \I__3022\ : CascadeMux
    port map (
            O => \N__17362\,
            I => \N__17356\
        );

    \I__3021\ : LocalMux
    port map (
            O => \N__17359\,
            I => \N__17353\
        );

    \I__3020\ : InMux
    port map (
            O => \N__17356\,
            I => \N__17350\
        );

    \I__3019\ : Span4Mux_v
    port map (
            O => \N__17353\,
            I => \N__17345\
        );

    \I__3018\ : LocalMux
    port map (
            O => \N__17350\,
            I => \N__17345\
        );

    \I__3017\ : Odrv4
    port map (
            O => \N__17345\,
            I => \eeprom.n2713\
        );

    \I__3016\ : CascadeMux
    port map (
            O => \N__17342\,
            I => \N__17339\
        );

    \I__3015\ : InMux
    port map (
            O => \N__17339\,
            I => \N__17336\
        );

    \I__3014\ : LocalMux
    port map (
            O => \N__17336\,
            I => \N__17333\
        );

    \I__3013\ : Odrv4
    port map (
            O => \N__17333\,
            I => \eeprom.n2780\
        );

    \I__3012\ : InMux
    port map (
            O => \N__17330\,
            I => \bfn_9_17_0_\
        );

    \I__3011\ : CascadeMux
    port map (
            O => \N__17327\,
            I => \N__17324\
        );

    \I__3010\ : InMux
    port map (
            O => \N__17324\,
            I => \N__17320\
        );

    \I__3009\ : InMux
    port map (
            O => \N__17323\,
            I => \N__17316\
        );

    \I__3008\ : LocalMux
    port map (
            O => \N__17320\,
            I => \N__17313\
        );

    \I__3007\ : InMux
    port map (
            O => \N__17319\,
            I => \N__17310\
        );

    \I__3006\ : LocalMux
    port map (
            O => \N__17316\,
            I => \eeprom.n2714\
        );

    \I__3005\ : Odrv4
    port map (
            O => \N__17313\,
            I => \eeprom.n2714\
        );

    \I__3004\ : LocalMux
    port map (
            O => \N__17310\,
            I => \eeprom.n2714\
        );

    \I__3003\ : InMux
    port map (
            O => \N__17303\,
            I => \N__17300\
        );

    \I__3002\ : LocalMux
    port map (
            O => \N__17300\,
            I => \eeprom.n2781\
        );

    \I__3001\ : InMux
    port map (
            O => \N__17297\,
            I => \eeprom.n3605\
        );

    \I__3000\ : InMux
    port map (
            O => \N__17294\,
            I => \eeprom.n3606\
        );

    \I__2999\ : InMux
    port map (
            O => \N__17291\,
            I => \eeprom.n3607\
        );

    \I__2998\ : InMux
    port map (
            O => \N__17288\,
            I => \bfn_7_22_0_\
        );

    \I__2997\ : InMux
    port map (
            O => \N__17285\,
            I => \eeprom.n3609\
        );

    \I__2996\ : InMux
    port map (
            O => \N__17282\,
            I => \eeprom.n3610\
        );

    \I__2995\ : InMux
    port map (
            O => \N__17279\,
            I => \eeprom.n3611\
        );

    \I__2994\ : InMux
    port map (
            O => \N__17276\,
            I => \eeprom.n3612\
        );

    \I__2993\ : InMux
    port map (
            O => \N__17273\,
            I => \N__17270\
        );

    \I__2992\ : LocalMux
    port map (
            O => \N__17270\,
            I => \N__17267\
        );

    \I__2991\ : Span4Mux_v
    port map (
            O => \N__17267\,
            I => \N__17264\
        );

    \I__2990\ : Span4Mux_h
    port map (
            O => \N__17264\,
            I => \N__17261\
        );

    \I__2989\ : Odrv4
    port map (
            O => \N__17261\,
            I => \eeprom.n28\
        );

    \I__2988\ : InMux
    port map (
            O => \N__17258\,
            I => \N__17255\
        );

    \I__2987\ : LocalMux
    port map (
            O => \N__17255\,
            I => \N__17251\
        );

    \I__2986\ : InMux
    port map (
            O => \N__17254\,
            I => \N__17248\
        );

    \I__2985\ : Span4Mux_h
    port map (
            O => \N__17251\,
            I => \N__17244\
        );

    \I__2984\ : LocalMux
    port map (
            O => \N__17248\,
            I => \N__17241\
        );

    \I__2983\ : InMux
    port map (
            O => \N__17247\,
            I => \N__17238\
        );

    \I__2982\ : Odrv4
    port map (
            O => \N__17244\,
            I => \eeprom.n2610\
        );

    \I__2981\ : Odrv12
    port map (
            O => \N__17241\,
            I => \eeprom.n2610\
        );

    \I__2980\ : LocalMux
    port map (
            O => \N__17238\,
            I => \eeprom.n2610\
        );

    \I__2979\ : CascadeMux
    port map (
            O => \N__17231\,
            I => \N__17228\
        );

    \I__2978\ : InMux
    port map (
            O => \N__17228\,
            I => \N__17225\
        );

    \I__2977\ : LocalMux
    port map (
            O => \N__17225\,
            I => \eeprom.n2677\
        );

    \I__2976\ : InMux
    port map (
            O => \N__17222\,
            I => \N__17214\
        );

    \I__2975\ : CascadeMux
    port map (
            O => \N__17221\,
            I => \N__17207\
        );

    \I__2974\ : CascadeMux
    port map (
            O => \N__17220\,
            I => \N__17204\
        );

    \I__2973\ : CascadeMux
    port map (
            O => \N__17219\,
            I => \N__17199\
        );

    \I__2972\ : CascadeMux
    port map (
            O => \N__17218\,
            I => \N__17195\
        );

    \I__2971\ : InMux
    port map (
            O => \N__17217\,
            I => \N__17191\
        );

    \I__2970\ : LocalMux
    port map (
            O => \N__17214\,
            I => \N__17188\
        );

    \I__2969\ : InMux
    port map (
            O => \N__17213\,
            I => \N__17185\
        );

    \I__2968\ : InMux
    port map (
            O => \N__17212\,
            I => \N__17180\
        );

    \I__2967\ : InMux
    port map (
            O => \N__17211\,
            I => \N__17180\
        );

    \I__2966\ : InMux
    port map (
            O => \N__17210\,
            I => \N__17171\
        );

    \I__2965\ : InMux
    port map (
            O => \N__17207\,
            I => \N__17171\
        );

    \I__2964\ : InMux
    port map (
            O => \N__17204\,
            I => \N__17171\
        );

    \I__2963\ : InMux
    port map (
            O => \N__17203\,
            I => \N__17171\
        );

    \I__2962\ : InMux
    port map (
            O => \N__17202\,
            I => \N__17160\
        );

    \I__2961\ : InMux
    port map (
            O => \N__17199\,
            I => \N__17160\
        );

    \I__2960\ : InMux
    port map (
            O => \N__17198\,
            I => \N__17160\
        );

    \I__2959\ : InMux
    port map (
            O => \N__17195\,
            I => \N__17160\
        );

    \I__2958\ : InMux
    port map (
            O => \N__17194\,
            I => \N__17160\
        );

    \I__2957\ : LocalMux
    port map (
            O => \N__17191\,
            I => \eeprom.n2638\
        );

    \I__2956\ : Odrv4
    port map (
            O => \N__17188\,
            I => \eeprom.n2638\
        );

    \I__2955\ : LocalMux
    port map (
            O => \N__17185\,
            I => \eeprom.n2638\
        );

    \I__2954\ : LocalMux
    port map (
            O => \N__17180\,
            I => \eeprom.n2638\
        );

    \I__2953\ : LocalMux
    port map (
            O => \N__17171\,
            I => \eeprom.n2638\
        );

    \I__2952\ : LocalMux
    port map (
            O => \N__17160\,
            I => \eeprom.n2638\
        );

    \I__2951\ : InMux
    port map (
            O => \N__17147\,
            I => \N__17144\
        );

    \I__2950\ : LocalMux
    port map (
            O => \N__17144\,
            I => \N__17141\
        );

    \I__2949\ : Odrv4
    port map (
            O => \N__17141\,
            I => \eeprom.n18\
        );

    \I__2948\ : CascadeMux
    port map (
            O => \N__17138\,
            I => \eeprom.n2709_cascade_\
        );

    \I__2947\ : InMux
    port map (
            O => \N__17135\,
            I => \N__17132\
        );

    \I__2946\ : LocalMux
    port map (
            O => \N__17132\,
            I => \eeprom.n13_adj_417\
        );

    \I__2945\ : CascadeMux
    port map (
            O => \N__17129\,
            I => \eeprom.n2737_cascade_\
        );

    \I__2944\ : InMux
    port map (
            O => \N__17126\,
            I => \N__17123\
        );

    \I__2943\ : LocalMux
    port map (
            O => \N__17123\,
            I => \N__17118\
        );

    \I__2942\ : InMux
    port map (
            O => \N__17122\,
            I => \N__17115\
        );

    \I__2941\ : InMux
    port map (
            O => \N__17121\,
            I => \N__17112\
        );

    \I__2940\ : Span4Mux_h
    port map (
            O => \N__17118\,
            I => \N__17109\
        );

    \I__2939\ : LocalMux
    port map (
            O => \N__17115\,
            I => \N__17104\
        );

    \I__2938\ : LocalMux
    port map (
            O => \N__17112\,
            I => \N__17104\
        );

    \I__2937\ : Span4Mux_h
    port map (
            O => \N__17109\,
            I => \N__17101\
        );

    \I__2936\ : Span12Mux_v
    port map (
            O => \N__17104\,
            I => \N__17098\
        );

    \I__2935\ : Odrv4
    port map (
            O => \N__17101\,
            I => \eeprom.n2719\
        );

    \I__2934\ : Odrv12
    port map (
            O => \N__17098\,
            I => \eeprom.n2719\
        );

    \I__2933\ : InMux
    port map (
            O => \N__17093\,
            I => \N__17090\
        );

    \I__2932\ : LocalMux
    port map (
            O => \N__17090\,
            I => \eeprom.n2786\
        );

    \I__2931\ : InMux
    port map (
            O => \N__17087\,
            I => \bfn_7_21_0_\
        );

    \I__2930\ : CascadeMux
    port map (
            O => \N__17084\,
            I => \N__17081\
        );

    \I__2929\ : InMux
    port map (
            O => \N__17081\,
            I => \N__17077\
        );

    \I__2928\ : InMux
    port map (
            O => \N__17080\,
            I => \N__17074\
        );

    \I__2927\ : LocalMux
    port map (
            O => \N__17077\,
            I => \N__17071\
        );

    \I__2926\ : LocalMux
    port map (
            O => \N__17074\,
            I => \eeprom.n2718\
        );

    \I__2925\ : Odrv4
    port map (
            O => \N__17071\,
            I => \eeprom.n2718\
        );

    \I__2924\ : InMux
    port map (
            O => \N__17066\,
            I => \N__17063\
        );

    \I__2923\ : LocalMux
    port map (
            O => \N__17063\,
            I => \eeprom.n2785\
        );

    \I__2922\ : InMux
    port map (
            O => \N__17060\,
            I => \eeprom.n3601\
        );

    \I__2921\ : InMux
    port map (
            O => \N__17057\,
            I => \eeprom.n3602\
        );

    \I__2920\ : CascadeMux
    port map (
            O => \N__17054\,
            I => \N__17051\
        );

    \I__2919\ : InMux
    port map (
            O => \N__17051\,
            I => \N__17047\
        );

    \I__2918\ : InMux
    port map (
            O => \N__17050\,
            I => \N__17043\
        );

    \I__2917\ : LocalMux
    port map (
            O => \N__17047\,
            I => \N__17040\
        );

    \I__2916\ : InMux
    port map (
            O => \N__17046\,
            I => \N__17037\
        );

    \I__2915\ : LocalMux
    port map (
            O => \N__17043\,
            I => \eeprom.n2716\
        );

    \I__2914\ : Odrv4
    port map (
            O => \N__17040\,
            I => \eeprom.n2716\
        );

    \I__2913\ : LocalMux
    port map (
            O => \N__17037\,
            I => \eeprom.n2716\
        );

    \I__2912\ : InMux
    port map (
            O => \N__17030\,
            I => \N__17027\
        );

    \I__2911\ : LocalMux
    port map (
            O => \N__17027\,
            I => \eeprom.n2783\
        );

    \I__2910\ : InMux
    port map (
            O => \N__17024\,
            I => \eeprom.n3603\
        );

    \I__2909\ : InMux
    port map (
            O => \N__17021\,
            I => \eeprom.n3604\
        );

    \I__2908\ : CascadeMux
    port map (
            O => \N__17018\,
            I => \N__17015\
        );

    \I__2907\ : InMux
    port map (
            O => \N__17015\,
            I => \N__17012\
        );

    \I__2906\ : LocalMux
    port map (
            O => \N__17012\,
            I => \eeprom.n2675\
        );

    \I__2905\ : InMux
    port map (
            O => \N__17009\,
            I => \N__17006\
        );

    \I__2904\ : LocalMux
    port map (
            O => \N__17006\,
            I => \eeprom.n2682\
        );

    \I__2903\ : InMux
    port map (
            O => \N__17003\,
            I => \N__16999\
        );

    \I__2902\ : CascadeMux
    port map (
            O => \N__17002\,
            I => \N__16996\
        );

    \I__2901\ : LocalMux
    port map (
            O => \N__16999\,
            I => \N__16993\
        );

    \I__2900\ : InMux
    port map (
            O => \N__16996\,
            I => \N__16990\
        );

    \I__2899\ : Odrv12
    port map (
            O => \N__16993\,
            I => \eeprom.n2615\
        );

    \I__2898\ : LocalMux
    port map (
            O => \N__16990\,
            I => \eeprom.n2615\
        );

    \I__2897\ : CascadeMux
    port map (
            O => \N__16985\,
            I => \N__16982\
        );

    \I__2896\ : InMux
    port map (
            O => \N__16982\,
            I => \N__16977\
        );

    \I__2895\ : InMux
    port map (
            O => \N__16981\,
            I => \N__16972\
        );

    \I__2894\ : InMux
    port map (
            O => \N__16980\,
            I => \N__16972\
        );

    \I__2893\ : LocalMux
    port map (
            O => \N__16977\,
            I => \eeprom.n2608\
        );

    \I__2892\ : LocalMux
    port map (
            O => \N__16972\,
            I => \eeprom.n2608\
        );

    \I__2891\ : InMux
    port map (
            O => \N__16967\,
            I => \N__16964\
        );

    \I__2890\ : LocalMux
    port map (
            O => \N__16964\,
            I => \N__16961\
        );

    \I__2889\ : Odrv4
    port map (
            O => \N__16961\,
            I => \eeprom.n12\
        );

    \I__2888\ : CascadeMux
    port map (
            O => \N__16958\,
            I => \N__16954\
        );

    \I__2887\ : CascadeMux
    port map (
            O => \N__16957\,
            I => \N__16950\
        );

    \I__2886\ : InMux
    port map (
            O => \N__16954\,
            I => \N__16947\
        );

    \I__2885\ : InMux
    port map (
            O => \N__16953\,
            I => \N__16942\
        );

    \I__2884\ : InMux
    port map (
            O => \N__16950\,
            I => \N__16942\
        );

    \I__2883\ : LocalMux
    port map (
            O => \N__16947\,
            I => \eeprom.n2607\
        );

    \I__2882\ : LocalMux
    port map (
            O => \N__16942\,
            I => \eeprom.n2607\
        );

    \I__2881\ : InMux
    port map (
            O => \N__16937\,
            I => \N__16934\
        );

    \I__2880\ : LocalMux
    port map (
            O => \N__16934\,
            I => \N__16931\
        );

    \I__2879\ : Span4Mux_v
    port map (
            O => \N__16931\,
            I => \N__16928\
        );

    \I__2878\ : Odrv4
    port map (
            O => \N__16928\,
            I => \eeprom.n16\
        );

    \I__2877\ : InMux
    port map (
            O => \N__16925\,
            I => \N__16922\
        );

    \I__2876\ : LocalMux
    port map (
            O => \N__16922\,
            I => \eeprom.n2683\
        );

    \I__2875\ : CascadeMux
    port map (
            O => \N__16919\,
            I => \eeprom.n2638_cascade_\
        );

    \I__2874\ : InMux
    port map (
            O => \N__16916\,
            I => \N__16912\
        );

    \I__2873\ : CascadeMux
    port map (
            O => \N__16915\,
            I => \N__16909\
        );

    \I__2872\ : LocalMux
    port map (
            O => \N__16912\,
            I => \N__16905\
        );

    \I__2871\ : InMux
    port map (
            O => \N__16909\,
            I => \N__16902\
        );

    \I__2870\ : InMux
    port map (
            O => \N__16908\,
            I => \N__16899\
        );

    \I__2869\ : Odrv4
    port map (
            O => \N__16905\,
            I => \eeprom.n2616\
        );

    \I__2868\ : LocalMux
    port map (
            O => \N__16902\,
            I => \eeprom.n2616\
        );

    \I__2867\ : LocalMux
    port map (
            O => \N__16899\,
            I => \eeprom.n2616\
        );

    \I__2866\ : InMux
    port map (
            O => \N__16892\,
            I => \N__16888\
        );

    \I__2865\ : CascadeMux
    port map (
            O => \N__16891\,
            I => \N__16885\
        );

    \I__2864\ : LocalMux
    port map (
            O => \N__16888\,
            I => \N__16881\
        );

    \I__2863\ : InMux
    port map (
            O => \N__16885\,
            I => \N__16878\
        );

    \I__2862\ : InMux
    port map (
            O => \N__16884\,
            I => \N__16875\
        );

    \I__2861\ : Odrv4
    port map (
            O => \N__16881\,
            I => \eeprom.n2617\
        );

    \I__2860\ : LocalMux
    port map (
            O => \N__16878\,
            I => \eeprom.n2617\
        );

    \I__2859\ : LocalMux
    port map (
            O => \N__16875\,
            I => \eeprom.n2617\
        );

    \I__2858\ : CascadeMux
    port map (
            O => \N__16868\,
            I => \N__16865\
        );

    \I__2857\ : InMux
    port map (
            O => \N__16865\,
            I => \N__16862\
        );

    \I__2856\ : LocalMux
    port map (
            O => \N__16862\,
            I => \eeprom.n2684\
        );

    \I__2855\ : CascadeMux
    port map (
            O => \N__16859\,
            I => \eeprom.n2815_cascade_\
        );

    \I__2854\ : InMux
    port map (
            O => \N__16856\,
            I => \N__16852\
        );

    \I__2853\ : CascadeMux
    port map (
            O => \N__16855\,
            I => \N__16849\
        );

    \I__2852\ : LocalMux
    port map (
            O => \N__16852\,
            I => \N__16846\
        );

    \I__2851\ : InMux
    port map (
            O => \N__16849\,
            I => \N__16843\
        );

    \I__2850\ : Span4Mux_h
    port map (
            O => \N__16846\,
            I => \N__16839\
        );

    \I__2849\ : LocalMux
    port map (
            O => \N__16843\,
            I => \N__16836\
        );

    \I__2848\ : InMux
    port map (
            O => \N__16842\,
            I => \N__16833\
        );

    \I__2847\ : Odrv4
    port map (
            O => \N__16839\,
            I => \eeprom.n2614\
        );

    \I__2846\ : Odrv4
    port map (
            O => \N__16836\,
            I => \eeprom.n2614\
        );

    \I__2845\ : LocalMux
    port map (
            O => \N__16833\,
            I => \eeprom.n2614\
        );

    \I__2844\ : InMux
    port map (
            O => \N__16826\,
            I => \N__16823\
        );

    \I__2843\ : LocalMux
    port map (
            O => \N__16823\,
            I => \eeprom.n2681\
        );

    \I__2842\ : CascadeMux
    port map (
            O => \N__16820\,
            I => \eeprom.n2713_cascade_\
        );

    \I__2841\ : CascadeMux
    port map (
            O => \N__16817\,
            I => \eeprom.n4695_cascade_\
        );

    \I__2840\ : CascadeMux
    port map (
            O => \N__16814\,
            I => \eeprom.n16_adj_416_cascade_\
        );

    \I__2839\ : CascadeMux
    port map (
            O => \N__16811\,
            I => \N__16806\
        );

    \I__2838\ : InMux
    port map (
            O => \N__16810\,
            I => \N__16803\
        );

    \I__2837\ : InMux
    port map (
            O => \N__16809\,
            I => \N__16800\
        );

    \I__2836\ : InMux
    port map (
            O => \N__16806\,
            I => \N__16797\
        );

    \I__2835\ : LocalMux
    port map (
            O => \N__16803\,
            I => \eeprom.n2618\
        );

    \I__2834\ : LocalMux
    port map (
            O => \N__16800\,
            I => \eeprom.n2618\
        );

    \I__2833\ : LocalMux
    port map (
            O => \N__16797\,
            I => \eeprom.n2618\
        );

    \I__2832\ : CascadeMux
    port map (
            O => \N__16790\,
            I => \N__16787\
        );

    \I__2831\ : InMux
    port map (
            O => \N__16787\,
            I => \N__16784\
        );

    \I__2830\ : LocalMux
    port map (
            O => \N__16784\,
            I => \eeprom.n2685\
        );

    \I__2829\ : InMux
    port map (
            O => \N__16781\,
            I => \N__16778\
        );

    \I__2828\ : LocalMux
    port map (
            O => \N__16778\,
            I => \eeprom.n2674\
        );

    \I__2827\ : InMux
    port map (
            O => \N__16775\,
            I => \N__16772\
        );

    \I__2826\ : LocalMux
    port map (
            O => \N__16772\,
            I => \N__16769\
        );

    \I__2825\ : Span4Mux_h
    port map (
            O => \N__16769\,
            I => \N__16766\
        );

    \I__2824\ : Odrv4
    port map (
            O => \N__16766\,
            I => \eeprom.n2686\
        );

    \I__2823\ : InMux
    port map (
            O => \N__16763\,
            I => \N__16758\
        );

    \I__2822\ : InMux
    port map (
            O => \N__16762\,
            I => \N__16755\
        );

    \I__2821\ : InMux
    port map (
            O => \N__16761\,
            I => \N__16752\
        );

    \I__2820\ : LocalMux
    port map (
            O => \N__16758\,
            I => \N__16747\
        );

    \I__2819\ : LocalMux
    port map (
            O => \N__16755\,
            I => \N__16747\
        );

    \I__2818\ : LocalMux
    port map (
            O => \N__16752\,
            I => \N__16744\
        );

    \I__2817\ : Span4Mux_h
    port map (
            O => \N__16747\,
            I => \N__16741\
        );

    \I__2816\ : Odrv4
    port map (
            O => \N__16744\,
            I => \eeprom.n2619\
        );

    \I__2815\ : Odrv4
    port map (
            O => \N__16741\,
            I => \eeprom.n2619\
        );

    \I__2814\ : CascadeMux
    port map (
            O => \N__16736\,
            I => \eeprom.n2718_cascade_\
        );

    \I__2813\ : InMux
    port map (
            O => \N__16733\,
            I => \N__16730\
        );

    \I__2812\ : LocalMux
    port map (
            O => \N__16730\,
            I => \eeprom.n4699\
        );

    \I__2811\ : CascadeMux
    port map (
            O => \N__16727\,
            I => \N__16724\
        );

    \I__2810\ : InMux
    port map (
            O => \N__16724\,
            I => \N__16721\
        );

    \I__2809\ : LocalMux
    port map (
            O => \N__16721\,
            I => \N__16718\
        );

    \I__2808\ : Span4Mux_h
    port map (
            O => \N__16718\,
            I => \N__16715\
        );

    \I__2807\ : Odrv4
    port map (
            O => \N__16715\,
            I => \eeprom.n2280\
        );

    \I__2806\ : InMux
    port map (
            O => \N__16712\,
            I => \eeprom.n3546\
        );

    \I__2805\ : CascadeMux
    port map (
            O => \N__16709\,
            I => \N__16704\
        );

    \I__2804\ : InMux
    port map (
            O => \N__16708\,
            I => \N__16701\
        );

    \I__2803\ : InMux
    port map (
            O => \N__16707\,
            I => \N__16698\
        );

    \I__2802\ : InMux
    port map (
            O => \N__16704\,
            I => \N__16695\
        );

    \I__2801\ : LocalMux
    port map (
            O => \N__16701\,
            I => \N__16692\
        );

    \I__2800\ : LocalMux
    port map (
            O => \N__16698\,
            I => \eeprom.n2212\
        );

    \I__2799\ : LocalMux
    port map (
            O => \N__16695\,
            I => \eeprom.n2212\
        );

    \I__2798\ : Odrv4
    port map (
            O => \N__16692\,
            I => \eeprom.n2212\
        );

    \I__2797\ : InMux
    port map (
            O => \N__16685\,
            I => \N__16682\
        );

    \I__2796\ : LocalMux
    port map (
            O => \N__16682\,
            I => \eeprom.n2279\
        );

    \I__2795\ : InMux
    port map (
            O => \N__16679\,
            I => \eeprom.n3547\
        );

    \I__2794\ : CascadeMux
    port map (
            O => \N__16676\,
            I => \N__16671\
        );

    \I__2793\ : InMux
    port map (
            O => \N__16675\,
            I => \N__16666\
        );

    \I__2792\ : InMux
    port map (
            O => \N__16674\,
            I => \N__16666\
        );

    \I__2791\ : InMux
    port map (
            O => \N__16671\,
            I => \N__16663\
        );

    \I__2790\ : LocalMux
    port map (
            O => \N__16666\,
            I => \N__16660\
        );

    \I__2789\ : LocalMux
    port map (
            O => \N__16663\,
            I => \eeprom.n2211\
        );

    \I__2788\ : Odrv4
    port map (
            O => \N__16660\,
            I => \eeprom.n2211\
        );

    \I__2787\ : CascadeMux
    port map (
            O => \N__16655\,
            I => \N__16652\
        );

    \I__2786\ : InMux
    port map (
            O => \N__16652\,
            I => \N__16649\
        );

    \I__2785\ : LocalMux
    port map (
            O => \N__16649\,
            I => \N__16646\
        );

    \I__2784\ : Span4Mux_h
    port map (
            O => \N__16646\,
            I => \N__16643\
        );

    \I__2783\ : Odrv4
    port map (
            O => \N__16643\,
            I => \eeprom.n2278\
        );

    \I__2782\ : InMux
    port map (
            O => \N__16640\,
            I => \bfn_6_27_0_\
        );

    \I__2781\ : InMux
    port map (
            O => \N__16637\,
            I => \N__16633\
        );

    \I__2780\ : CascadeMux
    port map (
            O => \N__16636\,
            I => \N__16630\
        );

    \I__2779\ : LocalMux
    port map (
            O => \N__16633\,
            I => \N__16626\
        );

    \I__2778\ : InMux
    port map (
            O => \N__16630\,
            I => \N__16621\
        );

    \I__2777\ : InMux
    port map (
            O => \N__16629\,
            I => \N__16621\
        );

    \I__2776\ : Odrv4
    port map (
            O => \N__16626\,
            I => \eeprom.n2210\
        );

    \I__2775\ : LocalMux
    port map (
            O => \N__16621\,
            I => \eeprom.n2210\
        );

    \I__2774\ : InMux
    port map (
            O => \N__16616\,
            I => \N__16613\
        );

    \I__2773\ : LocalMux
    port map (
            O => \N__16613\,
            I => \N__16610\
        );

    \I__2772\ : Odrv4
    port map (
            O => \N__16610\,
            I => \eeprom.n2277\
        );

    \I__2771\ : InMux
    port map (
            O => \N__16607\,
            I => \eeprom.n3549\
        );

    \I__2770\ : InMux
    port map (
            O => \N__16604\,
            I => \N__16594\
        );

    \I__2769\ : InMux
    port map (
            O => \N__16603\,
            I => \N__16588\
        );

    \I__2768\ : InMux
    port map (
            O => \N__16602\,
            I => \N__16583\
        );

    \I__2767\ : InMux
    port map (
            O => \N__16601\,
            I => \N__16583\
        );

    \I__2766\ : InMux
    port map (
            O => \N__16600\,
            I => \N__16580\
        );

    \I__2765\ : InMux
    port map (
            O => \N__16599\,
            I => \N__16575\
        );

    \I__2764\ : InMux
    port map (
            O => \N__16598\,
            I => \N__16575\
        );

    \I__2763\ : InMux
    port map (
            O => \N__16597\,
            I => \N__16572\
        );

    \I__2762\ : LocalMux
    port map (
            O => \N__16594\,
            I => \N__16569\
        );

    \I__2761\ : InMux
    port map (
            O => \N__16593\,
            I => \N__16562\
        );

    \I__2760\ : InMux
    port map (
            O => \N__16592\,
            I => \N__16562\
        );

    \I__2759\ : InMux
    port map (
            O => \N__16591\,
            I => \N__16562\
        );

    \I__2758\ : LocalMux
    port map (
            O => \N__16588\,
            I => \eeprom.n2242\
        );

    \I__2757\ : LocalMux
    port map (
            O => \N__16583\,
            I => \eeprom.n2242\
        );

    \I__2756\ : LocalMux
    port map (
            O => \N__16580\,
            I => \eeprom.n2242\
        );

    \I__2755\ : LocalMux
    port map (
            O => \N__16575\,
            I => \eeprom.n2242\
        );

    \I__2754\ : LocalMux
    port map (
            O => \N__16572\,
            I => \eeprom.n2242\
        );

    \I__2753\ : Odrv4
    port map (
            O => \N__16569\,
            I => \eeprom.n2242\
        );

    \I__2752\ : LocalMux
    port map (
            O => \N__16562\,
            I => \eeprom.n2242\
        );

    \I__2751\ : InMux
    port map (
            O => \N__16547\,
            I => \N__16543\
        );

    \I__2750\ : CascadeMux
    port map (
            O => \N__16546\,
            I => \N__16540\
        );

    \I__2749\ : LocalMux
    port map (
            O => \N__16543\,
            I => \N__16537\
        );

    \I__2748\ : InMux
    port map (
            O => \N__16540\,
            I => \N__16534\
        );

    \I__2747\ : Span4Mux_h
    port map (
            O => \N__16537\,
            I => \N__16531\
        );

    \I__2746\ : LocalMux
    port map (
            O => \N__16534\,
            I => \eeprom.n2209\
        );

    \I__2745\ : Odrv4
    port map (
            O => \N__16531\,
            I => \eeprom.n2209\
        );

    \I__2744\ : InMux
    port map (
            O => \N__16526\,
            I => \eeprom.n3550\
        );

    \I__2743\ : InMux
    port map (
            O => \N__16523\,
            I => \N__16519\
        );

    \I__2742\ : InMux
    port map (
            O => \N__16522\,
            I => \N__16516\
        );

    \I__2741\ : LocalMux
    port map (
            O => \N__16519\,
            I => \N__16513\
        );

    \I__2740\ : LocalMux
    port map (
            O => \N__16516\,
            I => \N__16510\
        );

    \I__2739\ : Span4Mux_h
    port map (
            O => \N__16513\,
            I => \N__16507\
        );

    \I__2738\ : Span4Mux_h
    port map (
            O => \N__16510\,
            I => \N__16504\
        );

    \I__2737\ : Odrv4
    port map (
            O => \N__16507\,
            I => \eeprom.n2308\
        );

    \I__2736\ : Odrv4
    port map (
            O => \N__16504\,
            I => \eeprom.n2308\
        );

    \I__2735\ : InMux
    port map (
            O => \N__16499\,
            I => \N__16495\
        );

    \I__2734\ : CascadeMux
    port map (
            O => \N__16498\,
            I => \N__16492\
        );

    \I__2733\ : LocalMux
    port map (
            O => \N__16495\,
            I => \N__16489\
        );

    \I__2732\ : InMux
    port map (
            O => \N__16492\,
            I => \N__16486\
        );

    \I__2731\ : Span4Mux_v
    port map (
            O => \N__16489\,
            I => \N__16482\
        );

    \I__2730\ : LocalMux
    port map (
            O => \N__16486\,
            I => \N__16479\
        );

    \I__2729\ : InMux
    port map (
            O => \N__16485\,
            I => \N__16476\
        );

    \I__2728\ : Odrv4
    port map (
            O => \N__16482\,
            I => \eeprom.n2612\
        );

    \I__2727\ : Odrv12
    port map (
            O => \N__16479\,
            I => \eeprom.n2612\
        );

    \I__2726\ : LocalMux
    port map (
            O => \N__16476\,
            I => \eeprom.n2612\
        );

    \I__2725\ : CascadeMux
    port map (
            O => \N__16469\,
            I => \N__16466\
        );

    \I__2724\ : InMux
    port map (
            O => \N__16466\,
            I => \N__16463\
        );

    \I__2723\ : LocalMux
    port map (
            O => \N__16463\,
            I => \eeprom.n2679\
        );

    \I__2722\ : InMux
    port map (
            O => \N__16460\,
            I => \N__16457\
        );

    \I__2721\ : LocalMux
    port map (
            O => \N__16457\,
            I => \N__16453\
        );

    \I__2720\ : InMux
    port map (
            O => \N__16456\,
            I => \N__16450\
        );

    \I__2719\ : Span4Mux_v
    port map (
            O => \N__16453\,
            I => \N__16447\
        );

    \I__2718\ : LocalMux
    port map (
            O => \N__16450\,
            I => \N__16444\
        );

    \I__2717\ : Odrv4
    port map (
            O => \N__16447\,
            I => \eeprom.n2606\
        );

    \I__2716\ : Odrv12
    port map (
            O => \N__16444\,
            I => \eeprom.n2606\
        );

    \I__2715\ : InMux
    port map (
            O => \N__16439\,
            I => \N__16436\
        );

    \I__2714\ : LocalMux
    port map (
            O => \N__16436\,
            I => \eeprom.n2673\
        );

    \I__2713\ : InMux
    port map (
            O => \N__16433\,
            I => \N__16430\
        );

    \I__2712\ : LocalMux
    port map (
            O => \N__16430\,
            I => \eeprom.n2680\
        );

    \I__2711\ : InMux
    port map (
            O => \N__16427\,
            I => \N__16423\
        );

    \I__2710\ : CascadeMux
    port map (
            O => \N__16426\,
            I => \N__16420\
        );

    \I__2709\ : LocalMux
    port map (
            O => \N__16423\,
            I => \N__16417\
        );

    \I__2708\ : InMux
    port map (
            O => \N__16420\,
            I => \N__16414\
        );

    \I__2707\ : Span4Mux_v
    port map (
            O => \N__16417\,
            I => \N__16410\
        );

    \I__2706\ : LocalMux
    port map (
            O => \N__16414\,
            I => \N__16407\
        );

    \I__2705\ : InMux
    port map (
            O => \N__16413\,
            I => \N__16404\
        );

    \I__2704\ : Odrv4
    port map (
            O => \N__16410\,
            I => \eeprom.n2613\
        );

    \I__2703\ : Odrv4
    port map (
            O => \N__16407\,
            I => \eeprom.n2613\
        );

    \I__2702\ : LocalMux
    port map (
            O => \N__16404\,
            I => \eeprom.n2613\
        );

    \I__2701\ : CascadeMux
    port map (
            O => \N__16397\,
            I => \N__16393\
        );

    \I__2700\ : InMux
    port map (
            O => \N__16396\,
            I => \N__16390\
        );

    \I__2699\ : InMux
    port map (
            O => \N__16393\,
            I => \N__16387\
        );

    \I__2698\ : LocalMux
    port map (
            O => \N__16390\,
            I => \N__16383\
        );

    \I__2697\ : LocalMux
    port map (
            O => \N__16387\,
            I => \N__16380\
        );

    \I__2696\ : InMux
    port map (
            O => \N__16386\,
            I => \N__16377\
        );

    \I__2695\ : Odrv4
    port map (
            O => \N__16383\,
            I => \eeprom.n2113\
        );

    \I__2694\ : Odrv12
    port map (
            O => \N__16380\,
            I => \eeprom.n2113\
        );

    \I__2693\ : LocalMux
    port map (
            O => \N__16377\,
            I => \eeprom.n2113\
        );

    \I__2692\ : CascadeMux
    port map (
            O => \N__16370\,
            I => \N__16361\
        );

    \I__2691\ : InMux
    port map (
            O => \N__16369\,
            I => \N__16358\
        );

    \I__2690\ : CascadeMux
    port map (
            O => \N__16368\,
            I => \N__16355\
        );

    \I__2689\ : CascadeMux
    port map (
            O => \N__16367\,
            I => \N__16350\
        );

    \I__2688\ : CascadeMux
    port map (
            O => \N__16366\,
            I => \N__16347\
        );

    \I__2687\ : CascadeMux
    port map (
            O => \N__16365\,
            I => \N__16343\
        );

    \I__2686\ : CascadeMux
    port map (
            O => \N__16364\,
            I => \N__16340\
        );

    \I__2685\ : InMux
    port map (
            O => \N__16361\,
            I => \N__16336\
        );

    \I__2684\ : LocalMux
    port map (
            O => \N__16358\,
            I => \N__16333\
        );

    \I__2683\ : InMux
    port map (
            O => \N__16355\,
            I => \N__16328\
        );

    \I__2682\ : InMux
    port map (
            O => \N__16354\,
            I => \N__16328\
        );

    \I__2681\ : InMux
    port map (
            O => \N__16353\,
            I => \N__16319\
        );

    \I__2680\ : InMux
    port map (
            O => \N__16350\,
            I => \N__16319\
        );

    \I__2679\ : InMux
    port map (
            O => \N__16347\,
            I => \N__16319\
        );

    \I__2678\ : InMux
    port map (
            O => \N__16346\,
            I => \N__16319\
        );

    \I__2677\ : InMux
    port map (
            O => \N__16343\,
            I => \N__16312\
        );

    \I__2676\ : InMux
    port map (
            O => \N__16340\,
            I => \N__16312\
        );

    \I__2675\ : InMux
    port map (
            O => \N__16339\,
            I => \N__16312\
        );

    \I__2674\ : LocalMux
    port map (
            O => \N__16336\,
            I => \N__16309\
        );

    \I__2673\ : Odrv4
    port map (
            O => \N__16333\,
            I => \eeprom.n2143\
        );

    \I__2672\ : LocalMux
    port map (
            O => \N__16328\,
            I => \eeprom.n2143\
        );

    \I__2671\ : LocalMux
    port map (
            O => \N__16319\,
            I => \eeprom.n2143\
        );

    \I__2670\ : LocalMux
    port map (
            O => \N__16312\,
            I => \eeprom.n2143\
        );

    \I__2669\ : Odrv4
    port map (
            O => \N__16309\,
            I => \eeprom.n2143\
        );

    \I__2668\ : InMux
    port map (
            O => \N__16298\,
            I => \N__16295\
        );

    \I__2667\ : LocalMux
    port map (
            O => \N__16295\,
            I => \N__16292\
        );

    \I__2666\ : Odrv4
    port map (
            O => \N__16292\,
            I => \eeprom.n2180\
        );

    \I__2665\ : InMux
    port map (
            O => \N__16289\,
            I => \N__16285\
        );

    \I__2664\ : InMux
    port map (
            O => \N__16288\,
            I => \N__16282\
        );

    \I__2663\ : LocalMux
    port map (
            O => \N__16285\,
            I => \N__16277\
        );

    \I__2662\ : LocalMux
    port map (
            O => \N__16282\,
            I => \N__16277\
        );

    \I__2661\ : Odrv4
    port map (
            O => \N__16277\,
            I => \eeprom.n2219\
        );

    \I__2660\ : InMux
    port map (
            O => \N__16274\,
            I => \N__16271\
        );

    \I__2659\ : LocalMux
    port map (
            O => \N__16271\,
            I => \N__16268\
        );

    \I__2658\ : Odrv12
    port map (
            O => \N__16268\,
            I => \eeprom.n2286\
        );

    \I__2657\ : InMux
    port map (
            O => \N__16265\,
            I => \bfn_6_26_0_\
        );

    \I__2656\ : CascadeMux
    port map (
            O => \N__16262\,
            I => \N__16259\
        );

    \I__2655\ : InMux
    port map (
            O => \N__16259\,
            I => \N__16255\
        );

    \I__2654\ : InMux
    port map (
            O => \N__16258\,
            I => \N__16252\
        );

    \I__2653\ : LocalMux
    port map (
            O => \N__16255\,
            I => \eeprom.n2218\
        );

    \I__2652\ : LocalMux
    port map (
            O => \N__16252\,
            I => \eeprom.n2218\
        );

    \I__2651\ : InMux
    port map (
            O => \N__16247\,
            I => \N__16244\
        );

    \I__2650\ : LocalMux
    port map (
            O => \N__16244\,
            I => \eeprom.n2285\
        );

    \I__2649\ : InMux
    port map (
            O => \N__16241\,
            I => \eeprom.n3541\
        );

    \I__2648\ : CascadeMux
    port map (
            O => \N__16238\,
            I => \N__16234\
        );

    \I__2647\ : CascadeMux
    port map (
            O => \N__16237\,
            I => \N__16231\
        );

    \I__2646\ : InMux
    port map (
            O => \N__16234\,
            I => \N__16227\
        );

    \I__2645\ : InMux
    port map (
            O => \N__16231\,
            I => \N__16224\
        );

    \I__2644\ : InMux
    port map (
            O => \N__16230\,
            I => \N__16221\
        );

    \I__2643\ : LocalMux
    port map (
            O => \N__16227\,
            I => \eeprom.n2217\
        );

    \I__2642\ : LocalMux
    port map (
            O => \N__16224\,
            I => \eeprom.n2217\
        );

    \I__2641\ : LocalMux
    port map (
            O => \N__16221\,
            I => \eeprom.n2217\
        );

    \I__2640\ : InMux
    port map (
            O => \N__16214\,
            I => \N__16211\
        );

    \I__2639\ : LocalMux
    port map (
            O => \N__16211\,
            I => \eeprom.n2284\
        );

    \I__2638\ : InMux
    port map (
            O => \N__16208\,
            I => \eeprom.n3542\
        );

    \I__2637\ : CascadeMux
    port map (
            O => \N__16205\,
            I => \N__16200\
        );

    \I__2636\ : CascadeMux
    port map (
            O => \N__16204\,
            I => \N__16197\
        );

    \I__2635\ : InMux
    port map (
            O => \N__16203\,
            I => \N__16194\
        );

    \I__2634\ : InMux
    port map (
            O => \N__16200\,
            I => \N__16191\
        );

    \I__2633\ : InMux
    port map (
            O => \N__16197\,
            I => \N__16188\
        );

    \I__2632\ : LocalMux
    port map (
            O => \N__16194\,
            I => \eeprom.n2216\
        );

    \I__2631\ : LocalMux
    port map (
            O => \N__16191\,
            I => \eeprom.n2216\
        );

    \I__2630\ : LocalMux
    port map (
            O => \N__16188\,
            I => \eeprom.n2216\
        );

    \I__2629\ : CascadeMux
    port map (
            O => \N__16181\,
            I => \N__16178\
        );

    \I__2628\ : InMux
    port map (
            O => \N__16178\,
            I => \N__16175\
        );

    \I__2627\ : LocalMux
    port map (
            O => \N__16175\,
            I => \eeprom.n2283\
        );

    \I__2626\ : InMux
    port map (
            O => \N__16172\,
            I => \eeprom.n3543\
        );

    \I__2625\ : CascadeMux
    port map (
            O => \N__16169\,
            I => \N__16166\
        );

    \I__2624\ : InMux
    port map (
            O => \N__16166\,
            I => \N__16162\
        );

    \I__2623\ : InMux
    port map (
            O => \N__16165\,
            I => \N__16159\
        );

    \I__2622\ : LocalMux
    port map (
            O => \N__16162\,
            I => \eeprom.n2215\
        );

    \I__2621\ : LocalMux
    port map (
            O => \N__16159\,
            I => \eeprom.n2215\
        );

    \I__2620\ : CascadeMux
    port map (
            O => \N__16154\,
            I => \N__16151\
        );

    \I__2619\ : InMux
    port map (
            O => \N__16151\,
            I => \N__16148\
        );

    \I__2618\ : LocalMux
    port map (
            O => \N__16148\,
            I => \N__16145\
        );

    \I__2617\ : Odrv4
    port map (
            O => \N__16145\,
            I => \eeprom.n2282\
        );

    \I__2616\ : InMux
    port map (
            O => \N__16142\,
            I => \eeprom.n3544\
        );

    \I__2615\ : CascadeMux
    port map (
            O => \N__16139\,
            I => \N__16136\
        );

    \I__2614\ : InMux
    port map (
            O => \N__16136\,
            I => \N__16132\
        );

    \I__2613\ : InMux
    port map (
            O => \N__16135\,
            I => \N__16129\
        );

    \I__2612\ : LocalMux
    port map (
            O => \N__16132\,
            I => \eeprom.n2214\
        );

    \I__2611\ : LocalMux
    port map (
            O => \N__16129\,
            I => \eeprom.n2214\
        );

    \I__2610\ : InMux
    port map (
            O => \N__16124\,
            I => \N__16121\
        );

    \I__2609\ : LocalMux
    port map (
            O => \N__16121\,
            I => \eeprom.n2281\
        );

    \I__2608\ : InMux
    port map (
            O => \N__16118\,
            I => \eeprom.n3545\
        );

    \I__2607\ : InMux
    port map (
            O => \N__16115\,
            I => \N__16111\
        );

    \I__2606\ : CascadeMux
    port map (
            O => \N__16114\,
            I => \N__16108\
        );

    \I__2605\ : LocalMux
    port map (
            O => \N__16111\,
            I => \N__16104\
        );

    \I__2604\ : InMux
    port map (
            O => \N__16108\,
            I => \N__16101\
        );

    \I__2603\ : InMux
    port map (
            O => \N__16107\,
            I => \N__16098\
        );

    \I__2602\ : Odrv4
    port map (
            O => \N__16104\,
            I => \eeprom.n2213\
        );

    \I__2601\ : LocalMux
    port map (
            O => \N__16101\,
            I => \eeprom.n2213\
        );

    \I__2600\ : LocalMux
    port map (
            O => \N__16098\,
            I => \eeprom.n2213\
        );

    \I__2599\ : InMux
    port map (
            O => \N__16091\,
            I => \N__16087\
        );

    \I__2598\ : CascadeMux
    port map (
            O => \N__16090\,
            I => \N__16084\
        );

    \I__2597\ : LocalMux
    port map (
            O => \N__16087\,
            I => \N__16080\
        );

    \I__2596\ : InMux
    port map (
            O => \N__16084\,
            I => \N__16077\
        );

    \I__2595\ : InMux
    port map (
            O => \N__16083\,
            I => \N__16074\
        );

    \I__2594\ : Odrv12
    port map (
            O => \N__16080\,
            I => \eeprom.n2413\
        );

    \I__2593\ : LocalMux
    port map (
            O => \N__16077\,
            I => \eeprom.n2413\
        );

    \I__2592\ : LocalMux
    port map (
            O => \N__16074\,
            I => \eeprom.n2413\
        );

    \I__2591\ : CascadeMux
    port map (
            O => \N__16067\,
            I => \N__16064\
        );

    \I__2590\ : InMux
    port map (
            O => \N__16064\,
            I => \N__16061\
        );

    \I__2589\ : LocalMux
    port map (
            O => \N__16061\,
            I => \N__16058\
        );

    \I__2588\ : Span4Mux_h
    port map (
            O => \N__16058\,
            I => \N__16055\
        );

    \I__2587\ : Odrv4
    port map (
            O => \N__16055\,
            I => \eeprom.n2480\
        );

    \I__2586\ : InMux
    port map (
            O => \N__16052\,
            I => \N__16047\
        );

    \I__2585\ : CascadeMux
    port map (
            O => \N__16051\,
            I => \N__16044\
        );

    \I__2584\ : InMux
    port map (
            O => \N__16050\,
            I => \N__16041\
        );

    \I__2583\ : LocalMux
    port map (
            O => \N__16047\,
            I => \N__16038\
        );

    \I__2582\ : InMux
    port map (
            O => \N__16044\,
            I => \N__16035\
        );

    \I__2581\ : LocalMux
    port map (
            O => \N__16041\,
            I => \N__16032\
        );

    \I__2580\ : Span4Mux_h
    port map (
            O => \N__16038\,
            I => \N__16025\
        );

    \I__2579\ : LocalMux
    port map (
            O => \N__16035\,
            I => \N__16025\
        );

    \I__2578\ : Span4Mux_h
    port map (
            O => \N__16032\,
            I => \N__16025\
        );

    \I__2577\ : Odrv4
    port map (
            O => \N__16025\,
            I => \eeprom.n2512\
        );

    \I__2576\ : InMux
    port map (
            O => \N__16022\,
            I => \N__16018\
        );

    \I__2575\ : InMux
    port map (
            O => \N__16021\,
            I => \N__16015\
        );

    \I__2574\ : LocalMux
    port map (
            O => \N__16018\,
            I => \N__16011\
        );

    \I__2573\ : LocalMux
    port map (
            O => \N__16015\,
            I => \N__16008\
        );

    \I__2572\ : InMux
    port map (
            O => \N__16014\,
            I => \N__16005\
        );

    \I__2571\ : Odrv12
    port map (
            O => \N__16011\,
            I => \eeprom.n2408\
        );

    \I__2570\ : Odrv4
    port map (
            O => \N__16008\,
            I => \eeprom.n2408\
        );

    \I__2569\ : LocalMux
    port map (
            O => \N__16005\,
            I => \eeprom.n2408\
        );

    \I__2568\ : CascadeMux
    port map (
            O => \N__15998\,
            I => \N__15995\
        );

    \I__2567\ : InMux
    port map (
            O => \N__15995\,
            I => \N__15992\
        );

    \I__2566\ : LocalMux
    port map (
            O => \N__15992\,
            I => \N__15989\
        );

    \I__2565\ : Span4Mux_v
    port map (
            O => \N__15989\,
            I => \N__15986\
        );

    \I__2564\ : Odrv4
    port map (
            O => \N__15986\,
            I => \eeprom.n2475\
        );

    \I__2563\ : CascadeMux
    port map (
            O => \N__15983\,
            I => \N__15979\
        );

    \I__2562\ : InMux
    port map (
            O => \N__15982\,
            I => \N__15974\
        );

    \I__2561\ : InMux
    port map (
            O => \N__15979\,
            I => \N__15967\
        );

    \I__2560\ : InMux
    port map (
            O => \N__15978\,
            I => \N__15967\
        );

    \I__2559\ : CascadeMux
    port map (
            O => \N__15977\,
            I => \N__15964\
        );

    \I__2558\ : LocalMux
    port map (
            O => \N__15974\,
            I => \N__15956\
        );

    \I__2557\ : InMux
    port map (
            O => \N__15973\,
            I => \N__15951\
        );

    \I__2556\ : InMux
    port map (
            O => \N__15972\,
            I => \N__15951\
        );

    \I__2555\ : LocalMux
    port map (
            O => \N__15967\,
            I => \N__15948\
        );

    \I__2554\ : InMux
    port map (
            O => \N__15964\,
            I => \N__15941\
        );

    \I__2553\ : InMux
    port map (
            O => \N__15963\,
            I => \N__15941\
        );

    \I__2552\ : InMux
    port map (
            O => \N__15962\,
            I => \N__15941\
        );

    \I__2551\ : InMux
    port map (
            O => \N__15961\,
            I => \N__15936\
        );

    \I__2550\ : InMux
    port map (
            O => \N__15960\,
            I => \N__15936\
        );

    \I__2549\ : CascadeMux
    port map (
            O => \N__15959\,
            I => \N__15932\
        );

    \I__2548\ : Span4Mux_h
    port map (
            O => \N__15956\,
            I => \N__15928\
        );

    \I__2547\ : LocalMux
    port map (
            O => \N__15951\,
            I => \N__15925\
        );

    \I__2546\ : Span4Mux_v
    port map (
            O => \N__15948\,
            I => \N__15920\
        );

    \I__2545\ : LocalMux
    port map (
            O => \N__15941\,
            I => \N__15920\
        );

    \I__2544\ : LocalMux
    port map (
            O => \N__15936\,
            I => \N__15917\
        );

    \I__2543\ : InMux
    port map (
            O => \N__15935\,
            I => \N__15910\
        );

    \I__2542\ : InMux
    port map (
            O => \N__15932\,
            I => \N__15910\
        );

    \I__2541\ : InMux
    port map (
            O => \N__15931\,
            I => \N__15910\
        );

    \I__2540\ : Odrv4
    port map (
            O => \N__15928\,
            I => \eeprom.n2440\
        );

    \I__2539\ : Odrv4
    port map (
            O => \N__15925\,
            I => \eeprom.n2440\
        );

    \I__2538\ : Odrv4
    port map (
            O => \N__15920\,
            I => \eeprom.n2440\
        );

    \I__2537\ : Odrv4
    port map (
            O => \N__15917\,
            I => \eeprom.n2440\
        );

    \I__2536\ : LocalMux
    port map (
            O => \N__15910\,
            I => \eeprom.n2440\
        );

    \I__2535\ : InMux
    port map (
            O => \N__15899\,
            I => \N__15894\
        );

    \I__2534\ : InMux
    port map (
            O => \N__15898\,
            I => \N__15891\
        );

    \I__2533\ : InMux
    port map (
            O => \N__15897\,
            I => \N__15888\
        );

    \I__2532\ : LocalMux
    port map (
            O => \N__15894\,
            I => \N__15885\
        );

    \I__2531\ : LocalMux
    port map (
            O => \N__15891\,
            I => \N__15878\
        );

    \I__2530\ : LocalMux
    port map (
            O => \N__15888\,
            I => \N__15878\
        );

    \I__2529\ : Span4Mux_h
    port map (
            O => \N__15885\,
            I => \N__15878\
        );

    \I__2528\ : Odrv4
    port map (
            O => \N__15878\,
            I => \eeprom.n2507\
        );

    \I__2527\ : InMux
    port map (
            O => \N__15875\,
            I => \N__15872\
        );

    \I__2526\ : LocalMux
    port map (
            O => \N__15872\,
            I => \eeprom.n4801\
        );

    \I__2525\ : InMux
    port map (
            O => \N__15869\,
            I => \N__15865\
        );

    \I__2524\ : CascadeMux
    port map (
            O => \N__15868\,
            I => \N__15862\
        );

    \I__2523\ : LocalMux
    port map (
            O => \N__15865\,
            I => \N__15859\
        );

    \I__2522\ : InMux
    port map (
            O => \N__15862\,
            I => \N__15855\
        );

    \I__2521\ : Span4Mux_v
    port map (
            O => \N__15859\,
            I => \N__15852\
        );

    \I__2520\ : InMux
    port map (
            O => \N__15858\,
            I => \N__15849\
        );

    \I__2519\ : LocalMux
    port map (
            O => \N__15855\,
            I => \N__15846\
        );

    \I__2518\ : Odrv4
    port map (
            O => \N__15852\,
            I => \eeprom.n2017\
        );

    \I__2517\ : LocalMux
    port map (
            O => \N__15849\,
            I => \eeprom.n2017\
        );

    \I__2516\ : Odrv4
    port map (
            O => \N__15846\,
            I => \eeprom.n2017\
        );

    \I__2515\ : CascadeMux
    port map (
            O => \N__15839\,
            I => \eeprom.n4799_cascade_\
        );

    \I__2514\ : InMux
    port map (
            O => \N__15836\,
            I => \N__15833\
        );

    \I__2513\ : LocalMux
    port map (
            O => \N__15833\,
            I => \eeprom.n4872\
        );

    \I__2512\ : CascadeMux
    port map (
            O => \N__15830\,
            I => \N__15826\
        );

    \I__2511\ : CascadeMux
    port map (
            O => \N__15829\,
            I => \N__15823\
        );

    \I__2510\ : InMux
    port map (
            O => \N__15826\,
            I => \N__15820\
        );

    \I__2509\ : InMux
    port map (
            O => \N__15823\,
            I => \N__15816\
        );

    \I__2508\ : LocalMux
    port map (
            O => \N__15820\,
            I => \N__15813\
        );

    \I__2507\ : CascadeMux
    port map (
            O => \N__15819\,
            I => \N__15810\
        );

    \I__2506\ : LocalMux
    port map (
            O => \N__15816\,
            I => \N__15807\
        );

    \I__2505\ : Span4Mux_h
    port map (
            O => \N__15813\,
            I => \N__15804\
        );

    \I__2504\ : InMux
    port map (
            O => \N__15810\,
            I => \N__15801\
        );

    \I__2503\ : Odrv4
    port map (
            O => \N__15807\,
            I => \eeprom.n2314\
        );

    \I__2502\ : Odrv4
    port map (
            O => \N__15804\,
            I => \eeprom.n2314\
        );

    \I__2501\ : LocalMux
    port map (
            O => \N__15801\,
            I => \eeprom.n2314\
        );

    \I__2500\ : CascadeMux
    port map (
            O => \N__15794\,
            I => \N__15790\
        );

    \I__2499\ : InMux
    port map (
            O => \N__15793\,
            I => \N__15787\
        );

    \I__2498\ : InMux
    port map (
            O => \N__15790\,
            I => \N__15784\
        );

    \I__2497\ : LocalMux
    port map (
            O => \N__15787\,
            I => \N__15781\
        );

    \I__2496\ : LocalMux
    port map (
            O => \N__15784\,
            I => \N__15777\
        );

    \I__2495\ : Span4Mux_h
    port map (
            O => \N__15781\,
            I => \N__15774\
        );

    \I__2494\ : InMux
    port map (
            O => \N__15780\,
            I => \N__15771\
        );

    \I__2493\ : Span4Mux_h
    port map (
            O => \N__15777\,
            I => \N__15768\
        );

    \I__2492\ : Odrv4
    port map (
            O => \N__15774\,
            I => \eeprom.n2316\
        );

    \I__2491\ : LocalMux
    port map (
            O => \N__15771\,
            I => \eeprom.n2316\
        );

    \I__2490\ : Odrv4
    port map (
            O => \N__15768\,
            I => \eeprom.n2316\
        );

    \I__2489\ : InMux
    port map (
            O => \N__15761\,
            I => \N__15758\
        );

    \I__2488\ : LocalMux
    port map (
            O => \N__15758\,
            I => \N__15755\
        );

    \I__2487\ : Odrv4
    port map (
            O => \N__15755\,
            I => \eeprom.n2186\
        );

    \I__2486\ : InMux
    port map (
            O => \N__15752\,
            I => \N__15747\
        );

    \I__2485\ : InMux
    port map (
            O => \N__15751\,
            I => \N__15744\
        );

    \I__2484\ : InMux
    port map (
            O => \N__15750\,
            I => \N__15741\
        );

    \I__2483\ : LocalMux
    port map (
            O => \N__15747\,
            I => \N__15738\
        );

    \I__2482\ : LocalMux
    port map (
            O => \N__15744\,
            I => \eeprom.n2119\
        );

    \I__2481\ : LocalMux
    port map (
            O => \N__15741\,
            I => \eeprom.n2119\
        );

    \I__2480\ : Odrv4
    port map (
            O => \N__15738\,
            I => \eeprom.n2119\
        );

    \I__2479\ : CascadeMux
    port map (
            O => \N__15731\,
            I => \eeprom.n2218_cascade_\
        );

    \I__2478\ : CascadeMux
    port map (
            O => \N__15728\,
            I => \N__15724\
        );

    \I__2477\ : InMux
    port map (
            O => \N__15727\,
            I => \N__15721\
        );

    \I__2476\ : InMux
    port map (
            O => \N__15724\,
            I => \N__15718\
        );

    \I__2475\ : LocalMux
    port map (
            O => \N__15721\,
            I => \N__15712\
        );

    \I__2474\ : LocalMux
    port map (
            O => \N__15718\,
            I => \N__15712\
        );

    \I__2473\ : InMux
    port map (
            O => \N__15717\,
            I => \N__15709\
        );

    \I__2472\ : Span4Mux_v
    port map (
            O => \N__15712\,
            I => \N__15706\
        );

    \I__2471\ : LocalMux
    port map (
            O => \N__15709\,
            I => \eeprom.n2317\
        );

    \I__2470\ : Odrv4
    port map (
            O => \N__15706\,
            I => \eeprom.n2317\
        );

    \I__2469\ : CascadeMux
    port map (
            O => \N__15701\,
            I => \eeprom.n4447_cascade_\
        );

    \I__2468\ : InMux
    port map (
            O => \N__15698\,
            I => \N__15695\
        );

    \I__2467\ : LocalMux
    port map (
            O => \N__15695\,
            I => \eeprom.n4218\
        );

    \I__2466\ : InMux
    port map (
            O => \N__15692\,
            I => \N__15689\
        );

    \I__2465\ : LocalMux
    port map (
            O => \N__15689\,
            I => \N__15686\
        );

    \I__2464\ : Span4Mux_h
    port map (
            O => \N__15686\,
            I => \N__15681\
        );

    \I__2463\ : InMux
    port map (
            O => \N__15685\,
            I => \N__15678\
        );

    \I__2462\ : InMux
    port map (
            O => \N__15684\,
            I => \N__15675\
        );

    \I__2461\ : Odrv4
    port map (
            O => \N__15681\,
            I => \eeprom.n2412\
        );

    \I__2460\ : LocalMux
    port map (
            O => \N__15678\,
            I => \eeprom.n2412\
        );

    \I__2459\ : LocalMux
    port map (
            O => \N__15675\,
            I => \eeprom.n2412\
        );

    \I__2458\ : CascadeMux
    port map (
            O => \N__15668\,
            I => \N__15665\
        );

    \I__2457\ : InMux
    port map (
            O => \N__15665\,
            I => \N__15662\
        );

    \I__2456\ : LocalMux
    port map (
            O => \N__15662\,
            I => \N__15659\
        );

    \I__2455\ : Span4Mux_h
    port map (
            O => \N__15659\,
            I => \N__15656\
        );

    \I__2454\ : Odrv4
    port map (
            O => \N__15656\,
            I => \eeprom.n2479\
        );

    \I__2453\ : InMux
    port map (
            O => \N__15653\,
            I => \N__15649\
        );

    \I__2452\ : CascadeMux
    port map (
            O => \N__15652\,
            I => \N__15646\
        );

    \I__2451\ : LocalMux
    port map (
            O => \N__15649\,
            I => \N__15643\
        );

    \I__2450\ : InMux
    port map (
            O => \N__15646\,
            I => \N__15640\
        );

    \I__2449\ : Odrv4
    port map (
            O => \N__15643\,
            I => \eeprom.n2511\
        );

    \I__2448\ : LocalMux
    port map (
            O => \N__15640\,
            I => \eeprom.n2511\
        );

    \I__2447\ : InMux
    port map (
            O => \N__15635\,
            I => \N__15632\
        );

    \I__2446\ : LocalMux
    port map (
            O => \N__15632\,
            I => \eeprom.n2578\
        );

    \I__2445\ : CascadeMux
    port map (
            O => \N__15629\,
            I => \eeprom.n2511_cascade_\
        );

    \I__2444\ : InMux
    port map (
            O => \N__15626\,
            I => \N__15623\
        );

    \I__2443\ : LocalMux
    port map (
            O => \N__15623\,
            I => \N__15620\
        );

    \I__2442\ : Odrv12
    port map (
            O => \N__15620\,
            I => \eeprom.n12_adj_351\
        );

    \I__2441\ : InMux
    port map (
            O => \N__15617\,
            I => \N__15613\
        );

    \I__2440\ : InMux
    port map (
            O => \N__15616\,
            I => \N__15610\
        );

    \I__2439\ : LocalMux
    port map (
            O => \N__15613\,
            I => \N__15606\
        );

    \I__2438\ : LocalMux
    port map (
            O => \N__15610\,
            I => \N__15603\
        );

    \I__2437\ : InMux
    port map (
            O => \N__15609\,
            I => \N__15600\
        );

    \I__2436\ : Span4Mux_v
    port map (
            O => \N__15606\,
            I => \N__15597\
        );

    \I__2435\ : Span4Mux_h
    port map (
            O => \N__15603\,
            I => \N__15594\
        );

    \I__2434\ : LocalMux
    port map (
            O => \N__15600\,
            I => \eeprom.delay_counter_21\
        );

    \I__2433\ : Odrv4
    port map (
            O => \N__15597\,
            I => \eeprom.delay_counter_21\
        );

    \I__2432\ : Odrv4
    port map (
            O => \N__15594\,
            I => \eeprom.delay_counter_21\
        );

    \I__2431\ : CascadeMux
    port map (
            O => \N__15587\,
            I => \eeprom.n2219_cascade_\
        );

    \I__2430\ : CascadeMux
    port map (
            O => \N__15584\,
            I => \N__15580\
        );

    \I__2429\ : InMux
    port map (
            O => \N__15583\,
            I => \N__15576\
        );

    \I__2428\ : InMux
    port map (
            O => \N__15580\,
            I => \N__15573\
        );

    \I__2427\ : InMux
    port map (
            O => \N__15579\,
            I => \N__15570\
        );

    \I__2426\ : LocalMux
    port map (
            O => \N__15576\,
            I => \N__15565\
        );

    \I__2425\ : LocalMux
    port map (
            O => \N__15573\,
            I => \N__15565\
        );

    \I__2424\ : LocalMux
    port map (
            O => \N__15570\,
            I => \eeprom.n2318\
        );

    \I__2423\ : Odrv4
    port map (
            O => \N__15565\,
            I => \eeprom.n2318\
        );

    \I__2422\ : InMux
    port map (
            O => \N__15560\,
            I => \N__15557\
        );

    \I__2421\ : LocalMux
    port map (
            O => \N__15557\,
            I => \N__15554\
        );

    \I__2420\ : Odrv4
    port map (
            O => \N__15554\,
            I => \eeprom.n2580\
        );

    \I__2419\ : CascadeMux
    port map (
            O => \N__15551\,
            I => \N__15548\
        );

    \I__2418\ : InMux
    port map (
            O => \N__15548\,
            I => \N__15544\
        );

    \I__2417\ : InMux
    port map (
            O => \N__15547\,
            I => \N__15541\
        );

    \I__2416\ : LocalMux
    port map (
            O => \N__15544\,
            I => \N__15538\
        );

    \I__2415\ : LocalMux
    port map (
            O => \N__15541\,
            I => \N__15534\
        );

    \I__2414\ : Span4Mux_h
    port map (
            O => \N__15538\,
            I => \N__15531\
        );

    \I__2413\ : InMux
    port map (
            O => \N__15537\,
            I => \N__15528\
        );

    \I__2412\ : Odrv4
    port map (
            O => \N__15534\,
            I => \eeprom.n2513\
        );

    \I__2411\ : Odrv4
    port map (
            O => \N__15531\,
            I => \eeprom.n2513\
        );

    \I__2410\ : LocalMux
    port map (
            O => \N__15528\,
            I => \eeprom.n2513\
        );

    \I__2409\ : CascadeMux
    port map (
            O => \N__15521\,
            I => \N__15514\
        );

    \I__2408\ : CascadeMux
    port map (
            O => \N__15520\,
            I => \N__15509\
        );

    \I__2407\ : CascadeMux
    port map (
            O => \N__15519\,
            I => \N__15506\
        );

    \I__2406\ : CascadeMux
    port map (
            O => \N__15518\,
            I => \N__15501\
        );

    \I__2405\ : CascadeMux
    port map (
            O => \N__15517\,
            I => \N__15495\
        );

    \I__2404\ : InMux
    port map (
            O => \N__15514\,
            I => \N__15489\
        );

    \I__2403\ : InMux
    port map (
            O => \N__15513\,
            I => \N__15489\
        );

    \I__2402\ : InMux
    port map (
            O => \N__15512\,
            I => \N__15484\
        );

    \I__2401\ : InMux
    port map (
            O => \N__15509\,
            I => \N__15484\
        );

    \I__2400\ : InMux
    port map (
            O => \N__15506\,
            I => \N__15479\
        );

    \I__2399\ : InMux
    port map (
            O => \N__15505\,
            I => \N__15479\
        );

    \I__2398\ : InMux
    port map (
            O => \N__15504\,
            I => \N__15472\
        );

    \I__2397\ : InMux
    port map (
            O => \N__15501\,
            I => \N__15472\
        );

    \I__2396\ : InMux
    port map (
            O => \N__15500\,
            I => \N__15472\
        );

    \I__2395\ : InMux
    port map (
            O => \N__15499\,
            I => \N__15469\
        );

    \I__2394\ : InMux
    port map (
            O => \N__15498\,
            I => \N__15462\
        );

    \I__2393\ : InMux
    port map (
            O => \N__15495\,
            I => \N__15462\
        );

    \I__2392\ : InMux
    port map (
            O => \N__15494\,
            I => \N__15462\
        );

    \I__2391\ : LocalMux
    port map (
            O => \N__15489\,
            I => \N__15457\
        );

    \I__2390\ : LocalMux
    port map (
            O => \N__15484\,
            I => \N__15457\
        );

    \I__2389\ : LocalMux
    port map (
            O => \N__15479\,
            I => \eeprom.n2539\
        );

    \I__2388\ : LocalMux
    port map (
            O => \N__15472\,
            I => \eeprom.n2539\
        );

    \I__2387\ : LocalMux
    port map (
            O => \N__15469\,
            I => \eeprom.n2539\
        );

    \I__2386\ : LocalMux
    port map (
            O => \N__15462\,
            I => \eeprom.n2539\
        );

    \I__2385\ : Odrv4
    port map (
            O => \N__15457\,
            I => \eeprom.n2539\
        );

    \I__2384\ : InMux
    port map (
            O => \N__15446\,
            I => \N__15443\
        );

    \I__2383\ : LocalMux
    port map (
            O => \N__15443\,
            I => \eeprom.n2574\
        );

    \I__2382\ : CascadeMux
    port map (
            O => \N__15440\,
            I => \eeprom.n2606_cascade_\
        );

    \I__2381\ : CascadeMux
    port map (
            O => \N__15437\,
            I => \N__15434\
        );

    \I__2380\ : InMux
    port map (
            O => \N__15434\,
            I => \N__15431\
        );

    \I__2379\ : LocalMux
    port map (
            O => \N__15431\,
            I => \N__15427\
        );

    \I__2378\ : InMux
    port map (
            O => \N__15430\,
            I => \N__15424\
        );

    \I__2377\ : Odrv4
    port map (
            O => \N__15427\,
            I => \eeprom.n2605\
        );

    \I__2376\ : LocalMux
    port map (
            O => \N__15424\,
            I => \eeprom.n2605\
        );

    \I__2375\ : CascadeMux
    port map (
            O => \N__15419\,
            I => \N__15415\
        );

    \I__2374\ : InMux
    port map (
            O => \N__15418\,
            I => \N__15412\
        );

    \I__2373\ : InMux
    port map (
            O => \N__15415\,
            I => \N__15409\
        );

    \I__2372\ : LocalMux
    port map (
            O => \N__15412\,
            I => \N__15406\
        );

    \I__2371\ : LocalMux
    port map (
            O => \N__15409\,
            I => \eeprom.n2611\
        );

    \I__2370\ : Odrv4
    port map (
            O => \N__15406\,
            I => \eeprom.n2611\
        );

    \I__2369\ : CascadeMux
    port map (
            O => \N__15401\,
            I => \eeprom.n10_adj_475_cascade_\
        );

    \I__2368\ : InMux
    port map (
            O => \N__15398\,
            I => \N__15395\
        );

    \I__2367\ : LocalMux
    port map (
            O => \N__15395\,
            I => \eeprom.n2581\
        );

    \I__2366\ : InMux
    port map (
            O => \N__15392\,
            I => \eeprom.n3578\
        );

    \I__2365\ : InMux
    port map (
            O => \N__15389\,
            I => \eeprom.n3579\
        );

    \I__2364\ : CascadeMux
    port map (
            O => \N__15386\,
            I => \N__15383\
        );

    \I__2363\ : InMux
    port map (
            O => \N__15383\,
            I => \N__15380\
        );

    \I__2362\ : LocalMux
    port map (
            O => \N__15380\,
            I => \eeprom.n2579\
        );

    \I__2361\ : InMux
    port map (
            O => \N__15377\,
            I => \eeprom.n3580\
        );

    \I__2360\ : InMux
    port map (
            O => \N__15374\,
            I => \bfn_6_22_0_\
        );

    \I__2359\ : CascadeMux
    port map (
            O => \N__15371\,
            I => \N__15366\
        );

    \I__2358\ : CascadeMux
    port map (
            O => \N__15370\,
            I => \N__15363\
        );

    \I__2357\ : InMux
    port map (
            O => \N__15369\,
            I => \N__15360\
        );

    \I__2356\ : InMux
    port map (
            O => \N__15366\,
            I => \N__15357\
        );

    \I__2355\ : InMux
    port map (
            O => \N__15363\,
            I => \N__15354\
        );

    \I__2354\ : LocalMux
    port map (
            O => \N__15360\,
            I => \eeprom.n2510\
        );

    \I__2353\ : LocalMux
    port map (
            O => \N__15357\,
            I => \eeprom.n2510\
        );

    \I__2352\ : LocalMux
    port map (
            O => \N__15354\,
            I => \eeprom.n2510\
        );

    \I__2351\ : InMux
    port map (
            O => \N__15347\,
            I => \N__15344\
        );

    \I__2350\ : LocalMux
    port map (
            O => \N__15344\,
            I => \N__15341\
        );

    \I__2349\ : Odrv4
    port map (
            O => \N__15341\,
            I => \eeprom.n2577\
        );

    \I__2348\ : InMux
    port map (
            O => \N__15338\,
            I => \eeprom.n3582\
        );

    \I__2347\ : InMux
    port map (
            O => \N__15335\,
            I => \N__15331\
        );

    \I__2346\ : CascadeMux
    port map (
            O => \N__15334\,
            I => \N__15328\
        );

    \I__2345\ : LocalMux
    port map (
            O => \N__15331\,
            I => \N__15324\
        );

    \I__2344\ : InMux
    port map (
            O => \N__15328\,
            I => \N__15321\
        );

    \I__2343\ : InMux
    port map (
            O => \N__15327\,
            I => \N__15318\
        );

    \I__2342\ : Span4Mux_h
    port map (
            O => \N__15324\,
            I => \N__15315\
        );

    \I__2341\ : LocalMux
    port map (
            O => \N__15321\,
            I => \N__15312\
        );

    \I__2340\ : LocalMux
    port map (
            O => \N__15318\,
            I => \N__15309\
        );

    \I__2339\ : Span4Mux_v
    port map (
            O => \N__15315\,
            I => \N__15306\
        );

    \I__2338\ : Span4Mux_h
    port map (
            O => \N__15312\,
            I => \N__15301\
        );

    \I__2337\ : Span4Mux_v
    port map (
            O => \N__15309\,
            I => \N__15301\
        );

    \I__2336\ : Odrv4
    port map (
            O => \N__15306\,
            I => \eeprom.n2509\
        );

    \I__2335\ : Odrv4
    port map (
            O => \N__15301\,
            I => \eeprom.n2509\
        );

    \I__2334\ : InMux
    port map (
            O => \N__15296\,
            I => \N__15293\
        );

    \I__2333\ : LocalMux
    port map (
            O => \N__15293\,
            I => \N__15290\
        );

    \I__2332\ : Odrv4
    port map (
            O => \N__15290\,
            I => \eeprom.n2576\
        );

    \I__2331\ : InMux
    port map (
            O => \N__15287\,
            I => \eeprom.n3583\
        );

    \I__2330\ : InMux
    port map (
            O => \N__15284\,
            I => \N__15280\
        );

    \I__2329\ : CascadeMux
    port map (
            O => \N__15283\,
            I => \N__15277\
        );

    \I__2328\ : LocalMux
    port map (
            O => \N__15280\,
            I => \N__15273\
        );

    \I__2327\ : InMux
    port map (
            O => \N__15277\,
            I => \N__15270\
        );

    \I__2326\ : CascadeMux
    port map (
            O => \N__15276\,
            I => \N__15267\
        );

    \I__2325\ : Span4Mux_v
    port map (
            O => \N__15273\,
            I => \N__15262\
        );

    \I__2324\ : LocalMux
    port map (
            O => \N__15270\,
            I => \N__15262\
        );

    \I__2323\ : InMux
    port map (
            O => \N__15267\,
            I => \N__15259\
        );

    \I__2322\ : Span4Mux_h
    port map (
            O => \N__15262\,
            I => \N__15256\
        );

    \I__2321\ : LocalMux
    port map (
            O => \N__15259\,
            I => \N__15253\
        );

    \I__2320\ : Span4Mux_v
    port map (
            O => \N__15256\,
            I => \N__15250\
        );

    \I__2319\ : Span4Mux_v
    port map (
            O => \N__15253\,
            I => \N__15247\
        );

    \I__2318\ : Odrv4
    port map (
            O => \N__15250\,
            I => \eeprom.n2508\
        );

    \I__2317\ : Odrv4
    port map (
            O => \N__15247\,
            I => \eeprom.n2508\
        );

    \I__2316\ : CascadeMux
    port map (
            O => \N__15242\,
            I => \N__15239\
        );

    \I__2315\ : InMux
    port map (
            O => \N__15239\,
            I => \N__15236\
        );

    \I__2314\ : LocalMux
    port map (
            O => \N__15236\,
            I => \N__15233\
        );

    \I__2313\ : Odrv4
    port map (
            O => \N__15233\,
            I => \eeprom.n2575\
        );

    \I__2312\ : InMux
    port map (
            O => \N__15230\,
            I => \eeprom.n3584\
        );

    \I__2311\ : InMux
    port map (
            O => \N__15227\,
            I => \eeprom.n3585\
        );

    \I__2310\ : InMux
    port map (
            O => \N__15224\,
            I => \N__15220\
        );

    \I__2309\ : InMux
    port map (
            O => \N__15223\,
            I => \N__15217\
        );

    \I__2308\ : LocalMux
    port map (
            O => \N__15220\,
            I => \N__15214\
        );

    \I__2307\ : LocalMux
    port map (
            O => \N__15217\,
            I => \N__15211\
        );

    \I__2306\ : Span4Mux_h
    port map (
            O => \N__15214\,
            I => \N__15206\
        );

    \I__2305\ : Span4Mux_v
    port map (
            O => \N__15211\,
            I => \N__15206\
        );

    \I__2304\ : Odrv4
    port map (
            O => \N__15206\,
            I => \eeprom.n2506\
        );

    \I__2303\ : InMux
    port map (
            O => \N__15203\,
            I => \eeprom.n3586\
        );

    \I__2302\ : InMux
    port map (
            O => \N__15200\,
            I => \N__15197\
        );

    \I__2301\ : LocalMux
    port map (
            O => \N__15197\,
            I => \eeprom.n2678\
        );

    \I__2300\ : CascadeMux
    port map (
            O => \N__15194\,
            I => \eeprom.n2611_cascade_\
        );

    \I__2299\ : InMux
    port map (
            O => \N__15191\,
            I => \N__15188\
        );

    \I__2298\ : LocalMux
    port map (
            O => \N__15188\,
            I => \N__15184\
        );

    \I__2297\ : InMux
    port map (
            O => \N__15187\,
            I => \N__15181\
        );

    \I__2296\ : Span4Mux_v
    port map (
            O => \N__15184\,
            I => \N__15175\
        );

    \I__2295\ : LocalMux
    port map (
            O => \N__15181\,
            I => \N__15175\
        );

    \I__2294\ : InMux
    port map (
            O => \N__15180\,
            I => \N__15172\
        );

    \I__2293\ : Span4Mux_h
    port map (
            O => \N__15175\,
            I => \N__15169\
        );

    \I__2292\ : LocalMux
    port map (
            O => \N__15172\,
            I => \eeprom.n2519\
        );

    \I__2291\ : Odrv4
    port map (
            O => \N__15169\,
            I => \eeprom.n2519\
        );

    \I__2290\ : InMux
    port map (
            O => \N__15164\,
            I => \N__15161\
        );

    \I__2289\ : LocalMux
    port map (
            O => \N__15161\,
            I => \N__15158\
        );

    \I__2288\ : Odrv4
    port map (
            O => \N__15158\,
            I => \eeprom.n2586\
        );

    \I__2287\ : InMux
    port map (
            O => \N__15155\,
            I => \bfn_6_21_0_\
        );

    \I__2286\ : CascadeMux
    port map (
            O => \N__15152\,
            I => \N__15149\
        );

    \I__2285\ : InMux
    port map (
            O => \N__15149\,
            I => \N__15145\
        );

    \I__2284\ : CascadeMux
    port map (
            O => \N__15148\,
            I => \N__15141\
        );

    \I__2283\ : LocalMux
    port map (
            O => \N__15145\,
            I => \N__15138\
        );

    \I__2282\ : InMux
    port map (
            O => \N__15144\,
            I => \N__15135\
        );

    \I__2281\ : InMux
    port map (
            O => \N__15141\,
            I => \N__15132\
        );

    \I__2280\ : Odrv4
    port map (
            O => \N__15138\,
            I => \eeprom.n2518\
        );

    \I__2279\ : LocalMux
    port map (
            O => \N__15135\,
            I => \eeprom.n2518\
        );

    \I__2278\ : LocalMux
    port map (
            O => \N__15132\,
            I => \eeprom.n2518\
        );

    \I__2277\ : InMux
    port map (
            O => \N__15125\,
            I => \N__15122\
        );

    \I__2276\ : LocalMux
    port map (
            O => \N__15122\,
            I => \N__15119\
        );

    \I__2275\ : Odrv4
    port map (
            O => \N__15119\,
            I => \eeprom.n2585\
        );

    \I__2274\ : InMux
    port map (
            O => \N__15116\,
            I => \eeprom.n3574\
        );

    \I__2273\ : CascadeMux
    port map (
            O => \N__15113\,
            I => \N__15109\
        );

    \I__2272\ : InMux
    port map (
            O => \N__15112\,
            I => \N__15106\
        );

    \I__2271\ : InMux
    port map (
            O => \N__15109\,
            I => \N__15103\
        );

    \I__2270\ : LocalMux
    port map (
            O => \N__15106\,
            I => \N__15100\
        );

    \I__2269\ : LocalMux
    port map (
            O => \N__15103\,
            I => \N__15097\
        );

    \I__2268\ : Span4Mux_v
    port map (
            O => \N__15100\,
            I => \N__15093\
        );

    \I__2267\ : Span4Mux_h
    port map (
            O => \N__15097\,
            I => \N__15090\
        );

    \I__2266\ : InMux
    port map (
            O => \N__15096\,
            I => \N__15087\
        );

    \I__2265\ : Odrv4
    port map (
            O => \N__15093\,
            I => \eeprom.n2517\
        );

    \I__2264\ : Odrv4
    port map (
            O => \N__15090\,
            I => \eeprom.n2517\
        );

    \I__2263\ : LocalMux
    port map (
            O => \N__15087\,
            I => \eeprom.n2517\
        );

    \I__2262\ : InMux
    port map (
            O => \N__15080\,
            I => \N__15077\
        );

    \I__2261\ : LocalMux
    port map (
            O => \N__15077\,
            I => \N__15074\
        );

    \I__2260\ : Odrv4
    port map (
            O => \N__15074\,
            I => \eeprom.n2584\
        );

    \I__2259\ : InMux
    port map (
            O => \N__15071\,
            I => \eeprom.n3575\
        );

    \I__2258\ : CascadeMux
    port map (
            O => \N__15068\,
            I => \N__15064\
        );

    \I__2257\ : InMux
    port map (
            O => \N__15067\,
            I => \N__15061\
        );

    \I__2256\ : InMux
    port map (
            O => \N__15064\,
            I => \N__15058\
        );

    \I__2255\ : LocalMux
    port map (
            O => \N__15061\,
            I => \N__15055\
        );

    \I__2254\ : LocalMux
    port map (
            O => \N__15058\,
            I => \N__15052\
        );

    \I__2253\ : Span4Mux_v
    port map (
            O => \N__15055\,
            I => \N__15048\
        );

    \I__2252\ : Span4Mux_h
    port map (
            O => \N__15052\,
            I => \N__15045\
        );

    \I__2251\ : InMux
    port map (
            O => \N__15051\,
            I => \N__15042\
        );

    \I__2250\ : Odrv4
    port map (
            O => \N__15048\,
            I => \eeprom.n2516\
        );

    \I__2249\ : Odrv4
    port map (
            O => \N__15045\,
            I => \eeprom.n2516\
        );

    \I__2248\ : LocalMux
    port map (
            O => \N__15042\,
            I => \eeprom.n2516\
        );

    \I__2247\ : CascadeMux
    port map (
            O => \N__15035\,
            I => \N__15032\
        );

    \I__2246\ : InMux
    port map (
            O => \N__15032\,
            I => \N__15029\
        );

    \I__2245\ : LocalMux
    port map (
            O => \N__15029\,
            I => \N__15026\
        );

    \I__2244\ : Odrv4
    port map (
            O => \N__15026\,
            I => \eeprom.n2583\
        );

    \I__2243\ : InMux
    port map (
            O => \N__15023\,
            I => \eeprom.n3576\
        );

    \I__2242\ : CascadeMux
    port map (
            O => \N__15020\,
            I => \N__15016\
        );

    \I__2241\ : CascadeMux
    port map (
            O => \N__15019\,
            I => \N__15013\
        );

    \I__2240\ : InMux
    port map (
            O => \N__15016\,
            I => \N__15010\
        );

    \I__2239\ : InMux
    port map (
            O => \N__15013\,
            I => \N__15007\
        );

    \I__2238\ : LocalMux
    port map (
            O => \N__15010\,
            I => \N__15003\
        );

    \I__2237\ : LocalMux
    port map (
            O => \N__15007\,
            I => \N__15000\
        );

    \I__2236\ : CascadeMux
    port map (
            O => \N__15006\,
            I => \N__14997\
        );

    \I__2235\ : Span4Mux_h
    port map (
            O => \N__15003\,
            I => \N__14994\
        );

    \I__2234\ : Span4Mux_h
    port map (
            O => \N__15000\,
            I => \N__14991\
        );

    \I__2233\ : InMux
    port map (
            O => \N__14997\,
            I => \N__14988\
        );

    \I__2232\ : Odrv4
    port map (
            O => \N__14994\,
            I => \eeprom.n2515\
        );

    \I__2231\ : Odrv4
    port map (
            O => \N__14991\,
            I => \eeprom.n2515\
        );

    \I__2230\ : LocalMux
    port map (
            O => \N__14988\,
            I => \eeprom.n2515\
        );

    \I__2229\ : InMux
    port map (
            O => \N__14981\,
            I => \N__14978\
        );

    \I__2228\ : LocalMux
    port map (
            O => \N__14978\,
            I => \eeprom.n2582\
        );

    \I__2227\ : InMux
    port map (
            O => \N__14975\,
            I => \eeprom.n3577\
        );

    \I__2226\ : CascadeMux
    port map (
            O => \N__14972\,
            I => \N__14969\
        );

    \I__2225\ : InMux
    port map (
            O => \N__14969\,
            I => \N__14965\
        );

    \I__2224\ : InMux
    port map (
            O => \N__14968\,
            I => \N__14962\
        );

    \I__2223\ : LocalMux
    port map (
            O => \N__14965\,
            I => \N__14959\
        );

    \I__2222\ : LocalMux
    port map (
            O => \N__14962\,
            I => \N__14955\
        );

    \I__2221\ : Span4Mux_h
    port map (
            O => \N__14959\,
            I => \N__14952\
        );

    \I__2220\ : InMux
    port map (
            O => \N__14958\,
            I => \N__14949\
        );

    \I__2219\ : Odrv4
    port map (
            O => \N__14955\,
            I => \eeprom.n2514\
        );

    \I__2218\ : Odrv4
    port map (
            O => \N__14952\,
            I => \eeprom.n2514\
        );

    \I__2217\ : LocalMux
    port map (
            O => \N__14949\,
            I => \eeprom.n2514\
        );

    \I__2216\ : InMux
    port map (
            O => \N__14942\,
            I => \eeprom.n3597\
        );

    \I__2215\ : InMux
    port map (
            O => \N__14939\,
            I => \eeprom.n3598\
        );

    \I__2214\ : InMux
    port map (
            O => \N__14936\,
            I => \eeprom.n3599\
        );

    \I__2213\ : InMux
    port map (
            O => \N__14933\,
            I => \eeprom.n3600\
        );

    \I__2212\ : InMux
    port map (
            O => \N__14930\,
            I => \N__14927\
        );

    \I__2211\ : LocalMux
    port map (
            O => \N__14927\,
            I => \N__14924\
        );

    \I__2210\ : Span4Mux_v
    port map (
            O => \N__14924\,
            I => \N__14921\
        );

    \I__2209\ : Odrv4
    port map (
            O => \N__14921\,
            I => \eeprom.n21\
        );

    \I__2208\ : InMux
    port map (
            O => \N__14918\,
            I => \N__14915\
        );

    \I__2207\ : LocalMux
    port map (
            O => \N__14915\,
            I => \N__14911\
        );

    \I__2206\ : InMux
    port map (
            O => \N__14914\,
            I => \N__14907\
        );

    \I__2205\ : Span4Mux_h
    port map (
            O => \N__14911\,
            I => \N__14904\
        );

    \I__2204\ : InMux
    port map (
            O => \N__14910\,
            I => \N__14901\
        );

    \I__2203\ : LocalMux
    port map (
            O => \N__14907\,
            I => \eeprom.delay_counter_12\
        );

    \I__2202\ : Odrv4
    port map (
            O => \N__14904\,
            I => \eeprom.delay_counter_12\
        );

    \I__2201\ : LocalMux
    port map (
            O => \N__14901\,
            I => \eeprom.delay_counter_12\
        );

    \I__2200\ : CascadeMux
    port map (
            O => \N__14894\,
            I => \N__14891\
        );

    \I__2199\ : InMux
    port map (
            O => \N__14891\,
            I => \N__14888\
        );

    \I__2198\ : LocalMux
    port map (
            O => \N__14888\,
            I => \N__14885\
        );

    \I__2197\ : Span4Mux_h
    port map (
            O => \N__14885\,
            I => \N__14882\
        );

    \I__2196\ : Odrv4
    port map (
            O => \N__14882\,
            I => \eeprom.n29_adj_460\
        );

    \I__2195\ : CascadeMux
    port map (
            O => \N__14879\,
            I => \N__14875\
        );

    \I__2194\ : InMux
    port map (
            O => \N__14878\,
            I => \N__14871\
        );

    \I__2193\ : InMux
    port map (
            O => \N__14875\,
            I => \N__14868\
        );

    \I__2192\ : InMux
    port map (
            O => \N__14874\,
            I => \N__14865\
        );

    \I__2191\ : LocalMux
    port map (
            O => \N__14871\,
            I => \eeprom.n2609\
        );

    \I__2190\ : LocalMux
    port map (
            O => \N__14868\,
            I => \eeprom.n2609\
        );

    \I__2189\ : LocalMux
    port map (
            O => \N__14865\,
            I => \eeprom.n2609\
        );

    \I__2188\ : CascadeMux
    port map (
            O => \N__14858\,
            I => \N__14855\
        );

    \I__2187\ : InMux
    port map (
            O => \N__14855\,
            I => \N__14852\
        );

    \I__2186\ : LocalMux
    port map (
            O => \N__14852\,
            I => \eeprom.n2676\
        );

    \I__2185\ : InMux
    port map (
            O => \N__14849\,
            I => \eeprom.n3588\
        );

    \I__2184\ : InMux
    port map (
            O => \N__14846\,
            I => \eeprom.n3589\
        );

    \I__2183\ : InMux
    port map (
            O => \N__14843\,
            I => \eeprom.n3590\
        );

    \I__2182\ : InMux
    port map (
            O => \N__14840\,
            I => \eeprom.n3591\
        );

    \I__2181\ : InMux
    port map (
            O => \N__14837\,
            I => \eeprom.n3592\
        );

    \I__2180\ : InMux
    port map (
            O => \N__14834\,
            I => \eeprom.n3593\
        );

    \I__2179\ : InMux
    port map (
            O => \N__14831\,
            I => \bfn_6_19_0_\
        );

    \I__2178\ : InMux
    port map (
            O => \N__14828\,
            I => \eeprom.n3595\
        );

    \I__2177\ : InMux
    port map (
            O => \N__14825\,
            I => \eeprom.n3596\
        );

    \I__2176\ : InMux
    port map (
            O => \N__14822\,
            I => \N__14819\
        );

    \I__2175\ : LocalMux
    port map (
            O => \N__14819\,
            I => n7
        );

    \I__2174\ : InMux
    port map (
            O => \N__14816\,
            I => n3503
        );

    \I__2173\ : InMux
    port map (
            O => \N__14813\,
            I => \N__14810\
        );

    \I__2172\ : LocalMux
    port map (
            O => \N__14810\,
            I => n6
        );

    \I__2171\ : InMux
    port map (
            O => \N__14807\,
            I => n3504
        );

    \I__2170\ : CascadeMux
    port map (
            O => \N__14804\,
            I => \N__14801\
        );

    \I__2169\ : InMux
    port map (
            O => \N__14801\,
            I => \N__14794\
        );

    \I__2168\ : InMux
    port map (
            O => \N__14800\,
            I => \N__14794\
        );

    \I__2167\ : InMux
    port map (
            O => \N__14799\,
            I => \N__14791\
        );

    \I__2166\ : LocalMux
    port map (
            O => \N__14794\,
            I => blink_counter_21
        );

    \I__2165\ : LocalMux
    port map (
            O => \N__14791\,
            I => blink_counter_21
        );

    \I__2164\ : InMux
    port map (
            O => \N__14786\,
            I => n3505
        );

    \I__2163\ : InMux
    port map (
            O => \N__14783\,
            I => \N__14776\
        );

    \I__2162\ : InMux
    port map (
            O => \N__14782\,
            I => \N__14776\
        );

    \I__2161\ : InMux
    port map (
            O => \N__14781\,
            I => \N__14773\
        );

    \I__2160\ : LocalMux
    port map (
            O => \N__14776\,
            I => blink_counter_22
        );

    \I__2159\ : LocalMux
    port map (
            O => \N__14773\,
            I => blink_counter_22
        );

    \I__2158\ : InMux
    port map (
            O => \N__14768\,
            I => n3506
        );

    \I__2157\ : CascadeMux
    port map (
            O => \N__14765\,
            I => \N__14761\
        );

    \I__2156\ : InMux
    port map (
            O => \N__14764\,
            I => \N__14755\
        );

    \I__2155\ : InMux
    port map (
            O => \N__14761\,
            I => \N__14755\
        );

    \I__2154\ : InMux
    port map (
            O => \N__14760\,
            I => \N__14752\
        );

    \I__2153\ : LocalMux
    port map (
            O => \N__14755\,
            I => blink_counter_23
        );

    \I__2152\ : LocalMux
    port map (
            O => \N__14752\,
            I => blink_counter_23
        );

    \I__2151\ : InMux
    port map (
            O => \N__14747\,
            I => n3507
        );

    \I__2150\ : InMux
    port map (
            O => \N__14744\,
            I => \N__14737\
        );

    \I__2149\ : InMux
    port map (
            O => \N__14743\,
            I => \N__14737\
        );

    \I__2148\ : InMux
    port map (
            O => \N__14742\,
            I => \N__14734\
        );

    \I__2147\ : LocalMux
    port map (
            O => \N__14737\,
            I => blink_counter_24
        );

    \I__2146\ : LocalMux
    port map (
            O => \N__14734\,
            I => blink_counter_24
        );

    \I__2145\ : InMux
    port map (
            O => \N__14729\,
            I => \bfn_5_32_0_\
        );

    \I__2144\ : InMux
    port map (
            O => \N__14726\,
            I => n3509
        );

    \I__2143\ : InMux
    port map (
            O => \N__14723\,
            I => \N__14719\
        );

    \I__2142\ : InMux
    port map (
            O => \N__14722\,
            I => \N__14716\
        );

    \I__2141\ : LocalMux
    port map (
            O => \N__14719\,
            I => blink_counter_25
        );

    \I__2140\ : LocalMux
    port map (
            O => \N__14716\,
            I => blink_counter_25
        );

    \I__2139\ : InMux
    port map (
            O => \N__14711\,
            I => \bfn_6_18_0_\
        );

    \I__2138\ : InMux
    port map (
            O => \N__14708\,
            I => \eeprom.n3587\
        );

    \I__2137\ : InMux
    port map (
            O => \N__14705\,
            I => \N__14702\
        );

    \I__2136\ : LocalMux
    port map (
            O => \N__14702\,
            I => n15
        );

    \I__2135\ : InMux
    port map (
            O => \N__14699\,
            I => n3495
        );

    \I__2134\ : InMux
    port map (
            O => \N__14696\,
            I => \N__14693\
        );

    \I__2133\ : LocalMux
    port map (
            O => \N__14693\,
            I => n14
        );

    \I__2132\ : InMux
    port map (
            O => \N__14690\,
            I => n3496
        );

    \I__2131\ : InMux
    port map (
            O => \N__14687\,
            I => \N__14684\
        );

    \I__2130\ : LocalMux
    port map (
            O => \N__14684\,
            I => n13
        );

    \I__2129\ : InMux
    port map (
            O => \N__14681\,
            I => n3497
        );

    \I__2128\ : InMux
    port map (
            O => \N__14678\,
            I => \N__14675\
        );

    \I__2127\ : LocalMux
    port map (
            O => \N__14675\,
            I => n12
        );

    \I__2126\ : InMux
    port map (
            O => \N__14672\,
            I => n3498
        );

    \I__2125\ : InMux
    port map (
            O => \N__14669\,
            I => \N__14666\
        );

    \I__2124\ : LocalMux
    port map (
            O => \N__14666\,
            I => n11
        );

    \I__2123\ : InMux
    port map (
            O => \N__14663\,
            I => n3499
        );

    \I__2122\ : InMux
    port map (
            O => \N__14660\,
            I => \N__14657\
        );

    \I__2121\ : LocalMux
    port map (
            O => \N__14657\,
            I => n10
        );

    \I__2120\ : InMux
    port map (
            O => \N__14654\,
            I => \bfn_5_31_0_\
        );

    \I__2119\ : InMux
    port map (
            O => \N__14651\,
            I => \N__14648\
        );

    \I__2118\ : LocalMux
    port map (
            O => \N__14648\,
            I => n9
        );

    \I__2117\ : InMux
    port map (
            O => \N__14645\,
            I => n3501
        );

    \I__2116\ : InMux
    port map (
            O => \N__14642\,
            I => \N__14639\
        );

    \I__2115\ : LocalMux
    port map (
            O => \N__14639\,
            I => n8
        );

    \I__2114\ : InMux
    port map (
            O => \N__14636\,
            I => n3502
        );

    \I__2113\ : InMux
    port map (
            O => \N__14633\,
            I => \N__14630\
        );

    \I__2112\ : LocalMux
    port map (
            O => \N__14630\,
            I => n23
        );

    \I__2111\ : InMux
    port map (
            O => \N__14627\,
            I => n3487
        );

    \I__2110\ : InMux
    port map (
            O => \N__14624\,
            I => \N__14621\
        );

    \I__2109\ : LocalMux
    port map (
            O => \N__14621\,
            I => n22
        );

    \I__2108\ : InMux
    port map (
            O => \N__14618\,
            I => n3488
        );

    \I__2107\ : InMux
    port map (
            O => \N__14615\,
            I => \N__14612\
        );

    \I__2106\ : LocalMux
    port map (
            O => \N__14612\,
            I => n21
        );

    \I__2105\ : InMux
    port map (
            O => \N__14609\,
            I => n3489
        );

    \I__2104\ : InMux
    port map (
            O => \N__14606\,
            I => \N__14603\
        );

    \I__2103\ : LocalMux
    port map (
            O => \N__14603\,
            I => n20
        );

    \I__2102\ : InMux
    port map (
            O => \N__14600\,
            I => n3490
        );

    \I__2101\ : InMux
    port map (
            O => \N__14597\,
            I => \N__14594\
        );

    \I__2100\ : LocalMux
    port map (
            O => \N__14594\,
            I => n19
        );

    \I__2099\ : InMux
    port map (
            O => \N__14591\,
            I => n3491
        );

    \I__2098\ : InMux
    port map (
            O => \N__14588\,
            I => \N__14585\
        );

    \I__2097\ : LocalMux
    port map (
            O => \N__14585\,
            I => n18
        );

    \I__2096\ : InMux
    port map (
            O => \N__14582\,
            I => \bfn_5_30_0_\
        );

    \I__2095\ : InMux
    port map (
            O => \N__14579\,
            I => \N__14576\
        );

    \I__2094\ : LocalMux
    port map (
            O => \N__14576\,
            I => n17
        );

    \I__2093\ : InMux
    port map (
            O => \N__14573\,
            I => n3493
        );

    \I__2092\ : InMux
    port map (
            O => \N__14570\,
            I => \N__14567\
        );

    \I__2091\ : LocalMux
    port map (
            O => \N__14567\,
            I => n16
        );

    \I__2090\ : InMux
    port map (
            O => \N__14564\,
            I => n3494
        );

    \I__2089\ : CascadeMux
    port map (
            O => \N__14561\,
            I => \N__14558\
        );

    \I__2088\ : InMux
    port map (
            O => \N__14558\,
            I => \N__14553\
        );

    \I__2087\ : InMux
    port map (
            O => \N__14557\,
            I => \N__14550\
        );

    \I__2086\ : CascadeMux
    port map (
            O => \N__14556\,
            I => \N__14547\
        );

    \I__2085\ : LocalMux
    port map (
            O => \N__14553\,
            I => \N__14544\
        );

    \I__2084\ : LocalMux
    port map (
            O => \N__14550\,
            I => \N__14541\
        );

    \I__2083\ : InMux
    port map (
            O => \N__14547\,
            I => \N__14538\
        );

    \I__2082\ : Odrv4
    port map (
            O => \N__14544\,
            I => \eeprom.n2115\
        );

    \I__2081\ : Odrv12
    port map (
            O => \N__14541\,
            I => \eeprom.n2115\
        );

    \I__2080\ : LocalMux
    port map (
            O => \N__14538\,
            I => \eeprom.n2115\
        );

    \I__2079\ : InMux
    port map (
            O => \N__14531\,
            I => \N__14528\
        );

    \I__2078\ : LocalMux
    port map (
            O => \N__14528\,
            I => \N__14525\
        );

    \I__2077\ : Odrv4
    port map (
            O => \N__14525\,
            I => \eeprom.n2182\
        );

    \I__2076\ : InMux
    port map (
            O => \N__14522\,
            I => \eeprom.n3535\
        );

    \I__2075\ : InMux
    port map (
            O => \N__14519\,
            I => \N__14516\
        );

    \I__2074\ : LocalMux
    port map (
            O => \N__14516\,
            I => \N__14512\
        );

    \I__2073\ : InMux
    port map (
            O => \N__14515\,
            I => \N__14509\
        );

    \I__2072\ : Span4Mux_v
    port map (
            O => \N__14512\,
            I => \N__14506\
        );

    \I__2071\ : LocalMux
    port map (
            O => \N__14509\,
            I => \N__14503\
        );

    \I__2070\ : Span4Mux_v
    port map (
            O => \N__14506\,
            I => \N__14500\
        );

    \I__2069\ : Span4Mux_v
    port map (
            O => \N__14503\,
            I => \N__14497\
        );

    \I__2068\ : Odrv4
    port map (
            O => \N__14500\,
            I => \eeprom.n2114\
        );

    \I__2067\ : Odrv4
    port map (
            O => \N__14497\,
            I => \eeprom.n2114\
        );

    \I__2066\ : InMux
    port map (
            O => \N__14492\,
            I => \N__14489\
        );

    \I__2065\ : LocalMux
    port map (
            O => \N__14489\,
            I => \eeprom.n2181\
        );

    \I__2064\ : InMux
    port map (
            O => \N__14486\,
            I => \eeprom.n3536\
        );

    \I__2063\ : InMux
    port map (
            O => \N__14483\,
            I => \eeprom.n3537\
        );

    \I__2062\ : CascadeMux
    port map (
            O => \N__14480\,
            I => \N__14475\
        );

    \I__2061\ : InMux
    port map (
            O => \N__14479\,
            I => \N__14470\
        );

    \I__2060\ : InMux
    port map (
            O => \N__14478\,
            I => \N__14470\
        );

    \I__2059\ : InMux
    port map (
            O => \N__14475\,
            I => \N__14467\
        );

    \I__2058\ : LocalMux
    port map (
            O => \N__14470\,
            I => \N__14462\
        );

    \I__2057\ : LocalMux
    port map (
            O => \N__14467\,
            I => \N__14462\
        );

    \I__2056\ : Span4Mux_v
    port map (
            O => \N__14462\,
            I => \N__14459\
        );

    \I__2055\ : Odrv4
    port map (
            O => \N__14459\,
            I => \eeprom.n2112\
        );

    \I__2054\ : CascadeMux
    port map (
            O => \N__14456\,
            I => \N__14453\
        );

    \I__2053\ : InMux
    port map (
            O => \N__14453\,
            I => \N__14450\
        );

    \I__2052\ : LocalMux
    port map (
            O => \N__14450\,
            I => \eeprom.n2179\
        );

    \I__2051\ : InMux
    port map (
            O => \N__14447\,
            I => \eeprom.n3538\
        );

    \I__2050\ : CascadeMux
    port map (
            O => \N__14444\,
            I => \N__14441\
        );

    \I__2049\ : InMux
    port map (
            O => \N__14441\,
            I => \N__14437\
        );

    \I__2048\ : InMux
    port map (
            O => \N__14440\,
            I => \N__14433\
        );

    \I__2047\ : LocalMux
    port map (
            O => \N__14437\,
            I => \N__14430\
        );

    \I__2046\ : InMux
    port map (
            O => \N__14436\,
            I => \N__14427\
        );

    \I__2045\ : LocalMux
    port map (
            O => \N__14433\,
            I => \N__14424\
        );

    \I__2044\ : Span4Mux_v
    port map (
            O => \N__14430\,
            I => \N__14419\
        );

    \I__2043\ : LocalMux
    port map (
            O => \N__14427\,
            I => \N__14419\
        );

    \I__2042\ : Odrv4
    port map (
            O => \N__14424\,
            I => \eeprom.n2111\
        );

    \I__2041\ : Odrv4
    port map (
            O => \N__14419\,
            I => \eeprom.n2111\
        );

    \I__2040\ : InMux
    port map (
            O => \N__14414\,
            I => \N__14411\
        );

    \I__2039\ : LocalMux
    port map (
            O => \N__14411\,
            I => \N__14408\
        );

    \I__2038\ : Odrv4
    port map (
            O => \N__14408\,
            I => \eeprom.n2178\
        );

    \I__2037\ : InMux
    port map (
            O => \N__14405\,
            I => \bfn_5_28_0_\
        );

    \I__2036\ : InMux
    port map (
            O => \N__14402\,
            I => \N__14399\
        );

    \I__2035\ : LocalMux
    port map (
            O => \N__14399\,
            I => \N__14395\
        );

    \I__2034\ : InMux
    port map (
            O => \N__14398\,
            I => \N__14392\
        );

    \I__2033\ : Span4Mux_v
    port map (
            O => \N__14395\,
            I => \N__14387\
        );

    \I__2032\ : LocalMux
    port map (
            O => \N__14392\,
            I => \N__14387\
        );

    \I__2031\ : Span4Mux_v
    port map (
            O => \N__14387\,
            I => \N__14384\
        );

    \I__2030\ : Odrv4
    port map (
            O => \N__14384\,
            I => \eeprom.n2110\
        );

    \I__2029\ : InMux
    port map (
            O => \N__14381\,
            I => \eeprom.n3540\
        );

    \I__2028\ : InMux
    port map (
            O => \N__14378\,
            I => \N__14375\
        );

    \I__2027\ : LocalMux
    port map (
            O => \N__14375\,
            I => n26
        );

    \I__2026\ : InMux
    port map (
            O => \N__14372\,
            I => \bfn_5_29_0_\
        );

    \I__2025\ : InMux
    port map (
            O => \N__14369\,
            I => \N__14366\
        );

    \I__2024\ : LocalMux
    port map (
            O => \N__14366\,
            I => n25
        );

    \I__2023\ : InMux
    port map (
            O => \N__14363\,
            I => n3485
        );

    \I__2022\ : InMux
    port map (
            O => \N__14360\,
            I => \N__14357\
        );

    \I__2021\ : LocalMux
    port map (
            O => \N__14357\,
            I => n24
        );

    \I__2020\ : InMux
    port map (
            O => \N__14354\,
            I => n3486
        );

    \I__2019\ : CascadeMux
    port map (
            O => \N__14351\,
            I => \eeprom.n2143_cascade_\
        );

    \I__2018\ : InMux
    port map (
            O => \N__14348\,
            I => \bfn_5_27_0_\
        );

    \I__2017\ : CascadeMux
    port map (
            O => \N__14345\,
            I => \N__14340\
        );

    \I__2016\ : InMux
    port map (
            O => \N__14344\,
            I => \N__14335\
        );

    \I__2015\ : InMux
    port map (
            O => \N__14343\,
            I => \N__14335\
        );

    \I__2014\ : InMux
    port map (
            O => \N__14340\,
            I => \N__14332\
        );

    \I__2013\ : LocalMux
    port map (
            O => \N__14335\,
            I => \N__14327\
        );

    \I__2012\ : LocalMux
    port map (
            O => \N__14332\,
            I => \N__14327\
        );

    \I__2011\ : Odrv12
    port map (
            O => \N__14327\,
            I => \eeprom.n2118\
        );

    \I__2010\ : InMux
    port map (
            O => \N__14324\,
            I => \N__14321\
        );

    \I__2009\ : LocalMux
    port map (
            O => \N__14321\,
            I => \eeprom.n2185\
        );

    \I__2008\ : InMux
    port map (
            O => \N__14318\,
            I => \eeprom.n3532\
        );

    \I__2007\ : CascadeMux
    port map (
            O => \N__14315\,
            I => \N__14311\
        );

    \I__2006\ : CascadeMux
    port map (
            O => \N__14314\,
            I => \N__14308\
        );

    \I__2005\ : InMux
    port map (
            O => \N__14311\,
            I => \N__14305\
        );

    \I__2004\ : InMux
    port map (
            O => \N__14308\,
            I => \N__14302\
        );

    \I__2003\ : LocalMux
    port map (
            O => \N__14305\,
            I => \N__14299\
        );

    \I__2002\ : LocalMux
    port map (
            O => \N__14302\,
            I => \N__14296\
        );

    \I__2001\ : Span4Mux_v
    port map (
            O => \N__14299\,
            I => \N__14290\
        );

    \I__2000\ : Span4Mux_v
    port map (
            O => \N__14296\,
            I => \N__14290\
        );

    \I__1999\ : InMux
    port map (
            O => \N__14295\,
            I => \N__14287\
        );

    \I__1998\ : Odrv4
    port map (
            O => \N__14290\,
            I => \eeprom.n2117\
        );

    \I__1997\ : LocalMux
    port map (
            O => \N__14287\,
            I => \eeprom.n2117\
        );

    \I__1996\ : InMux
    port map (
            O => \N__14282\,
            I => \N__14279\
        );

    \I__1995\ : LocalMux
    port map (
            O => \N__14279\,
            I => \eeprom.n2184\
        );

    \I__1994\ : InMux
    port map (
            O => \N__14276\,
            I => \eeprom.n3533\
        );

    \I__1993\ : CascadeMux
    port map (
            O => \N__14273\,
            I => \N__14269\
        );

    \I__1992\ : InMux
    port map (
            O => \N__14272\,
            I => \N__14266\
        );

    \I__1991\ : InMux
    port map (
            O => \N__14269\,
            I => \N__14263\
        );

    \I__1990\ : LocalMux
    port map (
            O => \N__14266\,
            I => \N__14257\
        );

    \I__1989\ : LocalMux
    port map (
            O => \N__14263\,
            I => \N__14257\
        );

    \I__1988\ : InMux
    port map (
            O => \N__14262\,
            I => \N__14254\
        );

    \I__1987\ : Odrv12
    port map (
            O => \N__14257\,
            I => \eeprom.n2116\
        );

    \I__1986\ : LocalMux
    port map (
            O => \N__14254\,
            I => \eeprom.n2116\
        );

    \I__1985\ : InMux
    port map (
            O => \N__14249\,
            I => \N__14246\
        );

    \I__1984\ : LocalMux
    port map (
            O => \N__14246\,
            I => \N__14242\
        );

    \I__1983\ : InMux
    port map (
            O => \N__14245\,
            I => \N__14239\
        );

    \I__1982\ : Odrv4
    port map (
            O => \N__14242\,
            I => \eeprom.n2183\
        );

    \I__1981\ : LocalMux
    port map (
            O => \N__14239\,
            I => \eeprom.n2183\
        );

    \I__1980\ : InMux
    port map (
            O => \N__14234\,
            I => \eeprom.n3534\
        );

    \I__1979\ : CascadeMux
    port map (
            O => \N__14231\,
            I => \eeprom.n2214_cascade_\
        );

    \I__1978\ : InMux
    port map (
            O => \N__14228\,
            I => \N__14225\
        );

    \I__1977\ : LocalMux
    port map (
            O => \N__14225\,
            I => \N__14221\
        );

    \I__1976\ : InMux
    port map (
            O => \N__14224\,
            I => \N__14218\
        );

    \I__1975\ : Span4Mux_v
    port map (
            O => \N__14221\,
            I => \N__14215\
        );

    \I__1974\ : LocalMux
    port map (
            O => \N__14218\,
            I => \eeprom.n2313\
        );

    \I__1973\ : Odrv4
    port map (
            O => \N__14215\,
            I => \eeprom.n2313\
        );

    \I__1972\ : CascadeMux
    port map (
            O => \N__14210\,
            I => \eeprom.n2313_cascade_\
        );

    \I__1971\ : InMux
    port map (
            O => \N__14207\,
            I => \N__14204\
        );

    \I__1970\ : LocalMux
    port map (
            O => \N__14204\,
            I => \eeprom.n4505\
        );

    \I__1969\ : InMux
    port map (
            O => \N__14201\,
            I => \N__14198\
        );

    \I__1968\ : LocalMux
    port map (
            O => \N__14198\,
            I => \N__14195\
        );

    \I__1967\ : Span4Mux_h
    port map (
            O => \N__14195\,
            I => \N__14192\
        );

    \I__1966\ : Odrv4
    port map (
            O => \N__14192\,
            I => \eeprom.n11\
        );

    \I__1965\ : InMux
    port map (
            O => \N__14189\,
            I => \N__14186\
        );

    \I__1964\ : LocalMux
    port map (
            O => \N__14186\,
            I => \N__14182\
        );

    \I__1963\ : InMux
    port map (
            O => \N__14185\,
            I => \N__14179\
        );

    \I__1962\ : Span4Mux_v
    port map (
            O => \N__14182\,
            I => \N__14175\
        );

    \I__1961\ : LocalMux
    port map (
            O => \N__14179\,
            I => \N__14172\
        );

    \I__1960\ : InMux
    port map (
            O => \N__14178\,
            I => \N__14169\
        );

    \I__1959\ : Span4Mux_h
    port map (
            O => \N__14175\,
            I => \N__14164\
        );

    \I__1958\ : Span4Mux_v
    port map (
            O => \N__14172\,
            I => \N__14164\
        );

    \I__1957\ : LocalMux
    port map (
            O => \N__14169\,
            I => \eeprom.delay_counter_22\
        );

    \I__1956\ : Odrv4
    port map (
            O => \N__14164\,
            I => \eeprom.delay_counter_22\
        );

    \I__1955\ : CascadeMux
    port map (
            O => \N__14159\,
            I => \N__14156\
        );

    \I__1954\ : InMux
    port map (
            O => \N__14156\,
            I => \N__14152\
        );

    \I__1953\ : CascadeMux
    port map (
            O => \N__14155\,
            I => \N__14149\
        );

    \I__1952\ : LocalMux
    port map (
            O => \N__14152\,
            I => \N__14146\
        );

    \I__1951\ : InMux
    port map (
            O => \N__14149\,
            I => \N__14142\
        );

    \I__1950\ : Span4Mux_h
    port map (
            O => \N__14146\,
            I => \N__14139\
        );

    \I__1949\ : InMux
    port map (
            O => \N__14145\,
            I => \N__14136\
        );

    \I__1948\ : LocalMux
    port map (
            O => \N__14142\,
            I => \eeprom.n2315\
        );

    \I__1947\ : Odrv4
    port map (
            O => \N__14139\,
            I => \eeprom.n2315\
        );

    \I__1946\ : LocalMux
    port map (
            O => \N__14136\,
            I => \eeprom.n2315\
        );

    \I__1945\ : CascadeMux
    port map (
            O => \N__14129\,
            I => \N__14124\
        );

    \I__1944\ : CascadeMux
    port map (
            O => \N__14128\,
            I => \N__14121\
        );

    \I__1943\ : InMux
    port map (
            O => \N__14127\,
            I => \N__14118\
        );

    \I__1942\ : InMux
    port map (
            O => \N__14124\,
            I => \N__14115\
        );

    \I__1941\ : InMux
    port map (
            O => \N__14121\,
            I => \N__14112\
        );

    \I__1940\ : LocalMux
    port map (
            O => \N__14118\,
            I => \N__14109\
        );

    \I__1939\ : LocalMux
    port map (
            O => \N__14115\,
            I => \N__14104\
        );

    \I__1938\ : LocalMux
    port map (
            O => \N__14112\,
            I => \N__14104\
        );

    \I__1937\ : Span4Mux_s3_h
    port map (
            O => \N__14109\,
            I => \N__14099\
        );

    \I__1936\ : Span4Mux_v
    port map (
            O => \N__14104\,
            I => \N__14099\
        );

    \I__1935\ : Odrv4
    port map (
            O => \N__14099\,
            I => \eeprom.n2311\
        );

    \I__1934\ : CascadeMux
    port map (
            O => \N__14096\,
            I => \N__14093\
        );

    \I__1933\ : InMux
    port map (
            O => \N__14093\,
            I => \N__14090\
        );

    \I__1932\ : LocalMux
    port map (
            O => \N__14090\,
            I => \N__14087\
        );

    \I__1931\ : Odrv4
    port map (
            O => \N__14087\,
            I => \eeprom.n4461\
        );

    \I__1930\ : InMux
    port map (
            O => \N__14084\,
            I => \N__14081\
        );

    \I__1929\ : LocalMux
    port map (
            O => \N__14081\,
            I => \N__14078\
        );

    \I__1928\ : Odrv12
    port map (
            O => \N__14078\,
            I => \eeprom.n4463\
        );

    \I__1927\ : CascadeMux
    port map (
            O => \N__14075\,
            I => \eeprom.n4225_cascade_\
        );

    \I__1926\ : InMux
    port map (
            O => \N__14072\,
            I => \N__14069\
        );

    \I__1925\ : LocalMux
    port map (
            O => \N__14069\,
            I => \N__14065\
        );

    \I__1924\ : InMux
    port map (
            O => \N__14068\,
            I => \N__14061\
        );

    \I__1923\ : Span12Mux_s10_v
    port map (
            O => \N__14065\,
            I => \N__14058\
        );

    \I__1922\ : InMux
    port map (
            O => \N__14064\,
            I => \N__14055\
        );

    \I__1921\ : LocalMux
    port map (
            O => \N__14061\,
            I => \N__14052\
        );

    \I__1920\ : Odrv12
    port map (
            O => \N__14058\,
            I => \eeprom.n2019\
        );

    \I__1919\ : LocalMux
    port map (
            O => \N__14055\,
            I => \eeprom.n2019\
        );

    \I__1918\ : Odrv12
    port map (
            O => \N__14052\,
            I => \eeprom.n2019\
        );

    \I__1917\ : CascadeMux
    port map (
            O => \N__14045\,
            I => \N__14042\
        );

    \I__1916\ : InMux
    port map (
            O => \N__14042\,
            I => \N__14039\
        );

    \I__1915\ : LocalMux
    port map (
            O => \N__14039\,
            I => \eeprom.n2086\
        );

    \I__1914\ : InMux
    port map (
            O => \N__14036\,
            I => \N__14031\
        );

    \I__1913\ : CascadeMux
    port map (
            O => \N__14035\,
            I => \N__14028\
        );

    \I__1912\ : InMux
    port map (
            O => \N__14034\,
            I => \N__14025\
        );

    \I__1911\ : LocalMux
    port map (
            O => \N__14031\,
            I => \N__14022\
        );

    \I__1910\ : InMux
    port map (
            O => \N__14028\,
            I => \N__14019\
        );

    \I__1909\ : LocalMux
    port map (
            O => \N__14025\,
            I => \eeprom.n2309\
        );

    \I__1908\ : Odrv4
    port map (
            O => \N__14022\,
            I => \eeprom.n2309\
        );

    \I__1907\ : LocalMux
    port map (
            O => \N__14019\,
            I => \eeprom.n2309\
        );

    \I__1906\ : InMux
    port map (
            O => \N__14012\,
            I => \N__14008\
        );

    \I__1905\ : InMux
    port map (
            O => \N__14011\,
            I => \N__14005\
        );

    \I__1904\ : LocalMux
    port map (
            O => \N__14008\,
            I => \N__14001\
        );

    \I__1903\ : LocalMux
    port map (
            O => \N__14005\,
            I => \N__13998\
        );

    \I__1902\ : InMux
    port map (
            O => \N__14004\,
            I => \N__13995\
        );

    \I__1901\ : Odrv4
    port map (
            O => \N__14001\,
            I => \eeprom.n2319\
        );

    \I__1900\ : Odrv4
    port map (
            O => \N__13998\,
            I => \eeprom.n2319\
        );

    \I__1899\ : LocalMux
    port map (
            O => \N__13995\,
            I => \eeprom.n2319\
        );

    \I__1898\ : CascadeMux
    port map (
            O => \N__13988\,
            I => \eeprom.n4509_cascade_\
        );

    \I__1897\ : InMux
    port map (
            O => \N__13985\,
            I => \N__13982\
        );

    \I__1896\ : LocalMux
    port map (
            O => \N__13982\,
            I => \eeprom.n8_adj_468\
        );

    \I__1895\ : InMux
    port map (
            O => \N__13979\,
            I => \N__13975\
        );

    \I__1894\ : InMux
    port map (
            O => \N__13978\,
            I => \N__13971\
        );

    \I__1893\ : LocalMux
    port map (
            O => \N__13975\,
            I => \N__13968\
        );

    \I__1892\ : InMux
    port map (
            O => \N__13974\,
            I => \N__13965\
        );

    \I__1891\ : LocalMux
    port map (
            O => \N__13971\,
            I => \eeprom.n2310\
        );

    \I__1890\ : Odrv4
    port map (
            O => \N__13968\,
            I => \eeprom.n2310\
        );

    \I__1889\ : LocalMux
    port map (
            O => \N__13965\,
            I => \eeprom.n2310\
        );

    \I__1888\ : CascadeMux
    port map (
            O => \N__13958\,
            I => \eeprom.n6_cascade_\
        );

    \I__1887\ : CascadeMux
    port map (
            O => \N__13955\,
            I => \eeprom.n2242_cascade_\
        );

    \I__1886\ : InMux
    port map (
            O => \N__13952\,
            I => \N__13946\
        );

    \I__1885\ : CascadeMux
    port map (
            O => \N__13951\,
            I => \N__13943\
        );

    \I__1884\ : CascadeMux
    port map (
            O => \N__13950\,
            I => \N__13940\
        );

    \I__1883\ : CascadeMux
    port map (
            O => \N__13949\,
            I => \N__13932\
        );

    \I__1882\ : LocalMux
    port map (
            O => \N__13946\,
            I => \N__13928\
        );

    \I__1881\ : InMux
    port map (
            O => \N__13943\,
            I => \N__13917\
        );

    \I__1880\ : InMux
    port map (
            O => \N__13940\,
            I => \N__13917\
        );

    \I__1879\ : InMux
    port map (
            O => \N__13939\,
            I => \N__13917\
        );

    \I__1878\ : InMux
    port map (
            O => \N__13938\,
            I => \N__13917\
        );

    \I__1877\ : InMux
    port map (
            O => \N__13937\,
            I => \N__13917\
        );

    \I__1876\ : InMux
    port map (
            O => \N__13936\,
            I => \N__13908\
        );

    \I__1875\ : InMux
    port map (
            O => \N__13935\,
            I => \N__13908\
        );

    \I__1874\ : InMux
    port map (
            O => \N__13932\,
            I => \N__13908\
        );

    \I__1873\ : InMux
    port map (
            O => \N__13931\,
            I => \N__13908\
        );

    \I__1872\ : Odrv4
    port map (
            O => \N__13928\,
            I => \eeprom.n2044\
        );

    \I__1871\ : LocalMux
    port map (
            O => \N__13917\,
            I => \eeprom.n2044\
        );

    \I__1870\ : LocalMux
    port map (
            O => \N__13908\,
            I => \eeprom.n2044\
        );

    \I__1869\ : InMux
    port map (
            O => \N__13901\,
            I => \N__13898\
        );

    \I__1868\ : LocalMux
    port map (
            O => \N__13898\,
            I => \N__13894\
        );

    \I__1867\ : InMux
    port map (
            O => \N__13897\,
            I => \N__13891\
        );

    \I__1866\ : Odrv4
    port map (
            O => \N__13894\,
            I => \eeprom.n2084\
        );

    \I__1865\ : LocalMux
    port map (
            O => \N__13891\,
            I => \eeprom.n2084\
        );

    \I__1864\ : CascadeMux
    port map (
            O => \N__13886\,
            I => \N__13881\
        );

    \I__1863\ : CascadeMux
    port map (
            O => \N__13885\,
            I => \N__13878\
        );

    \I__1862\ : InMux
    port map (
            O => \N__13884\,
            I => \N__13875\
        );

    \I__1861\ : InMux
    port map (
            O => \N__13881\,
            I => \N__13872\
        );

    \I__1860\ : InMux
    port map (
            O => \N__13878\,
            I => \N__13869\
        );

    \I__1859\ : LocalMux
    port map (
            O => \N__13875\,
            I => \eeprom.n2013\
        );

    \I__1858\ : LocalMux
    port map (
            O => \N__13872\,
            I => \eeprom.n2013\
        );

    \I__1857\ : LocalMux
    port map (
            O => \N__13869\,
            I => \eeprom.n2013\
        );

    \I__1856\ : CascadeMux
    port map (
            O => \N__13862\,
            I => \N__13859\
        );

    \I__1855\ : InMux
    port map (
            O => \N__13859\,
            I => \N__13856\
        );

    \I__1854\ : LocalMux
    port map (
            O => \N__13856\,
            I => \eeprom.n2080\
        );

    \I__1853\ : InMux
    port map (
            O => \N__13853\,
            I => \eeprom.n3529\
        );

    \I__1852\ : InMux
    port map (
            O => \N__13850\,
            I => \eeprom.n3530\
        );

    \I__1851\ : InMux
    port map (
            O => \N__13847\,
            I => \N__13844\
        );

    \I__1850\ : LocalMux
    port map (
            O => \N__13844\,
            I => \N__13840\
        );

    \I__1849\ : InMux
    port map (
            O => \N__13843\,
            I => \N__13837\
        );

    \I__1848\ : Span4Mux_v
    port map (
            O => \N__13840\,
            I => \N__13834\
        );

    \I__1847\ : LocalMux
    port map (
            O => \N__13837\,
            I => \N__13831\
        );

    \I__1846\ : Odrv4
    port map (
            O => \N__13834\,
            I => \eeprom.n2011\
        );

    \I__1845\ : Odrv4
    port map (
            O => \N__13831\,
            I => \eeprom.n2011\
        );

    \I__1844\ : InMux
    port map (
            O => \N__13826\,
            I => \bfn_5_23_0_\
        );

    \I__1843\ : InMux
    port map (
            O => \N__13823\,
            I => \N__13820\
        );

    \I__1842\ : LocalMux
    port map (
            O => \N__13820\,
            I => \eeprom.n2081\
        );

    \I__1841\ : CascadeMux
    port map (
            O => \N__13817\,
            I => \N__13814\
        );

    \I__1840\ : InMux
    port map (
            O => \N__13814\,
            I => \N__13810\
        );

    \I__1839\ : CascadeMux
    port map (
            O => \N__13813\,
            I => \N__13807\
        );

    \I__1838\ : LocalMux
    port map (
            O => \N__13810\,
            I => \N__13804\
        );

    \I__1837\ : InMux
    port map (
            O => \N__13807\,
            I => \N__13801\
        );

    \I__1836\ : Odrv4
    port map (
            O => \N__13804\,
            I => \eeprom.n2014\
        );

    \I__1835\ : LocalMux
    port map (
            O => \N__13801\,
            I => \eeprom.n2014\
        );

    \I__1834\ : InMux
    port map (
            O => \N__13796\,
            I => \N__13793\
        );

    \I__1833\ : LocalMux
    port map (
            O => \N__13793\,
            I => \N__13788\
        );

    \I__1832\ : InMux
    port map (
            O => \N__13792\,
            I => \N__13785\
        );

    \I__1831\ : InMux
    port map (
            O => \N__13791\,
            I => \N__13782\
        );

    \I__1830\ : Span4Mux_h
    port map (
            O => \N__13788\,
            I => \N__13777\
        );

    \I__1829\ : LocalMux
    port map (
            O => \N__13785\,
            I => \N__13777\
        );

    \I__1828\ : LocalMux
    port map (
            O => \N__13782\,
            I => \eeprom.n2012\
        );

    \I__1827\ : Odrv4
    port map (
            O => \N__13777\,
            I => \eeprom.n2012\
        );

    \I__1826\ : InMux
    port map (
            O => \N__13772\,
            I => \N__13769\
        );

    \I__1825\ : LocalMux
    port map (
            O => \N__13769\,
            I => \eeprom.n2079\
        );

    \I__1824\ : InMux
    port map (
            O => \N__13766\,
            I => \N__13763\
        );

    \I__1823\ : LocalMux
    port map (
            O => \N__13763\,
            I => \eeprom.n2083\
        );

    \I__1822\ : CascadeMux
    port map (
            O => \N__13760\,
            I => \N__13757\
        );

    \I__1821\ : InMux
    port map (
            O => \N__13757\,
            I => \N__13753\
        );

    \I__1820\ : CascadeMux
    port map (
            O => \N__13756\,
            I => \N__13750\
        );

    \I__1819\ : LocalMux
    port map (
            O => \N__13753\,
            I => \N__13747\
        );

    \I__1818\ : InMux
    port map (
            O => \N__13750\,
            I => \N__13744\
        );

    \I__1817\ : Span4Mux_v
    port map (
            O => \N__13747\,
            I => \N__13738\
        );

    \I__1816\ : LocalMux
    port map (
            O => \N__13744\,
            I => \N__13738\
        );

    \I__1815\ : InMux
    port map (
            O => \N__13743\,
            I => \N__13735\
        );

    \I__1814\ : Odrv4
    port map (
            O => \N__13738\,
            I => \eeprom.n2016\
        );

    \I__1813\ : LocalMux
    port map (
            O => \N__13735\,
            I => \eeprom.n2016\
        );

    \I__1812\ : InMux
    port map (
            O => \N__13730\,
            I => \N__13727\
        );

    \I__1811\ : LocalMux
    port map (
            O => \N__13727\,
            I => \eeprom.n7_adj_470\
        );

    \I__1810\ : InMux
    port map (
            O => \N__13724\,
            I => \N__13721\
        );

    \I__1809\ : LocalMux
    port map (
            O => \N__13721\,
            I => \N__13716\
        );

    \I__1808\ : InMux
    port map (
            O => \N__13720\,
            I => \N__13713\
        );

    \I__1807\ : InMux
    port map (
            O => \N__13719\,
            I => \N__13710\
        );

    \I__1806\ : Span4Mux_v
    port map (
            O => \N__13716\,
            I => \N__13705\
        );

    \I__1805\ : LocalMux
    port map (
            O => \N__13713\,
            I => \N__13705\
        );

    \I__1804\ : LocalMux
    port map (
            O => \N__13710\,
            I => \N__13702\
        );

    \I__1803\ : Span4Mux_h
    port map (
            O => \N__13705\,
            I => \N__13699\
        );

    \I__1802\ : Odrv4
    port map (
            O => \N__13702\,
            I => \eeprom.n2419\
        );

    \I__1801\ : Odrv4
    port map (
            O => \N__13699\,
            I => \eeprom.n2419\
        );

    \I__1800\ : InMux
    port map (
            O => \N__13694\,
            I => \N__13691\
        );

    \I__1799\ : LocalMux
    port map (
            O => \N__13691\,
            I => \N__13688\
        );

    \I__1798\ : Span4Mux_v
    port map (
            O => \N__13688\,
            I => \N__13685\
        );

    \I__1797\ : Odrv4
    port map (
            O => \N__13685\,
            I => \eeprom.n2486\
        );

    \I__1796\ : InMux
    port map (
            O => \N__13682\,
            I => \bfn_5_22_0_\
        );

    \I__1795\ : CascadeMux
    port map (
            O => \N__13679\,
            I => \N__13675\
        );

    \I__1794\ : InMux
    port map (
            O => \N__13678\,
            I => \N__13671\
        );

    \I__1793\ : InMux
    port map (
            O => \N__13675\,
            I => \N__13668\
        );

    \I__1792\ : InMux
    port map (
            O => \N__13674\,
            I => \N__13665\
        );

    \I__1791\ : LocalMux
    port map (
            O => \N__13671\,
            I => \eeprom.n2018\
        );

    \I__1790\ : LocalMux
    port map (
            O => \N__13668\,
            I => \eeprom.n2018\
        );

    \I__1789\ : LocalMux
    port map (
            O => \N__13665\,
            I => \eeprom.n2018\
        );

    \I__1788\ : CascadeMux
    port map (
            O => \N__13658\,
            I => \N__13655\
        );

    \I__1787\ : InMux
    port map (
            O => \N__13655\,
            I => \N__13652\
        );

    \I__1786\ : LocalMux
    port map (
            O => \N__13652\,
            I => \eeprom.n2085\
        );

    \I__1785\ : InMux
    port map (
            O => \N__13649\,
            I => \eeprom.n3524\
        );

    \I__1784\ : InMux
    port map (
            O => \N__13646\,
            I => \eeprom.n3525\
        );

    \I__1783\ : InMux
    port map (
            O => \N__13643\,
            I => \eeprom.n3526\
        );

    \I__1782\ : CascadeMux
    port map (
            O => \N__13640\,
            I => \N__13637\
        );

    \I__1781\ : InMux
    port map (
            O => \N__13637\,
            I => \N__13633\
        );

    \I__1780\ : InMux
    port map (
            O => \N__13636\,
            I => \N__13629\
        );

    \I__1779\ : LocalMux
    port map (
            O => \N__13633\,
            I => \N__13626\
        );

    \I__1778\ : InMux
    port map (
            O => \N__13632\,
            I => \N__13623\
        );

    \I__1777\ : LocalMux
    port map (
            O => \N__13629\,
            I => \eeprom.n2015\
        );

    \I__1776\ : Odrv4
    port map (
            O => \N__13626\,
            I => \eeprom.n2015\
        );

    \I__1775\ : LocalMux
    port map (
            O => \N__13623\,
            I => \eeprom.n2015\
        );

    \I__1774\ : CascadeMux
    port map (
            O => \N__13616\,
            I => \N__13613\
        );

    \I__1773\ : InMux
    port map (
            O => \N__13613\,
            I => \N__13610\
        );

    \I__1772\ : LocalMux
    port map (
            O => \N__13610\,
            I => \eeprom.n2082\
        );

    \I__1771\ : InMux
    port map (
            O => \N__13607\,
            I => \eeprom.n3527\
        );

    \I__1770\ : InMux
    port map (
            O => \N__13604\,
            I => \eeprom.n3528\
        );

    \I__1769\ : CascadeMux
    port map (
            O => \N__13601\,
            I => \eeprom.n13_adj_474_cascade_\
        );

    \I__1768\ : InMux
    port map (
            O => \N__13598\,
            I => \N__13595\
        );

    \I__1767\ : LocalMux
    port map (
            O => \N__13595\,
            I => \eeprom.n11_adj_473\
        );

    \I__1766\ : CascadeMux
    port map (
            O => \N__13592\,
            I => \eeprom.n2539_cascade_\
        );

    \I__1765\ : InMux
    port map (
            O => \N__13589\,
            I => \N__13586\
        );

    \I__1764\ : LocalMux
    port map (
            O => \N__13586\,
            I => \N__13581\
        );

    \I__1763\ : InMux
    port map (
            O => \N__13585\,
            I => \N__13578\
        );

    \I__1762\ : InMux
    port map (
            O => \N__13584\,
            I => \N__13575\
        );

    \I__1761\ : Span4Mux_h
    port map (
            O => \N__13581\,
            I => \N__13570\
        );

    \I__1760\ : LocalMux
    port map (
            O => \N__13578\,
            I => \N__13570\
        );

    \I__1759\ : LocalMux
    port map (
            O => \N__13575\,
            I => \N__13565\
        );

    \I__1758\ : Span4Mux_v
    port map (
            O => \N__13570\,
            I => \N__13565\
        );

    \I__1757\ : Odrv4
    port map (
            O => \N__13565\,
            I => \eeprom.delay_counter_14\
        );

    \I__1756\ : CascadeMux
    port map (
            O => \N__13562\,
            I => \N__13559\
        );

    \I__1755\ : InMux
    port map (
            O => \N__13559\,
            I => \N__13556\
        );

    \I__1754\ : LocalMux
    port map (
            O => \N__13556\,
            I => \N__13553\
        );

    \I__1753\ : Span4Mux_h
    port map (
            O => \N__13553\,
            I => \N__13550\
        );

    \I__1752\ : Odrv4
    port map (
            O => \N__13550\,
            I => \eeprom.n19_adj_429\
        );

    \I__1751\ : InMux
    port map (
            O => \N__13547\,
            I => \N__13544\
        );

    \I__1750\ : LocalMux
    port map (
            O => \N__13544\,
            I => \N__13541\
        );

    \I__1749\ : Odrv12
    port map (
            O => \N__13541\,
            I => \eeprom.n30\
        );

    \I__1748\ : CascadeMux
    port map (
            O => \N__13538\,
            I => \eeprom.n2114_cascade_\
        );

    \I__1747\ : InMux
    port map (
            O => \N__13535\,
            I => \N__13532\
        );

    \I__1746\ : LocalMux
    port map (
            O => \N__13532\,
            I => \N__13528\
        );

    \I__1745\ : InMux
    port map (
            O => \N__13531\,
            I => \N__13525\
        );

    \I__1744\ : Span4Mux_v
    port map (
            O => \N__13528\,
            I => \N__13520\
        );

    \I__1743\ : LocalMux
    port map (
            O => \N__13525\,
            I => \N__13520\
        );

    \I__1742\ : Odrv4
    port map (
            O => \N__13520\,
            I => \eeprom.n2411\
        );

    \I__1741\ : InMux
    port map (
            O => \N__13517\,
            I => \N__13514\
        );

    \I__1740\ : LocalMux
    port map (
            O => \N__13514\,
            I => \N__13511\
        );

    \I__1739\ : Span4Mux_v
    port map (
            O => \N__13511\,
            I => \N__13508\
        );

    \I__1738\ : Odrv4
    port map (
            O => \N__13508\,
            I => \eeprom.n2478\
        );

    \I__1737\ : InMux
    port map (
            O => \N__13505\,
            I => \N__13502\
        );

    \I__1736\ : LocalMux
    port map (
            O => \N__13502\,
            I => n4826
        );

    \I__1735\ : CascadeMux
    port map (
            O => \N__13499\,
            I => \n4825_cascade_\
        );

    \I__1734\ : IoInMux
    port map (
            O => \N__13496\,
            I => \N__13493\
        );

    \I__1733\ : LocalMux
    port map (
            O => \N__13493\,
            I => \N__13490\
        );

    \I__1732\ : Odrv4
    port map (
            O => \N__13490\,
            I => \LED_c\
        );

    \I__1731\ : InMux
    port map (
            O => \N__13487\,
            I => \N__13484\
        );

    \I__1730\ : LocalMux
    port map (
            O => \N__13484\,
            I => \N__13481\
        );

    \I__1729\ : Span4Mux_h
    port map (
            O => \N__13481\,
            I => \N__13478\
        );

    \I__1728\ : Odrv4
    port map (
            O => \N__13478\,
            I => \eeprom.n23_adj_464\
        );

    \I__1727\ : InMux
    port map (
            O => \N__13475\,
            I => \N__13471\
        );

    \I__1726\ : InMux
    port map (
            O => \N__13474\,
            I => \N__13467\
        );

    \I__1725\ : LocalMux
    port map (
            O => \N__13471\,
            I => \N__13464\
        );

    \I__1724\ : InMux
    port map (
            O => \N__13470\,
            I => \N__13461\
        );

    \I__1723\ : LocalMux
    port map (
            O => \N__13467\,
            I => \eeprom.delay_counter_10\
        );

    \I__1722\ : Odrv4
    port map (
            O => \N__13464\,
            I => \eeprom.delay_counter_10\
        );

    \I__1721\ : LocalMux
    port map (
            O => \N__13461\,
            I => \eeprom.delay_counter_10\
        );

    \I__1720\ : CascadeMux
    port map (
            O => \N__13454\,
            I => \eeprom.n2615_cascade_\
        );

    \I__1719\ : CascadeMux
    port map (
            O => \N__13451\,
            I => \eeprom.n4497_cascade_\
        );

    \I__1718\ : CascadeMux
    port map (
            O => \N__13448\,
            I => \eeprom.n4501_cascade_\
        );

    \I__1717\ : InMux
    port map (
            O => \N__13445\,
            I => \bfn_4_26_0_\
        );

    \I__1716\ : InMux
    port map (
            O => \N__13442\,
            I => \eeprom.n3570\
        );

    \I__1715\ : InMux
    port map (
            O => \N__13439\,
            I => \eeprom.n3571\
        );

    \I__1714\ : InMux
    port map (
            O => \N__13436\,
            I => \eeprom.n3572\
        );

    \I__1713\ : InMux
    port map (
            O => \N__13433\,
            I => \N__13430\
        );

    \I__1712\ : LocalMux
    port map (
            O => \N__13430\,
            I => \N__13426\
        );

    \I__1711\ : InMux
    port map (
            O => \N__13429\,
            I => \N__13423\
        );

    \I__1710\ : Odrv4
    port map (
            O => \N__13426\,
            I => \eeprom.n2407\
        );

    \I__1709\ : LocalMux
    port map (
            O => \N__13423\,
            I => \eeprom.n2407\
        );

    \I__1708\ : InMux
    port map (
            O => \N__13418\,
            I => \eeprom.n3573\
        );

    \I__1707\ : InMux
    port map (
            O => \N__13415\,
            I => \N__13408\
        );

    \I__1706\ : InMux
    port map (
            O => \N__13414\,
            I => \N__13408\
        );

    \I__1705\ : InMux
    port map (
            O => \N__13413\,
            I => \N__13405\
        );

    \I__1704\ : LocalMux
    port map (
            O => \N__13408\,
            I => \eeprom.n2410\
        );

    \I__1703\ : LocalMux
    port map (
            O => \N__13405\,
            I => \eeprom.n2410\
        );

    \I__1702\ : CascadeMux
    port map (
            O => \N__13400\,
            I => \N__13397\
        );

    \I__1701\ : InMux
    port map (
            O => \N__13397\,
            I => \N__13394\
        );

    \I__1700\ : LocalMux
    port map (
            O => \N__13394\,
            I => \eeprom.n2477\
        );

    \I__1699\ : InMux
    port map (
            O => \N__13391\,
            I => \N__13388\
        );

    \I__1698\ : LocalMux
    port map (
            O => \N__13388\,
            I => \eeprom.n2476\
        );

    \I__1697\ : CascadeMux
    port map (
            O => \N__13385\,
            I => \N__13382\
        );

    \I__1696\ : InMux
    port map (
            O => \N__13382\,
            I => \N__13376\
        );

    \I__1695\ : InMux
    port map (
            O => \N__13381\,
            I => \N__13376\
        );

    \I__1694\ : LocalMux
    port map (
            O => \N__13376\,
            I => \N__13372\
        );

    \I__1693\ : InMux
    port map (
            O => \N__13375\,
            I => \N__13369\
        );

    \I__1692\ : Odrv4
    port map (
            O => \N__13372\,
            I => \eeprom.n2409\
        );

    \I__1691\ : LocalMux
    port map (
            O => \N__13369\,
            I => \eeprom.n2409\
        );

    \I__1690\ : InMux
    port map (
            O => \N__13364\,
            I => \bfn_4_25_0_\
        );

    \I__1689\ : CascadeMux
    port map (
            O => \N__13361\,
            I => \N__13356\
        );

    \I__1688\ : InMux
    port map (
            O => \N__13360\,
            I => \N__13351\
        );

    \I__1687\ : InMux
    port map (
            O => \N__13359\,
            I => \N__13351\
        );

    \I__1686\ : InMux
    port map (
            O => \N__13356\,
            I => \N__13348\
        );

    \I__1685\ : LocalMux
    port map (
            O => \N__13351\,
            I => \eeprom.n2418\
        );

    \I__1684\ : LocalMux
    port map (
            O => \N__13348\,
            I => \eeprom.n2418\
        );

    \I__1683\ : CascadeMux
    port map (
            O => \N__13343\,
            I => \N__13340\
        );

    \I__1682\ : InMux
    port map (
            O => \N__13340\,
            I => \N__13337\
        );

    \I__1681\ : LocalMux
    port map (
            O => \N__13337\,
            I => \N__13334\
        );

    \I__1680\ : Odrv4
    port map (
            O => \N__13334\,
            I => \eeprom.n2485\
        );

    \I__1679\ : InMux
    port map (
            O => \N__13331\,
            I => \eeprom.n3562\
        );

    \I__1678\ : CascadeMux
    port map (
            O => \N__13328\,
            I => \N__13325\
        );

    \I__1677\ : InMux
    port map (
            O => \N__13325\,
            I => \N__13321\
        );

    \I__1676\ : InMux
    port map (
            O => \N__13324\,
            I => \N__13317\
        );

    \I__1675\ : LocalMux
    port map (
            O => \N__13321\,
            I => \N__13314\
        );

    \I__1674\ : InMux
    port map (
            O => \N__13320\,
            I => \N__13311\
        );

    \I__1673\ : LocalMux
    port map (
            O => \N__13317\,
            I => \eeprom.n2417\
        );

    \I__1672\ : Odrv4
    port map (
            O => \N__13314\,
            I => \eeprom.n2417\
        );

    \I__1671\ : LocalMux
    port map (
            O => \N__13311\,
            I => \eeprom.n2417\
        );

    \I__1670\ : CascadeMux
    port map (
            O => \N__13304\,
            I => \N__13301\
        );

    \I__1669\ : InMux
    port map (
            O => \N__13301\,
            I => \N__13298\
        );

    \I__1668\ : LocalMux
    port map (
            O => \N__13298\,
            I => \N__13295\
        );

    \I__1667\ : Odrv4
    port map (
            O => \N__13295\,
            I => \eeprom.n2484\
        );

    \I__1666\ : InMux
    port map (
            O => \N__13292\,
            I => \eeprom.n3563\
        );

    \I__1665\ : CascadeMux
    port map (
            O => \N__13289\,
            I => \N__13285\
        );

    \I__1664\ : CascadeMux
    port map (
            O => \N__13288\,
            I => \N__13281\
        );

    \I__1663\ : InMux
    port map (
            O => \N__13285\,
            I => \N__13278\
        );

    \I__1662\ : InMux
    port map (
            O => \N__13284\,
            I => \N__13273\
        );

    \I__1661\ : InMux
    port map (
            O => \N__13281\,
            I => \N__13273\
        );

    \I__1660\ : LocalMux
    port map (
            O => \N__13278\,
            I => \eeprom.n2416\
        );

    \I__1659\ : LocalMux
    port map (
            O => \N__13273\,
            I => \eeprom.n2416\
        );

    \I__1658\ : InMux
    port map (
            O => \N__13268\,
            I => \N__13265\
        );

    \I__1657\ : LocalMux
    port map (
            O => \N__13265\,
            I => \N__13262\
        );

    \I__1656\ : Odrv4
    port map (
            O => \N__13262\,
            I => \eeprom.n2483\
        );

    \I__1655\ : InMux
    port map (
            O => \N__13259\,
            I => \eeprom.n3564\
        );

    \I__1654\ : InMux
    port map (
            O => \N__13256\,
            I => \N__13251\
        );

    \I__1653\ : CascadeMux
    port map (
            O => \N__13255\,
            I => \N__13248\
        );

    \I__1652\ : InMux
    port map (
            O => \N__13254\,
            I => \N__13245\
        );

    \I__1651\ : LocalMux
    port map (
            O => \N__13251\,
            I => \N__13242\
        );

    \I__1650\ : InMux
    port map (
            O => \N__13248\,
            I => \N__13239\
        );

    \I__1649\ : LocalMux
    port map (
            O => \N__13245\,
            I => \eeprom.n2415\
        );

    \I__1648\ : Odrv4
    port map (
            O => \N__13242\,
            I => \eeprom.n2415\
        );

    \I__1647\ : LocalMux
    port map (
            O => \N__13239\,
            I => \eeprom.n2415\
        );

    \I__1646\ : CascadeMux
    port map (
            O => \N__13232\,
            I => \N__13229\
        );

    \I__1645\ : InMux
    port map (
            O => \N__13229\,
            I => \N__13226\
        );

    \I__1644\ : LocalMux
    port map (
            O => \N__13226\,
            I => \N__13223\
        );

    \I__1643\ : Odrv4
    port map (
            O => \N__13223\,
            I => \eeprom.n2482\
        );

    \I__1642\ : InMux
    port map (
            O => \N__13220\,
            I => \eeprom.n3565\
        );

    \I__1641\ : CascadeMux
    port map (
            O => \N__13217\,
            I => \N__13213\
        );

    \I__1640\ : CascadeMux
    port map (
            O => \N__13216\,
            I => \N__13210\
        );

    \I__1639\ : InMux
    port map (
            O => \N__13213\,
            I => \N__13206\
        );

    \I__1638\ : InMux
    port map (
            O => \N__13210\,
            I => \N__13201\
        );

    \I__1637\ : InMux
    port map (
            O => \N__13209\,
            I => \N__13201\
        );

    \I__1636\ : LocalMux
    port map (
            O => \N__13206\,
            I => \eeprom.n2414\
        );

    \I__1635\ : LocalMux
    port map (
            O => \N__13201\,
            I => \eeprom.n2414\
        );

    \I__1634\ : InMux
    port map (
            O => \N__13196\,
            I => \N__13193\
        );

    \I__1633\ : LocalMux
    port map (
            O => \N__13193\,
            I => \N__13190\
        );

    \I__1632\ : Odrv4
    port map (
            O => \N__13190\,
            I => \eeprom.n2481\
        );

    \I__1631\ : InMux
    port map (
            O => \N__13187\,
            I => \eeprom.n3566\
        );

    \I__1630\ : InMux
    port map (
            O => \N__13184\,
            I => \eeprom.n3567\
        );

    \I__1629\ : InMux
    port map (
            O => \N__13181\,
            I => \eeprom.n3568\
        );

    \I__1628\ : InMux
    port map (
            O => \N__13178\,
            I => \N__13175\
        );

    \I__1627\ : LocalMux
    port map (
            O => \N__13175\,
            I => \eeprom.n2376\
        );

    \I__1626\ : InMux
    port map (
            O => \N__13172\,
            I => \N__13168\
        );

    \I__1625\ : InMux
    port map (
            O => \N__13171\,
            I => \N__13165\
        );

    \I__1624\ : LocalMux
    port map (
            O => \N__13168\,
            I => \eeprom.n2312\
        );

    \I__1623\ : LocalMux
    port map (
            O => \N__13165\,
            I => \eeprom.n2312\
        );

    \I__1622\ : CascadeMux
    port map (
            O => \N__13160\,
            I => \eeprom.n2312_cascade_\
        );

    \I__1621\ : InMux
    port map (
            O => \N__13157\,
            I => \N__13154\
        );

    \I__1620\ : LocalMux
    port map (
            O => \N__13154\,
            I => \eeprom.n2379\
        );

    \I__1619\ : CascadeMux
    port map (
            O => \N__13151\,
            I => \eeprom.n2411_cascade_\
        );

    \I__1618\ : InMux
    port map (
            O => \N__13148\,
            I => \N__13145\
        );

    \I__1617\ : LocalMux
    port map (
            O => \N__13145\,
            I => \eeprom.n4133\
        );

    \I__1616\ : CascadeMux
    port map (
            O => \N__13142\,
            I => \eeprom.n12_adj_472_cascade_\
        );

    \I__1615\ : InMux
    port map (
            O => \N__13139\,
            I => \N__13136\
        );

    \I__1614\ : LocalMux
    port map (
            O => \N__13136\,
            I => \eeprom.n2382\
        );

    \I__1613\ : InMux
    port map (
            O => \N__13133\,
            I => \N__13130\
        );

    \I__1612\ : LocalMux
    port map (
            O => \N__13130\,
            I => \eeprom.n2377\
        );

    \I__1611\ : CascadeMux
    port map (
            O => \N__13127\,
            I => \N__13124\
        );

    \I__1610\ : InMux
    port map (
            O => \N__13124\,
            I => \N__13121\
        );

    \I__1609\ : LocalMux
    port map (
            O => \N__13121\,
            I => \eeprom.n2380\
        );

    \I__1608\ : InMux
    port map (
            O => \N__13118\,
            I => \N__13110\
        );

    \I__1607\ : CascadeMux
    port map (
            O => \N__13117\,
            I => \N__13107\
        );

    \I__1606\ : CascadeMux
    port map (
            O => \N__13116\,
            I => \N__13104\
        );

    \I__1605\ : CascadeMux
    port map (
            O => \N__13115\,
            I => \N__13097\
        );

    \I__1604\ : CascadeMux
    port map (
            O => \N__13114\,
            I => \N__13094\
        );

    \I__1603\ : CascadeMux
    port map (
            O => \N__13113\,
            I => \N__13091\
        );

    \I__1602\ : LocalMux
    port map (
            O => \N__13110\,
            I => \N__13087\
        );

    \I__1601\ : InMux
    port map (
            O => \N__13107\,
            I => \N__13076\
        );

    \I__1600\ : InMux
    port map (
            O => \N__13104\,
            I => \N__13076\
        );

    \I__1599\ : InMux
    port map (
            O => \N__13103\,
            I => \N__13076\
        );

    \I__1598\ : InMux
    port map (
            O => \N__13102\,
            I => \N__13076\
        );

    \I__1597\ : InMux
    port map (
            O => \N__13101\,
            I => \N__13076\
        );

    \I__1596\ : InMux
    port map (
            O => \N__13100\,
            I => \N__13073\
        );

    \I__1595\ : InMux
    port map (
            O => \N__13097\,
            I => \N__13064\
        );

    \I__1594\ : InMux
    port map (
            O => \N__13094\,
            I => \N__13064\
        );

    \I__1593\ : InMux
    port map (
            O => \N__13091\,
            I => \N__13064\
        );

    \I__1592\ : InMux
    port map (
            O => \N__13090\,
            I => \N__13064\
        );

    \I__1591\ : Odrv4
    port map (
            O => \N__13087\,
            I => \eeprom.n2341\
        );

    \I__1590\ : LocalMux
    port map (
            O => \N__13076\,
            I => \eeprom.n2341\
        );

    \I__1589\ : LocalMux
    port map (
            O => \N__13073\,
            I => \eeprom.n2341\
        );

    \I__1588\ : LocalMux
    port map (
            O => \N__13064\,
            I => \eeprom.n2341\
        );

    \I__1587\ : InMux
    port map (
            O => \N__13055\,
            I => \N__13052\
        );

    \I__1586\ : LocalMux
    port map (
            O => \N__13052\,
            I => \N__13047\
        );

    \I__1585\ : InMux
    port map (
            O => \N__13051\,
            I => \N__13044\
        );

    \I__1584\ : InMux
    port map (
            O => \N__13050\,
            I => \N__13041\
        );

    \I__1583\ : Span4Mux_h
    port map (
            O => \N__13047\,
            I => \N__13036\
        );

    \I__1582\ : LocalMux
    port map (
            O => \N__13044\,
            I => \N__13036\
        );

    \I__1581\ : LocalMux
    port map (
            O => \N__13041\,
            I => \eeprom.delay_counter_20\
        );

    \I__1580\ : Odrv4
    port map (
            O => \N__13036\,
            I => \eeprom.delay_counter_20\
        );

    \I__1579\ : CascadeMux
    port map (
            O => \N__13031\,
            I => \eeprom.n4479_cascade_\
        );

    \I__1578\ : InMux
    port map (
            O => \N__13028\,
            I => \N__13025\
        );

    \I__1577\ : LocalMux
    port map (
            O => \N__13025\,
            I => \eeprom.n4477\
        );

    \I__1576\ : InMux
    port map (
            O => \N__13022\,
            I => \N__13019\
        );

    \I__1575\ : LocalMux
    port map (
            O => \N__13019\,
            I => \eeprom.n2385\
        );

    \I__1574\ : CascadeMux
    port map (
            O => \N__13016\,
            I => \eeprom.n2341_cascade_\
        );

    \I__1573\ : InMux
    port map (
            O => \N__13013\,
            I => \N__13010\
        );

    \I__1572\ : LocalMux
    port map (
            O => \N__13010\,
            I => \N__13006\
        );

    \I__1571\ : InMux
    port map (
            O => \N__13009\,
            I => \N__13003\
        );

    \I__1570\ : Odrv12
    port map (
            O => \N__13006\,
            I => \eeprom.n1915\
        );

    \I__1569\ : LocalMux
    port map (
            O => \N__13003\,
            I => \eeprom.n1915\
        );

    \I__1568\ : CascadeMux
    port map (
            O => \N__12998\,
            I => \N__12995\
        );

    \I__1567\ : InMux
    port map (
            O => \N__12995\,
            I => \N__12992\
        );

    \I__1566\ : LocalMux
    port map (
            O => \N__12992\,
            I => \N__12989\
        );

    \I__1565\ : Odrv4
    port map (
            O => \N__12989\,
            I => \eeprom.n1982\
        );

    \I__1564\ : CascadeMux
    port map (
            O => \N__12986\,
            I => \eeprom.n2014_cascade_\
        );

    \I__1563\ : InMux
    port map (
            O => \N__12983\,
            I => \N__12980\
        );

    \I__1562\ : LocalMux
    port map (
            O => \N__12980\,
            I => \eeprom.n4415\
        );

    \I__1561\ : InMux
    port map (
            O => \N__12977\,
            I => \N__12972\
        );

    \I__1560\ : InMux
    port map (
            O => \N__12976\,
            I => \N__12969\
        );

    \I__1559\ : InMux
    port map (
            O => \N__12975\,
            I => \N__12966\
        );

    \I__1558\ : LocalMux
    port map (
            O => \N__12972\,
            I => \eeprom.n1919\
        );

    \I__1557\ : LocalMux
    port map (
            O => \N__12969\,
            I => \eeprom.n1919\
        );

    \I__1556\ : LocalMux
    port map (
            O => \N__12966\,
            I => \eeprom.n1919\
        );

    \I__1555\ : CascadeMux
    port map (
            O => \N__12959\,
            I => \N__12956\
        );

    \I__1554\ : InMux
    port map (
            O => \N__12956\,
            I => \N__12953\
        );

    \I__1553\ : LocalMux
    port map (
            O => \N__12953\,
            I => \N__12950\
        );

    \I__1552\ : Odrv4
    port map (
            O => \N__12950\,
            I => \eeprom.n1986\
        );

    \I__1551\ : InMux
    port map (
            O => \N__12947\,
            I => \N__12943\
        );

    \I__1550\ : CascadeMux
    port map (
            O => \N__12946\,
            I => \N__12940\
        );

    \I__1549\ : LocalMux
    port map (
            O => \N__12943\,
            I => \N__12937\
        );

    \I__1548\ : InMux
    port map (
            O => \N__12940\,
            I => \N__12934\
        );

    \I__1547\ : Odrv4
    port map (
            O => \N__12937\,
            I => \eeprom.n1913\
        );

    \I__1546\ : LocalMux
    port map (
            O => \N__12934\,
            I => \eeprom.n1913\
        );

    \I__1545\ : CascadeMux
    port map (
            O => \N__12929\,
            I => \N__12923\
        );

    \I__1544\ : CascadeMux
    port map (
            O => \N__12928\,
            I => \N__12920\
        );

    \I__1543\ : CascadeMux
    port map (
            O => \N__12927\,
            I => \N__12917\
        );

    \I__1542\ : CascadeMux
    port map (
            O => \N__12926\,
            I => \N__12912\
        );

    \I__1541\ : InMux
    port map (
            O => \N__12923\,
            I => \N__12908\
        );

    \I__1540\ : InMux
    port map (
            O => \N__12920\,
            I => \N__12899\
        );

    \I__1539\ : InMux
    port map (
            O => \N__12917\,
            I => \N__12899\
        );

    \I__1538\ : InMux
    port map (
            O => \N__12916\,
            I => \N__12899\
        );

    \I__1537\ : InMux
    port map (
            O => \N__12915\,
            I => \N__12899\
        );

    \I__1536\ : InMux
    port map (
            O => \N__12912\,
            I => \N__12894\
        );

    \I__1535\ : InMux
    port map (
            O => \N__12911\,
            I => \N__12894\
        );

    \I__1534\ : LocalMux
    port map (
            O => \N__12908\,
            I => \eeprom.n1945\
        );

    \I__1533\ : LocalMux
    port map (
            O => \N__12899\,
            I => \eeprom.n1945\
        );

    \I__1532\ : LocalMux
    port map (
            O => \N__12894\,
            I => \eeprom.n1945\
        );

    \I__1531\ : InMux
    port map (
            O => \N__12887\,
            I => \N__12884\
        );

    \I__1530\ : LocalMux
    port map (
            O => \N__12884\,
            I => \N__12881\
        );

    \I__1529\ : Odrv4
    port map (
            O => \N__12881\,
            I => \eeprom.n1980\
        );

    \I__1528\ : InMux
    port map (
            O => \N__12878\,
            I => \N__12875\
        );

    \I__1527\ : LocalMux
    port map (
            O => \N__12875\,
            I => \eeprom.n4419\
        );

    \I__1526\ : CascadeMux
    port map (
            O => \N__12872\,
            I => \eeprom.n4575_cascade_\
        );

    \I__1525\ : InMux
    port map (
            O => \N__12869\,
            I => \N__12866\
        );

    \I__1524\ : LocalMux
    port map (
            O => \N__12866\,
            I => \eeprom.n4579\
        );

    \I__1523\ : InMux
    port map (
            O => \N__12863\,
            I => \N__12860\
        );

    \I__1522\ : LocalMux
    port map (
            O => \N__12860\,
            I => \N__12857\
        );

    \I__1521\ : Span4Mux_h
    port map (
            O => \N__12857\,
            I => \N__12854\
        );

    \I__1520\ : Odrv4
    port map (
            O => \N__12854\,
            I => \eeprom.n13\
        );

    \I__1519\ : InMux
    port map (
            O => \N__12851\,
            I => \eeprom.n3523\
        );

    \I__1518\ : InMux
    port map (
            O => \N__12848\,
            I => \N__12845\
        );

    \I__1517\ : LocalMux
    port map (
            O => \N__12845\,
            I => \N__12842\
        );

    \I__1516\ : Span4Mux_v
    port map (
            O => \N__12842\,
            I => \N__12839\
        );

    \I__1515\ : Odrv4
    port map (
            O => \N__12839\,
            I => \eeprom.n26_adj_469\
        );

    \I__1514\ : InMux
    port map (
            O => \N__12836\,
            I => \N__12833\
        );

    \I__1513\ : LocalMux
    port map (
            O => \N__12833\,
            I => \N__12829\
        );

    \I__1512\ : InMux
    port map (
            O => \N__12832\,
            I => \N__12825\
        );

    \I__1511\ : Span4Mux_v
    port map (
            O => \N__12829\,
            I => \N__12822\
        );

    \I__1510\ : InMux
    port map (
            O => \N__12828\,
            I => \N__12819\
        );

    \I__1509\ : LocalMux
    port map (
            O => \N__12825\,
            I => \eeprom.delay_counter_7\
        );

    \I__1508\ : Odrv4
    port map (
            O => \N__12822\,
            I => \eeprom.delay_counter_7\
        );

    \I__1507\ : LocalMux
    port map (
            O => \N__12819\,
            I => \eeprom.delay_counter_7\
        );

    \I__1506\ : CascadeMux
    port map (
            O => \N__12812\,
            I => \N__12809\
        );

    \I__1505\ : InMux
    port map (
            O => \N__12809\,
            I => \N__12806\
        );

    \I__1504\ : LocalMux
    port map (
            O => \N__12806\,
            I => \eeprom.n1984\
        );

    \I__1503\ : InMux
    port map (
            O => \N__12803\,
            I => \N__12800\
        );

    \I__1502\ : LocalMux
    port map (
            O => \N__12800\,
            I => \eeprom.n1985\
        );

    \I__1501\ : CascadeMux
    port map (
            O => \N__12797\,
            I => \eeprom.n2017_cascade_\
        );

    \I__1500\ : CascadeMux
    port map (
            O => \N__12794\,
            I => \N__12789\
        );

    \I__1499\ : InMux
    port map (
            O => \N__12793\,
            I => \N__12784\
        );

    \I__1498\ : InMux
    port map (
            O => \N__12792\,
            I => \N__12784\
        );

    \I__1497\ : InMux
    port map (
            O => \N__12789\,
            I => \N__12781\
        );

    \I__1496\ : LocalMux
    port map (
            O => \N__12784\,
            I => \eeprom.n1917\
        );

    \I__1495\ : LocalMux
    port map (
            O => \N__12781\,
            I => \eeprom.n1917\
        );

    \I__1494\ : InMux
    port map (
            O => \N__12776\,
            I => \N__12773\
        );

    \I__1493\ : LocalMux
    port map (
            O => \N__12773\,
            I => \N__12770\
        );

    \I__1492\ : Odrv4
    port map (
            O => \N__12770\,
            I => \eeprom.n4437\
        );

    \I__1491\ : CascadeMux
    port map (
            O => \N__12767\,
            I => \N__12762\
        );

    \I__1490\ : InMux
    port map (
            O => \N__12766\,
            I => \N__12759\
        );

    \I__1489\ : InMux
    port map (
            O => \N__12765\,
            I => \N__12756\
        );

    \I__1488\ : InMux
    port map (
            O => \N__12762\,
            I => \N__12753\
        );

    \I__1487\ : LocalMux
    port map (
            O => \N__12759\,
            I => \eeprom.n1918\
        );

    \I__1486\ : LocalMux
    port map (
            O => \N__12756\,
            I => \eeprom.n1918\
        );

    \I__1485\ : LocalMux
    port map (
            O => \N__12753\,
            I => \eeprom.n1918\
        );

    \I__1484\ : CascadeMux
    port map (
            O => \N__12746\,
            I => \eeprom.n4441_cascade_\
        );

    \I__1483\ : InMux
    port map (
            O => \N__12743\,
            I => \N__12739\
        );

    \I__1482\ : InMux
    port map (
            O => \N__12742\,
            I => \N__12736\
        );

    \I__1481\ : LocalMux
    port map (
            O => \N__12739\,
            I => \N__12733\
        );

    \I__1480\ : LocalMux
    port map (
            O => \N__12736\,
            I => \eeprom.n1912\
        );

    \I__1479\ : Odrv4
    port map (
            O => \N__12733\,
            I => \eeprom.n1912\
        );

    \I__1478\ : CascadeMux
    port map (
            O => \N__12728\,
            I => \N__12723\
        );

    \I__1477\ : CascadeMux
    port map (
            O => \N__12727\,
            I => \N__12720\
        );

    \I__1476\ : InMux
    port map (
            O => \N__12726\,
            I => \N__12715\
        );

    \I__1475\ : InMux
    port map (
            O => \N__12723\,
            I => \N__12715\
        );

    \I__1474\ : InMux
    port map (
            O => \N__12720\,
            I => \N__12712\
        );

    \I__1473\ : LocalMux
    port map (
            O => \N__12715\,
            I => \N__12709\
        );

    \I__1472\ : LocalMux
    port map (
            O => \N__12712\,
            I => \eeprom.n1916\
        );

    \I__1471\ : Odrv4
    port map (
            O => \N__12709\,
            I => \eeprom.n1916\
        );

    \I__1470\ : CascadeMux
    port map (
            O => \N__12704\,
            I => \eeprom.n1945_cascade_\
        );

    \I__1469\ : InMux
    port map (
            O => \N__12701\,
            I => \N__12698\
        );

    \I__1468\ : LocalMux
    port map (
            O => \N__12698\,
            I => \eeprom.n1983\
        );

    \I__1467\ : InMux
    port map (
            O => \N__12695\,
            I => \N__12692\
        );

    \I__1466\ : LocalMux
    port map (
            O => \N__12692\,
            I => \N__12689\
        );

    \I__1465\ : Odrv4
    port map (
            O => \N__12689\,
            I => \eeprom.n1981\
        );

    \I__1464\ : CascadeMux
    port map (
            O => \N__12686\,
            I => \N__12682\
        );

    \I__1463\ : InMux
    port map (
            O => \N__12685\,
            I => \N__12678\
        );

    \I__1462\ : InMux
    port map (
            O => \N__12682\,
            I => \N__12675\
        );

    \I__1461\ : InMux
    port map (
            O => \N__12681\,
            I => \N__12672\
        );

    \I__1460\ : LocalMux
    port map (
            O => \N__12678\,
            I => \eeprom.n1914\
        );

    \I__1459\ : LocalMux
    port map (
            O => \N__12675\,
            I => \eeprom.n1914\
        );

    \I__1458\ : LocalMux
    port map (
            O => \N__12672\,
            I => \eeprom.n1914\
        );

    \I__1457\ : InMux
    port map (
            O => \N__12665\,
            I => \N__12662\
        );

    \I__1456\ : LocalMux
    port map (
            O => \N__12662\,
            I => \N__12657\
        );

    \I__1455\ : InMux
    port map (
            O => \N__12661\,
            I => \N__12654\
        );

    \I__1454\ : InMux
    port map (
            O => \N__12660\,
            I => \N__12651\
        );

    \I__1453\ : Span4Mux_v
    port map (
            O => \N__12657\,
            I => \N__12648\
        );

    \I__1452\ : LocalMux
    port map (
            O => \N__12654\,
            I => \N__12645\
        );

    \I__1451\ : LocalMux
    port map (
            O => \N__12651\,
            I => \N__12638\
        );

    \I__1450\ : Span4Mux_h
    port map (
            O => \N__12648\,
            I => \N__12638\
        );

    \I__1449\ : Span4Mux_v
    port map (
            O => \N__12645\,
            I => \N__12638\
        );

    \I__1448\ : Odrv4
    port map (
            O => \N__12638\,
            I => \eeprom.delay_counter_17\
        );

    \I__1447\ : InMux
    port map (
            O => \N__12635\,
            I => \N__12632\
        );

    \I__1446\ : LocalMux
    port map (
            O => \N__12632\,
            I => \N__12629\
        );

    \I__1445\ : Span4Mux_v
    port map (
            O => \N__12629\,
            I => \N__12626\
        );

    \I__1444\ : Span4Mux_v
    port map (
            O => \N__12626\,
            I => \N__12623\
        );

    \I__1443\ : Odrv4
    port map (
            O => \N__12623\,
            I => \eeprom.n16_adj_377\
        );

    \I__1442\ : CascadeMux
    port map (
            O => \N__12620\,
            I => \N__12617\
        );

    \I__1441\ : InMux
    port map (
            O => \N__12617\,
            I => \N__12611\
        );

    \I__1440\ : InMux
    port map (
            O => \N__12616\,
            I => \N__12611\
        );

    \I__1439\ : LocalMux
    port map (
            O => \N__12611\,
            I => \eeprom.n4734\
        );

    \I__1438\ : InMux
    port map (
            O => \N__12608\,
            I => \N__12602\
        );

    \I__1437\ : CascadeMux
    port map (
            O => \N__12607\,
            I => \N__12595\
        );

    \I__1436\ : InMux
    port map (
            O => \N__12606\,
            I => \N__12590\
        );

    \I__1435\ : InMux
    port map (
            O => \N__12605\,
            I => \N__12590\
        );

    \I__1434\ : LocalMux
    port map (
            O => \N__12602\,
            I => \N__12587\
        );

    \I__1433\ : InMux
    port map (
            O => \N__12601\,
            I => \N__12578\
        );

    \I__1432\ : InMux
    port map (
            O => \N__12600\,
            I => \N__12578\
        );

    \I__1431\ : InMux
    port map (
            O => \N__12599\,
            I => \N__12578\
        );

    \I__1430\ : InMux
    port map (
            O => \N__12598\,
            I => \N__12578\
        );

    \I__1429\ : InMux
    port map (
            O => \N__12595\,
            I => \N__12575\
        );

    \I__1428\ : LocalMux
    port map (
            O => \N__12590\,
            I => \eeprom.n1256\
        );

    \I__1427\ : Odrv4
    port map (
            O => \N__12587\,
            I => \eeprom.n1256\
        );

    \I__1426\ : LocalMux
    port map (
            O => \N__12578\,
            I => \eeprom.n1256\
        );

    \I__1425\ : LocalMux
    port map (
            O => \N__12575\,
            I => \eeprom.n1256\
        );

    \I__1424\ : InMux
    port map (
            O => \N__12566\,
            I => \bfn_4_19_0_\
        );

    \I__1423\ : InMux
    port map (
            O => \N__12563\,
            I => \eeprom.n3517\
        );

    \I__1422\ : InMux
    port map (
            O => \N__12560\,
            I => \eeprom.n3518\
        );

    \I__1421\ : InMux
    port map (
            O => \N__12557\,
            I => \eeprom.n3519\
        );

    \I__1420\ : InMux
    port map (
            O => \N__12554\,
            I => \eeprom.n3520\
        );

    \I__1419\ : InMux
    port map (
            O => \N__12551\,
            I => \eeprom.n3521\
        );

    \I__1418\ : InMux
    port map (
            O => \N__12548\,
            I => \eeprom.n3522\
        );

    \I__1417\ : InMux
    port map (
            O => \N__12545\,
            I => \N__12542\
        );

    \I__1416\ : LocalMux
    port map (
            O => \N__12542\,
            I => \eeprom.n2381\
        );

    \I__1415\ : InMux
    port map (
            O => \N__12539\,
            I => \N__12536\
        );

    \I__1414\ : LocalMux
    port map (
            O => \N__12536\,
            I => \eeprom.n2384\
        );

    \I__1413\ : CascadeMux
    port map (
            O => \N__12533\,
            I => \N__12530\
        );

    \I__1412\ : InMux
    port map (
            O => \N__12530\,
            I => \N__12527\
        );

    \I__1411\ : LocalMux
    port map (
            O => \N__12527\,
            I => \eeprom.n2378\
        );

    \I__1410\ : InMux
    port map (
            O => \N__12524\,
            I => \N__12521\
        );

    \I__1409\ : LocalMux
    port map (
            O => \N__12521\,
            I => \eeprom.n4733\
        );

    \I__1408\ : InMux
    port map (
            O => \N__12518\,
            I => \N__12515\
        );

    \I__1407\ : LocalMux
    port map (
            O => \N__12515\,
            I => \eeprom.n1340\
        );

    \I__1406\ : InMux
    port map (
            O => \N__12512\,
            I => \N__12508\
        );

    \I__1405\ : InMux
    port map (
            O => \N__12511\,
            I => \N__12504\
        );

    \I__1404\ : LocalMux
    port map (
            O => \N__12508\,
            I => \N__12501\
        );

    \I__1403\ : InMux
    port map (
            O => \N__12507\,
            I => \N__12498\
        );

    \I__1402\ : LocalMux
    port map (
            O => \N__12504\,
            I => \eeprom.n1138\
        );

    \I__1401\ : Odrv4
    port map (
            O => \N__12501\,
            I => \eeprom.n1138\
        );

    \I__1400\ : LocalMux
    port map (
            O => \N__12498\,
            I => \eeprom.n1138\
        );

    \I__1399\ : CascadeMux
    port map (
            O => \N__12491\,
            I => \eeprom.n1915_cascade_\
        );

    \I__1398\ : CascadeMux
    port map (
            O => \N__12488\,
            I => \N__12484\
        );

    \I__1397\ : InMux
    port map (
            O => \N__12487\,
            I => \N__12481\
        );

    \I__1396\ : InMux
    port map (
            O => \N__12484\,
            I => \N__12478\
        );

    \I__1395\ : LocalMux
    port map (
            O => \N__12481\,
            I => \eeprom.n1135\
        );

    \I__1394\ : LocalMux
    port map (
            O => \N__12478\,
            I => \eeprom.n1135\
        );

    \I__1393\ : CascadeMux
    port map (
            O => \N__12473\,
            I => \N__12467\
        );

    \I__1392\ : CascadeMux
    port map (
            O => \N__12472\,
            I => \N__12463\
        );

    \I__1391\ : CascadeMux
    port map (
            O => \N__12471\,
            I => \N__12460\
        );

    \I__1390\ : InMux
    port map (
            O => \N__12470\,
            I => \N__12456\
        );

    \I__1389\ : InMux
    port map (
            O => \N__12467\,
            I => \N__12453\
        );

    \I__1388\ : InMux
    port map (
            O => \N__12466\,
            I => \N__12450\
        );

    \I__1387\ : InMux
    port map (
            O => \N__12463\,
            I => \N__12443\
        );

    \I__1386\ : InMux
    port map (
            O => \N__12460\,
            I => \N__12443\
        );

    \I__1385\ : InMux
    port map (
            O => \N__12459\,
            I => \N__12443\
        );

    \I__1384\ : LocalMux
    port map (
            O => \N__12456\,
            I => \eeprom.n4405\
        );

    \I__1383\ : LocalMux
    port map (
            O => \N__12453\,
            I => \eeprom.n4405\
        );

    \I__1382\ : LocalMux
    port map (
            O => \N__12450\,
            I => \eeprom.n4405\
        );

    \I__1381\ : LocalMux
    port map (
            O => \N__12443\,
            I => \eeprom.n4405\
        );

    \I__1380\ : InMux
    port map (
            O => \N__12434\,
            I => \N__12431\
        );

    \I__1379\ : LocalMux
    port map (
            O => \N__12431\,
            I => \eeprom.n1337\
        );

    \I__1378\ : CascadeMux
    port map (
            O => \N__12428\,
            I => \N__12425\
        );

    \I__1377\ : InMux
    port map (
            O => \N__12425\,
            I => \N__12422\
        );

    \I__1376\ : LocalMux
    port map (
            O => \N__12422\,
            I => \N__12419\
        );

    \I__1375\ : Span4Mux_v
    port map (
            O => \N__12419\,
            I => \N__12416\
        );

    \I__1374\ : Span4Mux_v
    port map (
            O => \N__12416\,
            I => \N__12413\
        );

    \I__1373\ : Odrv4
    port map (
            O => \N__12413\,
            I => \eeprom.n12_adj_411\
        );

    \I__1372\ : InMux
    port map (
            O => \N__12410\,
            I => \N__12407\
        );

    \I__1371\ : LocalMux
    port map (
            O => \N__12407\,
            I => \N__12404\
        );

    \I__1370\ : Span12Mux_h
    port map (
            O => \N__12404\,
            I => \N__12401\
        );

    \I__1369\ : Odrv12
    port map (
            O => \N__12401\,
            I => \eeprom.n25_adj_471\
        );

    \I__1368\ : InMux
    port map (
            O => \N__12398\,
            I => \N__12394\
        );

    \I__1367\ : InMux
    port map (
            O => \N__12397\,
            I => \N__12390\
        );

    \I__1366\ : LocalMux
    port map (
            O => \N__12394\,
            I => \N__12387\
        );

    \I__1365\ : InMux
    port map (
            O => \N__12393\,
            I => \N__12384\
        );

    \I__1364\ : LocalMux
    port map (
            O => \N__12390\,
            I => \eeprom.delay_counter_8\
        );

    \I__1363\ : Odrv4
    port map (
            O => \N__12387\,
            I => \eeprom.delay_counter_8\
        );

    \I__1362\ : LocalMux
    port map (
            O => \N__12384\,
            I => \eeprom.delay_counter_8\
        );

    \I__1361\ : InMux
    port map (
            O => \N__12377\,
            I => \eeprom.n3554\
        );

    \I__1360\ : InMux
    port map (
            O => \N__12374\,
            I => \eeprom.n3555\
        );

    \I__1359\ : InMux
    port map (
            O => \N__12371\,
            I => \eeprom.n3556\
        );

    \I__1358\ : InMux
    port map (
            O => \N__12368\,
            I => \eeprom.n3557\
        );

    \I__1357\ : InMux
    port map (
            O => \N__12365\,
            I => \bfn_3_24_0_\
        );

    \I__1356\ : InMux
    port map (
            O => \N__12362\,
            I => \eeprom.n3559\
        );

    \I__1355\ : InMux
    port map (
            O => \N__12359\,
            I => \eeprom.n3560\
        );

    \I__1354\ : InMux
    port map (
            O => \N__12356\,
            I => \eeprom.n3561\
        );

    \I__1353\ : InMux
    port map (
            O => \N__12353\,
            I => \N__12350\
        );

    \I__1352\ : LocalMux
    port map (
            O => \N__12350\,
            I => \N__12347\
        );

    \I__1351\ : Odrv4
    port map (
            O => \N__12347\,
            I => \eeprom.n2386\
        );

    \I__1350\ : InMux
    port map (
            O => \N__12344\,
            I => \N__12341\
        );

    \I__1349\ : LocalMux
    port map (
            O => \N__12341\,
            I => \eeprom.n19_adj_428\
        );

    \I__1348\ : InMux
    port map (
            O => \N__12338\,
            I => \N__12335\
        );

    \I__1347\ : LocalMux
    port map (
            O => \N__12335\,
            I => \N__12331\
        );

    \I__1346\ : InMux
    port map (
            O => \N__12334\,
            I => \N__12327\
        );

    \I__1345\ : Span4Mux_v
    port map (
            O => \N__12331\,
            I => \N__12324\
        );

    \I__1344\ : InMux
    port map (
            O => \N__12330\,
            I => \N__12321\
        );

    \I__1343\ : LocalMux
    port map (
            O => \N__12327\,
            I => \eeprom.delay_counter_18\
        );

    \I__1342\ : Odrv4
    port map (
            O => \N__12324\,
            I => \eeprom.delay_counter_18\
        );

    \I__1341\ : LocalMux
    port map (
            O => \N__12321\,
            I => \eeprom.delay_counter_18\
        );

    \I__1340\ : InMux
    port map (
            O => \N__12314\,
            I => \N__12311\
        );

    \I__1339\ : LocalMux
    port map (
            O => \N__12311\,
            I => \eeprom.n15_adj_414\
        );

    \I__1338\ : InMux
    port map (
            O => \N__12308\,
            I => \N__12303\
        );

    \I__1337\ : InMux
    port map (
            O => \N__12307\,
            I => \N__12300\
        );

    \I__1336\ : InMux
    port map (
            O => \N__12306\,
            I => \N__12297\
        );

    \I__1335\ : LocalMux
    port map (
            O => \N__12303\,
            I => \N__12292\
        );

    \I__1334\ : LocalMux
    port map (
            O => \N__12300\,
            I => \N__12292\
        );

    \I__1333\ : LocalMux
    port map (
            O => \N__12297\,
            I => \eeprom.delay_counter_23\
        );

    \I__1332\ : Odrv4
    port map (
            O => \N__12292\,
            I => \eeprom.delay_counter_23\
        );

    \I__1331\ : InMux
    port map (
            O => \N__12287\,
            I => \N__12284\
        );

    \I__1330\ : LocalMux
    port map (
            O => \N__12284\,
            I => \eeprom.n10\
        );

    \I__1329\ : InMux
    port map (
            O => \N__12281\,
            I => \N__12278\
        );

    \I__1328\ : LocalMux
    port map (
            O => \N__12278\,
            I => \eeprom.n18_adj_426\
        );

    \I__1327\ : InMux
    port map (
            O => \N__12275\,
            I => \N__12272\
        );

    \I__1326\ : LocalMux
    port map (
            O => \N__12272\,
            I => \N__12268\
        );

    \I__1325\ : InMux
    port map (
            O => \N__12271\,
            I => \N__12264\
        );

    \I__1324\ : Span12Mux_v
    port map (
            O => \N__12268\,
            I => \N__12261\
        );

    \I__1323\ : InMux
    port map (
            O => \N__12267\,
            I => \N__12258\
        );

    \I__1322\ : LocalMux
    port map (
            O => \N__12264\,
            I => \eeprom.delay_counter_15\
        );

    \I__1321\ : Odrv12
    port map (
            O => \N__12261\,
            I => \eeprom.delay_counter_15\
        );

    \I__1320\ : LocalMux
    port map (
            O => \N__12258\,
            I => \eeprom.delay_counter_15\
        );

    \I__1319\ : InMux
    port map (
            O => \N__12251\,
            I => \bfn_3_23_0_\
        );

    \I__1318\ : InMux
    port map (
            O => \N__12248\,
            I => \eeprom.n3551\
        );

    \I__1317\ : InMux
    port map (
            O => \N__12245\,
            I => \eeprom.n3552\
        );

    \I__1316\ : CascadeMux
    port map (
            O => \N__12242\,
            I => \N__12239\
        );

    \I__1315\ : InMux
    port map (
            O => \N__12239\,
            I => \N__12236\
        );

    \I__1314\ : LocalMux
    port map (
            O => \N__12236\,
            I => \eeprom.n2383\
        );

    \I__1313\ : InMux
    port map (
            O => \N__12233\,
            I => \eeprom.n3553\
        );

    \I__1312\ : CascadeMux
    port map (
            O => \N__12230\,
            I => \N__12225\
        );

    \I__1311\ : InMux
    port map (
            O => \N__12229\,
            I => \N__12222\
        );

    \I__1310\ : InMux
    port map (
            O => \N__12228\,
            I => \N__12219\
        );

    \I__1309\ : InMux
    port map (
            O => \N__12225\,
            I => \N__12216\
        );

    \I__1308\ : LocalMux
    port map (
            O => \N__12222\,
            I => \eeprom.delay_counter_26\
        );

    \I__1307\ : LocalMux
    port map (
            O => \N__12219\,
            I => \eeprom.delay_counter_26\
        );

    \I__1306\ : LocalMux
    port map (
            O => \N__12216\,
            I => \eeprom.delay_counter_26\
        );

    \I__1305\ : CascadeMux
    port map (
            O => \N__12209\,
            I => \N__12206\
        );

    \I__1304\ : InMux
    port map (
            O => \N__12206\,
            I => \N__12202\
        );

    \I__1303\ : InMux
    port map (
            O => \N__12205\,
            I => \N__12199\
        );

    \I__1302\ : LocalMux
    port map (
            O => \N__12202\,
            I => \N__12194\
        );

    \I__1301\ : LocalMux
    port map (
            O => \N__12199\,
            I => \N__12194\
        );

    \I__1300\ : Span4Mux_v
    port map (
            O => \N__12194\,
            I => \N__12191\
        );

    \I__1299\ : Odrv4
    port map (
            O => \N__12191\,
            I => \eeprom.n7\
        );

    \I__1298\ : CascadeMux
    port map (
            O => \N__12188\,
            I => \N__12184\
        );

    \I__1297\ : InMux
    port map (
            O => \N__12187\,
            I => \N__12181\
        );

    \I__1296\ : InMux
    port map (
            O => \N__12184\,
            I => \N__12178\
        );

    \I__1295\ : LocalMux
    port map (
            O => \N__12181\,
            I => \N__12175\
        );

    \I__1294\ : LocalMux
    port map (
            O => \N__12178\,
            I => \N__12172\
        );

    \I__1293\ : Odrv4
    port map (
            O => \N__12175\,
            I => \eeprom.n1140\
        );

    \I__1292\ : Odrv4
    port map (
            O => \N__12172\,
            I => \eeprom.n1140\
        );

    \I__1291\ : InMux
    port map (
            O => \N__12167\,
            I => \N__12162\
        );

    \I__1290\ : InMux
    port map (
            O => \N__12166\,
            I => \N__12159\
        );

    \I__1289\ : InMux
    port map (
            O => \N__12165\,
            I => \N__12156\
        );

    \I__1288\ : LocalMux
    port map (
            O => \N__12162\,
            I => \eeprom.delay_counter_29\
        );

    \I__1287\ : LocalMux
    port map (
            O => \N__12159\,
            I => \eeprom.delay_counter_29\
        );

    \I__1286\ : LocalMux
    port map (
            O => \N__12156\,
            I => \eeprom.delay_counter_29\
        );

    \I__1285\ : InMux
    port map (
            O => \N__12149\,
            I => \N__12146\
        );

    \I__1284\ : LocalMux
    port map (
            O => \N__12146\,
            I => \N__12143\
        );

    \I__1283\ : Span4Mux_h
    port map (
            O => \N__12143\,
            I => \N__12140\
        );

    \I__1282\ : Odrv4
    port map (
            O => \N__12140\,
            I => \eeprom.n4\
        );

    \I__1281\ : CascadeMux
    port map (
            O => \N__12137\,
            I => \N__12134\
        );

    \I__1280\ : InMux
    port map (
            O => \N__12134\,
            I => \N__12131\
        );

    \I__1279\ : LocalMux
    port map (
            O => \N__12131\,
            I => \N__12127\
        );

    \I__1278\ : InMux
    port map (
            O => \N__12130\,
            I => \N__12124\
        );

    \I__1277\ : Odrv4
    port map (
            O => \N__12127\,
            I => \eeprom.n1137\
        );

    \I__1276\ : LocalMux
    port map (
            O => \N__12124\,
            I => \eeprom.n1137\
        );

    \I__1275\ : InMux
    port map (
            O => \N__12119\,
            I => \N__12116\
        );

    \I__1274\ : LocalMux
    port map (
            O => \N__12116\,
            I => \N__12113\
        );

    \I__1273\ : Odrv4
    port map (
            O => \N__12113\,
            I => \eeprom.n1339\
        );

    \I__1272\ : CascadeMux
    port map (
            O => \N__12110\,
            I => \eeprom.n1137_cascade_\
        );

    \I__1271\ : InMux
    port map (
            O => \N__12107\,
            I => \N__12104\
        );

    \I__1270\ : LocalMux
    port map (
            O => \N__12104\,
            I => \N__12101\
        );

    \I__1269\ : Span4Mux_h
    port map (
            O => \N__12101\,
            I => \N__12098\
        );

    \I__1268\ : Odrv4
    port map (
            O => \N__12098\,
            I => \eeprom.n24_adj_467\
        );

    \I__1267\ : InMux
    port map (
            O => \N__12095\,
            I => \N__12091\
        );

    \I__1266\ : InMux
    port map (
            O => \N__12094\,
            I => \N__12087\
        );

    \I__1265\ : LocalMux
    port map (
            O => \N__12091\,
            I => \N__12084\
        );

    \I__1264\ : InMux
    port map (
            O => \N__12090\,
            I => \N__12081\
        );

    \I__1263\ : LocalMux
    port map (
            O => \N__12087\,
            I => \eeprom.delay_counter_9\
        );

    \I__1262\ : Odrv4
    port map (
            O => \N__12084\,
            I => \eeprom.delay_counter_9\
        );

    \I__1261\ : LocalMux
    port map (
            O => \N__12081\,
            I => \eeprom.delay_counter_9\
        );

    \I__1260\ : InMux
    port map (
            O => \N__12074\,
            I => \N__12071\
        );

    \I__1259\ : LocalMux
    port map (
            O => \N__12071\,
            I => \eeprom.n33_adj_483\
        );

    \I__1258\ : CascadeMux
    port map (
            O => \N__12068\,
            I => \N__12065\
        );

    \I__1257\ : InMux
    port map (
            O => \N__12065\,
            I => \N__12062\
        );

    \I__1256\ : LocalMux
    port map (
            O => \N__12062\,
            I => \N__12059\
        );

    \I__1255\ : Odrv4
    port map (
            O => \N__12059\,
            I => \eeprom.n13_adj_412\
        );

    \I__1254\ : CascadeMux
    port map (
            O => \N__12056\,
            I => \N__12053\
        );

    \I__1253\ : InMux
    port map (
            O => \N__12053\,
            I => \N__12050\
        );

    \I__1252\ : LocalMux
    port map (
            O => \N__12050\,
            I => \N__12047\
        );

    \I__1251\ : Odrv4
    port map (
            O => \N__12047\,
            I => \eeprom.n10_adj_409\
        );

    \I__1250\ : InMux
    port map (
            O => \N__12044\,
            I => \N__12040\
        );

    \I__1249\ : InMux
    port map (
            O => \N__12043\,
            I => \N__12037\
        );

    \I__1248\ : LocalMux
    port map (
            O => \N__12040\,
            I => \N__12034\
        );

    \I__1247\ : LocalMux
    port map (
            O => \N__12037\,
            I => \N__12031\
        );

    \I__1246\ : Span4Mux_v
    port map (
            O => \N__12034\,
            I => \N__12028\
        );

    \I__1245\ : Span4Mux_v
    port map (
            O => \N__12031\,
            I => \N__12025\
        );

    \I__1244\ : Odrv4
    port map (
            O => \N__12028\,
            I => \eeprom.n2_adj_395\
        );

    \I__1243\ : Odrv4
    port map (
            O => \N__12025\,
            I => \eeprom.n2_adj_395\
        );

    \I__1242\ : CascadeMux
    port map (
            O => \N__12020\,
            I => \eeprom.n4399_cascade_\
        );

    \I__1241\ : InMux
    port map (
            O => \N__12017\,
            I => \N__12014\
        );

    \I__1240\ : LocalMux
    port map (
            O => \N__12014\,
            I => \N__12011\
        );

    \I__1239\ : Odrv4
    port map (
            O => \N__12011\,
            I => \eeprom.n1343\
        );

    \I__1238\ : CascadeMux
    port map (
            O => \N__12008\,
            I => \N__12005\
        );

    \I__1237\ : InMux
    port map (
            O => \N__12005\,
            I => \N__12001\
        );

    \I__1236\ : InMux
    port map (
            O => \N__12004\,
            I => \N__11998\
        );

    \I__1235\ : LocalMux
    port map (
            O => \N__12001\,
            I => \N__11995\
        );

    \I__1234\ : LocalMux
    port map (
            O => \N__11998\,
            I => \eeprom.n1141\
        );

    \I__1233\ : Odrv4
    port map (
            O => \N__11995\,
            I => \eeprom.n1141\
        );

    \I__1232\ : CascadeMux
    port map (
            O => \N__11990\,
            I => \eeprom.n4405_cascade_\
        );

    \I__1231\ : InMux
    port map (
            O => \N__11987\,
            I => \N__11984\
        );

    \I__1230\ : LocalMux
    port map (
            O => \N__11984\,
            I => \N__11979\
        );

    \I__1229\ : InMux
    port map (
            O => \N__11983\,
            I => \N__11976\
        );

    \I__1228\ : InMux
    port map (
            O => \N__11982\,
            I => \N__11973\
        );

    \I__1227\ : Span4Mux_v
    port map (
            O => \N__11979\,
            I => \N__11970\
        );

    \I__1226\ : LocalMux
    port map (
            O => \N__11976\,
            I => \N__11967\
        );

    \I__1225\ : LocalMux
    port map (
            O => \N__11973\,
            I => \eeprom.delay_counter_28\
        );

    \I__1224\ : Odrv4
    port map (
            O => \N__11970\,
            I => \eeprom.delay_counter_28\
        );

    \I__1223\ : Odrv4
    port map (
            O => \N__11967\,
            I => \eeprom.delay_counter_28\
        );

    \I__1222\ : InMux
    port map (
            O => \N__11960\,
            I => \N__11957\
        );

    \I__1221\ : LocalMux
    port map (
            O => \N__11957\,
            I => \N__11954\
        );

    \I__1220\ : Span4Mux_v
    port map (
            O => \N__11954\,
            I => \N__11951\
        );

    \I__1219\ : Odrv4
    port map (
            O => \N__11951\,
            I => \eeprom.n5\
        );

    \I__1218\ : InMux
    port map (
            O => \N__11948\,
            I => \N__11945\
        );

    \I__1217\ : LocalMux
    port map (
            O => \N__11945\,
            I => \N__11942\
        );

    \I__1216\ : Odrv4
    port map (
            O => \N__11942\,
            I => \eeprom.n1342\
        );

    \I__1215\ : CascadeMux
    port map (
            O => \N__11939\,
            I => \N__11936\
        );

    \I__1214\ : InMux
    port map (
            O => \N__11936\,
            I => \N__11930\
        );

    \I__1213\ : InMux
    port map (
            O => \N__11935\,
            I => \N__11930\
        );

    \I__1212\ : LocalMux
    port map (
            O => \N__11930\,
            I => \N__11927\
        );

    \I__1211\ : Span4Mux_v
    port map (
            O => \N__11927\,
            I => \N__11924\
        );

    \I__1210\ : Odrv4
    port map (
            O => \N__11924\,
            I => \eeprom.n6_adj_402\
        );

    \I__1209\ : InMux
    port map (
            O => \N__11921\,
            I => \N__11916\
        );

    \I__1208\ : InMux
    port map (
            O => \N__11920\,
            I => \N__11913\
        );

    \I__1207\ : InMux
    port map (
            O => \N__11919\,
            I => \N__11910\
        );

    \I__1206\ : LocalMux
    port map (
            O => \N__11916\,
            I => \eeprom.delay_counter_27\
        );

    \I__1205\ : LocalMux
    port map (
            O => \N__11913\,
            I => \eeprom.delay_counter_27\
        );

    \I__1204\ : LocalMux
    port map (
            O => \N__11910\,
            I => \eeprom.delay_counter_27\
        );

    \I__1203\ : InMux
    port map (
            O => \N__11903\,
            I => \N__11899\
        );

    \I__1202\ : InMux
    port map (
            O => \N__11902\,
            I => \N__11896\
        );

    \I__1201\ : LocalMux
    port map (
            O => \N__11899\,
            I => \N__11893\
        );

    \I__1200\ : LocalMux
    port map (
            O => \N__11896\,
            I => \eeprom.n1139\
        );

    \I__1199\ : Odrv4
    port map (
            O => \N__11893\,
            I => \eeprom.n1139\
        );

    \I__1198\ : InMux
    port map (
            O => \N__11888\,
            I => \N__11885\
        );

    \I__1197\ : LocalMux
    port map (
            O => \N__11885\,
            I => \N__11882\
        );

    \I__1196\ : Odrv4
    port map (
            O => \N__11882\,
            I => \eeprom.n25\
        );

    \I__1195\ : CascadeMux
    port map (
            O => \N__11879\,
            I => \N__11876\
        );

    \I__1194\ : InMux
    port map (
            O => \N__11876\,
            I => \N__11873\
        );

    \I__1193\ : LocalMux
    port map (
            O => \N__11873\,
            I => \N__11870\
        );

    \I__1192\ : Span4Mux_h
    port map (
            O => \N__11870\,
            I => \N__11867\
        );

    \I__1191\ : Odrv4
    port map (
            O => \N__11867\,
            I => \eeprom.n9\
        );

    \I__1190\ : CascadeMux
    port map (
            O => \N__11864\,
            I => \N__11859\
        );

    \I__1189\ : InMux
    port map (
            O => \N__11863\,
            I => \N__11856\
        );

    \I__1188\ : InMux
    port map (
            O => \N__11862\,
            I => \N__11851\
        );

    \I__1187\ : InMux
    port map (
            O => \N__11859\,
            I => \N__11851\
        );

    \I__1186\ : LocalMux
    port map (
            O => \N__11856\,
            I => \eeprom.delay_counter_24\
        );

    \I__1185\ : LocalMux
    port map (
            O => \N__11851\,
            I => \eeprom.delay_counter_24\
        );

    \I__1184\ : CascadeMux
    port map (
            O => \N__11846\,
            I => \N__11843\
        );

    \I__1183\ : InMux
    port map (
            O => \N__11843\,
            I => \N__11840\
        );

    \I__1182\ : LocalMux
    port map (
            O => \N__11840\,
            I => \N__11837\
        );

    \I__1181\ : Span4Mux_v
    port map (
            O => \N__11837\,
            I => \N__11834\
        );

    \I__1180\ : Odrv4
    port map (
            O => \N__11834\,
            I => \eeprom.n9_adj_408\
        );

    \I__1179\ : CascadeMux
    port map (
            O => \N__11831\,
            I => \N__11828\
        );

    \I__1178\ : InMux
    port map (
            O => \N__11828\,
            I => \N__11825\
        );

    \I__1177\ : LocalMux
    port map (
            O => \N__11825\,
            I => \eeprom.n32\
        );

    \I__1176\ : InMux
    port map (
            O => \N__11822\,
            I => \N__11819\
        );

    \I__1175\ : LocalMux
    port map (
            O => \N__11819\,
            I => \N__11816\
        );

    \I__1174\ : Odrv4
    port map (
            O => \N__11816\,
            I => \eeprom.n26\
        );

    \I__1173\ : InMux
    port map (
            O => \N__11813\,
            I => \N__11809\
        );

    \I__1172\ : InMux
    port map (
            O => \N__11812\,
            I => \N__11805\
        );

    \I__1171\ : LocalMux
    port map (
            O => \N__11809\,
            I => \N__11802\
        );

    \I__1170\ : InMux
    port map (
            O => \N__11808\,
            I => \N__11799\
        );

    \I__1169\ : LocalMux
    port map (
            O => \N__11805\,
            I => \eeprom.delay_counter_30\
        );

    \I__1168\ : Odrv4
    port map (
            O => \N__11802\,
            I => \eeprom.delay_counter_30\
        );

    \I__1167\ : LocalMux
    port map (
            O => \N__11799\,
            I => \eeprom.delay_counter_30\
        );

    \I__1166\ : InMux
    port map (
            O => \N__11792\,
            I => \N__11789\
        );

    \I__1165\ : LocalMux
    port map (
            O => \N__11789\,
            I => \N__11786\
        );

    \I__1164\ : Span4Mux_v
    port map (
            O => \N__11786\,
            I => \N__11783\
        );

    \I__1163\ : Odrv4
    port map (
            O => \N__11783\,
            I => \eeprom.n3\
        );

    \I__1162\ : InMux
    port map (
            O => \N__11780\,
            I => \N__11777\
        );

    \I__1161\ : LocalMux
    port map (
            O => \N__11777\,
            I => \eeprom.n1341\
        );

    \I__1160\ : CascadeMux
    port map (
            O => \N__11774\,
            I => \eeprom.n1256_cascade_\
        );

    \I__1159\ : CascadeMux
    port map (
            O => \N__11771\,
            I => \N__11768\
        );

    \I__1158\ : InMux
    port map (
            O => \N__11768\,
            I => \N__11765\
        );

    \I__1157\ : LocalMux
    port map (
            O => \N__11765\,
            I => \N__11762\
        );

    \I__1156\ : Span4Mux_v
    port map (
            O => \N__11762\,
            I => \N__11759\
        );

    \I__1155\ : Odrv4
    port map (
            O => \N__11759\,
            I => \eeprom.n5_adj_400\
        );

    \I__1154\ : CascadeMux
    port map (
            O => \N__11756\,
            I => \N__11753\
        );

    \I__1153\ : InMux
    port map (
            O => \N__11753\,
            I => \N__11750\
        );

    \I__1152\ : LocalMux
    port map (
            O => \N__11750\,
            I => \N__11747\
        );

    \I__1151\ : Span4Mux_v
    port map (
            O => \N__11747\,
            I => \N__11744\
        );

    \I__1150\ : Odrv4
    port map (
            O => \N__11744\,
            I => \eeprom.n15_adj_415\
        );

    \I__1149\ : InMux
    port map (
            O => \N__11741\,
            I => \N__11738\
        );

    \I__1148\ : LocalMux
    port map (
            O => \N__11738\,
            I => \N__11735\
        );

    \I__1147\ : Odrv4
    port map (
            O => \N__11735\,
            I => \eeprom.n33\
        );

    \I__1146\ : CascadeMux
    port map (
            O => \N__11732\,
            I => \N__11728\
        );

    \I__1145\ : InMux
    port map (
            O => \N__11731\,
            I => \N__11724\
        );

    \I__1144\ : InMux
    port map (
            O => \N__11728\,
            I => \N__11721\
        );

    \I__1143\ : InMux
    port map (
            O => \N__11727\,
            I => \N__11718\
        );

    \I__1142\ : LocalMux
    port map (
            O => \N__11724\,
            I => \eeprom.delay_counter_25\
        );

    \I__1141\ : LocalMux
    port map (
            O => \N__11721\,
            I => \eeprom.delay_counter_25\
        );

    \I__1140\ : LocalMux
    port map (
            O => \N__11718\,
            I => \eeprom.delay_counter_25\
        );

    \I__1139\ : InMux
    port map (
            O => \N__11711\,
            I => \N__11708\
        );

    \I__1138\ : LocalMux
    port map (
            O => \N__11708\,
            I => \N__11705\
        );

    \I__1137\ : Span4Mux_v
    port map (
            O => \N__11705\,
            I => \N__11702\
        );

    \I__1136\ : Odrv4
    port map (
            O => \N__11702\,
            I => \eeprom.n8\
        );

    \I__1135\ : CascadeMux
    port map (
            O => \N__11699\,
            I => \eeprom.n1141_cascade_\
        );

    \I__1134\ : CascadeMux
    port map (
            O => \N__11696\,
            I => \N__11693\
        );

    \I__1133\ : InMux
    port map (
            O => \N__11693\,
            I => \N__11690\
        );

    \I__1132\ : LocalMux
    port map (
            O => \N__11690\,
            I => \N__11687\
        );

    \I__1131\ : Odrv4
    port map (
            O => \N__11687\,
            I => \eeprom.n11_adj_410\
        );

    \I__1130\ : InMux
    port map (
            O => \N__11684\,
            I => \bfn_3_17_0_\
        );

    \I__1129\ : InMux
    port map (
            O => \N__11681\,
            I => \eeprom.n3448\
        );

    \I__1128\ : InMux
    port map (
            O => \N__11678\,
            I => \eeprom.n3449\
        );

    \I__1127\ : InMux
    port map (
            O => \N__11675\,
            I => \eeprom.n3450\
        );

    \I__1126\ : InMux
    port map (
            O => \N__11672\,
            I => \eeprom.n3451\
        );

    \I__1125\ : InMux
    port map (
            O => \N__11669\,
            I => \eeprom.n3452\
        );

    \I__1124\ : InMux
    port map (
            O => \N__11666\,
            I => \eeprom.n3453\
        );

    \I__1123\ : CascadeMux
    port map (
            O => \N__11663\,
            I => \N__11660\
        );

    \I__1122\ : InMux
    port map (
            O => \N__11660\,
            I => \N__11657\
        );

    \I__1121\ : LocalMux
    port map (
            O => \N__11657\,
            I => \N__11654\
        );

    \I__1120\ : Span4Mux_v
    port map (
            O => \N__11654\,
            I => \N__11651\
        );

    \I__1119\ : Odrv4
    port map (
            O => \N__11651\,
            I => \eeprom.n30_adj_458\
        );

    \I__1118\ : InMux
    port map (
            O => \N__11648\,
            I => \bfn_2_24_0_\
        );

    \I__1117\ : CascadeMux
    port map (
            O => \N__11645\,
            I => \N__11642\
        );

    \I__1116\ : InMux
    port map (
            O => \N__11642\,
            I => \N__11639\
        );

    \I__1115\ : LocalMux
    port map (
            O => \N__11639\,
            I => \N__11636\
        );

    \I__1114\ : Span4Mux_v
    port map (
            O => \N__11636\,
            I => \N__11633\
        );

    \I__1113\ : Odrv4
    port map (
            O => \N__11633\,
            I => \eeprom.n8_adj_407\
        );

    \I__1112\ : InMux
    port map (
            O => \N__11630\,
            I => \eeprom.n3810\
        );

    \I__1111\ : CascadeMux
    port map (
            O => \N__11627\,
            I => \N__11624\
        );

    \I__1110\ : InMux
    port map (
            O => \N__11624\,
            I => \N__11621\
        );

    \I__1109\ : LocalMux
    port map (
            O => \N__11621\,
            I => \N__11618\
        );

    \I__1108\ : Span4Mux_v
    port map (
            O => \N__11618\,
            I => \N__11615\
        );

    \I__1107\ : Odrv4
    port map (
            O => \N__11615\,
            I => \eeprom.n7_adj_405\
        );

    \I__1106\ : InMux
    port map (
            O => \N__11612\,
            I => \eeprom.n3811\
        );

    \I__1105\ : CascadeMux
    port map (
            O => \N__11609\,
            I => \N__11606\
        );

    \I__1104\ : InMux
    port map (
            O => \N__11606\,
            I => \N__11603\
        );

    \I__1103\ : LocalMux
    port map (
            O => \N__11603\,
            I => \N__11600\
        );

    \I__1102\ : Span4Mux_v
    port map (
            O => \N__11600\,
            I => \N__11597\
        );

    \I__1101\ : Odrv4
    port map (
            O => \N__11597\,
            I => \eeprom.n6_adj_403\
        );

    \I__1100\ : InMux
    port map (
            O => \N__11594\,
            I => \eeprom.n3812\
        );

    \I__1099\ : InMux
    port map (
            O => \N__11591\,
            I => \eeprom.n3813\
        );

    \I__1098\ : CascadeMux
    port map (
            O => \N__11588\,
            I => \N__11585\
        );

    \I__1097\ : InMux
    port map (
            O => \N__11585\,
            I => \N__11582\
        );

    \I__1096\ : LocalMux
    port map (
            O => \N__11582\,
            I => \N__11579\
        );

    \I__1095\ : Span4Mux_v
    port map (
            O => \N__11579\,
            I => \N__11576\
        );

    \I__1094\ : Odrv4
    port map (
            O => \N__11576\,
            I => \eeprom.n4_adj_397\
        );

    \I__1093\ : InMux
    port map (
            O => \N__11573\,
            I => \eeprom.n3814\
        );

    \I__1092\ : CascadeMux
    port map (
            O => \N__11570\,
            I => \N__11567\
        );

    \I__1091\ : InMux
    port map (
            O => \N__11567\,
            I => \N__11564\
        );

    \I__1090\ : LocalMux
    port map (
            O => \N__11564\,
            I => \N__11561\
        );

    \I__1089\ : Span4Mux_v
    port map (
            O => \N__11561\,
            I => \N__11558\
        );

    \I__1088\ : Odrv4
    port map (
            O => \N__11558\,
            I => \eeprom.n3_adj_396\
        );

    \I__1087\ : InMux
    port map (
            O => \N__11555\,
            I => \eeprom.n3815\
        );

    \I__1086\ : InMux
    port map (
            O => \N__11552\,
            I => \eeprom.n3816\
        );

    \I__1085\ : InMux
    port map (
            O => \N__11549\,
            I => \N__11546\
        );

    \I__1084\ : LocalMux
    port map (
            O => \N__11546\,
            I => \N__11543\
        );

    \I__1083\ : Odrv12
    port map (
            O => \N__11543\,
            I => \eeprom.n14\
        );

    \I__1082\ : InMux
    port map (
            O => \N__11540\,
            I => \N__11537\
        );

    \I__1081\ : LocalMux
    port map (
            O => \N__11537\,
            I => \N__11532\
        );

    \I__1080\ : InMux
    port map (
            O => \N__11536\,
            I => \N__11529\
        );

    \I__1079\ : InMux
    port map (
            O => \N__11535\,
            I => \N__11526\
        );

    \I__1078\ : Span4Mux_v
    port map (
            O => \N__11532\,
            I => \N__11521\
        );

    \I__1077\ : LocalMux
    port map (
            O => \N__11529\,
            I => \N__11521\
        );

    \I__1076\ : LocalMux
    port map (
            O => \N__11526\,
            I => \eeprom.delay_counter_19\
        );

    \I__1075\ : Odrv4
    port map (
            O => \N__11521\,
            I => \eeprom.delay_counter_19\
        );

    \I__1074\ : InMux
    port map (
            O => \N__11516\,
            I => \eeprom.n3800\
        );

    \I__1073\ : InMux
    port map (
            O => \N__11513\,
            I => \N__11510\
        );

    \I__1072\ : LocalMux
    port map (
            O => \N__11510\,
            I => \eeprom.n17_adj_425\
        );

    \I__1071\ : InMux
    port map (
            O => \N__11507\,
            I => \N__11504\
        );

    \I__1070\ : LocalMux
    port map (
            O => \N__11504\,
            I => \eeprom.n17\
        );

    \I__1069\ : InMux
    port map (
            O => \N__11501\,
            I => \bfn_2_23_0_\
        );

    \I__1068\ : CascadeMux
    port map (
            O => \N__11498\,
            I => \N__11495\
        );

    \I__1067\ : InMux
    port map (
            O => \N__11495\,
            I => \N__11492\
        );

    \I__1066\ : LocalMux
    port map (
            O => \N__11492\,
            I => \eeprom.n16_adj_424\
        );

    \I__1065\ : InMux
    port map (
            O => \N__11489\,
            I => \eeprom.n3802\
        );

    \I__1064\ : InMux
    port map (
            O => \N__11486\,
            I => \eeprom.n3803\
        );

    \I__1063\ : CascadeMux
    port map (
            O => \N__11483\,
            I => \N__11480\
        );

    \I__1062\ : InMux
    port map (
            O => \N__11480\,
            I => \N__11477\
        );

    \I__1061\ : LocalMux
    port map (
            O => \N__11477\,
            I => \eeprom.n14_adj_413\
        );

    \I__1060\ : InMux
    port map (
            O => \N__11474\,
            I => \eeprom.n3804\
        );

    \I__1059\ : InMux
    port map (
            O => \N__11471\,
            I => \eeprom.n3805\
        );

    \I__1058\ : InMux
    port map (
            O => \N__11468\,
            I => \eeprom.n3806\
        );

    \I__1057\ : InMux
    port map (
            O => \N__11465\,
            I => \eeprom.n3807\
        );

    \I__1056\ : InMux
    port map (
            O => \N__11462\,
            I => \eeprom.n3808\
        );

    \I__1055\ : InMux
    port map (
            O => \N__11459\,
            I => \eeprom.n3792\
        );

    \I__1054\ : InMux
    port map (
            O => \N__11456\,
            I => \bfn_2_22_0_\
        );

    \I__1053\ : CascadeMux
    port map (
            O => \N__11453\,
            I => \N__11450\
        );

    \I__1052\ : InMux
    port map (
            O => \N__11450\,
            I => \N__11447\
        );

    \I__1051\ : LocalMux
    port map (
            O => \N__11447\,
            I => \N__11444\
        );

    \I__1050\ : Span4Mux_v
    port map (
            O => \N__11444\,
            I => \N__11441\
        );

    \I__1049\ : Odrv4
    port map (
            O => \N__11441\,
            I => \eeprom.n24_adj_463\
        );

    \I__1048\ : InMux
    port map (
            O => \N__11438\,
            I => \eeprom.n3794\
        );

    \I__1047\ : CascadeMux
    port map (
            O => \N__11435\,
            I => \N__11432\
        );

    \I__1046\ : InMux
    port map (
            O => \N__11432\,
            I => \N__11429\
        );

    \I__1045\ : LocalMux
    port map (
            O => \N__11429\,
            I => \N__11426\
        );

    \I__1044\ : Span4Mux_v
    port map (
            O => \N__11426\,
            I => \N__11423\
        );

    \I__1043\ : Odrv4
    port map (
            O => \N__11423\,
            I => \eeprom.n23\
        );

    \I__1042\ : InMux
    port map (
            O => \N__11420\,
            I => \eeprom.n3795\
        );

    \I__1041\ : CascadeMux
    port map (
            O => \N__11417\,
            I => \N__11414\
        );

    \I__1040\ : InMux
    port map (
            O => \N__11414\,
            I => \N__11411\
        );

    \I__1039\ : LocalMux
    port map (
            O => \N__11411\,
            I => \N__11408\
        );

    \I__1038\ : Span4Mux_v
    port map (
            O => \N__11408\,
            I => \N__11405\
        );

    \I__1037\ : Odrv4
    port map (
            O => \N__11405\,
            I => \eeprom.n22_adj_448\
        );

    \I__1036\ : InMux
    port map (
            O => \N__11402\,
            I => \N__11399\
        );

    \I__1035\ : LocalMux
    port map (
            O => \N__11399\,
            I => \N__11396\
        );

    \I__1034\ : Sp12to4
    port map (
            O => \N__11396\,
            I => \N__11393\
        );

    \I__1033\ : Odrv12
    port map (
            O => \N__11393\,
            I => \eeprom.n22_adj_447\
        );

    \I__1032\ : InMux
    port map (
            O => \N__11390\,
            I => \eeprom.n3796\
        );

    \I__1031\ : CascadeMux
    port map (
            O => \N__11387\,
            I => \N__11384\
        );

    \I__1030\ : InMux
    port map (
            O => \N__11384\,
            I => \N__11381\
        );

    \I__1029\ : LocalMux
    port map (
            O => \N__11381\,
            I => \N__11378\
        );

    \I__1028\ : Span4Mux_v
    port map (
            O => \N__11378\,
            I => \N__11375\
        );

    \I__1027\ : Odrv4
    port map (
            O => \N__11375\,
            I => \eeprom.n21_adj_440\
        );

    \I__1026\ : InMux
    port map (
            O => \N__11372\,
            I => \eeprom.n3797\
        );

    \I__1025\ : CascadeMux
    port map (
            O => \N__11369\,
            I => \N__11366\
        );

    \I__1024\ : InMux
    port map (
            O => \N__11366\,
            I => \N__11363\
        );

    \I__1023\ : LocalMux
    port map (
            O => \N__11363\,
            I => \eeprom.n20_adj_431\
        );

    \I__1022\ : InMux
    port map (
            O => \N__11360\,
            I => \N__11357\
        );

    \I__1021\ : LocalMux
    port map (
            O => \N__11357\,
            I => \N__11354\
        );

    \I__1020\ : Span4Mux_s1_h
    port map (
            O => \N__11354\,
            I => \N__11351\
        );

    \I__1019\ : Odrv4
    port map (
            O => \N__11351\,
            I => \eeprom.n20_adj_430\
        );

    \I__1018\ : InMux
    port map (
            O => \N__11348\,
            I => \eeprom.n3798\
        );

    \I__1017\ : InMux
    port map (
            O => \N__11345\,
            I => \eeprom.n3799\
        );

    \I__1016\ : CascadeMux
    port map (
            O => \N__11342\,
            I => \N__11339\
        );

    \I__1015\ : InMux
    port map (
            O => \N__11339\,
            I => \N__11336\
        );

    \I__1014\ : LocalMux
    port map (
            O => \N__11336\,
            I => \N__11333\
        );

    \I__1013\ : Span4Mux_v
    port map (
            O => \N__11333\,
            I => \N__11330\
        );

    \I__1012\ : Odrv4
    port map (
            O => \N__11330\,
            I => \eeprom.n18_adj_427\
        );

    \I__1011\ : InMux
    port map (
            O => \N__11327\,
            I => \eeprom.n3483\
        );

    \I__1010\ : InMux
    port map (
            O => \N__11324\,
            I => \eeprom.n3484\
        );

    \I__1009\ : InMux
    port map (
            O => \N__11321\,
            I => \bfn_2_21_0_\
        );

    \I__1008\ : InMux
    port map (
            O => \N__11318\,
            I => \eeprom.n3786\
        );

    \I__1007\ : CascadeMux
    port map (
            O => \N__11315\,
            I => \N__11312\
        );

    \I__1006\ : InMux
    port map (
            O => \N__11312\,
            I => \N__11309\
        );

    \I__1005\ : LocalMux
    port map (
            O => \N__11309\,
            I => \N__11306\
        );

    \I__1004\ : Odrv4
    port map (
            O => \N__11306\,
            I => \eeprom.n31_adj_457\
        );

    \I__1003\ : InMux
    port map (
            O => \N__11303\,
            I => \eeprom.n3787\
        );

    \I__1002\ : InMux
    port map (
            O => \N__11300\,
            I => \eeprom.n3788\
        );

    \I__1001\ : InMux
    port map (
            O => \N__11297\,
            I => \eeprom.n3789\
        );

    \I__1000\ : CascadeMux
    port map (
            O => \N__11294\,
            I => \N__11291\
        );

    \I__999\ : InMux
    port map (
            O => \N__11291\,
            I => \N__11288\
        );

    \I__998\ : LocalMux
    port map (
            O => \N__11288\,
            I => \N__11285\
        );

    \I__997\ : Odrv4
    port map (
            O => \N__11285\,
            I => \eeprom.n28_adj_461\
        );

    \I__996\ : InMux
    port map (
            O => \N__11282\,
            I => \eeprom.n3790\
        );

    \I__995\ : CascadeMux
    port map (
            O => \N__11279\,
            I => \N__11276\
        );

    \I__994\ : InMux
    port map (
            O => \N__11276\,
            I => \N__11273\
        );

    \I__993\ : LocalMux
    port map (
            O => \N__11273\,
            I => \N__11270\
        );

    \I__992\ : Span4Mux_v
    port map (
            O => \N__11270\,
            I => \N__11267\
        );

    \I__991\ : Odrv4
    port map (
            O => \N__11267\,
            I => \eeprom.n27_adj_462\
        );

    \I__990\ : InMux
    port map (
            O => \N__11264\,
            I => \eeprom.n3791\
        );

    \I__989\ : InMux
    port map (
            O => \N__11261\,
            I => \eeprom.n3474\
        );

    \I__988\ : InMux
    port map (
            O => \N__11258\,
            I => \eeprom.n3475\
        );

    \I__987\ : InMux
    port map (
            O => \N__11255\,
            I => \eeprom.n3476\
        );

    \I__986\ : InMux
    port map (
            O => \N__11252\,
            I => \bfn_2_20_0_\
        );

    \I__985\ : InMux
    port map (
            O => \N__11249\,
            I => \eeprom.n3478\
        );

    \I__984\ : InMux
    port map (
            O => \N__11246\,
            I => \eeprom.n3479\
        );

    \I__983\ : InMux
    port map (
            O => \N__11243\,
            I => \eeprom.n3480\
        );

    \I__982\ : InMux
    port map (
            O => \N__11240\,
            I => \eeprom.n3481\
        );

    \I__981\ : InMux
    port map (
            O => \N__11237\,
            I => \eeprom.n3482\
        );

    \I__980\ : InMux
    port map (
            O => \N__11234\,
            I => \eeprom.n3465\
        );

    \I__979\ : InMux
    port map (
            O => \N__11231\,
            I => \N__11227\
        );

    \I__978\ : InMux
    port map (
            O => \N__11230\,
            I => \N__11223\
        );

    \I__977\ : LocalMux
    port map (
            O => \N__11227\,
            I => \N__11220\
        );

    \I__976\ : InMux
    port map (
            O => \N__11226\,
            I => \N__11217\
        );

    \I__975\ : LocalMux
    port map (
            O => \N__11223\,
            I => \N__11212\
        );

    \I__974\ : Span4Mux_v
    port map (
            O => \N__11220\,
            I => \N__11212\
        );

    \I__973\ : LocalMux
    port map (
            O => \N__11217\,
            I => \eeprom.delay_counter_13\
        );

    \I__972\ : Odrv4
    port map (
            O => \N__11212\,
            I => \eeprom.delay_counter_13\
        );

    \I__971\ : InMux
    port map (
            O => \N__11207\,
            I => \eeprom.n3466\
        );

    \I__970\ : InMux
    port map (
            O => \N__11204\,
            I => \eeprom.n3467\
        );

    \I__969\ : InMux
    port map (
            O => \N__11201\,
            I => \eeprom.n3468\
        );

    \I__968\ : InMux
    port map (
            O => \N__11198\,
            I => \N__11192\
        );

    \I__967\ : InMux
    port map (
            O => \N__11197\,
            I => \N__11192\
        );

    \I__966\ : LocalMux
    port map (
            O => \N__11192\,
            I => \N__11188\
        );

    \I__965\ : InMux
    port map (
            O => \N__11191\,
            I => \N__11185\
        );

    \I__964\ : Span4Mux_v
    port map (
            O => \N__11188\,
            I => \N__11182\
        );

    \I__963\ : LocalMux
    port map (
            O => \N__11185\,
            I => \eeprom.delay_counter_16\
        );

    \I__962\ : Odrv4
    port map (
            O => \N__11182\,
            I => \eeprom.delay_counter_16\
        );

    \I__961\ : InMux
    port map (
            O => \N__11177\,
            I => \bfn_2_19_0_\
        );

    \I__960\ : InMux
    port map (
            O => \N__11174\,
            I => \eeprom.n3470\
        );

    \I__959\ : InMux
    port map (
            O => \N__11171\,
            I => \eeprom.n3471\
        );

    \I__958\ : InMux
    port map (
            O => \N__11168\,
            I => \eeprom.n3472\
        );

    \I__957\ : InMux
    port map (
            O => \N__11165\,
            I => \eeprom.n3473\
        );

    \I__956\ : InMux
    port map (
            O => \N__11162\,
            I => \eeprom.n3456\
        );

    \I__955\ : InMux
    port map (
            O => \N__11159\,
            I => \eeprom.n3457\
        );

    \I__954\ : InMux
    port map (
            O => \N__11156\,
            I => \eeprom.n3458\
        );

    \I__953\ : InMux
    port map (
            O => \N__11153\,
            I => \eeprom.n3459\
        );

    \I__952\ : InMux
    port map (
            O => \N__11150\,
            I => \eeprom.n3460\
        );

    \I__951\ : InMux
    port map (
            O => \N__11147\,
            I => \bfn_2_18_0_\
        );

    \I__950\ : InMux
    port map (
            O => \N__11144\,
            I => \eeprom.n3462\
        );

    \I__949\ : InMux
    port map (
            O => \N__11141\,
            I => \eeprom.n3463\
        );

    \I__948\ : InMux
    port map (
            O => \N__11138\,
            I => \N__11133\
        );

    \I__947\ : InMux
    port map (
            O => \N__11137\,
            I => \N__11128\
        );

    \I__946\ : InMux
    port map (
            O => \N__11136\,
            I => \N__11128\
        );

    \I__945\ : LocalMux
    port map (
            O => \N__11133\,
            I => \eeprom.delay_counter_11\
        );

    \I__944\ : LocalMux
    port map (
            O => \N__11128\,
            I => \eeprom.delay_counter_11\
        );

    \I__943\ : InMux
    port map (
            O => \N__11123\,
            I => \eeprom.n3464\
        );

    \I__942\ : InMux
    port map (
            O => \N__11120\,
            I => \bfn_2_17_0_\
        );

    \I__941\ : InMux
    port map (
            O => \N__11117\,
            I => \eeprom.n3454\
        );

    \I__940\ : InMux
    port map (
            O => \N__11114\,
            I => \eeprom.n3455\
        );

    \I__939\ : IoInMux
    port map (
            O => \N__11111\,
            I => \N__11108\
        );

    \I__938\ : LocalMux
    port map (
            O => \N__11108\,
            I => \N__11105\
        );

    \I__937\ : IoSpan4Mux
    port map (
            O => \N__11105\,
            I => \N__11102\
        );

    \I__936\ : IoSpan4Mux
    port map (
            O => \N__11102\,
            I => \N__11099\
        );

    \I__935\ : IoSpan4Mux
    port map (
            O => \N__11099\,
            I => \N__11096\
        );

    \I__934\ : Odrv4
    port map (
            O => \N__11096\,
            I => \CLK_pad_gb_input\
        );

    \IN_MUX_bfv_2_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_2_21_0_\
        );

    \IN_MUX_bfv_2_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \eeprom.n3793\,
            carryinitout => \bfn_2_22_0_\
        );

    \IN_MUX_bfv_2_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \eeprom.n3801\,
            carryinitout => \bfn_2_23_0_\
        );

    \IN_MUX_bfv_2_24_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \eeprom.n3809\,
            carryinitout => \bfn_2_24_0_\
        );

    \IN_MUX_bfv_15_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_15_20_0_\
        );

    \IN_MUX_bfv_15_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \eeprom.n3779\,
            carryinitout => \bfn_15_21_0_\
        );

    \IN_MUX_bfv_16_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_16_17_0_\
        );

    \IN_MUX_bfv_16_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \eeprom.n3756\,
            carryinitout => \bfn_16_18_0_\
        );

    \IN_MUX_bfv_16_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \eeprom.n3764\,
            carryinitout => \bfn_16_19_0_\
        );

    \IN_MUX_bfv_14_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_14_17_0_\
        );

    \IN_MUX_bfv_14_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \eeprom.n3734\,
            carryinitout => \bfn_14_18_0_\
        );

    \IN_MUX_bfv_14_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \eeprom.n3742\,
            carryinitout => \bfn_14_19_0_\
        );

    \IN_MUX_bfv_9_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_17_0_\
        );

    \IN_MUX_bfv_9_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \eeprom.n3713\,
            carryinitout => \bfn_9_18_0_\
        );

    \IN_MUX_bfv_9_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \eeprom.n3721\,
            carryinitout => \bfn_9_19_0_\
        );

    \IN_MUX_bfv_9_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_20_0_\
        );

    \IN_MUX_bfv_9_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \eeprom.n3693\,
            carryinitout => \bfn_9_21_0_\
        );

    \IN_MUX_bfv_9_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \eeprom.n3701\,
            carryinitout => \bfn_9_22_0_\
        );

    \IN_MUX_bfv_12_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_12_22_0_\
        );

    \IN_MUX_bfv_12_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \eeprom.n3674\,
            carryinitout => \bfn_12_23_0_\
        );

    \IN_MUX_bfv_12_24_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \eeprom.n3682\,
            carryinitout => \bfn_12_24_0_\
        );

    \IN_MUX_bfv_16_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_16_23_0_\
        );

    \IN_MUX_bfv_16_24_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \eeprom.n3656\,
            carryinitout => \bfn_16_24_0_\
        );

    \IN_MUX_bfv_16_25_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \eeprom.n3664\,
            carryinitout => \bfn_16_25_0_\
        );

    \IN_MUX_bfv_11_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_21_0_\
        );

    \IN_MUX_bfv_11_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \eeprom.n3639\,
            carryinitout => \bfn_11_22_0_\
        );

    \IN_MUX_bfv_11_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \eeprom.n3647\,
            carryinitout => \bfn_11_23_0_\
        );

    \IN_MUX_bfv_9_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_23_0_\
        );

    \IN_MUX_bfv_9_24_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \eeprom.n3623\,
            carryinitout => \bfn_9_24_0_\
        );

    \IN_MUX_bfv_9_25_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \eeprom.n3631\,
            carryinitout => \bfn_9_25_0_\
        );

    \IN_MUX_bfv_7_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_21_0_\
        );

    \IN_MUX_bfv_7_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \eeprom.n3608\,
            carryinitout => \bfn_7_22_0_\
        );

    \IN_MUX_bfv_6_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_6_18_0_\
        );

    \IN_MUX_bfv_6_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \eeprom.n3594\,
            carryinitout => \bfn_6_19_0_\
        );

    \IN_MUX_bfv_6_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_6_21_0_\
        );

    \IN_MUX_bfv_6_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \eeprom.n3581\,
            carryinitout => \bfn_6_22_0_\
        );

    \IN_MUX_bfv_4_25_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_4_25_0_\
        );

    \IN_MUX_bfv_4_26_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \eeprom.n3569\,
            carryinitout => \bfn_4_26_0_\
        );

    \IN_MUX_bfv_3_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_3_23_0_\
        );

    \IN_MUX_bfv_3_24_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \eeprom.n3558\,
            carryinitout => \bfn_3_24_0_\
        );

    \IN_MUX_bfv_6_26_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_6_26_0_\
        );

    \IN_MUX_bfv_6_27_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \eeprom.n3548\,
            carryinitout => \bfn_6_27_0_\
        );

    \IN_MUX_bfv_5_27_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_5_27_0_\
        );

    \IN_MUX_bfv_5_28_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \eeprom.n3539\,
            carryinitout => \bfn_5_28_0_\
        );

    \IN_MUX_bfv_5_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_5_22_0_\
        );

    \IN_MUX_bfv_5_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \eeprom.n3531\,
            carryinitout => \bfn_5_23_0_\
        );

    \IN_MUX_bfv_4_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_4_19_0_\
        );

    \IN_MUX_bfv_2_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_2_17_0_\
        );

    \IN_MUX_bfv_2_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \eeprom.n3461\,
            carryinitout => \bfn_2_18_0_\
        );

    \IN_MUX_bfv_2_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \eeprom.n3469\,
            carryinitout => \bfn_2_19_0_\
        );

    \IN_MUX_bfv_2_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \eeprom.n3477\,
            carryinitout => \bfn_2_20_0_\
        );

    \IN_MUX_bfv_16_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_16_20_0_\
        );

    \IN_MUX_bfv_3_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_3_17_0_\
        );

    \IN_MUX_bfv_5_29_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_5_29_0_\
        );

    \IN_MUX_bfv_5_30_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n3492,
            carryinitout => \bfn_5_30_0_\
        );

    \IN_MUX_bfv_5_31_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n3500,
            carryinitout => \bfn_5_31_0_\
        );

    \IN_MUX_bfv_5_32_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n3508,
            carryinitout => \bfn_5_32_0_\
        );

    \CLK_pad_gb\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__11111\,
            GLOBALBUFFEROUTPUT => \CLK_N\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \eeprom.rem_4_unary_minus_2_inv_0_i10_1_lut_LC_1_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12090\,
            lcout => \eeprom.n24_adj_463\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_unary_minus_2_inv_0_i7_1_lut_LC_1_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23595\,
            lcout => \eeprom.n27_adj_462\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_unary_minus_2_inv_0_i11_1_lut_LC_1_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13470\,
            lcout => \eeprom.n23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_mux_3_i12_3_lut_LC_1_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__11137\,
            in1 => \N__11402\,
            in2 => \_gnd_net_\,
            in3 => \N__22970\,
            lcout => \eeprom.n3219\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_unary_minus_2_inv_0_i12_1_lut_LC_1_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11136\,
            lcout => \eeprom.n22_adj_448\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_unary_minus_2_inv_0_i16_1_lut_LC_1_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12267\,
            lcout => \eeprom.n18_adj_427\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_unary_minus_2_inv_0_i13_1_lut_LC_1_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14910\,
            lcout => \eeprom.n21_adj_440\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_unary_minus_2_inv_0_i26_1_lut_LC_1_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11727\,
            lcout => \eeprom.n8_adj_407\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_unary_minus_2_inv_0_i27_1_lut_LC_1_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__12230\,
            in3 => \_gnd_net_\,
            lcout => \eeprom.n7_adj_405\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_unary_minus_2_inv_0_i28_1_lut_LC_1_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11919\,
            lcout => \eeprom.n6_adj_403\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_unary_minus_2_inv_0_i30_1_lut_LC_1_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12165\,
            lcout => \eeprom.n4_adj_397\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_unary_minus_2_inv_0_i31_1_lut_LC_1_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11808\,
            lcout => \eeprom.n3_adj_396\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_unary_minus_2_inv_0_i3_1_lut_LC_1_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__23838\,
            in3 => \_gnd_net_\,
            lcout => \eeprom.n31_adj_457\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_unary_minus_2_inv_0_i6_1_lut_LC_1_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__23658\,
            in3 => \_gnd_net_\,
            lcout => \eeprom.n28_adj_461\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_mux_3_i14_3_lut_LC_1_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__11360\,
            in1 => \N__22888\,
            in2 => \_gnd_net_\,
            in3 => \N__11230\,
            lcout => \eeprom.n3019\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_unary_minus_2_inv_0_i14_1_lut_LC_1_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11231\,
            lcout => \eeprom.n20_adj_431\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_mux_3_i17_3_lut_LC_1_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__11198\,
            in1 => \N__11507\,
            in2 => \_gnd_net_\,
            in3 => \N__22938\,
            lcout => \eeprom.n2719\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_unary_minus_2_inv_0_i17_1_lut_LC_1_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11197\,
            lcout => \eeprom.n17_adj_425\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_unary_minus_2_inv_0_i18_1_lut_LC_1_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12661\,
            lcout => \eeprom.n16_adj_424\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_unary_minus_2_inv_0_i20_1_lut_LC_1_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11536\,
            lcout => \eeprom.n14_adj_413\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.delay_counter_288__i0_LC_2_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23481\,
            in2 => \_gnd_net_\,
            in3 => \N__11120\,
            lcout => \eeprom.delay_counter_0\,
            ltout => OPEN,
            carryin => \bfn_2_17_0_\,
            carryout => \eeprom.n3454\,
            clk => \N__24342\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.delay_counter_288__i1_LC_2_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23891\,
            in2 => \_gnd_net_\,
            in3 => \N__11117\,
            lcout => \eeprom.delay_counter_1\,
            ltout => OPEN,
            carryin => \eeprom.n3454\,
            carryout => \eeprom.n3455\,
            clk => \N__24342\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.delay_counter_288__i2_LC_2_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23828\,
            in2 => \_gnd_net_\,
            in3 => \N__11114\,
            lcout => \eeprom.delay_counter_2\,
            ltout => OPEN,
            carryin => \eeprom.n3455\,
            carryout => \eeprom.n3456\,
            clk => \N__24342\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.delay_counter_288__i3_LC_2_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23772\,
            in2 => \_gnd_net_\,
            in3 => \N__11162\,
            lcout => \eeprom.delay_counter_3\,
            ltout => OPEN,
            carryin => \eeprom.n3456\,
            carryout => \eeprom.n3457\,
            clk => \N__24342\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.delay_counter_288__i4_LC_2_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23703\,
            in2 => \_gnd_net_\,
            in3 => \N__11159\,
            lcout => \eeprom.delay_counter_4\,
            ltout => OPEN,
            carryin => \eeprom.n3457\,
            carryout => \eeprom.n3458\,
            clk => \N__24342\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.delay_counter_288__i5_LC_2_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23649\,
            in2 => \_gnd_net_\,
            in3 => \N__11156\,
            lcout => \eeprom.delay_counter_5\,
            ltout => OPEN,
            carryin => \eeprom.n3458\,
            carryout => \eeprom.n3459\,
            clk => \N__24342\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.delay_counter_288__i6_LC_2_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23599\,
            in2 => \_gnd_net_\,
            in3 => \N__11153\,
            lcout => \eeprom.delay_counter_6\,
            ltout => OPEN,
            carryin => \eeprom.n3459\,
            carryout => \eeprom.n3460\,
            clk => \N__24342\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.delay_counter_288__i7_LC_2_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12832\,
            in2 => \_gnd_net_\,
            in3 => \N__11150\,
            lcout => \eeprom.delay_counter_7\,
            ltout => OPEN,
            carryin => \eeprom.n3460\,
            carryout => \eeprom.n3461\,
            clk => \N__24342\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.delay_counter_288__i8_LC_2_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12397\,
            in2 => \_gnd_net_\,
            in3 => \N__11147\,
            lcout => \eeprom.delay_counter_8\,
            ltout => OPEN,
            carryin => \bfn_2_18_0_\,
            carryout => \eeprom.n3462\,
            clk => \N__24343\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.delay_counter_288__i9_LC_2_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12094\,
            in2 => \_gnd_net_\,
            in3 => \N__11144\,
            lcout => \eeprom.delay_counter_9\,
            ltout => OPEN,
            carryin => \eeprom.n3462\,
            carryout => \eeprom.n3463\,
            clk => \N__24343\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.delay_counter_288__i10_LC_2_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13474\,
            in2 => \_gnd_net_\,
            in3 => \N__11141\,
            lcout => \eeprom.delay_counter_10\,
            ltout => OPEN,
            carryin => \eeprom.n3463\,
            carryout => \eeprom.n3464\,
            clk => \N__24343\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.delay_counter_288__i11_LC_2_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11138\,
            in2 => \_gnd_net_\,
            in3 => \N__11123\,
            lcout => \eeprom.delay_counter_11\,
            ltout => OPEN,
            carryin => \eeprom.n3464\,
            carryout => \eeprom.n3465\,
            clk => \N__24343\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.delay_counter_288__i12_LC_2_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14914\,
            in2 => \_gnd_net_\,
            in3 => \N__11234\,
            lcout => \eeprom.delay_counter_12\,
            ltout => OPEN,
            carryin => \eeprom.n3465\,
            carryout => \eeprom.n3466\,
            clk => \N__24343\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.delay_counter_288__i13_LC_2_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11226\,
            in2 => \_gnd_net_\,
            in3 => \N__11207\,
            lcout => \eeprom.delay_counter_13\,
            ltout => OPEN,
            carryin => \eeprom.n3466\,
            carryout => \eeprom.n3467\,
            clk => \N__24343\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.delay_counter_288__i14_LC_2_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13584\,
            in2 => \_gnd_net_\,
            in3 => \N__11204\,
            lcout => \eeprom.delay_counter_14\,
            ltout => OPEN,
            carryin => \eeprom.n3467\,
            carryout => \eeprom.n3468\,
            clk => \N__24343\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.delay_counter_288__i15_LC_2_18_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12271\,
            in2 => \_gnd_net_\,
            in3 => \N__11201\,
            lcout => \eeprom.delay_counter_15\,
            ltout => OPEN,
            carryin => \eeprom.n3468\,
            carryout => \eeprom.n3469\,
            clk => \N__24343\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.delay_counter_288__i16_LC_2_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11191\,
            in2 => \_gnd_net_\,
            in3 => \N__11177\,
            lcout => \eeprom.delay_counter_16\,
            ltout => OPEN,
            carryin => \bfn_2_19_0_\,
            carryout => \eeprom.n3470\,
            clk => \N__24344\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.delay_counter_288__i17_LC_2_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12660\,
            in2 => \_gnd_net_\,
            in3 => \N__11174\,
            lcout => \eeprom.delay_counter_17\,
            ltout => OPEN,
            carryin => \eeprom.n3470\,
            carryout => \eeprom.n3471\,
            clk => \N__24344\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.delay_counter_288__i18_LC_2_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12334\,
            in2 => \_gnd_net_\,
            in3 => \N__11171\,
            lcout => \eeprom.delay_counter_18\,
            ltout => OPEN,
            carryin => \eeprom.n3471\,
            carryout => \eeprom.n3472\,
            clk => \N__24344\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.delay_counter_288__i19_LC_2_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11535\,
            in2 => \_gnd_net_\,
            in3 => \N__11168\,
            lcout => \eeprom.delay_counter_19\,
            ltout => OPEN,
            carryin => \eeprom.n3472\,
            carryout => \eeprom.n3473\,
            clk => \N__24344\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.delay_counter_288__i20_LC_2_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13050\,
            in2 => \_gnd_net_\,
            in3 => \N__11165\,
            lcout => \eeprom.delay_counter_20\,
            ltout => OPEN,
            carryin => \eeprom.n3473\,
            carryout => \eeprom.n3474\,
            clk => \N__24344\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.delay_counter_288__i21_LC_2_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15609\,
            in2 => \_gnd_net_\,
            in3 => \N__11261\,
            lcout => \eeprom.delay_counter_21\,
            ltout => OPEN,
            carryin => \eeprom.n3474\,
            carryout => \eeprom.n3475\,
            clk => \N__24344\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.delay_counter_288__i22_LC_2_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14178\,
            in2 => \_gnd_net_\,
            in3 => \N__11258\,
            lcout => \eeprom.delay_counter_22\,
            ltout => OPEN,
            carryin => \eeprom.n3475\,
            carryout => \eeprom.n3476\,
            clk => \N__24344\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.delay_counter_288__i23_LC_2_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12306\,
            in2 => \_gnd_net_\,
            in3 => \N__11255\,
            lcout => \eeprom.delay_counter_23\,
            ltout => OPEN,
            carryin => \eeprom.n3476\,
            carryout => \eeprom.n3477\,
            clk => \N__24344\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.delay_counter_288__i24_LC_2_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11863\,
            in2 => \_gnd_net_\,
            in3 => \N__11252\,
            lcout => \eeprom.delay_counter_24\,
            ltout => OPEN,
            carryin => \bfn_2_20_0_\,
            carryout => \eeprom.n3478\,
            clk => \N__24345\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.delay_counter_288__i25_LC_2_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11731\,
            in2 => \_gnd_net_\,
            in3 => \N__11249\,
            lcout => \eeprom.delay_counter_25\,
            ltout => OPEN,
            carryin => \eeprom.n3478\,
            carryout => \eeprom.n3479\,
            clk => \N__24345\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.delay_counter_288__i26_LC_2_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12229\,
            in2 => \_gnd_net_\,
            in3 => \N__11246\,
            lcout => \eeprom.delay_counter_26\,
            ltout => OPEN,
            carryin => \eeprom.n3479\,
            carryout => \eeprom.n3480\,
            clk => \N__24345\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.delay_counter_288__i27_LC_2_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11921\,
            in2 => \_gnd_net_\,
            in3 => \N__11243\,
            lcout => \eeprom.delay_counter_27\,
            ltout => OPEN,
            carryin => \eeprom.n3480\,
            carryout => \eeprom.n3481\,
            clk => \N__24345\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.delay_counter_288__i28_LC_2_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11982\,
            in2 => \_gnd_net_\,
            in3 => \N__11240\,
            lcout => \eeprom.delay_counter_28\,
            ltout => OPEN,
            carryin => \eeprom.n3481\,
            carryout => \eeprom.n3482\,
            clk => \N__24345\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.delay_counter_288__i29_LC_2_20_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12167\,
            in2 => \_gnd_net_\,
            in3 => \N__11237\,
            lcout => \eeprom.delay_counter_29\,
            ltout => OPEN,
            carryin => \eeprom.n3482\,
            carryout => \eeprom.n3483\,
            clk => \N__24345\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.delay_counter_288__i30_LC_2_20_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11812\,
            in2 => \_gnd_net_\,
            in3 => \N__11327\,
            lcout => \eeprom.delay_counter_30\,
            ltout => OPEN,
            carryin => \eeprom.n3483\,
            carryout => \eeprom.n3484\,
            clk => \N__24345\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.delay_counter_288__i31_LC_2_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22906\,
            in2 => \_gnd_net_\,
            in3 => \N__11324\,
            lcout => \eeprom.delay_counter_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24345\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_unary_minus_2_add_3_2_lut_LC_2_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11741\,
            in2 => \_gnd_net_\,
            in3 => \N__11321\,
            lcout => \eeprom.n33_adj_483\,
            ltout => OPEN,
            carryin => \bfn_2_21_0_\,
            carryout => \eeprom.n3786\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_unary_minus_2_add_3_3_lut_LC_2_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__11831\,
            in3 => \N__11318\,
            lcout => \eeprom.n32_adj_480\,
            ltout => OPEN,
            carryin => \eeprom.n3786\,
            carryout => \eeprom.n3787\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_unary_minus_2_add_3_4_lut_LC_2_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__11315\,
            in3 => \N__11303\,
            lcout => \eeprom.n31_adj_476\,
            ltout => OPEN,
            carryin => \eeprom.n3787\,
            carryout => \eeprom.n3788\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_unary_minus_2_add_3_5_lut_LC_2_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__11663\,
            in3 => \N__11300\,
            lcout => \eeprom.n30\,
            ltout => OPEN,
            carryin => \eeprom.n3788\,
            carryout => \eeprom.n3789\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_unary_minus_2_add_3_6_lut_LC_2_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__14894\,
            in3 => \N__11297\,
            lcout => \eeprom.n29\,
            ltout => OPEN,
            carryin => \eeprom.n3789\,
            carryout => \eeprom.n3790\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_unary_minus_2_add_3_7_lut_LC_2_21_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__11294\,
            in3 => \N__11282\,
            lcout => \eeprom.n28\,
            ltout => OPEN,
            carryin => \eeprom.n3790\,
            carryout => \eeprom.n3791\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_unary_minus_2_add_3_8_lut_LC_2_21_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__11279\,
            in3 => \N__11264\,
            lcout => \eeprom.n27\,
            ltout => OPEN,
            carryin => \eeprom.n3791\,
            carryout => \eeprom.n3792\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_unary_minus_2_add_3_9_lut_LC_2_21_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11822\,
            in2 => \_gnd_net_\,
            in3 => \N__11459\,
            lcout => \eeprom.n26_adj_469\,
            ltout => OPEN,
            carryin => \eeprom.n3792\,
            carryout => \eeprom.n3793\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_unary_minus_2_add_3_10_lut_LC_2_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11888\,
            in2 => \_gnd_net_\,
            in3 => \N__11456\,
            lcout => \eeprom.n25_adj_471\,
            ltout => OPEN,
            carryin => \bfn_2_22_0_\,
            carryout => \eeprom.n3794\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_unary_minus_2_add_3_11_lut_LC_2_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__11453\,
            in3 => \N__11438\,
            lcout => \eeprom.n24_adj_467\,
            ltout => OPEN,
            carryin => \eeprom.n3794\,
            carryout => \eeprom.n3795\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_unary_minus_2_add_3_12_lut_LC_2_22_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__11435\,
            in3 => \N__11420\,
            lcout => \eeprom.n23_adj_464\,
            ltout => OPEN,
            carryin => \eeprom.n3795\,
            carryout => \eeprom.n3796\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_unary_minus_2_add_3_13_lut_LC_2_22_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__11417\,
            in3 => \N__11390\,
            lcout => \eeprom.n22_adj_447\,
            ltout => OPEN,
            carryin => \eeprom.n3796\,
            carryout => \eeprom.n3797\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_unary_minus_2_add_3_14_lut_LC_2_22_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__11387\,
            in3 => \N__11372\,
            lcout => \eeprom.n21\,
            ltout => OPEN,
            carryin => \eeprom.n3797\,
            carryout => \eeprom.n3798\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_unary_minus_2_add_3_15_lut_LC_2_22_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__11369\,
            in3 => \N__11348\,
            lcout => \eeprom.n20_adj_430\,
            ltout => OPEN,
            carryin => \eeprom.n3798\,
            carryout => \eeprom.n3799\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_unary_minus_2_add_3_16_lut_LC_2_22_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__13562\,
            in3 => \N__11345\,
            lcout => \eeprom.n19_adj_428\,
            ltout => OPEN,
            carryin => \eeprom.n3799\,
            carryout => \eeprom.n3800\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_unary_minus_2_add_3_17_lut_LC_2_22_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__11342\,
            in3 => \N__11516\,
            lcout => \eeprom.n18_adj_426\,
            ltout => OPEN,
            carryin => \eeprom.n3800\,
            carryout => \eeprom.n3801\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_unary_minus_2_add_3_18_lut_LC_2_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11513\,
            in2 => \_gnd_net_\,
            in3 => \N__11501\,
            lcout => \eeprom.n17\,
            ltout => OPEN,
            carryin => \bfn_2_23_0_\,
            carryout => \eeprom.n3802\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_unary_minus_2_add_3_19_lut_LC_2_23_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__11498\,
            in3 => \N__11489\,
            lcout => \eeprom.n16_adj_377\,
            ltout => OPEN,
            carryin => \eeprom.n3802\,
            carryout => \eeprom.n3803\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_unary_minus_2_add_3_20_lut_LC_2_23_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__11756\,
            in3 => \N__11486\,
            lcout => \eeprom.n15_adj_414\,
            ltout => OPEN,
            carryin => \eeprom.n3803\,
            carryout => \eeprom.n3804\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_unary_minus_2_add_3_21_lut_LC_2_23_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__11483\,
            in3 => \N__11474\,
            lcout => \eeprom.n14\,
            ltout => OPEN,
            carryin => \eeprom.n3804\,
            carryout => \eeprom.n3805\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_unary_minus_2_add_3_22_lut_LC_2_23_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__12068\,
            in3 => \N__11471\,
            lcout => \eeprom.n13\,
            ltout => OPEN,
            carryin => \eeprom.n3805\,
            carryout => \eeprom.n3806\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_unary_minus_2_add_3_23_lut_LC_2_23_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__12428\,
            in3 => \N__11468\,
            lcout => \eeprom.n12_adj_351\,
            ltout => OPEN,
            carryin => \eeprom.n3806\,
            carryout => \eeprom.n3807\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_unary_minus_2_add_3_24_lut_LC_2_23_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__11696\,
            in3 => \N__11465\,
            lcout => \eeprom.n11\,
            ltout => OPEN,
            carryin => \eeprom.n3807\,
            carryout => \eeprom.n3808\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_unary_minus_2_add_3_25_lut_LC_2_23_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__12056\,
            in3 => \N__11462\,
            lcout => \eeprom.n10\,
            ltout => OPEN,
            carryin => \eeprom.n3808\,
            carryout => \eeprom.n3809\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_unary_minus_2_add_3_26_lut_LC_2_24_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__11846\,
            in3 => \N__11648\,
            lcout => \eeprom.n9\,
            ltout => OPEN,
            carryin => \bfn_2_24_0_\,
            carryout => \eeprom.n3810\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_unary_minus_2_add_3_27_lut_LC_2_24_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__11645\,
            in3 => \N__11630\,
            lcout => \eeprom.n8\,
            ltout => OPEN,
            carryin => \eeprom.n3810\,
            carryout => \eeprom.n3811\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_unary_minus_2_add_3_28_lut_LC_2_24_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__11627\,
            in3 => \N__11612\,
            lcout => \eeprom.n7\,
            ltout => OPEN,
            carryin => \eeprom.n3811\,
            carryout => \eeprom.n3812\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_unary_minus_2_add_3_29_lut_LC_2_24_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__11609\,
            in3 => \N__11594\,
            lcout => \eeprom.n6_adj_402\,
            ltout => OPEN,
            carryin => \eeprom.n3812\,
            carryout => \eeprom.n3813\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_unary_minus_2_add_3_30_lut_LC_2_24_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__11771\,
            in3 => \N__11591\,
            lcout => \eeprom.n5\,
            ltout => OPEN,
            carryin => \eeprom.n3813\,
            carryout => \eeprom.n3814\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_unary_minus_2_add_3_31_lut_LC_2_24_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__11588\,
            in3 => \N__11573\,
            lcout => \eeprom.n4\,
            ltout => OPEN,
            carryin => \eeprom.n3814\,
            carryout => \eeprom.n3815\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_unary_minus_2_add_3_32_lut_LC_2_24_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__11570\,
            in3 => \N__11555\,
            lcout => \eeprom.n3\,
            ltout => OPEN,
            carryin => \eeprom.n3815\,
            carryout => \eeprom.n3816\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_unary_minus_2_add_3_33_lut_LC_2_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24004\,
            in2 => \_gnd_net_\,
            in3 => \N__11552\,
            lcout => \eeprom.n2_adj_395\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_mux_3_i20_3_lut_LC_2_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__11549\,
            in1 => \N__22969\,
            in2 => \_gnd_net_\,
            in3 => \N__11540\,
            lcout => \eeprom.n2419\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_unary_minus_2_inv_0_i23_1_lut_LC_2_26_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14185\,
            lcout => \eeprom.n11_adj_410\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.add_937_2_lut_LC_3_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__12008\,
            in3 => \N__11684\,
            lcout => \eeprom.n1343\,
            ltout => OPEN,
            carryin => \bfn_3_17_0_\,
            carryout => \eeprom.n3448\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.add_937_3_lut_LC_3_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27731\,
            in2 => \N__12188\,
            in3 => \N__11681\,
            lcout => \eeprom.n1342\,
            ltout => OPEN,
            carryin => \eeprom.n3448\,
            carryout => \eeprom.n3449\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.add_937_4_lut_LC_3_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11903\,
            in2 => \_gnd_net_\,
            in3 => \N__11678\,
            lcout => \eeprom.n1341\,
            ltout => OPEN,
            carryin => \eeprom.n3449\,
            carryout => \eeprom.n3450\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.add_937_5_lut_LC_3_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12512\,
            in2 => \_gnd_net_\,
            in3 => \N__11675\,
            lcout => \eeprom.n1340\,
            ltout => OPEN,
            carryin => \eeprom.n3450\,
            carryout => \eeprom.n3451\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.add_937_6_lut_LC_3_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__12137\,
            in3 => \N__11672\,
            lcout => \eeprom.n1339\,
            ltout => OPEN,
            carryin => \eeprom.n3451\,
            carryout => \eeprom.n3452\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.add_937_7_lut_LC_3_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101110111110"
        )
    port map (
            in0 => \N__12524\,
            in1 => \_gnd_net_\,
            in2 => \N__12607\,
            in3 => \N__11669\,
            lcout => \eeprom.n4734\,
            ltout => OPEN,
            carryin => \eeprom.n3452\,
            carryout => \eeprom.n3453\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.add_937_8_lut_LC_3_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__12488\,
            in3 => \N__11666\,
            lcout => \eeprom.n1337\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_unary_minus_2_inv_0_i4_1_lut_LC_3_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23768\,
            lcout => \eeprom.n30_adj_458\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i520_2_lut_LC_3_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22955\,
            in2 => \_gnd_net_\,
            in3 => \N__12044\,
            lcout => \eeprom.n1135\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_unary_minus_2_inv_0_i8_1_lut_LC_3_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12828\,
            lcout => \eeprom.n26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_mux_3_i31_3_lut_LC_3_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__11813\,
            in1 => \N__22954\,
            in2 => \_gnd_net_\,
            in3 => \N__11792\,
            lcout => \eeprom.n1256\,
            ltout => \eeprom.n1256_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1224_3_lut_4_lut_LC_3_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110011001100"
        )
    port map (
            in0 => \N__11780\,
            in1 => \N__11902\,
            in2 => \N__11774\,
            in3 => \N__12466\,
            lcout => \eeprom.n1916\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_unary_minus_2_inv_0_i29_1_lut_LC_3_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11983\,
            lcout => \eeprom.n5_adj_400\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_unary_minus_2_inv_0_i19_1_lut_LC_3_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12330\,
            lcout => \eeprom.n15_adj_415\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_unary_minus_2_inv_0_i1_1_lut_LC_3_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23475\,
            lcout => \eeprom.n33\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_mux_3_i26_3_lut_LC_3_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22852\,
            in2 => \N__11732\,
            in3 => \N__11711\,
            lcout => \eeprom.n1141\,
            ltout => \eeprom.n1141_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i1_4_lut_adj_48_LC_3_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010000000"
        )
    port map (
            in0 => \N__22853\,
            in1 => \N__11935\,
            in2 => \N__11699\,
            in3 => \N__12205\,
            lcout => OPEN,
            ltout => \eeprom.n4399_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i1_4_lut_adj_49_LC_3_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__12043\,
            in1 => \N__12507\,
            in2 => \N__12020\,
            in3 => \N__12130\,
            lcout => \eeprom.n4405\,
            ltout => \eeprom.n4405_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1226_3_lut_4_lut_LC_3_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110011001100"
        )
    port map (
            in0 => \N__12017\,
            in1 => \N__12004\,
            in2 => \N__11990\,
            in3 => \N__12605\,
            lcout => \eeprom.n1918\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_mux_3_i29_3_lut_LC_3_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__11987\,
            in1 => \N__22851\,
            in2 => \_gnd_net_\,
            in3 => \N__11960\,
            lcout => \eeprom.n1138\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1225_3_lut_4_lut_LC_3_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101000101010"
        )
    port map (
            in0 => \N__12187\,
            in1 => \N__12606\,
            in2 => \N__12473\,
            in3 => \N__11948\,
            lcout => \eeprom.n1917\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_mux_3_i28_3_lut_LC_3_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22854\,
            in2 => \N__11939\,
            in3 => \N__11920\,
            lcout => \eeprom.n1139\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_unary_minus_2_inv_0_i9_1_lut_LC_3_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12393\,
            lcout => \eeprom.n25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_mux_3_i25_3_lut_LC_3_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22849\,
            in2 => \N__11879\,
            in3 => \N__11862\,
            lcout => \eeprom.n1919\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_unary_minus_2_inv_0_i25_1_lut_LC_3_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__11864\,
            in3 => \_gnd_net_\,
            lcout => \eeprom.n9_adj_408\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_unary_minus_2_inv_0_i2_1_lut_LC_3_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23901\,
            lcout => \eeprom.n32\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_mux_3_i27_3_lut_LC_3_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__12228\,
            in1 => \_gnd_net_\,
            in2 => \N__12209\,
            in3 => \N__22848\,
            lcout => \eeprom.n1140\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_mux_3_i30_3_lut_LC_3_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__22847\,
            in1 => \N__12166\,
            in2 => \_gnd_net_\,
            in3 => \N__12149\,
            lcout => \eeprom.n1137\,
            ltout => \eeprom.n1137_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i4030_3_lut_4_lut_LC_3_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100011110000"
        )
    port map (
            in0 => \N__12608\,
            in1 => \N__12119\,
            in2 => \N__12110\,
            in3 => \N__12470\,
            lcout => \eeprom.n1914\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_mux_3_i10_3_lut_LC_3_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__22850\,
            in1 => \N__12107\,
            in2 => \_gnd_net_\,
            in3 => \N__12095\,
            lcout => \eeprom.n3419\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_mux_3_i1_3_lut_LC_3_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010001110111"
        )
    port map (
            in0 => \N__12074\,
            in1 => \N__22846\,
            in2 => \_gnd_net_\,
            in3 => \N__23488\,
            lcout => \eeprom.n1166\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_unary_minus_2_inv_0_i21_1_lut_LC_3_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13051\,
            lcout => \eeprom.n13_adj_412\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_unary_minus_2_inv_0_i32_1_lut_LC_3_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22845\,
            lcout => \eeprom.n2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_unary_minus_2_inv_0_i24_1_lut_LC_3_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12307\,
            lcout => \eeprom.n10_adj_409\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_mux_3_i15_3_lut_LC_3_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__12344\,
            in1 => \N__22923\,
            in2 => \_gnd_net_\,
            in3 => \N__13589\,
            lcout => \eeprom.n2919\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i4037_3_lut_LC_3_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15793\,
            in2 => \N__12242\,
            in3 => \N__13100\,
            lcout => \eeprom.n2415\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_mux_3_i19_3_lut_LC_3_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__22921\,
            in1 => \N__12338\,
            in2 => \_gnd_net_\,
            in3 => \N__12314\,
            lcout => \eeprom.n2519\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_mux_3_i24_3_lut_LC_3_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__12308\,
            in1 => \N__12287\,
            in2 => \_gnd_net_\,
            in3 => \N__22920\,
            lcout => \eeprom.n2019\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_mux_3_i16_3_lut_LC_3_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__22922\,
            in1 => \N__12281\,
            in2 => \_gnd_net_\,
            in3 => \N__12275\,
            lcout => \eeprom.n2819\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1553_2_lut_LC_3_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14004\,
            in2 => \_gnd_net_\,
            in3 => \N__12251\,
            lcout => \eeprom.n2386\,
            ltout => OPEN,
            carryin => \bfn_3_23_0_\,
            carryout => \eeprom.n3551\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1553_3_lut_LC_3_23_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27582\,
            in2 => \N__15584\,
            in3 => \N__12248\,
            lcout => \eeprom.n2385\,
            ltout => OPEN,
            carryin => \eeprom.n3551\,
            carryout => \eeprom.n3552\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1553_4_lut_LC_3_23_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__15728\,
            in3 => \N__12245\,
            lcout => \eeprom.n2384\,
            ltout => OPEN,
            carryin => \eeprom.n3552\,
            carryout => \eeprom.n3553\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1553_5_lut_LC_3_23_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__15794\,
            in3 => \N__12233\,
            lcout => \eeprom.n2383\,
            ltout => OPEN,
            carryin => \eeprom.n3553\,
            carryout => \eeprom.n3554\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1553_6_lut_LC_3_23_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__14159\,
            in3 => \N__12377\,
            lcout => \eeprom.n2382\,
            ltout => OPEN,
            carryin => \eeprom.n3554\,
            carryout => \eeprom.n3555\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1553_7_lut_LC_3_23_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__15830\,
            in3 => \N__12374\,
            lcout => \eeprom.n2381\,
            ltout => OPEN,
            carryin => \eeprom.n3555\,
            carryout => \eeprom.n3556\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1553_8_lut_LC_3_23_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14228\,
            in2 => \_gnd_net_\,
            in3 => \N__12371\,
            lcout => \eeprom.n2380\,
            ltout => OPEN,
            carryin => \eeprom.n3556\,
            carryout => \eeprom.n3557\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1553_9_lut_LC_3_23_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13172\,
            in2 => \N__27784\,
            in3 => \N__12368\,
            lcout => \eeprom.n2379\,
            ltout => OPEN,
            carryin => \eeprom.n3557\,
            carryout => \eeprom.n3558\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1553_10_lut_LC_3_24_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27732\,
            in2 => \N__14129\,
            in3 => \N__12365\,
            lcout => \eeprom.n2378\,
            ltout => OPEN,
            carryin => \bfn_3_24_0_\,
            carryout => \eeprom.n3559\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1553_11_lut_LC_3_24_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13979\,
            in2 => \N__27783\,
            in3 => \N__12362\,
            lcout => \eeprom.n2377\,
            ltout => OPEN,
            carryin => \eeprom.n3559\,
            carryout => \eeprom.n3560\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1553_12_lut_LC_3_24_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14036\,
            in2 => \N__27785\,
            in3 => \N__12359\,
            lcout => \eeprom.n2376\,
            ltout => OPEN,
            carryin => \eeprom.n3560\,
            carryout => \eeprom.n3561\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1553_13_lut_LC_3_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001000001100000"
        )
    port map (
            in0 => \N__16523\,
            in1 => \N__27742\,
            in2 => \N__13115\,
            in3 => \N__12356\,
            lcout => \eeprom.n2407\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1566_3_lut_LC_3_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__14012\,
            in1 => \_gnd_net_\,
            in2 => \N__13114\,
            in3 => \N__12353\,
            lcout => \eeprom.n2418\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i4035_3_lut_LC_3_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12545\,
            in2 => \N__15829\,
            in3 => \N__13090\,
            lcout => \eeprom.n2413\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1564_3_lut_LC_3_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12539\,
            in2 => \N__13113\,
            in3 => \N__15727\,
            lcout => \eeprom.n2416\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1558_3_lut_LC_3_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14127\,
            in2 => \N__12533\,
            in3 => \N__13118\,
            lcout => \eeprom.n2410\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i3948_1_lut_LC_4_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12459\,
            lcout => \eeprom.n4733\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1223_3_lut_4_lut_LC_4_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111110000000"
        )
    port map (
            in0 => \N__12518\,
            in1 => \N__12598\,
            in2 => \N__12471\,
            in3 => \N__12511\,
            lcout => \eeprom.n1915\,
            ltout => \eeprom.n1915_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i1_2_lut_3_lut_LC_4_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000000000000"
        )
    port map (
            in0 => \N__12599\,
            in1 => \_gnd_net_\,
            in2 => \N__12491\,
            in3 => \N__12616\,
            lcout => \eeprom.n4437\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1220_3_lut_4_lut_LC_4_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101000101010"
        )
    port map (
            in0 => \N__12487\,
            in1 => \N__12600\,
            in2 => \N__12472\,
            in3 => \N__12434\,
            lcout => \eeprom.n1912\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_unary_minus_2_inv_0_i22_1_lut_LC_4_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15616\,
            lcout => \eeprom.n12_adj_411\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_mux_3_i9_3_lut_LC_4_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__22957\,
            in1 => \N__12410\,
            in2 => \_gnd_net_\,
            in3 => \N__12398\,
            lcout => \eeprom.n3519_adj_379\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_mux_3_i18_3_lut_LC_4_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__12665\,
            in1 => \N__12635\,
            in2 => \_gnd_net_\,
            in3 => \N__22956\,
            lcout => \eeprom.n2619\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i3950_2_lut_LC_4_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__12620\,
            in3 => \N__12601\,
            lcout => \eeprom.n1913\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1285_2_lut_LC_4_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12975\,
            in2 => \_gnd_net_\,
            in3 => \N__12566\,
            lcout => \eeprom.n1986\,
            ltout => OPEN,
            carryin => \bfn_4_19_0_\,
            carryout => \eeprom.n3517\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1285_3_lut_LC_4_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27730\,
            in2 => \N__12767\,
            in3 => \N__12563\,
            lcout => \eeprom.n1985\,
            ltout => OPEN,
            carryin => \eeprom.n3517\,
            carryout => \eeprom.n3518\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1285_4_lut_LC_4_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__12794\,
            in3 => \N__12560\,
            lcout => \eeprom.n1984\,
            ltout => OPEN,
            carryin => \eeprom.n3518\,
            carryout => \eeprom.n3519\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1285_5_lut_LC_4_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__12727\,
            in3 => \N__12557\,
            lcout => \eeprom.n1983\,
            ltout => OPEN,
            carryin => \eeprom.n3519\,
            carryout => \eeprom.n3520\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1285_6_lut_LC_4_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13009\,
            in2 => \_gnd_net_\,
            in3 => \N__12554\,
            lcout => \eeprom.n1982\,
            ltout => OPEN,
            carryin => \eeprom.n3520\,
            carryout => \eeprom.n3521\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1285_7_lut_LC_4_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__12686\,
            in3 => \N__12551\,
            lcout => \eeprom.n1981\,
            ltout => OPEN,
            carryin => \eeprom.n3521\,
            carryout => \eeprom.n3522\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1285_8_lut_LC_4_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__12946\,
            in3 => \N__12548\,
            lcout => \eeprom.n1980\,
            ltout => OPEN,
            carryin => \eeprom.n3522\,
            carryout => \eeprom.n3523\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1285_9_lut_LC_4_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001000001100000"
        )
    port map (
            in0 => \N__27383\,
            in1 => \N__12742\,
            in2 => \N__12929\,
            in3 => \N__12851\,
            lcout => \eeprom.n2011\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_mux_3_i8_3_lut_LC_4_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__22943\,
            in1 => \N__12848\,
            in2 => \_gnd_net_\,
            in3 => \N__12836\,
            lcout => \eeprom.n3619_adj_352\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1292_3_lut_LC_4_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__12793\,
            in1 => \_gnd_net_\,
            in2 => \N__12812\,
            in3 => \N__12911\,
            lcout => \eeprom.n2016\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1293_3_lut_LC_4_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__12803\,
            in1 => \_gnd_net_\,
            in2 => \N__12926\,
            in3 => \N__12766\,
            lcout => \eeprom.n2017\,
            ltout => \eeprom.n2017_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i1_3_lut_adj_68_LC_4_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13632\,
            in2 => \N__12797\,
            in3 => \N__13743\,
            lcout => \eeprom.n4415\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i1_4_lut_adj_65_LC_4_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__12792\,
            in1 => \N__12681\,
            in2 => \N__12728\,
            in3 => \N__12776\,
            lcout => OPEN,
            ltout => \eeprom.n4441_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i3028_4_lut_LC_4_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111100000"
        )
    port map (
            in0 => \N__12765\,
            in1 => \N__12976\,
            in2 => \N__12746\,
            in3 => \N__12743\,
            lcout => \eeprom.n1945\,
            ltout => \eeprom.n1945_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1291_3_lut_LC_4_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__12726\,
            in1 => \_gnd_net_\,
            in2 => \N__12704\,
            in3 => \N__12701\,
            lcout => \eeprom.n2015\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i4031_3_lut_LC_4_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12695\,
            in2 => \N__12928\,
            in3 => \N__12685\,
            lcout => \eeprom.n2013\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1290_3_lut_LC_4_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13013\,
            in2 => \N__12998\,
            in3 => \N__12916\,
            lcout => \eeprom.n2014\,
            ltout => \eeprom.n2014_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i1_4_lut_adj_70_LC_4_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000000000000"
        )
    port map (
            in0 => \N__14064\,
            in1 => \N__13674\,
            in2 => \N__12986\,
            in3 => \N__12983\,
            lcout => \eeprom.n4419\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1294_3_lut_LC_4_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12977\,
            in2 => \N__12959\,
            in3 => \N__12915\,
            lcout => \eeprom.n2018\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i3_4_lut_adj_80_LC_4_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011110000"
        )
    port map (
            in0 => \N__15180\,
            in1 => \N__15144\,
            in2 => \N__15370\,
            in3 => \N__12869\,
            lcout => \eeprom.n11_adj_473\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1288_3_lut_LC_4_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__12947\,
            in1 => \_gnd_net_\,
            in2 => \N__12927\,
            in3 => \N__12887\,
            lcout => \eeprom.n2012\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i1_4_lut_adj_71_LC_4_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011101110"
        )
    port map (
            in0 => \N__13843\,
            in1 => \N__13792\,
            in2 => \N__13885\,
            in3 => \N__12878\,
            lcout => \eeprom.n2044\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i1_2_lut_adj_78_LC_4_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__15006\,
            in3 => \N__15537\,
            lcout => OPEN,
            ltout => \eeprom.n4575_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i1_4_lut_adj_79_LC_4_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__15096\,
            in1 => \N__15051\,
            in2 => \N__12872\,
            in3 => \N__14958\,
            lcout => \eeprom.n4579\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_mux_3_i21_3_lut_LC_4_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__12863\,
            in1 => \N__13055\,
            in2 => \_gnd_net_\,
            in3 => \N__22959\,
            lcout => \eeprom.n2319\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1632_3_lut_LC_4_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13324\,
            in2 => \N__13304\,
            in3 => \N__15961\,
            lcout => \eeprom.n2516\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1630_3_lut_LC_4_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13254\,
            in2 => \N__13232\,
            in3 => \N__15960\,
            lcout => \eeprom.n2514\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i1_3_lut_adj_74_LC_4_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13320\,
            in2 => \N__13288\,
            in3 => \N__13209\,
            lcout => OPEN,
            ltout => \eeprom.n4479_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i1_4_lut_adj_75_LC_4_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000000000000"
        )
    port map (
            in0 => \N__13720\,
            in1 => \N__13359\,
            in2 => \N__13031\,
            in3 => \N__13028\,
            lcout => \eeprom.n4133\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i1_2_lut_adj_73_LC_4_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__13255\,
            in3 => \N__16083\,
            lcout => \eeprom.n4477\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i5_4_lut_LC_4_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__13171\,
            in1 => \N__13730\,
            in2 => \N__14128\,
            in3 => \N__13985\,
            lcout => \eeprom.n2341\,
            ltout => \eeprom.n2341_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1565_3_lut_LC_4_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__13022\,
            in1 => \_gnd_net_\,
            in2 => \N__13016\,
            in3 => \N__15583\,
            lcout => \eeprom.n2417\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1629_3_lut_LC_4_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13196\,
            in2 => \N__13216\,
            in3 => \N__15931\,
            lcout => \eeprom.n2513\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1631_3_lut_LC_4_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__13284\,
            in1 => \_gnd_net_\,
            in2 => \N__15959\,
            in3 => \N__13268\,
            lcout => \eeprom.n2515\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1633_3_lut_LC_4_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13360\,
            in2 => \N__13343\,
            in3 => \N__15935\,
            lcout => \eeprom.n2517\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1556_3_lut_LC_4_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13178\,
            in2 => \N__13117\,
            in3 => \N__14034\,
            lcout => \eeprom.n2408\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1492_3_lut_LC_4_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16115\,
            in2 => \N__16727\,
            in3 => \N__16603\,
            lcout => \eeprom.n2312\,
            ltout => \eeprom.n2312_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1559_3_lut_LC_4_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__13102\,
            in1 => \_gnd_net_\,
            in2 => \N__13160\,
            in3 => \N__13157\,
            lcout => \eeprom.n2411\,
            ltout => \eeprom.n2411_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i5_4_lut_adj_76_LC_4_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__13375\,
            in1 => \N__13413\,
            in2 => \N__13151\,
            in3 => \N__13148\,
            lcout => OPEN,
            ltout => \eeprom.n12_adj_472_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i6_4_lut_adj_77_LC_4_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__16014\,
            in1 => \N__13429\,
            in2 => \N__13142\,
            in3 => \N__15685\,
            lcout => \eeprom.n2440\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1562_3_lut_LC_4_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13139\,
            in2 => \N__14155\,
            in3 => \N__13101\,
            lcout => \eeprom.n2414\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1557_3_lut_LC_4_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13133\,
            in2 => \N__13116\,
            in3 => \N__13978\,
            lcout => \eeprom.n2409\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1560_3_lut_LC_4_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14224\,
            in2 => \N__13127\,
            in3 => \N__13103\,
            lcout => \eeprom.n2412\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1620_2_lut_LC_4_25_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13719\,
            in2 => \_gnd_net_\,
            in3 => \N__13364\,
            lcout => \eeprom.n2486\,
            ltout => OPEN,
            carryin => \bfn_4_25_0_\,
            carryout => \eeprom.n3562\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1620_3_lut_LC_4_25_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27371\,
            in2 => \N__13361\,
            in3 => \N__13331\,
            lcout => \eeprom.n2485\,
            ltout => OPEN,
            carryin => \eeprom.n3562\,
            carryout => \eeprom.n3563\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1620_4_lut_LC_4_25_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__13328\,
            in3 => \N__13292\,
            lcout => \eeprom.n2484\,
            ltout => OPEN,
            carryin => \eeprom.n3563\,
            carryout => \eeprom.n3564\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1620_5_lut_LC_4_25_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__13289\,
            in3 => \N__13259\,
            lcout => \eeprom.n2483\,
            ltout => OPEN,
            carryin => \eeprom.n3564\,
            carryout => \eeprom.n3565\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1620_6_lut_LC_4_25_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13256\,
            in2 => \_gnd_net_\,
            in3 => \N__13220\,
            lcout => \eeprom.n2482\,
            ltout => OPEN,
            carryin => \eeprom.n3565\,
            carryout => \eeprom.n3566\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1620_7_lut_LC_4_25_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__13217\,
            in3 => \N__13187\,
            lcout => \eeprom.n2481\,
            ltout => OPEN,
            carryin => \eeprom.n3566\,
            carryout => \eeprom.n3567\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1620_8_lut_LC_4_25_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__16090\,
            in3 => \N__13184\,
            lcout => \eeprom.n2480\,
            ltout => OPEN,
            carryin => \eeprom.n3567\,
            carryout => \eeprom.n3568\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1620_9_lut_LC_4_25_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15684\,
            in2 => \N__27581\,
            in3 => \N__13181\,
            lcout => \eeprom.n2479\,
            ltout => OPEN,
            carryin => \eeprom.n3568\,
            carryout => \eeprom.n3569\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1620_10_lut_LC_4_26_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13531\,
            in2 => \N__27744\,
            in3 => \N__13445\,
            lcout => \eeprom.n2478\,
            ltout => OPEN,
            carryin => \bfn_4_26_0_\,
            carryout => \eeprom.n3570\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1620_11_lut_LC_4_26_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13414\,
            in2 => \N__27746\,
            in3 => \N__13442\,
            lcout => \eeprom.n2477\,
            ltout => OPEN,
            carryin => \eeprom.n3570\,
            carryout => \eeprom.n3571\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1620_12_lut_LC_4_26_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13381\,
            in2 => \N__27745\,
            in3 => \N__13439\,
            lcout => \eeprom.n2476\,
            ltout => OPEN,
            carryin => \eeprom.n3571\,
            carryout => \eeprom.n3572\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1620_13_lut_LC_4_26_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16021\,
            in2 => \N__27747\,
            in3 => \N__13436\,
            lcout => \eeprom.n2475\,
            ltout => OPEN,
            carryin => \eeprom.n3572\,
            carryout => \eeprom.n3573\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1620_14_lut_LC_4_26_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001000001100000"
        )
    port map (
            in0 => \N__27620\,
            in1 => \N__13433\,
            in2 => \N__15977\,
            in3 => \N__13418\,
            lcout => \eeprom.n2506\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1625_3_lut_LC_4_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13415\,
            in2 => \N__13400\,
            in3 => \N__15963\,
            lcout => \eeprom.n2509\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1624_3_lut_LC_4_26_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13391\,
            in2 => \N__13385\,
            in3 => \N__15962\,
            lcout => \eeprom.n2508\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i3982_4_lut_LC_4_31_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110111100000"
        )
    port map (
            in0 => \N__14783\,
            in1 => \N__14744\,
            in2 => \N__14804\,
            in3 => \N__14764\,
            lcout => n4826,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i3981_4_lut_LC_4_31_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110101000000"
        )
    port map (
            in0 => \N__14743\,
            in1 => \N__14782\,
            in2 => \N__14765\,
            in3 => \N__14800\,
            lcout => OPEN,
            ltout => \n4825_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i3983_3_lut_LC_4_31_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13505\,
            in2 => \N__13499\,
            in3 => \N__14723\,
            lcout => \LED_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_mux_3_i11_3_lut_LC_5_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__13487\,
            in1 => \N__22958\,
            in2 => \_gnd_net_\,
            in3 => \N__13475\,
            lcout => \eeprom.n3319\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1700_3_lut_LC_5_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15080\,
            in2 => \N__15518\,
            in3 => \N__15112\,
            lcout => \eeprom.n2616\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1699_3_lut_LC_5_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15504\,
            in2 => \N__15035\,
            in3 => \N__15067\,
            lcout => \eeprom.n2615\,
            ltout => \eeprom.n2615_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i1_2_lut_adj_83_LC_5_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__13454\,
            in3 => \N__16413\,
            lcout => OPEN,
            ltout => \eeprom.n4497_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i1_4_lut_adj_84_LC_5_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__16884\,
            in1 => \N__16842\,
            in2 => \N__13451\,
            in3 => \N__16908\,
            lcout => OPEN,
            ltout => \eeprom.n4501_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i3_4_lut_adj_86_LC_5_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011101100"
        )
    port map (
            in0 => \N__16762\,
            in1 => \N__14874\,
            in2 => \N__13448\,
            in3 => \N__16809\,
            lcout => \eeprom.n12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1701_3_lut_LC_5_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15125\,
            in2 => \N__15152\,
            in3 => \N__15500\,
            lcout => \eeprom.n2617\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1698_3_lut_LC_5_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14981\,
            in2 => \N__15020\,
            in3 => \N__15505\,
            lcout => \eeprom.n2614\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1693_3_lut_LC_5_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15347\,
            in2 => \N__15519\,
            in3 => \N__15369\,
            lcout => \eeprom.n2609\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i5_4_lut_adj_81_LC_5_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__15327\,
            in1 => \N__15223\,
            in2 => \N__15276\,
            in3 => \N__15899\,
            lcout => OPEN,
            ltout => \eeprom.n13_adj_474_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i7_4_lut_adj_82_LC_5_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__15653\,
            in1 => \N__16050\,
            in2 => \N__13601\,
            in3 => \N__13598\,
            lcout => \eeprom.n2539\,
            ltout => \eeprom.n2539_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1697_3_lut_LC_5_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14968\,
            in2 => \N__13592\,
            in3 => \N__15398\,
            lcout => \eeprom.n2613\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_unary_minus_2_inv_0_i15_1_lut_LC_5_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13585\,
            lcout => \eeprom.n19_adj_429\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_mux_3_i4_3_lut_LC_5_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010011100100111"
        )
    port map (
            in0 => \N__22983\,
            in1 => \N__13547\,
            in2 => \N__23788\,
            in3 => \_gnd_net_\,
            lcout => \eeprom.n3722_adj_433\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1358_3_lut_LC_5_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13636\,
            in2 => \N__13616\,
            in3 => \N__13935\,
            lcout => \eeprom.n2114\,
            ltout => \eeprom.n2114_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i1_3_lut_LC_5_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14262\,
            in2 => \N__13538\,
            in3 => \N__14295\,
            lcout => \eeprom.n4463\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1356_3_lut_LC_5_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13884\,
            in2 => \N__13862\,
            in3 => \N__13936\,
            lcout => \eeprom.n2112\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1626_3_lut_LC_5_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13535\,
            in2 => \N__15983\,
            in3 => \N__13517\,
            lcout => \eeprom.n2510\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1361_3_lut_LC_5_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13678\,
            in2 => \N__13658\,
            in3 => \N__13931\,
            lcout => \eeprom.n2117\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1360_3_lut_LC_5_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13897\,
            in2 => \N__13949\,
            in3 => \N__15858\,
            lcout => \eeprom.n2116\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1634_3_lut_LC_5_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__13724\,
            in1 => \N__13694\,
            in2 => \_gnd_net_\,
            in3 => \N__15978\,
            lcout => \eeprom.n2518\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1352_2_lut_LC_5_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14068\,
            in2 => \_gnd_net_\,
            in3 => \N__13682\,
            lcout => \eeprom.n2086\,
            ltout => OPEN,
            carryin => \bfn_5_22_0_\,
            carryout => \eeprom.n3524\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1352_3_lut_LC_5_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27181\,
            in2 => \N__13679\,
            in3 => \N__13649\,
            lcout => \eeprom.n2085\,
            ltout => OPEN,
            carryin => \eeprom.n3524\,
            carryout => \eeprom.n3525\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1352_4_lut_LC_5_22_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__15868\,
            in3 => \N__13646\,
            lcout => \eeprom.n2084\,
            ltout => OPEN,
            carryin => \eeprom.n3525\,
            carryout => \eeprom.n3526\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1352_5_lut_LC_5_22_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__13756\,
            in3 => \N__13643\,
            lcout => \eeprom.n2083\,
            ltout => OPEN,
            carryin => \eeprom.n3526\,
            carryout => \eeprom.n3527\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1352_6_lut_LC_5_22_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__13640\,
            in3 => \N__13607\,
            lcout => \eeprom.n2082\,
            ltout => OPEN,
            carryin => \eeprom.n3527\,
            carryout => \eeprom.n3528\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1352_7_lut_LC_5_22_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__13813\,
            in3 => \N__13604\,
            lcout => \eeprom.n2081\,
            ltout => OPEN,
            carryin => \eeprom.n3528\,
            carryout => \eeprom.n3529\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1352_8_lut_LC_5_22_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__13886\,
            in3 => \N__13853\,
            lcout => \eeprom.n2080\,
            ltout => OPEN,
            carryin => \eeprom.n3529\,
            carryout => \eeprom.n3530\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1352_9_lut_LC_5_22_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13791\,
            in2 => \N__27729\,
            in3 => \N__13850\,
            lcout => \eeprom.n2079\,
            ltout => OPEN,
            carryin => \eeprom.n3530\,
            carryout => \eeprom.n3531\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1352_10_lut_LC_5_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001000001100000"
        )
    port map (
            in0 => \N__27629\,
            in1 => \N__13847\,
            in2 => \N__13950\,
            in3 => \N__13826\,
            lcout => \eeprom.n2110\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1357_3_lut_LC_5_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__13823\,
            in1 => \_gnd_net_\,
            in2 => \N__13817\,
            in3 => \N__13937\,
            lcout => \eeprom.n2113\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1355_3_lut_LC_5_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101011001010"
        )
    port map (
            in0 => \N__13796\,
            in1 => \N__13772\,
            in2 => \N__13951\,
            in3 => \_gnd_net_\,
            lcout => \eeprom.n2111\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i1_2_lut_LC_5_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__14556\,
            in3 => \N__16386\,
            lcout => \eeprom.n4461\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1359_3_lut_LC_5_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13766\,
            in2 => \N__13760\,
            in3 => \N__13938\,
            lcout => \eeprom.n2115\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i1_2_lut_adj_72_LC_5_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__14035\,
            in3 => \N__16522\,
            lcout => \eeprom.n7_adj_470\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1362_3_lut_LC_5_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__14072\,
            in1 => \_gnd_net_\,
            in2 => \N__14045\,
            in3 => \N__13939\,
            lcout => \eeprom.n2118\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1489_3_lut_LC_5_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16616\,
            in2 => \N__16636\,
            in3 => \N__16601\,
            lcout => \eeprom.n2309\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i1_4_lut_adj_50_LC_5_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__15780\,
            in1 => \N__15717\,
            in2 => \N__15819\,
            in3 => \N__14207\,
            lcout => OPEN,
            ltout => \eeprom.n4509_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2_4_lut_LC_5_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111100000"
        )
    port map (
            in0 => \N__14011\,
            in1 => \N__15579\,
            in2 => \N__13988\,
            in3 => \N__13974\,
            lcout => \eeprom.n8_adj_468\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1490_3_lut_LC_5_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16602\,
            in2 => \N__16655\,
            in3 => \N__16675\,
            lcout => \eeprom.n2310\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i1_2_lut_adj_25_LC_5_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16629\,
            in2 => \_gnd_net_\,
            in3 => \N__16547\,
            lcout => OPEN,
            ltout => \eeprom.n6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i4_4_lut_LC_5_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__16708\,
            in1 => \N__16674\,
            in2 => \N__13958\,
            in3 => \N__15698\,
            lcout => \eeprom.n2242\,
            ltout => \eeprom.n2242_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i4028_3_lut_LC_5_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16369\,
            in2 => \N__13955\,
            in3 => \N__13952\,
            lcout => \eeprom.n4872\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1360_rep_36_3_lut_LC_5_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13901\,
            in2 => \N__16365\,
            in3 => \N__14249\,
            lcout => \eeprom.n4801\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1426_3_lut_LC_5_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14531\,
            in2 => \N__14561\,
            in3 => \N__16339\,
            lcout => \eeprom.n2214\,
            ltout => \eeprom.n2214_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1493_3_lut_LC_5_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__16592\,
            in1 => \_gnd_net_\,
            in2 => \N__14231\,
            in3 => \N__16124\,
            lcout => \eeprom.n2313\,
            ltout => \eeprom.n2313_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i1_2_lut_adj_46_LC_5_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__14210\,
            in3 => \N__14145\,
            lcout => \eeprom.n4505\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_mux_3_i23_3_lut_LC_5_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__14201\,
            in1 => \N__22978\,
            in2 => \_gnd_net_\,
            in3 => \N__14189\,
            lcout => \eeprom.n2119\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1495_3_lut_LC_5_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16203\,
            in2 => \N__16181\,
            in3 => \N__16591\,
            lcout => \eeprom.n2315\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1422_3_lut_LC_5_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110010101100"
        )
    port map (
            in0 => \N__14414\,
            in1 => \N__14440\,
            in2 => \N__16364\,
            in3 => \_gnd_net_\,
            lcout => \eeprom.n2210\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1491_3_lut_LC_5_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__16685\,
            in1 => \N__16707\,
            in2 => \_gnd_net_\,
            in3 => \N__16593\,
            lcout => \eeprom.n2311\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i1_4_lut_LC_5_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000000000000"
        )
    port map (
            in0 => \N__14343\,
            in1 => \N__15750\,
            in2 => \N__14096\,
            in3 => \N__14084\,
            lcout => OPEN,
            ltout => \eeprom.n4225_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i3_4_lut_LC_5_26_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__14436\,
            in1 => \N__14478\,
            in2 => \N__14075\,
            in3 => \N__14398\,
            lcout => \eeprom.n2143\,
            ltout => \eeprom.n2143_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i4033_3_lut_LC_5_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__14272\,
            in1 => \_gnd_net_\,
            in2 => \N__14351\,
            in3 => \N__14245\,
            lcout => \eeprom.n2215\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1425_3_lut_LC_5_26_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__14492\,
            in1 => \_gnd_net_\,
            in2 => \N__16367\,
            in3 => \N__14519\,
            lcout => \eeprom.n2213\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1428_3_lut_LC_5_26_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14282\,
            in2 => \N__14315\,
            in3 => \N__16346\,
            lcout => \eeprom.n2216\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1423_3_lut_LC_5_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010011100100"
        )
    port map (
            in0 => \N__16353\,
            in1 => \N__14479\,
            in2 => \N__14456\,
            in3 => \_gnd_net_\,
            lcout => \eeprom.n2211\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1429_rep_30_3_lut_LC_5_26_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14324\,
            in2 => \N__16366\,
            in3 => \N__14344\,
            lcout => \eeprom.n2217\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1419_2_lut_LC_5_27_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15752\,
            in2 => \_gnd_net_\,
            in3 => \N__14348\,
            lcout => \eeprom.n2186\,
            ltout => OPEN,
            carryin => \bfn_5_27_0_\,
            carryout => \eeprom.n3532\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1419_3_lut_LC_5_27_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27627\,
            in2 => \N__14345\,
            in3 => \N__14318\,
            lcout => \eeprom.n2185\,
            ltout => OPEN,
            carryin => \eeprom.n3532\,
            carryout => \eeprom.n3533\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1419_4_lut_LC_5_27_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__14314\,
            in3 => \N__14276\,
            lcout => \eeprom.n2184\,
            ltout => OPEN,
            carryin => \eeprom.n3533\,
            carryout => \eeprom.n3534\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1419_5_lut_LC_5_27_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__14273\,
            in3 => \N__14234\,
            lcout => \eeprom.n2183\,
            ltout => OPEN,
            carryin => \eeprom.n3534\,
            carryout => \eeprom.n3535\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1419_6_lut_LC_5_27_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14557\,
            in2 => \_gnd_net_\,
            in3 => \N__14522\,
            lcout => \eeprom.n2182\,
            ltout => OPEN,
            carryin => \eeprom.n3535\,
            carryout => \eeprom.n3536\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1419_7_lut_LC_5_27_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14515\,
            in2 => \_gnd_net_\,
            in3 => \N__14486\,
            lcout => \eeprom.n2181\,
            ltout => OPEN,
            carryin => \eeprom.n3536\,
            carryout => \eeprom.n3537\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1419_8_lut_LC_5_27_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__16397\,
            in3 => \N__14483\,
            lcout => \eeprom.n2180\,
            ltout => OPEN,
            carryin => \eeprom.n3537\,
            carryout => \eeprom.n3538\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1419_9_lut_LC_5_27_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27628\,
            in2 => \N__14480\,
            in3 => \N__14447\,
            lcout => \eeprom.n2179\,
            ltout => OPEN,
            carryin => \eeprom.n3538\,
            carryout => \eeprom.n3539\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1419_10_lut_LC_5_28_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27612\,
            in2 => \N__14444\,
            in3 => \N__14405\,
            lcout => \eeprom.n2178\,
            ltout => OPEN,
            carryin => \bfn_5_28_0_\,
            carryout => \eeprom.n3540\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1419_11_lut_LC_5_28_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001000001100000"
        )
    port map (
            in0 => \N__27613\,
            in1 => \N__14402\,
            in2 => \N__16370\,
            in3 => \N__14381\,
            lcout => \eeprom.n2209\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_287__i0_LC_5_29_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14378\,
            in2 => \_gnd_net_\,
            in3 => \N__14372\,
            lcout => n26,
            ltout => OPEN,
            carryin => \bfn_5_29_0_\,
            carryout => n3485,
            clk => \N__24346\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_287__i1_LC_5_29_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14369\,
            in2 => \_gnd_net_\,
            in3 => \N__14363\,
            lcout => n25,
            ltout => OPEN,
            carryin => n3485,
            carryout => n3486,
            clk => \N__24346\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_287__i2_LC_5_29_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14360\,
            in2 => \_gnd_net_\,
            in3 => \N__14354\,
            lcout => n24,
            ltout => OPEN,
            carryin => n3486,
            carryout => n3487,
            clk => \N__24346\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_287__i3_LC_5_29_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14633\,
            in2 => \_gnd_net_\,
            in3 => \N__14627\,
            lcout => n23,
            ltout => OPEN,
            carryin => n3487,
            carryout => n3488,
            clk => \N__24346\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_287__i4_LC_5_29_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14624\,
            in2 => \_gnd_net_\,
            in3 => \N__14618\,
            lcout => n22,
            ltout => OPEN,
            carryin => n3488,
            carryout => n3489,
            clk => \N__24346\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_287__i5_LC_5_29_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14615\,
            in2 => \_gnd_net_\,
            in3 => \N__14609\,
            lcout => n21,
            ltout => OPEN,
            carryin => n3489,
            carryout => n3490,
            clk => \N__24346\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_287__i6_LC_5_29_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14606\,
            in2 => \_gnd_net_\,
            in3 => \N__14600\,
            lcout => n20,
            ltout => OPEN,
            carryin => n3490,
            carryout => n3491,
            clk => \N__24346\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_287__i7_LC_5_29_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14597\,
            in2 => \_gnd_net_\,
            in3 => \N__14591\,
            lcout => n19,
            ltout => OPEN,
            carryin => n3491,
            carryout => n3492,
            clk => \N__24346\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_287__i8_LC_5_30_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14588\,
            in2 => \_gnd_net_\,
            in3 => \N__14582\,
            lcout => n18,
            ltout => OPEN,
            carryin => \bfn_5_30_0_\,
            carryout => n3493,
            clk => \N__24347\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_287__i9_LC_5_30_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14579\,
            in2 => \_gnd_net_\,
            in3 => \N__14573\,
            lcout => n17,
            ltout => OPEN,
            carryin => n3493,
            carryout => n3494,
            clk => \N__24347\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_287__i10_LC_5_30_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14570\,
            in2 => \_gnd_net_\,
            in3 => \N__14564\,
            lcout => n16,
            ltout => OPEN,
            carryin => n3494,
            carryout => n3495,
            clk => \N__24347\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_287__i11_LC_5_30_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14705\,
            in2 => \_gnd_net_\,
            in3 => \N__14699\,
            lcout => n15,
            ltout => OPEN,
            carryin => n3495,
            carryout => n3496,
            clk => \N__24347\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_287__i12_LC_5_30_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14696\,
            in2 => \_gnd_net_\,
            in3 => \N__14690\,
            lcout => n14,
            ltout => OPEN,
            carryin => n3496,
            carryout => n3497,
            clk => \N__24347\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_287__i13_LC_5_30_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14687\,
            in2 => \_gnd_net_\,
            in3 => \N__14681\,
            lcout => n13,
            ltout => OPEN,
            carryin => n3497,
            carryout => n3498,
            clk => \N__24347\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_287__i14_LC_5_30_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14678\,
            in2 => \_gnd_net_\,
            in3 => \N__14672\,
            lcout => n12,
            ltout => OPEN,
            carryin => n3498,
            carryout => n3499,
            clk => \N__24347\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_287__i15_LC_5_30_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14669\,
            in2 => \_gnd_net_\,
            in3 => \N__14663\,
            lcout => n11,
            ltout => OPEN,
            carryin => n3499,
            carryout => n3500,
            clk => \N__24347\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_287__i16_LC_5_31_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14660\,
            in2 => \_gnd_net_\,
            in3 => \N__14654\,
            lcout => n10,
            ltout => OPEN,
            carryin => \bfn_5_31_0_\,
            carryout => n3501,
            clk => \N__24348\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_287__i17_LC_5_31_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14651\,
            in2 => \_gnd_net_\,
            in3 => \N__14645\,
            lcout => n9,
            ltout => OPEN,
            carryin => n3501,
            carryout => n3502,
            clk => \N__24348\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_287__i18_LC_5_31_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14642\,
            in2 => \_gnd_net_\,
            in3 => \N__14636\,
            lcout => n8,
            ltout => OPEN,
            carryin => n3502,
            carryout => n3503,
            clk => \N__24348\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_287__i19_LC_5_31_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14822\,
            in2 => \_gnd_net_\,
            in3 => \N__14816\,
            lcout => n7,
            ltout => OPEN,
            carryin => n3503,
            carryout => n3504,
            clk => \N__24348\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_287__i20_LC_5_31_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14813\,
            in2 => \_gnd_net_\,
            in3 => \N__14807\,
            lcout => n6,
            ltout => OPEN,
            carryin => n3504,
            carryout => n3505,
            clk => \N__24348\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_287__i21_LC_5_31_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14799\,
            in2 => \_gnd_net_\,
            in3 => \N__14786\,
            lcout => blink_counter_21,
            ltout => OPEN,
            carryin => n3505,
            carryout => n3506,
            clk => \N__24348\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_287__i22_LC_5_31_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14781\,
            in2 => \_gnd_net_\,
            in3 => \N__14768\,
            lcout => blink_counter_22,
            ltout => OPEN,
            carryin => n3506,
            carryout => n3507,
            clk => \N__24348\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_287__i23_LC_5_31_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14760\,
            in2 => \_gnd_net_\,
            in3 => \N__14747\,
            lcout => blink_counter_23,
            ltout => OPEN,
            carryin => n3507,
            carryout => n3508,
            clk => \N__24348\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_287__i24_LC_5_32_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14742\,
            in2 => \_gnd_net_\,
            in3 => \N__14729\,
            lcout => blink_counter_24,
            ltout => OPEN,
            carryin => \bfn_5_32_0_\,
            carryout => n3509,
            clk => \N__24350\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_287__i25_LC_5_32_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14722\,
            in2 => \_gnd_net_\,
            in3 => \N__14726\,
            lcout => blink_counter_25,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24350\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1754_2_lut_LC_6_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16761\,
            in2 => \_gnd_net_\,
            in3 => \N__14711\,
            lcout => \eeprom.n2686\,
            ltout => OPEN,
            carryin => \bfn_6_18_0_\,
            carryout => \eeprom.n3587\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1754_3_lut_LC_6_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27779\,
            in2 => \N__16811\,
            in3 => \N__14708\,
            lcout => \eeprom.n2685\,
            ltout => OPEN,
            carryin => \eeprom.n3587\,
            carryout => \eeprom.n3588\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1754_4_lut_LC_6_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__16891\,
            in3 => \N__14849\,
            lcout => \eeprom.n2684\,
            ltout => OPEN,
            carryin => \eeprom.n3588\,
            carryout => \eeprom.n3589\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1754_5_lut_LC_6_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__16915\,
            in3 => \N__14846\,
            lcout => \eeprom.n2683\,
            ltout => OPEN,
            carryin => \eeprom.n3589\,
            carryout => \eeprom.n3590\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1754_6_lut_LC_6_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__17002\,
            in3 => \N__14843\,
            lcout => \eeprom.n2682\,
            ltout => OPEN,
            carryin => \eeprom.n3590\,
            carryout => \eeprom.n3591\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1754_7_lut_LC_6_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__16855\,
            in3 => \N__14840\,
            lcout => \eeprom.n2681\,
            ltout => OPEN,
            carryin => \eeprom.n3591\,
            carryout => \eeprom.n3592\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1754_8_lut_LC_6_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__16426\,
            in3 => \N__14837\,
            lcout => \eeprom.n2680\,
            ltout => OPEN,
            carryin => \eeprom.n3592\,
            carryout => \eeprom.n3593\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1754_9_lut_LC_6_18_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27780\,
            in2 => \N__16498\,
            in3 => \N__14834\,
            lcout => \eeprom.n2679\,
            ltout => OPEN,
            carryin => \eeprom.n3593\,
            carryout => \eeprom.n3594\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1754_10_lut_LC_6_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27756\,
            in2 => \N__15419\,
            in3 => \N__14831\,
            lcout => \eeprom.n2678\,
            ltout => OPEN,
            carryin => \bfn_6_19_0_\,
            carryout => \eeprom.n3595\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1754_11_lut_LC_6_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17254\,
            in2 => \N__27786\,
            in3 => \N__14828\,
            lcout => \eeprom.n2677\,
            ltout => OPEN,
            carryin => \eeprom.n3595\,
            carryout => \eeprom.n3596\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1754_12_lut_LC_6_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27760\,
            in2 => \N__14879\,
            in3 => \N__14825\,
            lcout => \eeprom.n2676\,
            ltout => OPEN,
            carryin => \eeprom.n3596\,
            carryout => \eeprom.n3597\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1754_13_lut_LC_6_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27748\,
            in2 => \N__16985\,
            in3 => \N__14942\,
            lcout => \eeprom.n2675\,
            ltout => OPEN,
            carryin => \eeprom.n3597\,
            carryout => \eeprom.n3598\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1754_14_lut_LC_6_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27761\,
            in2 => \N__16958\,
            in3 => \N__14939\,
            lcout => \eeprom.n2674\,
            ltout => OPEN,
            carryin => \eeprom.n3598\,
            carryout => \eeprom.n3599\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1754_15_lut_LC_6_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16456\,
            in2 => \N__27787\,
            in3 => \N__14936\,
            lcout => \eeprom.n2673\,
            ltout => OPEN,
            carryin => \eeprom.n3599\,
            carryout => \eeprom.n3600\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1754_16_lut_LC_6_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000010001001000"
        )
    port map (
            in0 => \N__27749\,
            in1 => \N__17213\,
            in2 => \N__15437\,
            in3 => \N__14933\,
            lcout => \eeprom.n2704\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1702_3_lut_LC_6_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__15164\,
            in1 => \N__15191\,
            in2 => \_gnd_net_\,
            in3 => \N__15499\,
            lcout => \eeprom.n2618\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_mux_3_i13_3_lut_LC_6_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__14930\,
            in1 => \N__22942\,
            in2 => \_gnd_net_\,
            in3 => \N__14918\,
            lcout => \eeprom.n3119\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_unary_minus_2_inv_0_i5_1_lut_LC_6_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23710\,
            lcout => \eeprom.n29_adj_460\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1760_3_lut_LC_6_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14878\,
            in2 => \N__14858\,
            in3 => \N__17212\,
            lcout => \eeprom.n2708\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1695_3_lut_LC_6_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__16052\,
            in1 => \_gnd_net_\,
            in2 => \N__15386\,
            in3 => \N__15494\,
            lcout => \eeprom.n2611\,
            ltout => \eeprom.n2611_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1762_3_lut_LC_6_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15200\,
            in2 => \N__15194\,
            in3 => \N__17211\,
            lcout => \eeprom.n2710\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1691_3_lut_LC_6_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15284\,
            in2 => \N__15242\,
            in3 => \N__15498\,
            lcout => \eeprom.n2607\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1692_3_lut_LC_6_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15296\,
            in2 => \N__15517\,
            in3 => \N__15335\,
            lcout => \eeprom.n2608\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1687_2_lut_LC_6_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15187\,
            in2 => \_gnd_net_\,
            in3 => \N__15155\,
            lcout => \eeprom.n2586\,
            ltout => OPEN,
            carryin => \bfn_6_21_0_\,
            carryout => \eeprom.n3574\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1687_3_lut_LC_6_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27754\,
            in2 => \N__15148\,
            in3 => \N__15116\,
            lcout => \eeprom.n2585\,
            ltout => OPEN,
            carryin => \eeprom.n3574\,
            carryout => \eeprom.n3575\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1687_4_lut_LC_6_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__15113\,
            in3 => \N__15071\,
            lcout => \eeprom.n2584\,
            ltout => OPEN,
            carryin => \eeprom.n3575\,
            carryout => \eeprom.n3576\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1687_5_lut_LC_6_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__15068\,
            in3 => \N__15023\,
            lcout => \eeprom.n2583\,
            ltout => OPEN,
            carryin => \eeprom.n3576\,
            carryout => \eeprom.n3577\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1687_6_lut_LC_6_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__15019\,
            in3 => \N__14975\,
            lcout => \eeprom.n2582\,
            ltout => OPEN,
            carryin => \eeprom.n3577\,
            carryout => \eeprom.n3578\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1687_7_lut_LC_6_21_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__14972\,
            in3 => \N__15392\,
            lcout => \eeprom.n2581\,
            ltout => OPEN,
            carryin => \eeprom.n3578\,
            carryout => \eeprom.n3579\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1687_8_lut_LC_6_21_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__15551\,
            in3 => \N__15389\,
            lcout => \eeprom.n2580\,
            ltout => OPEN,
            carryin => \eeprom.n3579\,
            carryout => \eeprom.n3580\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1687_9_lut_LC_6_21_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27755\,
            in2 => \N__16051\,
            in3 => \N__15377\,
            lcout => \eeprom.n2579\,
            ltout => OPEN,
            carryin => \eeprom.n3580\,
            carryout => \eeprom.n3581\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1687_10_lut_LC_6_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27179\,
            in2 => \N__15652\,
            in3 => \N__15374\,
            lcout => \eeprom.n2578\,
            ltout => OPEN,
            carryin => \bfn_6_22_0_\,
            carryout => \eeprom.n3582\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1687_11_lut_LC_6_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27648\,
            in2 => \N__15371\,
            in3 => \N__15338\,
            lcout => \eeprom.n2577\,
            ltout => OPEN,
            carryin => \eeprom.n3582\,
            carryout => \eeprom.n3583\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1687_12_lut_LC_6_22_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27180\,
            in2 => \N__15334\,
            in3 => \N__15287\,
            lcout => \eeprom.n2576\,
            ltout => OPEN,
            carryin => \eeprom.n3583\,
            carryout => \eeprom.n3584\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1687_13_lut_LC_6_22_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27649\,
            in2 => \N__15283\,
            in3 => \N__15230\,
            lcout => \eeprom.n2575\,
            ltout => OPEN,
            carryin => \eeprom.n3584\,
            carryout => \eeprom.n3585\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1687_14_lut_LC_6_22_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15897\,
            in2 => \N__27753\,
            in3 => \N__15227\,
            lcout => \eeprom.n2574\,
            ltout => OPEN,
            carryin => \eeprom.n3585\,
            carryout => \eeprom.n3586\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1687_15_lut_LC_6_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001000001100000"
        )
    port map (
            in0 => \N__15224\,
            in1 => \N__27653\,
            in2 => \N__15520\,
            in3 => \N__15203\,
            lcout => \eeprom.n2605\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1627_3_lut_LC_6_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15692\,
            in2 => \N__15668\,
            in3 => \N__15982\,
            lcout => \eeprom.n2511\,
            ltout => \eeprom.n2511_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1694_3_lut_LC_6_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100011011000"
        )
    port map (
            in0 => \N__15512\,
            in1 => \N__15635\,
            in2 => \N__15629\,
            in3 => \_gnd_net_\,
            lcout => \eeprom.n2610\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_mux_3_i22_3_lut_LC_6_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__15626\,
            in1 => \N__22979\,
            in2 => \_gnd_net_\,
            in3 => \N__15617\,
            lcout => \eeprom.n2219\,
            ltout => \eeprom.n2219_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1498_3_lut_LC_6_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16274\,
            in2 => \N__15587\,
            in3 => \N__16600\,
            lcout => \eeprom.n2318\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1696_3_lut_LC_6_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__15560\,
            in1 => \N__15547\,
            in2 => \_gnd_net_\,
            in3 => \N__15513\,
            lcout => \eeprom.n2612\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1690_3_lut_LC_6_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15898\,
            in2 => \N__15521\,
            in3 => \N__15446\,
            lcout => \eeprom.n2606\,
            ltout => \eeprom.n2606_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i1_2_lut_adj_85_LC_6_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__15440\,
            in3 => \N__15430\,
            lcout => OPEN,
            ltout => \eeprom.n10_adj_475_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i7_4_lut_adj_87_LC_6_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__17247\,
            in1 => \N__15418\,
            in2 => \N__15401\,
            in3 => \N__16485\,
            lcout => \eeprom.n16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1628_3_lut_LC_6_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16091\,
            in2 => \N__16067\,
            in3 => \N__15973\,
            lcout => \eeprom.n2512\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1623_3_lut_LC_6_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16022\,
            in2 => \N__15998\,
            in3 => \N__15972\,
            lcout => \eeprom.n2507\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1427_rep_34_3_lut_LC_6_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15875\,
            in2 => \N__16154\,
            in3 => \N__16597\,
            lcout => OPEN,
            ltout => \eeprom.n4799_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1494_3_lut_LC_6_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__15869\,
            in1 => \_gnd_net_\,
            in2 => \N__15839\,
            in3 => \N__15836\,
            lcout => \eeprom.n2314\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i4036_3_lut_LC_6_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16214\,
            in2 => \N__16238\,
            in3 => \N__16599\,
            lcout => \eeprom.n2316\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1430_3_lut_LC_6_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__15761\,
            in1 => \N__15751\,
            in2 => \_gnd_net_\,
            in3 => \N__16354\,
            lcout => \eeprom.n2218\,
            ltout => \eeprom.n2218_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1497_3_lut_LC_6_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__16247\,
            in1 => \_gnd_net_\,
            in2 => \N__15731\,
            in3 => \N__16598\,
            lcout => \eeprom.n2317\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i1_4_lut_adj_24_LC_6_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__16165\,
            in1 => \N__16135\,
            in2 => \N__16204\,
            in3 => \N__16230\,
            lcout => OPEN,
            ltout => \eeprom.n4447_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i1_4_lut_adj_26_LC_6_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010000000"
        )
    port map (
            in0 => \N__16289\,
            in1 => \N__16107\,
            in2 => \N__15701\,
            in3 => \N__16258\,
            lcout => \eeprom.n4218\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1424_3_lut_LC_6_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16396\,
            in2 => \N__16368\,
            in3 => \N__16298\,
            lcout => \eeprom.n2212\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1486_2_lut_LC_6_26_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16288\,
            in2 => \_gnd_net_\,
            in3 => \N__16265\,
            lcout => \eeprom.n2286\,
            ltout => OPEN,
            carryin => \bfn_6_26_0_\,
            carryout => \eeprom.n3541\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1486_3_lut_LC_6_26_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27421\,
            in2 => \N__16262\,
            in3 => \N__16241\,
            lcout => \eeprom.n2285\,
            ltout => OPEN,
            carryin => \eeprom.n3541\,
            carryout => \eeprom.n3542\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1486_4_lut_LC_6_26_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__16237\,
            in3 => \N__16208\,
            lcout => \eeprom.n2284\,
            ltout => OPEN,
            carryin => \eeprom.n3542\,
            carryout => \eeprom.n3543\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1486_5_lut_LC_6_26_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__16205\,
            in3 => \N__16172\,
            lcout => \eeprom.n2283\,
            ltout => OPEN,
            carryin => \eeprom.n3543\,
            carryout => \eeprom.n3544\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1486_6_lut_LC_6_26_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__16169\,
            in3 => \N__16142\,
            lcout => \eeprom.n2282\,
            ltout => OPEN,
            carryin => \eeprom.n3544\,
            carryout => \eeprom.n3545\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1486_7_lut_LC_6_26_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__16139\,
            in3 => \N__16118\,
            lcout => \eeprom.n2281\,
            ltout => OPEN,
            carryin => \eeprom.n3545\,
            carryout => \eeprom.n3546\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1486_8_lut_LC_6_26_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__16114\,
            in3 => \N__16712\,
            lcout => \eeprom.n2280\,
            ltout => OPEN,
            carryin => \eeprom.n3546\,
            carryout => \eeprom.n3547\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1486_9_lut_LC_6_26_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27422\,
            in2 => \N__16709\,
            in3 => \N__16679\,
            lcout => \eeprom.n2279\,
            ltout => OPEN,
            carryin => \eeprom.n3547\,
            carryout => \eeprom.n3548\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1486_10_lut_LC_6_27_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27607\,
            in2 => \N__16676\,
            in3 => \N__16640\,
            lcout => \eeprom.n2278\,
            ltout => OPEN,
            carryin => \bfn_6_27_0_\,
            carryout => \eeprom.n3549\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1486_11_lut_LC_6_27_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16637\,
            in2 => \N__27743\,
            in3 => \N__16607\,
            lcout => \eeprom.n2277\,
            ltout => OPEN,
            carryin => \eeprom.n3549\,
            carryout => \eeprom.n3550\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1486_12_lut_LC_6_27_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000010001001000"
        )
    port map (
            in0 => \N__27611\,
            in1 => \N__16604\,
            in2 => \N__16546\,
            in3 => \N__16526\,
            lcout => \eeprom.n2308\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1763_3_lut_LC_7_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16499\,
            in2 => \N__16469\,
            in3 => \N__17222\,
            lcout => \eeprom.n2711\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1757_3_lut_LC_7_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__16460\,
            in1 => \_gnd_net_\,
            in2 => \N__17220\,
            in3 => \N__16439\,
            lcout => \eeprom.n2705\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1764_3_lut_LC_7_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__16433\,
            in1 => \N__16427\,
            in2 => \_gnd_net_\,
            in3 => \N__17210\,
            lcout => \eeprom.n2712\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1765_3_lut_LC_7_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16856\,
            in2 => \N__17221\,
            in3 => \N__16826\,
            lcout => \eeprom.n2713\,
            ltout => \eeprom.n2713_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i1_2_lut_adj_29_LC_7_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__16820\,
            in3 => \N__17376\,
            lcout => OPEN,
            ltout => \eeprom.n4695_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i1_4_lut_adj_30_LC_7_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__17046\,
            in1 => \N__17430\,
            in2 => \N__16817\,
            in3 => \N__17319\,
            lcout => \eeprom.n4699\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i6_4_lut_LC_7_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__18132\,
            in1 => \N__17706\,
            in2 => \N__17518\,
            in3 => \N__18459\,
            lcout => OPEN,
            ltout => \eeprom.n16_adj_416_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i8_3_lut_LC_7_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18504\,
            in2 => \N__16814\,
            in3 => \N__17487\,
            lcout => \eeprom.n18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1769_3_lut_LC_7_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16810\,
            in2 => \N__16790\,
            in3 => \N__17203\,
            lcout => \eeprom.n2717\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1758_3_lut_LC_7_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110010101100"
        )
    port map (
            in0 => \N__16781\,
            in1 => \N__16953\,
            in2 => \N__17219\,
            in3 => \_gnd_net_\,
            lcout => \eeprom.n2706\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1770_3_lut_LC_7_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__16775\,
            in1 => \N__16763\,
            in2 => \_gnd_net_\,
            in3 => \N__17194\,
            lcout => \eeprom.n2718\,
            ltout => \eeprom.n2718_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i3_4_lut_adj_31_LC_7_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011001100"
        )
    port map (
            in0 => \N__17126\,
            in1 => \N__18369\,
            in2 => \N__16736\,
            in3 => \N__16733\,
            lcout => \eeprom.n13_adj_417\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1759_3_lut_LC_7_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__16981\,
            in1 => \_gnd_net_\,
            in2 => \N__17018\,
            in3 => \N__17202\,
            lcout => \eeprom.n2707\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1766_3_lut_LC_7_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17009\,
            in2 => \N__17218\,
            in3 => \N__17003\,
            lcout => \eeprom.n2714\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i8_4_lut_LC_7_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__16980\,
            in1 => \N__16967\,
            in2 => \N__16957\,
            in3 => \N__16937\,
            lcout => \eeprom.n2638\,
            ltout => \eeprom.n2638_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1767_3_lut_LC_7_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__16925\,
            in1 => \_gnd_net_\,
            in2 => \N__16919\,
            in3 => \N__16916\,
            lcout => \eeprom.n2715\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1768_3_lut_LC_7_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16892\,
            in2 => \N__16868\,
            in3 => \N__17198\,
            lcout => \eeprom.n2716\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1837_3_lut_LC_7_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110010101100"
        )
    port map (
            in0 => \N__17066\,
            in1 => \N__17080\,
            in2 => \N__18313\,
            in3 => \_gnd_net_\,
            lcout => \eeprom.n2817\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1838_3_lut_LC_7_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__17122\,
            in1 => \N__17093\,
            in2 => \_gnd_net_\,
            in3 => \N__18278\,
            lcout => \eeprom.n2818\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1835_3_lut_LC_7_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17050\,
            in2 => \N__18314\,
            in3 => \N__17030\,
            lcout => \eeprom.n2815\,
            ltout => \eeprom.n2815_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i1_2_lut_adj_32_LC_7_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__16859\,
            in3 => \N__19615\,
            lcout => \eeprom.n4529\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_mux_3_i6_3_lut_LC_7_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001001110111"
        )
    port map (
            in0 => \N__22990\,
            in1 => \N__17273\,
            in2 => \_gnd_net_\,
            in3 => \N__23665\,
            lcout => \eeprom.n3720_adj_435\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1761_3_lut_LC_7_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17258\,
            in2 => \N__17231\,
            in3 => \N__17217\,
            lcout => \eeprom.n2709\,
            ltout => \eeprom.n2709_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i9_4_lut_LC_7_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__17458\,
            in1 => \N__17147\,
            in2 => \N__17138\,
            in3 => \N__17135\,
            lcout => \eeprom.n2737\,
            ltout => \eeprom.n2737_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1833_3_lut_LC_7_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__17303\,
            in1 => \_gnd_net_\,
            in2 => \N__17129\,
            in3 => \N__17323\,
            lcout => \eeprom.n2813\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1821_2_lut_LC_7_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17121\,
            in2 => \_gnd_net_\,
            in3 => \N__17087\,
            lcout => \eeprom.n2786\,
            ltout => OPEN,
            carryin => \bfn_7_21_0_\,
            carryout => \eeprom.n3601\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1821_3_lut_LC_7_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27589\,
            in2 => \N__17084\,
            in3 => \N__17060\,
            lcout => \eeprom.n2785\,
            ltout => OPEN,
            carryin => \eeprom.n3601\,
            carryout => \eeprom.n3602\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1821_4_lut_LC_7_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__17437\,
            in3 => \N__17057\,
            lcout => \eeprom.n2784\,
            ltout => OPEN,
            carryin => \eeprom.n3602\,
            carryout => \eeprom.n3603\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1821_5_lut_LC_7_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__17054\,
            in3 => \N__17024\,
            lcout => \eeprom.n2783\,
            ltout => OPEN,
            carryin => \eeprom.n3603\,
            carryout => \eeprom.n3604\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1821_6_lut_LC_7_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__17389\,
            in3 => \N__17021\,
            lcout => \eeprom.n2782\,
            ltout => OPEN,
            carryin => \eeprom.n3604\,
            carryout => \eeprom.n3605\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1821_7_lut_LC_7_21_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__17327\,
            in3 => \N__17297\,
            lcout => \eeprom.n2781\,
            ltout => OPEN,
            carryin => \eeprom.n3605\,
            carryout => \eeprom.n3606\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1821_8_lut_LC_7_21_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__17362\,
            in3 => \N__17294\,
            lcout => \eeprom.n2780\,
            ltout => OPEN,
            carryin => \eeprom.n3606\,
            carryout => \eeprom.n3607\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1821_9_lut_LC_7_21_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27590\,
            in2 => \N__18511\,
            in3 => \N__17291\,
            lcout => \eeprom.n2779\,
            ltout => OPEN,
            carryin => \eeprom.n3607\,
            carryout => \eeprom.n3608\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1821_10_lut_LC_7_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17457\,
            in2 => \N__27381\,
            in3 => \N__17288\,
            lcout => \eeprom.n2778\,
            ltout => OPEN,
            carryin => \bfn_7_22_0_\,
            carryout => \eeprom.n3609\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1821_11_lut_LC_7_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27174\,
            in2 => \N__17492\,
            in3 => \N__17285\,
            lcout => \eeprom.n2777\,
            ltout => OPEN,
            carryin => \eeprom.n3609\,
            carryout => \eeprom.n3610\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1821_12_lut_LC_7_22_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27642\,
            in2 => \N__17680\,
            in3 => \N__17282\,
            lcout => \eeprom.n2776\,
            ltout => OPEN,
            carryin => \eeprom.n3610\,
            carryout => \eeprom.n3611\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1821_13_lut_LC_7_22_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27175\,
            in2 => \N__18382\,
            in3 => \N__17279\,
            lcout => \eeprom.n2775\,
            ltout => OPEN,
            carryin => \eeprom.n3611\,
            carryout => \eeprom.n3612\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1821_14_lut_LC_7_22_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27643\,
            in2 => \N__18472\,
            in3 => \N__17276\,
            lcout => \eeprom.n2774\,
            ltout => OPEN,
            carryin => \eeprom.n3612\,
            carryout => \eeprom.n3613\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1821_15_lut_LC_7_22_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17713\,
            in2 => \N__27752\,
            in3 => \N__17528\,
            lcout => \eeprom.n2773\,
            ltout => OPEN,
            carryin => \eeprom.n3613\,
            carryout => \eeprom.n3614\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1821_16_lut_LC_7_22_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18139\,
            in2 => \N__27382\,
            in3 => \N__17525\,
            lcout => \eeprom.n2772\,
            ltout => OPEN,
            carryin => \eeprom.n3614\,
            carryout => \eeprom.n3615\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1821_17_lut_LC_7_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000010001001000"
        )
    port map (
            in0 => \N__27647\,
            in1 => \N__18326\,
            in2 => \N__17522\,
            in3 => \N__17501\,
            lcout => \eeprom.n2803\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1829_3_lut_LC_7_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17498\,
            in2 => \N__18339\,
            in3 => \N__17491\,
            lcout => \eeprom.n2809\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1830_3_lut_LC_7_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__17465\,
            in1 => \_gnd_net_\,
            in2 => \N__18338\,
            in3 => \N__17459\,
            lcout => \eeprom.n2810\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1836_3_lut_LC_7_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17438\,
            in2 => \N__17411\,
            in3 => \N__18315\,
            lcout => \eeprom.n2816\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1834_3_lut_LC_7_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17399\,
            in2 => \N__18337\,
            in3 => \N__17390\,
            lcout => \eeprom.n2814\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1832_3_lut_LC_7_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17363\,
            in2 => \N__17342\,
            in3 => \N__18319\,
            lcout => \eeprom.n2812\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2223_2_lut_LC_9_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20274\,
            in2 => \_gnd_net_\,
            in3 => \N__17330\,
            lcout => \eeprom.n3386\,
            ltout => OPEN,
            carryin => \bfn_9_17_0_\,
            carryout => \eeprom.n3706\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2223_3_lut_LC_9_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27727\,
            in2 => \N__18809\,
            in3 => \N__17555\,
            lcout => \eeprom.n3385\,
            ltout => OPEN,
            carryin => \eeprom.n3706\,
            carryout => \eeprom.n3707\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2223_4_lut_LC_9_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__19064\,
            in3 => \N__17552\,
            lcout => \eeprom.n3384\,
            ltout => OPEN,
            carryin => \eeprom.n3707\,
            carryout => \eeprom.n3708\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2223_5_lut_LC_9_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__20249\,
            in3 => \N__17549\,
            lcout => \eeprom.n3383\,
            ltout => OPEN,
            carryin => \eeprom.n3708\,
            carryout => \eeprom.n3709\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2223_6_lut_LC_9_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__19787\,
            in3 => \N__17546\,
            lcout => \eeprom.n3382\,
            ltout => OPEN,
            carryin => \eeprom.n3709\,
            carryout => \eeprom.n3710\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2223_7_lut_LC_9_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__20206\,
            in3 => \N__17543\,
            lcout => \eeprom.n3381\,
            ltout => OPEN,
            carryin => \eeprom.n3710\,
            carryout => \eeprom.n3711\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2223_8_lut_LC_9_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__20353\,
            in3 => \N__17540\,
            lcout => \eeprom.n3380\,
            ltout => OPEN,
            carryin => \eeprom.n3711\,
            carryout => \eeprom.n3712\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2223_9_lut_LC_9_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27728\,
            in2 => \N__17950\,
            in3 => \N__17537\,
            lcout => \eeprom.n3379\,
            ltout => OPEN,
            carryin => \eeprom.n3712\,
            carryout => \eeprom.n3713\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2223_10_lut_LC_9_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27769\,
            in2 => \N__20155\,
            in3 => \N__17534\,
            lcout => \eeprom.n3378\,
            ltout => OPEN,
            carryin => \bfn_9_18_0_\,
            carryout => \eeprom.n3714\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2223_11_lut_LC_9_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20385\,
            in2 => \N__27788\,
            in3 => \N__17531\,
            lcout => \eeprom.n3377\,
            ltout => OPEN,
            carryin => \eeprom.n3714\,
            carryout => \eeprom.n3715\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2223_12_lut_LC_9_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27773\,
            in2 => \N__18910\,
            in3 => \N__17582\,
            lcout => \eeprom.n3376\,
            ltout => OPEN,
            carryin => \eeprom.n3715\,
            carryout => \eeprom.n3716\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2223_13_lut_LC_9_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27776\,
            in2 => \N__19021\,
            in3 => \N__17579\,
            lcout => \eeprom.n3375\,
            ltout => OPEN,
            carryin => \eeprom.n3716\,
            carryout => \eeprom.n3717\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2223_14_lut_LC_9_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27774\,
            in2 => \N__17915\,
            in3 => \N__17576\,
            lcout => \eeprom.n3374\,
            ltout => OPEN,
            carryin => \eeprom.n3717\,
            carryout => \eeprom.n3718\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2223_15_lut_LC_9_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27777\,
            in2 => \N__18980\,
            in3 => \N__17573\,
            lcout => \eeprom.n3373\,
            ltout => OPEN,
            carryin => \eeprom.n3718\,
            carryout => \eeprom.n3719\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2223_16_lut_LC_9_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27775\,
            in2 => \N__18947\,
            in3 => \N__17570\,
            lcout => \eeprom.n3372\,
            ltout => OPEN,
            carryin => \eeprom.n3719\,
            carryout => \eeprom.n3720\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2223_17_lut_LC_9_18_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27778\,
            in2 => \N__18782\,
            in3 => \N__17567\,
            lcout => \eeprom.n3371\,
            ltout => OPEN,
            carryin => \eeprom.n3720\,
            carryout => \eeprom.n3721\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2223_18_lut_LC_9_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27560\,
            in2 => \N__20693\,
            in3 => \N__17564\,
            lcout => \eeprom.n3370\,
            ltout => OPEN,
            carryin => \bfn_9_19_0_\,
            carryout => \eeprom.n3722\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2223_19_lut_LC_9_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18756\,
            in2 => \N__27725\,
            in3 => \N__17561\,
            lcout => \eeprom.n3369\,
            ltout => OPEN,
            carryin => \eeprom.n3722\,
            carryout => \eeprom.n3723\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2223_20_lut_LC_9_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19309\,
            in2 => \N__27726\,
            in3 => \N__17558\,
            lcout => \eeprom.n3368\,
            ltout => OPEN,
            carryin => \eeprom.n3723\,
            carryout => \eeprom.n3724\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2223_21_lut_LC_9_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27569\,
            in2 => \N__19360\,
            in3 => \N__17615\,
            lcout => \eeprom.n3367\,
            ltout => OPEN,
            carryin => \eeprom.n3724\,
            carryout => \eeprom.n3725\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2223_22_lut_LC_9_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27564\,
            in2 => \N__20647\,
            in3 => \N__17612\,
            lcout => \eeprom.n3366\,
            ltout => OPEN,
            carryin => \eeprom.n3725\,
            carryout => \eeprom.n3726\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2223_23_lut_LC_9_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001000001100000"
        )
    port map (
            in0 => \N__27565\,
            in1 => \N__19336\,
            in2 => \N__20615\,
            in3 => \N__17609\,
            lcout => \eeprom.n3397\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2173_3_lut_LC_9_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20804\,
            in2 => \N__17591\,
            in3 => \N__19211\,
            lcout => \eeprom.n3313\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2156_2_lut_LC_9_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__19445\,
            in3 => \N__17606\,
            lcout => \eeprom.n3286\,
            ltout => OPEN,
            carryin => \bfn_9_20_0_\,
            carryout => \eeprom.n3686\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2156_3_lut_LC_9_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27556\,
            in2 => \N__19399\,
            in3 => \N__17603\,
            lcout => \eeprom.n3285\,
            ltout => OPEN,
            carryin => \eeprom.n3686\,
            carryout => \eeprom.n3687\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2156_4_lut_LC_9_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__20426\,
            in3 => \N__17600\,
            lcout => \eeprom.n3284\,
            ltout => OPEN,
            carryin => \eeprom.n3687\,
            carryout => \eeprom.n3688\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2156_5_lut_LC_9_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__20482\,
            in3 => \N__17597\,
            lcout => \eeprom.n3283\,
            ltout => OPEN,
            carryin => \eeprom.n3688\,
            carryout => \eeprom.n3689\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2156_6_lut_LC_9_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__19519\,
            in3 => \N__17594\,
            lcout => \eeprom.n3282\,
            ltout => OPEN,
            carryin => \eeprom.n3689\,
            carryout => \eeprom.n3690\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2156_7_lut_LC_9_20_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__20803\,
            in3 => \N__17645\,
            lcout => \eeprom.n3281\,
            ltout => OPEN,
            carryin => \eeprom.n3690\,
            carryout => \eeprom.n3691\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2156_8_lut_LC_9_20_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__19550\,
            in3 => \N__17642\,
            lcout => \eeprom.n3280\,
            ltout => OPEN,
            carryin => \eeprom.n3691\,
            carryout => \eeprom.n3692\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2156_9_lut_LC_9_20_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19112\,
            in2 => \N__27724\,
            in3 => \N__17639\,
            lcout => \eeprom.n3279\,
            ltout => OPEN,
            carryin => \eeprom.n3692\,
            carryout => \eeprom.n3693\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2156_10_lut_LC_9_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27670\,
            in2 => \N__21264\,
            in3 => \N__17636\,
            lcout => \eeprom.n3278\,
            ltout => OPEN,
            carryin => \bfn_9_21_0_\,
            carryout => \eeprom.n3694\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2156_11_lut_LC_9_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19139\,
            in2 => \N__27765\,
            in3 => \N__17633\,
            lcout => \eeprom.n3277\,
            ltout => OPEN,
            carryin => \eeprom.n3694\,
            carryout => \eeprom.n3695\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2156_12_lut_LC_9_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18035\,
            in2 => \N__27721\,
            in3 => \N__17630\,
            lcout => \eeprom.n3276\,
            ltout => OPEN,
            carryin => \eeprom.n3695\,
            carryout => \eeprom.n3696\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2156_13_lut_LC_9_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19090\,
            in2 => \N__27766\,
            in3 => \N__17627\,
            lcout => \eeprom.n3275\,
            ltout => OPEN,
            carryin => \eeprom.n3696\,
            carryout => \eeprom.n3697\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2156_14_lut_LC_9_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21559\,
            in2 => \N__27722\,
            in3 => \N__17624\,
            lcout => \eeprom.n3274\,
            ltout => OPEN,
            carryin => \eeprom.n3697\,
            carryout => \eeprom.n3698\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2156_15_lut_LC_9_21_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20830\,
            in2 => \N__27767\,
            in3 => \N__17621\,
            lcout => \eeprom.n3273\,
            ltout => OPEN,
            carryin => \eeprom.n3698\,
            carryout => \eeprom.n3699\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2156_16_lut_LC_9_21_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21676\,
            in2 => \N__27723\,
            in3 => \N__17618\,
            lcout => \eeprom.n3272\,
            ltout => OPEN,
            carryin => \eeprom.n3699\,
            carryout => \eeprom.n3700\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2156_17_lut_LC_9_21_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21306\,
            in2 => \N__27768\,
            in3 => \N__17735\,
            lcout => \eeprom.n3271\,
            ltout => OPEN,
            carryin => \eeprom.n3700\,
            carryout => \eeprom.n3701\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2156_18_lut_LC_9_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20449\,
            in2 => \N__27750\,
            in3 => \N__17732\,
            lcout => \eeprom.n3270\,
            ltout => OPEN,
            carryin => \bfn_9_22_0_\,
            carryout => \eeprom.n3702\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2156_19_lut_LC_9_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21925\,
            in2 => \N__27333\,
            in3 => \N__17729\,
            lcout => \eeprom.n3269\,
            ltout => OPEN,
            carryin => \eeprom.n3702\,
            carryout => \eeprom.n3703\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2156_20_lut_LC_9_22_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21580\,
            in2 => \N__27751\,
            in3 => \N__17726\,
            lcout => \eeprom.n3268\,
            ltout => OPEN,
            carryin => \eeprom.n3703\,
            carryout => \eeprom.n3704\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2156_21_lut_LC_9_22_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21889\,
            in2 => \N__27334\,
            in3 => \N__17723\,
            lcout => \eeprom.n3267\,
            ltout => OPEN,
            carryin => \eeprom.n3704\,
            carryout => \eeprom.n3705\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2156_22_lut_LC_9_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001000001100000"
        )
    port map (
            in0 => \N__27641\,
            in1 => \N__21650\,
            in2 => \N__19268\,
            in3 => \N__17720\,
            lcout => \eeprom.n3298\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1825_3_lut_LC_9_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17717\,
            in2 => \N__18340\,
            in3 => \N__17690\,
            lcout => \eeprom.n2805\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1828_3_lut_LC_9_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17681\,
            in2 => \N__17657\,
            in3 => \N__18327\,
            lcout => \eeprom.n2808\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1888_2_lut_LC_9_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18693\,
            in2 => \_gnd_net_\,
            in3 => \N__17765\,
            lcout => \eeprom.n2886\,
            ltout => OPEN,
            carryin => \bfn_9_23_0_\,
            carryout => \eeprom.n3616\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1888_3_lut_LC_9_23_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27459\,
            in2 => \N__18550\,
            in3 => \N__17762\,
            lcout => \eeprom.n2885\,
            ltout => OPEN,
            carryin => \eeprom.n3616\,
            carryout => \eeprom.n3617\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1888_4_lut_LC_9_23_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__20131\,
            in3 => \N__17759\,
            lcout => \eeprom.n2884\,
            ltout => OPEN,
            carryin => \eeprom.n3617\,
            carryout => \eeprom.n3618\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1888_5_lut_LC_9_23_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__18654\,
            in3 => \N__17756\,
            lcout => \eeprom.n2883\,
            ltout => OPEN,
            carryin => \eeprom.n3618\,
            carryout => \eeprom.n3619\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1888_6_lut_LC_9_23_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__18202\,
            in3 => \N__17753\,
            lcout => \eeprom.n2882\,
            ltout => OPEN,
            carryin => \eeprom.n3619\,
            carryout => \eeprom.n3620\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1888_7_lut_LC_9_23_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__18719\,
            in3 => \N__17750\,
            lcout => \eeprom.n2881\,
            ltout => OPEN,
            carryin => \eeprom.n3620\,
            carryout => \eeprom.n3621\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1888_8_lut_LC_9_23_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__19633\,
            in3 => \N__17747\,
            lcout => \eeprom.n2880\,
            ltout => OPEN,
            carryin => \eeprom.n3621\,
            carryout => \eeprom.n3622\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1888_9_lut_LC_9_23_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19668\,
            in2 => \N__27546\,
            in3 => \N__17744\,
            lcout => \eeprom.n2879\,
            ltout => OPEN,
            carryin => \eeprom.n3622\,
            carryout => \eeprom.n3623\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1888_10_lut_LC_9_24_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27411\,
            in2 => \N__19996\,
            in3 => \N__17741\,
            lcout => \eeprom.n2878\,
            ltout => OPEN,
            carryin => \bfn_9_24_0_\,
            carryout => \eeprom.n3624\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1888_11_lut_LC_9_24_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20071\,
            in2 => \N__27604\,
            in3 => \N__17738\,
            lcout => \eeprom.n2877\,
            ltout => OPEN,
            carryin => \eeprom.n3624\,
            carryout => \eeprom.n3625\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1888_12_lut_LC_9_24_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18621\,
            in2 => \N__27586\,
            in3 => \N__17801\,
            lcout => \eeprom.n2876\,
            ltout => OPEN,
            carryin => \eeprom.n3625\,
            carryout => \eeprom.n3626\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1888_13_lut_LC_9_24_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18862\,
            in2 => \N__27605\,
            in3 => \N__17798\,
            lcout => \eeprom.n2875\,
            ltout => OPEN,
            carryin => \eeprom.n3626\,
            carryout => \eeprom.n3627\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1888_14_lut_LC_9_24_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18251\,
            in2 => \N__27587\,
            in3 => \N__17795\,
            lcout => \eeprom.n2874\,
            ltout => OPEN,
            carryin => \eeprom.n3627\,
            carryout => \eeprom.n3628\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1888_15_lut_LC_9_24_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27393\,
            in2 => \N__18433\,
            in3 => \N__17792\,
            lcout => \eeprom.n2873\,
            ltout => OPEN,
            carryin => \eeprom.n3628\,
            carryout => \eeprom.n3629\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1888_16_lut_LC_9_24_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18409\,
            in2 => \N__27588\,
            in3 => \N__17789\,
            lcout => \eeprom.n2872\,
            ltout => OPEN,
            carryin => \eeprom.n3629\,
            carryout => \eeprom.n3630\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1888_17_lut_LC_9_24_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18587\,
            in2 => \N__27606\,
            in3 => \N__17786\,
            lcout => \eeprom.n2871\,
            ltout => OPEN,
            carryin => \eeprom.n3630\,
            carryout => \eeprom.n3631\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1888_18_lut_LC_9_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000010001001000"
        )
    port map (
            in0 => \N__27410\,
            in1 => \N__19959\,
            in2 => \N__18101\,
            in3 => \N__17783\,
            lcout => \eeprom.n2902\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1893_3_lut_LC_9_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18434\,
            in2 => \N__19967\,
            in3 => \N__17780\,
            lcout => \eeprom.n2905\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1892_3_lut_LC_9_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18410\,
            in2 => \N__17774\,
            in3 => \N__19963\,
            lcout => \eeprom.n2904\,
            ltout => \eeprom.n2904_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i7_4_lut_adj_37_LC_9_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__19703\,
            in1 => \N__19747\,
            in2 => \N__17870\,
            in3 => \N__21481\,
            lcout => \eeprom.n19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2178_3_lut_LC_10_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__19431\,
            in1 => \_gnd_net_\,
            in2 => \N__17867\,
            in3 => \N__19239\,
            lcout => \eeprom.n3318\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2177_3_lut_LC_10_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17852\,
            in2 => \N__19403\,
            in3 => \N__19240\,
            lcout => \eeprom.n3317\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2231_3_lut_LC_10_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18781\,
            in2 => \N__17843\,
            in3 => \N__20596\,
            lcout => \eeprom.n3403\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2174_3_lut_LC_10_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19520\,
            in2 => \N__19262\,
            in3 => \N__17834\,
            lcout => \eeprom.n3314\,
            ltout => \eeprom.n3314_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i1_3_lut_adj_96_LC_10_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19062\,
            in2 => \N__17825\,
            in3 => \N__20248\,
            lcout => \eeprom.n4721\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2164_3_lut_LC_10_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21680\,
            in2 => \N__19256\,
            in3 => \N__17822\,
            lcout => \eeprom.n3304\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i12_4_lut_adj_98_LC_10_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__17914\,
            in1 => \N__19017\,
            in2 => \N__17951\,
            in3 => \N__18906\,
            lcout => \eeprom.n28_adj_484\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2166_3_lut_LC_10_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__17810\,
            in1 => \_gnd_net_\,
            in2 => \N__19257\,
            in3 => \N__21563\,
            lcout => \eeprom.n3306\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2165_3_lut_LC_10_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17969\,
            in2 => \N__20840\,
            in3 => \N__19224\,
            lcout => \eeprom.n3305\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2172_3_lut_LC_10_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110010101100"
        )
    port map (
            in0 => \N__17960\,
            in1 => \N__19549\,
            in2 => \N__19254\,
            in3 => \_gnd_net_\,
            lcout => \eeprom.n3312\,
            ltout => \eeprom.n3312_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2239_3_lut_LC_10_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17933\,
            in2 => \N__17927\,
            in3 => \N__20607\,
            lcout => \eeprom.n3411\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2167_3_lut_LC_10_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19094\,
            in2 => \N__19255\,
            in3 => \N__17924\,
            lcout => \eeprom.n3307\,
            ltout => \eeprom.n3307_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2234_3_lut_LC_10_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__17900\,
            in1 => \_gnd_net_\,
            in2 => \N__17894\,
            in3 => \N__20606\,
            lcout => \eeprom.n3406\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i13_4_lut_adj_94_LC_10_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__19110\,
            in1 => \N__18033\,
            in2 => \N__19073\,
            in3 => \N__19373\,
            lcout => OPEN,
            ltout => \eeprom.n28_adj_482_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i14_4_lut_LC_10_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__21533\,
            in1 => \N__21265\,
            in2 => \N__17891\,
            in3 => \N__21632\,
            lcout => \eeprom.n3232\,
            ltout => \eeprom.n3232_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2170_3_lut_LC_10_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__17888\,
            in1 => \_gnd_net_\,
            in2 => \N__17879\,
            in3 => \N__21269\,
            lcout => \eeprom.n3310\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2227_3_lut_LC_10_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17876\,
            in2 => \N__19361\,
            in3 => \N__20578\,
            lcout => \eeprom.n3399\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2168_3_lut_LC_10_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18074\,
            in2 => \N__19258\,
            in3 => \N__18034\,
            lcout => \eeprom.n3308\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2171_3_lut_LC_10_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19111\,
            in2 => \N__18065\,
            in3 => \N__19225\,
            lcout => \eeprom.n3311\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2163_3_lut_LC_10_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__18056\,
            in1 => \_gnd_net_\,
            in2 => \N__19259\,
            in3 => \N__21311\,
            lcout => \eeprom.n3303\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2169_rep_54_3_lut_LC_10_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19135\,
            in2 => \N__18047\,
            in3 => \N__19226\,
            lcout => \eeprom.n3309\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2101_3_lut_LC_10_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24215\,
            in2 => \N__20873\,
            in3 => \N__21793\,
            lcout => \eeprom.n3209\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2229_3_lut_LC_10_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18020\,
            in2 => \N__20611\,
            in3 => \N__18757\,
            lcout => \eeprom.n3401\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_mux_3_i7_3_lut_LC_10_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010001110111"
        )
    port map (
            in0 => \N__18014\,
            in1 => \N__22950\,
            in2 => \_gnd_net_\,
            in3 => \N__23611\,
            lcout => \eeprom.n3719_adj_436\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2160_3_lut_LC_10_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21584\,
            in2 => \N__19260\,
            in3 => \N__17996\,
            lcout => \eeprom.n3300\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_mux_3_i2_3_lut_LC_10_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010001110111"
        )
    port map (
            in0 => \N__17987\,
            in1 => \N__22949\,
            in2 => \_gnd_net_\,
            in3 => \N__23908\,
            lcout => \eeprom.n3724_adj_335\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2161_3_lut_LC_10_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18212\,
            in2 => \N__19261\,
            in3 => \N__21926\,
            lcout => \eeprom.n3301\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1902_3_lut_LC_10_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18203\,
            in2 => \N__18179\,
            in3 => \N__19954\,
            lcout => \eeprom.n2914\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2110_3_lut_LC_10_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__20767\,
            in1 => \N__20726\,
            in2 => \_gnd_net_\,
            in3 => \N__21789\,
            lcout => \eeprom.n3218\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1906_3_lut_LC_10_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__18698\,
            in1 => \_gnd_net_\,
            in2 => \N__19966\,
            in3 => \N__18167\,
            lcout => \eeprom.n2918\,
            ltout => \eeprom.n2918_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1973_3_lut_LC_10_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19466\,
            in2 => \N__18155\,
            in3 => \N__24735\,
            lcout => \eeprom.n3017\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2100_3_lut_LC_10_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24248\,
            in2 => \N__21053\,
            in3 => \N__21790\,
            lcout => \eeprom.n3208\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2159_3_lut_LC_10_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21890\,
            in2 => \N__18152\,
            in3 => \N__19267\,
            lcout => \eeprom.n3299\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1824_3_lut_LC_10_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18143\,
            in2 => \N__18116\,
            in3 => \N__18336\,
            lcout => \eeprom.n2804\,
            ltout => \eeprom.n2804_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i9_4_lut_adj_34_LC_10_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__18094\,
            in1 => \N__19983\,
            in2 => \N__18077\,
            in3 => \N__18389\,
            lcout => \eeprom.n20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2162_3_lut_LC_10_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18521\,
            in2 => \N__20453\,
            in3 => \N__19266\,
            lcout => \eeprom.n3302\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1831_3_lut_LC_10_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18515\,
            in2 => \N__18341\,
            in3 => \N__18485\,
            lcout => \eeprom.n2811\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1826_3_lut_LC_10_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18473\,
            in2 => \N__18446\,
            in3 => \N__18332\,
            lcout => \eeprom.n2806\,
            ltout => \eeprom.n2806_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i7_4_lut_LC_10_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__18247\,
            in1 => \N__18855\,
            in2 => \N__18413\,
            in3 => \N__18402\,
            lcout => \eeprom.n18_adj_418\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1827_3_lut_LC_10_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18383\,
            in2 => \N__18353\,
            in3 => \N__18331\,
            lcout => \eeprom.n2807\,
            ltout => \eeprom.n2807_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1894_3_lut_LC_10_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18236\,
            in2 => \N__18227\,
            in3 => \N__19935\,
            lcout => \eeprom.n2906\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1901_3_lut_LC_10_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18718\,
            in2 => \N__18224\,
            in3 => \N__19930\,
            lcout => \eeprom.n2913\,
            ltout => \eeprom.n2913_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i1_2_lut_adj_27_LC_10_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__18215\,
            in3 => \N__19869\,
            lcout => \eeprom.n4703\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i1_4_lut_adj_33_LC_10_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__18731\,
            in1 => \N__18655\,
            in2 => \N__20132\,
            in3 => \N__18717\,
            lcout => OPEN,
            ltout => \eeprom.n4533_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i4_4_lut_adj_35_LC_10_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111100000"
        )
    port map (
            in0 => \N__18546\,
            in1 => \N__18694\,
            in2 => \N__18668\,
            in3 => \N__18622\,
            lcout => OPEN,
            ltout => \eeprom.n15_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i10_4_lut_LC_10_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__20070\,
            in1 => \N__18665\,
            in2 => \N__18659\,
            in3 => \N__19669\,
            lcout => \eeprom.n2836\,
            ltout => \eeprom.n2836_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1903_3_lut_LC_10_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__18656\,
            in1 => \_gnd_net_\,
            in2 => \N__18632\,
            in3 => \N__18629\,
            lcout => \eeprom.n2915\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1896_3_lut_LC_10_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__18623\,
            in1 => \_gnd_net_\,
            in2 => \N__18596\,
            in3 => \N__19934\,
            lcout => \eeprom.n2908\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1891_3_lut_LC_10_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18586\,
            in2 => \N__19958\,
            in3 => \N__18572\,
            lcout => \eeprom.n2903\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i10_4_lut_adj_38_LC_10_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__23178\,
            in1 => \N__18566\,
            in2 => \N__22125\,
            in3 => \N__18875\,
            lcout => OPEN,
            ltout => \eeprom.n22_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i11_4_lut_LC_10_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__20022\,
            in1 => \N__19842\,
            in2 => \N__18560\,
            in3 => \N__20042\,
            lcout => \eeprom.n2935\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1905_3_lut_LC_10_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18557\,
            in2 => \N__18551\,
            in3 => \N__19948\,
            lcout => \eeprom.n2917\,
            ltout => \eeprom.n2917_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i1_4_lut_adj_28_LC_10_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__21831\,
            in1 => \N__18887\,
            in2 => \N__18881\,
            in3 => \N__22080\,
            lcout => OPEN,
            ltout => \eeprom.n4707_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i3_4_lut_adj_36_LC_10_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011101010"
        )
    port map (
            in0 => \N__19733\,
            in1 => \N__24825\,
            in2 => \N__18878\,
            in3 => \N__19483\,
            lcout => \eeprom.n15_adj_419\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1895_3_lut_LC_10_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18869\,
            in2 => \N__19965\,
            in3 => \N__18863\,
            lcout => \eeprom.n2907\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2245_3_lut_LC_11_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18805\,
            in2 => \N__18839\,
            in3 => \N__20580\,
            lcout => \eeprom.n3417\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2175_3_lut_LC_11_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20483\,
            in2 => \N__18827\,
            in3 => \N__19253\,
            lcout => \eeprom.n3315\,
            ltout => \eeprom.n3315_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i1_2_lut_adj_95_LC_11_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__18812\,
            in3 => \N__20354\,
            lcout => OPEN,
            ltout => \eeprom.n4719_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i1_4_lut_adj_97_LC_11_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000000000000"
        )
    port map (
            in0 => \N__20281\,
            in1 => \N__18804\,
            in2 => \N__18791\,
            in3 => \N__18788\,
            lcout => OPEN,
            ltout => \eeprom.n4151_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i10_4_lut_adj_99_LC_11_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__18777\,
            in1 => \N__20688\,
            in2 => \N__18761\,
            in3 => \N__18758\,
            lcout => \eeprom.n26_adj_485\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2244_3_lut_LC_11_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19063\,
            in2 => \N__19043\,
            in3 => \N__20579\,
            lcout => \eeprom.n3416\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2235_3_lut_LC_11_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19031\,
            in2 => \N__20610\,
            in3 => \N__19022\,
            lcout => \eeprom.n3407\,
            ltout => \eeprom.n3407_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i12_4_lut_adj_108_LC_11_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__22155\,
            in1 => \N__22297\,
            in2 => \N__18998\,
            in3 => \N__22230\,
            lcout => \eeprom.n29_adj_491\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i11_4_lut_adj_100_LC_11_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__20386\,
            in1 => \N__18945\,
            in2 => \N__18979\,
            in3 => \N__20151\,
            lcout => OPEN,
            ltout => \eeprom.n27_adj_486_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i15_4_lut_LC_11_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__19316\,
            in1 => \N__18995\,
            in2 => \N__18989\,
            in3 => \N__18986\,
            lcout => \eeprom.n3331\,
            ltout => \eeprom.n3331_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2233_3_lut_LC_11_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__18975\,
            in1 => \_gnd_net_\,
            in2 => \N__18959\,
            in3 => \N__18956\,
            lcout => \eeprom.n3405\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2232_3_lut_LC_11_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__18946\,
            in1 => \_gnd_net_\,
            in2 => \N__20609\,
            in3 => \N__18929\,
            lcout => \eeprom.n3404\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i4038_3_lut_LC_11_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18920\,
            in2 => \N__18911\,
            in3 => \N__20588\,
            lcout => \eeprom.n3408\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i1_4_lut_adj_89_LC_11_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__20415\,
            in1 => \N__20469\,
            in2 => \N__20796\,
            in3 => \N__19367\,
            lcout => OPEN,
            ltout => \eeprom.n4615_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i6_4_lut_adj_90_LC_11_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011101100"
        )
    port map (
            in0 => \N__19438\,
            in1 => \N__19131\,
            in2 => \N__19406\,
            in3 => \N__19395\,
            lcout => \eeprom.n21_adj_477\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i1_2_lut_adj_88_LC_11_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__19512\,
            in3 => \N__19539\,
            lcout => \eeprom.n4611\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i9_4_lut_adj_101_LC_11_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__19353\,
            in1 => \N__19337\,
            in2 => \N__19310\,
            in3 => \N__20643\,
            lcout => \eeprom.n25_adj_487\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2228_3_lut_LC_11_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19308\,
            in2 => \N__19292\,
            in3 => \N__20595\,
            lcout => \eeprom.n3400\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2176_3_lut_LC_11_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19280\,
            in2 => \N__20425\,
            in3 => \N__19193\,
            lcout => \eeprom.n3316\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2102_3_lut_LC_11_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20888\,
            in2 => \N__21777\,
            in3 => \N__24283\,
            lcout => \eeprom.n3210\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2037_3_lut_LC_11_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26146\,
            in2 => \N__26117\,
            in3 => \N__27911\,
            lcout => \eeprom.n3113\,
            ltout => \eeprom.n3113_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2104_3_lut_LC_11_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__21746\,
            in1 => \_gnd_net_\,
            in2 => \N__19115\,
            in3 => \N__20906\,
            lcout => \eeprom.n3212\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i10_4_lut_adj_91_LC_11_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__20437\,
            in1 => \N__19089\,
            in2 => \N__20829\,
            in3 => \N__21310\,
            lcout => \eeprom.n25_adj_478\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2105_3_lut_LC_11_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21521\,
            in2 => \N__20939\,
            in3 => \N__21741\,
            lcout => \eeprom.n3213\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2040_3_lut_LC_11_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26283\,
            in2 => \N__27919\,
            in3 => \N__26267\,
            lcout => \eeprom.n3116\,
            ltout => \eeprom.n3116_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2107_3_lut_LC_11_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20960\,
            in2 => \N__19523\,
            in3 => \N__21742\,
            lcout => \eeprom.n3215\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1955_2_lut_LC_11_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24832\,
            in2 => \_gnd_net_\,
            in3 => \N__19487\,
            lcout => \eeprom.n2986\,
            ltout => OPEN,
            carryin => \bfn_11_21_0_\,
            carryout => \eeprom.n3632\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1955_3_lut_LC_11_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27325\,
            in2 => \N__19484\,
            in3 => \N__19460\,
            lcout => \eeprom.n2985\,
            ltout => OPEN,
            carryin => \eeprom.n3632\,
            carryout => \eeprom.n3633\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1955_4_lut_LC_11_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__19805\,
            in3 => \N__19457\,
            lcout => \eeprom.n2984\,
            ltout => OPEN,
            carryin => \eeprom.n3633\,
            carryout => \eeprom.n3634\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1955_5_lut_LC_11_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__21844\,
            in3 => \N__19454\,
            lcout => \eeprom.n2983\,
            ltout => OPEN,
            carryin => \eeprom.n3634\,
            carryout => \eeprom.n3635\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1955_6_lut_LC_11_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__19877\,
            in3 => \N__19451\,
            lcout => \eeprom.n2982\,
            ltout => OPEN,
            carryin => \eeprom.n3635\,
            carryout => \eeprom.n3636\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1955_7_lut_LC_11_21_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__22081\,
            in3 => \N__19448\,
            lcout => \eeprom.n2981\,
            ltout => OPEN,
            carryin => \eeprom.n3636\,
            carryout => \eeprom.n3637\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1955_8_lut_LC_11_21_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19604\,
            in2 => \_gnd_net_\,
            in3 => \N__19577\,
            lcout => \eeprom.n2980\,
            ltout => OPEN,
            carryin => \eeprom.n3637\,
            carryout => \eeprom.n3638\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1955_9_lut_LC_11_21_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27326\,
            in2 => \N__23188\,
            in3 => \N__19574\,
            lcout => \eeprom.n2979\,
            ltout => OPEN,
            carryin => \eeprom.n3638\,
            carryout => \eeprom.n3639\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1955_10_lut_LC_11_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19843\,
            in2 => \N__27543\,
            in3 => \N__19571\,
            lcout => \eeprom.n2978\,
            ltout => OPEN,
            carryin => \bfn_11_22_0_\,
            carryout => \eeprom.n3640\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1955_11_lut_LC_11_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27318\,
            in2 => \N__21080\,
            in3 => \N__19568\,
            lcout => \eeprom.n2977\,
            ltout => OPEN,
            carryin => \eeprom.n3640\,
            carryout => \eeprom.n3641\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1955_12_lut_LC_11_22_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27126\,
            in2 => \N__24797\,
            in3 => \N__19565\,
            lcout => \eeprom.n2976\,
            ltout => OPEN,
            carryin => \eeprom.n3641\,
            carryout => \eeprom.n3642\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1955_13_lut_LC_11_22_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20023\,
            in2 => \N__27330\,
            in3 => \N__19562\,
            lcout => \eeprom.n2975\,
            ltout => OPEN,
            carryin => \eeprom.n3642\,
            carryout => \eeprom.n3643\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1955_14_lut_LC_11_22_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22126\,
            in2 => \N__27544\,
            in3 => \N__19559\,
            lcout => \eeprom.n2974\,
            ltout => OPEN,
            carryin => \eeprom.n3643\,
            carryout => \eeprom.n3644\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1955_15_lut_LC_11_22_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19731\,
            in2 => \N__27331\,
            in3 => \N__19556\,
            lcout => \eeprom.n2973\,
            ltout => OPEN,
            carryin => \eeprom.n3644\,
            carryout => \eeprom.n3645\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1955_16_lut_LC_11_22_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21493\,
            in2 => \N__27545\,
            in3 => \N__19553\,
            lcout => \eeprom.n2972\,
            ltout => OPEN,
            carryin => \eeprom.n3645\,
            carryout => \eeprom.n3646\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1955_17_lut_LC_11_22_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21106\,
            in2 => \N__27332\,
            in3 => \N__19760\,
            lcout => \eeprom.n2971\,
            ltout => OPEN,
            carryin => \eeprom.n3646\,
            carryout => \eeprom.n3647\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1955_18_lut_LC_11_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19701\,
            in2 => \N__27541\,
            in3 => \N__19757\,
            lcout => \eeprom.n2970\,
            ltout => OPEN,
            carryin => \bfn_11_23_0_\,
            carryout => \eeprom.n3648\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1955_19_lut_LC_11_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001000001100000"
        )
    port map (
            in0 => \N__19754\,
            in1 => \N__27310\,
            in2 => \N__24758\,
            in3 => \N__19736\,
            lcout => \eeprom.n3001\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1961_3_lut_LC_11_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19732\,
            in2 => \N__19712\,
            in3 => \N__24727\,
            lcout => \eeprom.n3005\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1958_3_lut_LC_11_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__19702\,
            in1 => \_gnd_net_\,
            in2 => \N__24757\,
            in3 => \N__19685\,
            lcout => \eeprom.n3002\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1899_3_lut_LC_11_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19679\,
            in2 => \N__19964\,
            in3 => \N__19670\,
            lcout => \eeprom.n2911\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1900_3_lut_LC_11_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19646\,
            in2 => \N__19637\,
            in3 => \N__19944\,
            lcout => \eeprom.n2912\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1968_3_lut_LC_11_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19603\,
            in2 => \N__19589\,
            in3 => \N__24728\,
            lcout => \eeprom.n3012\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1904_3_lut_LC_11_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__20130\,
            in1 => \_gnd_net_\,
            in2 => \N__20096\,
            in3 => \N__19943\,
            lcout => \eeprom.n2916\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1897_3_lut_LC_11_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__19953\,
            in1 => \_gnd_net_\,
            in2 => \N__20084\,
            in3 => \N__20072\,
            lcout => \eeprom.n2909\,
            ltout => \eeprom.n2909_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i6_2_lut_LC_11_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__20045\,
            in3 => \N__21072\,
            lcout => \eeprom.n18_adj_420\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1963_3_lut_LC_11_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__24705\,
            in1 => \_gnd_net_\,
            in2 => \N__20036\,
            in3 => \N__20024\,
            lcout => \eeprom.n3007\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1898_3_lut_LC_11_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20006\,
            in2 => \N__19997\,
            in3 => \N__19952\,
            lcout => \eeprom.n2910\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1970_3_lut_LC_11_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__19873\,
            in1 => \_gnd_net_\,
            in2 => \N__24736\,
            in3 => \N__19853\,
            lcout => \eeprom.n3014\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1966_3_lut_LC_11_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19844\,
            in2 => \N__19826\,
            in3 => \N__24706\,
            lcout => \eeprom.n3010\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1972_3_lut_LC_11_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__19814\,
            in1 => \N__19801\,
            in2 => \_gnd_net_\,
            in3 => \N__24701\,
            lcout => \eeprom.n3016\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2242_3_lut_LC_12_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19783\,
            in2 => \N__20599\,
            in3 => \N__19769\,
            lcout => \eeprom.n3414\,
            ltout => \eeprom.n3414_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i1_3_lut_adj_104_LC_12_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23106\,
            in2 => \N__20303\,
            in3 => \N__23031\,
            lcout => OPEN,
            ltout => \eeprom.n4689_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i1_4_lut_adj_105_LC_12_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000000000000"
        )
    port map (
            in0 => \N__23421\,
            in1 => \N__23073\,
            in2 => \N__20300\,
            in3 => \N__20177\,
            lcout => OPEN,
            ltout => \eeprom.n4144_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i11_4_lut_adj_107_LC_12_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__23244\,
            in1 => \N__22674\,
            in2 => \N__20297\,
            in3 => \N__22635\,
            lcout => \eeprom.n28_adj_490\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2246_3_lut_LC_12_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20294\,
            in2 => \N__20597\,
            in3 => \N__20282\,
            lcout => \eeprom.n3418\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2243_3_lut_LC_12_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20244\,
            in2 => \N__20219\,
            in3 => \N__20557\,
            lcout => \eeprom.n3415\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2241_3_lut_LC_12_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20207\,
            in2 => \N__20598\,
            in3 => \N__20189\,
            lcout => \eeprom.n3413\,
            ltout => \eeprom.n3413_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i1_2_lut_adj_103_LC_12_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__20180\,
            in3 => \N__22002\,
            lcout => \eeprom.n4687\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2238_3_lut_LC_12_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20171\,
            in2 => \N__20162\,
            in3 => \N__20586\,
            lcout => \eeprom.n3410\,
            ltout => \eeprom.n3410_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2305_3_lut_LC_12_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22286\,
            in2 => \N__20399\,
            in3 => \N__23345\,
            lcout => \eeprom.n3509\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2373_3_lut_LC_12_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25013\,
            in2 => \N__25033\,
            in3 => \N__25659\,
            lcout => \eeprom.n3609_adj_445\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2301_3_lut_LC_12_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__23347\,
            in1 => \_gnd_net_\,
            in2 => \N__22142\,
            in3 => \N__22165\,
            lcout => \eeprom.n3505\,
            ltout => \eeprom.n3505_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i13_4_lut_adj_117_LC_12_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__24984\,
            in1 => \N__25026\,
            in2 => \N__20396\,
            in3 => \N__24870\,
            lcout => \eeprom.n31_adj_496\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2237_3_lut_LC_12_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20393\,
            in2 => \N__20369\,
            in3 => \N__20587\,
            lcout => \eeprom.n3409\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2302_3_lut_LC_12_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22178\,
            in2 => \N__22198\,
            in3 => \N__23346\,
            lcout => \eeprom.n3506\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2372_3_lut_LC_12_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24968\,
            in2 => \N__24994\,
            in3 => \N__25678\,
            lcout => OPEN,
            ltout => \eeprom.n3608_adj_451_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i1_4_lut_adj_54_LC_12_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011110100"
        )
    port map (
            in0 => \N__25679\,
            in1 => \N__25072\,
            in2 => \N__20357\,
            in3 => \N__25052\,
            lcout => \eeprom.n4581\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2240_3_lut_LC_12_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20352\,
            in2 => \N__20321\,
            in3 => \N__20581\,
            lcout => \eeprom.n3412\,
            ltout => \eeprom.n3412_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2307_3_lut_LC_12_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22355\,
            in2 => \N__20306\,
            in3 => \N__23353\,
            lcout => \eeprom.n3511_adj_362\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2230_3_lut_LC_12_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20692\,
            in2 => \N__20608\,
            in3 => \N__20666\,
            lcout => \eeprom.n3402\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2226_3_lut_LC_12_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20657\,
            in2 => \N__20648\,
            in3 => \N__20585\,
            lcout => \eeprom.n3398\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2296_3_lut_LC_12_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22544\,
            in2 => \N__22570\,
            in3 => \N__23362\,
            lcout => \eeprom.n3500\,
            ltout => \eeprom.n3500_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i11_4_lut_adj_118_LC_12_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__25393\,
            in1 => \N__25341\,
            in2 => \N__20486\,
            in3 => \N__25308\,
            lcout => \eeprom.n29_adj_497\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i10_4_lut_adj_109_LC_12_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__22563\,
            in1 => \N__22605\,
            in2 => \N__22524\,
            in3 => \N__22479\,
            lcout => \eeprom.n27_adj_492\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2108_3_lut_LC_12_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21391\,
            in2 => \N__20993\,
            in3 => \N__21772\,
            lcout => \eeprom.n3216\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2297_3_lut_LC_12_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22606\,
            in2 => \N__22592\,
            in3 => \N__23361\,
            lcout => \eeprom.n3501\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2095_3_lut_LC_12_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__21953\,
            in1 => \_gnd_net_\,
            in2 => \N__21791\,
            in3 => \N__21014\,
            lcout => \eeprom.n3203\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2109_3_lut_LC_12_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__21458\,
            in1 => \_gnd_net_\,
            in2 => \N__20708\,
            in3 => \N__21771\,
            lcout => \eeprom.n3217\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i4_4_lut_adj_47_LC_12_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011001100"
        )
    port map (
            in0 => \N__20768\,
            in1 => \N__21818\,
            in2 => \N__21454\,
            in3 => \N__20846\,
            lcout => OPEN,
            ltout => \eeprom.n18_adj_432_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i12_4_lut_adj_69_LC_12_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__21952\,
            in1 => \N__21340\,
            in2 => \N__20855\,
            in3 => \N__22772\,
            lcout => OPEN,
            ltout => \eeprom.n26_adj_466_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i13_4_lut_LC_12_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__23222\,
            in1 => \N__21370\,
            in2 => \N__20852\,
            in3 => \N__21413\,
            lcout => \eeprom.n3133\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i1_2_lut_adj_44_LC_12_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__21615\,
            in3 => \N__20917\,
            lcout => OPEN,
            ltout => \eeprom.n4711_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i1_4_lut_adj_45_LC_12_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__21390\,
            in1 => \N__21510\,
            in2 => \N__20849\,
            in3 => \N__20974\,
            lcout => \eeprom.n4715\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2098_3_lut_LC_12_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21032\,
            in2 => \N__24185\,
            in3 => \N__21762\,
            lcout => \eeprom.n3206\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2106_3_lut_LC_12_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20948\,
            in2 => \N__21616\,
            in3 => \N__21761\,
            lcout => \eeprom.n3214\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2089_2_lut_LC_12_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20763\,
            in2 => \_gnd_net_\,
            in3 => \N__20711\,
            lcout => \eeprom.n3186\,
            ltout => OPEN,
            carryin => \bfn_12_22_0_\,
            carryout => \eeprom.n3667\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2089_3_lut_LC_12_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27311\,
            in2 => \N__21453\,
            in3 => \N__20696\,
            lcout => \eeprom.n3185\,
            ltout => OPEN,
            carryin => \eeprom.n3667\,
            carryout => \eeprom.n3668\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2089_4_lut_LC_12_22_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__21392\,
            in3 => \N__20981\,
            lcout => \eeprom.n3184\,
            ltout => OPEN,
            carryin => \eeprom.n3668\,
            carryout => \eeprom.n3669\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2089_5_lut_LC_12_22_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__20978\,
            in3 => \N__20951\,
            lcout => \eeprom.n3183\,
            ltout => OPEN,
            carryin => \eeprom.n3669\,
            carryout => \eeprom.n3670\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2089_6_lut_LC_12_22_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__21617\,
            in3 => \N__20942\,
            lcout => \eeprom.n3182\,
            ltout => OPEN,
            carryin => \eeprom.n3670\,
            carryout => \eeprom.n3671\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2089_7_lut_LC_12_22_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__21517\,
            in3 => \N__20927\,
            lcout => \eeprom.n3181\,
            ltout => OPEN,
            carryin => \eeprom.n3671\,
            carryout => \eeprom.n3672\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2089_8_lut_LC_12_22_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__20924\,
            in3 => \N__20894\,
            lcout => \eeprom.n3180\,
            ltout => OPEN,
            carryin => \eeprom.n3672\,
            carryout => \eeprom.n3673\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2089_9_lut_LC_12_22_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23220\,
            in2 => \N__27542\,
            in3 => \N__20891\,
            lcout => \eeprom.n3179\,
            ltout => OPEN,
            carryin => \eeprom.n3673\,
            carryout => \eeprom.n3674\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2089_10_lut_LC_12_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27080\,
            in2 => \N__24284\,
            in3 => \N__20876\,
            lcout => \eeprom.n3178\,
            ltout => OPEN,
            carryin => \bfn_12_23_0_\,
            carryout => \eeprom.n3675\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2089_11_lut_LC_12_23_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24208\,
            in2 => \N__27302\,
            in3 => \N__20858\,
            lcout => \eeprom.n3177\,
            ltout => OPEN,
            carryin => \eeprom.n3675\,
            carryout => \eeprom.n3676\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2089_12_lut_LC_12_23_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27084\,
            in2 => \N__24244\,
            in3 => \N__21038\,
            lcout => \eeprom.n3176\,
            ltout => OPEN,
            carryin => \eeprom.n3676\,
            carryout => \eeprom.n3677\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2089_13_lut_LC_12_23_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21371\,
            in2 => \N__27303\,
            in3 => \N__21035\,
            lcout => \eeprom.n3175\,
            ltout => OPEN,
            carryin => \eeprom.n3677\,
            carryout => \eeprom.n3678\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2089_14_lut_LC_12_23_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24178\,
            in2 => \N__27306\,
            in3 => \N__21023\,
            lcout => \eeprom.n3174\,
            ltout => OPEN,
            carryin => \eeprom.n3678\,
            carryout => \eeprom.n3679\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2089_15_lut_LC_12_23_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21817\,
            in2 => \N__27304\,
            in3 => \N__21020\,
            lcout => \eeprom.n3173\,
            ltout => OPEN,
            carryin => \eeprom.n3679\,
            carryout => \eeprom.n3680\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2089_16_lut_LC_12_23_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27091\,
            in2 => \N__21344\,
            in3 => \N__21017\,
            lcout => \eeprom.n3172\,
            ltout => OPEN,
            carryin => \eeprom.n3680\,
            carryout => \eeprom.n3681\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2089_17_lut_LC_12_23_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21951\,
            in2 => \N__27305\,
            in3 => \N__21005\,
            lcout => \eeprom.n3171\,
            ltout => OPEN,
            carryin => \eeprom.n3681\,
            carryout => \eeprom.n3682\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2089_18_lut_LC_12_24_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23144\,
            in2 => \N__27384\,
            in3 => \N__21002\,
            lcout => \eeprom.n3170\,
            ltout => OPEN,
            carryin => \bfn_12_24_0_\,
            carryout => \eeprom.n3683\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2089_19_lut_LC_12_24_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21427\,
            in2 => \N__27386\,
            in3 => \N__20999\,
            lcout => \eeprom.n3169\,
            ltout => OPEN,
            carryin => \eeprom.n3683\,
            carryout => \eeprom.n3684\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2089_20_lut_LC_12_24_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22042\,
            in2 => \N__27385\,
            in3 => \N__20996\,
            lcout => \eeprom.n3168\,
            ltout => OPEN,
            carryin => \eeprom.n3684\,
            carryout => \eeprom.n3685\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2089_21_lut_LC_12_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001000001100000"
        )
    port map (
            in0 => \N__27205\,
            in1 => \N__27806\,
            in2 => \N__21792\,
            in3 => \N__21125\,
            lcout => \eeprom.n3199\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1959_3_lut_LC_12_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21122\,
            in2 => \N__21113\,
            in3 => \N__24753\,
            lcout => \eeprom.n3003\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1965_3_lut_LC_12_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__21089\,
            in1 => \_gnd_net_\,
            in2 => \N__24764\,
            in3 => \N__21076\,
            lcout => \eeprom.n3009\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2309_3_lut_LC_13_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21976\,
            in2 => \N__23363\,
            in3 => \N__21962\,
            lcout => \eeprom.n3513_adj_366\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2310_3_lut_LC_13_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__21986\,
            in1 => \_gnd_net_\,
            in2 => \N__22012\,
            in3 => \N__23324\,
            lcout => \eeprom.n3514_adj_368\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2308_3_lut_LC_13_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22385\,
            in2 => \N__22406\,
            in3 => \N__23331\,
            lcout => \eeprom.n3512_adj_364\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2294_3_lut_LC_13_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22489\,
            in2 => \N__23364\,
            in3 => \N__22457\,
            lcout => \eeprom.n3498\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2293_3_lut_LC_13_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22445\,
            in2 => \N__22418\,
            in3 => \N__23332\,
            lcout => \eeprom.n3497\,
            ltout => \eeprom.n3497_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i10_4_lut_adj_110_LC_13_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__25723\,
            in1 => \N__25240\,
            in2 => \N__21056\,
            in3 => \N__25186\,
            lcout => OPEN,
            ltout => \eeprom.n28_adj_493_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i14_3_lut_LC_13_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24946\,
            in2 => \N__21170\,
            in3 => \N__25113\,
            lcout => \eeprom.n32_adj_494\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i4039_3_lut_LC_13_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22240\,
            in2 => \N__22214\,
            in3 => \N__23352\,
            lcout => \eeprom.n3507\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2300_3_lut_LC_13_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22684\,
            in2 => \N__23371\,
            in3 => \N__22661\,
            lcout => \eeprom.n3504\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2306_3_lut_LC_13_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22339\,
            in2 => \N__22316\,
            in3 => \N__23348\,
            lcout => \eeprom.n3510_adj_360\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i1_2_lut_adj_102_LC_13_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__22443\,
            in3 => \N__22732\,
            lcout => OPEN,
            ltout => \eeprom.n18_adj_488_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i13_4_lut_adj_106_LC_13_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__22338\,
            in1 => \N__22369\,
            in2 => \N__21167\,
            in3 => \N__22269\,
            lcout => OPEN,
            ltout => \eeprom.n30_adj_489_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i16_4_lut_LC_13_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__21164\,
            in1 => \N__21155\,
            in2 => \N__21149\,
            in3 => \N__21146\,
            lcout => \eeprom.n3430\,
            ltout => \eeprom.n3430_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2304_3_lut_LC_13_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22270\,
            in2 => \N__21137\,
            in3 => \N__22253\,
            lcout => \eeprom.n3508\,
            ltout => \eeprom.n3508_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i1_4_lut_adj_52_LC_13_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011111010"
        )
    port map (
            in0 => \N__21134\,
            in1 => \N__24935\,
            in2 => \N__21128\,
            in3 => \N__25660\,
            lcout => \eeprom.n4429\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2298_3_lut_LC_13_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22619\,
            in2 => \N__23370\,
            in3 => \N__22645\,
            lcout => \eeprom.n3502\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i12_4_lut_adj_116_LC_13_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__25425\,
            in1 => \N__25071\,
            in2 => \N__24922\,
            in3 => \N__23126\,
            lcout => OPEN,
            ltout => \eeprom.n30_adj_495_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i17_4_lut_LC_13_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__21233\,
            in1 => \N__21227\,
            in2 => \N__21221\,
            in3 => \N__21218\,
            lcout => \eeprom.n3529_adj_336\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2295_3_lut_LC_13_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22528\,
            in2 => \N__22502\,
            in3 => \N__23341\,
            lcout => \eeprom.n3499\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2370_3_lut_LC_13_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24918\,
            in2 => \N__24902\,
            in3 => \N__25680\,
            lcout => OPEN,
            ltout => \eeprom.n3606_adj_446_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i1_4_lut_adj_51_LC_13_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110111111000"
        )
    port map (
            in0 => \N__25681\,
            in1 => \N__25409\,
            in2 => \N__21209\,
            in3 => \N__25429\,
            lcout => OPEN,
            ltout => \eeprom.n4451_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i1_4_lut_adj_53_LC_13_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111100"
        )
    port map (
            in0 => \N__25361\,
            in1 => \N__25394\,
            in2 => \N__21206\,
            in3 => \N__25682\,
            lcout => \eeprom.n4453\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2363_3_lut_LC_13_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25256\,
            in2 => \N__25276\,
            in3 => \N__25632\,
            lcout => OPEN,
            ltout => \eeprom.n3599_adj_450_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i1_4_lut_adj_57_LC_13_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__21404\,
            in1 => \N__21203\,
            in2 => \N__21197\,
            in3 => \N__21194\,
            lcout => \eeprom.n4433\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_mux_3_i5_3_lut_LC_13_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001001110111"
        )
    port map (
            in0 => \N__22977\,
            in1 => \N__21185\,
            in2 => \_gnd_net_\,
            in3 => \N__23722\,
            lcout => \eeprom.n3721_adj_434\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2364_3_lut_LC_13_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25292\,
            in2 => \N__25672\,
            in3 => \N__25312\,
            lcout => \eeprom.n3600_adj_449\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2377_3_lut_LC_13_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24487\,
            in2 => \N__24461\,
            in3 => \N__25628\,
            lcout => \eeprom.n3613_adj_342\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i1_4_lut_adj_55_LC_13_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011101110"
        )
    port map (
            in0 => \N__21398\,
            in1 => \N__25123\,
            in2 => \N__25097\,
            in3 => \N__25633\,
            lcout => \eeprom.n4583\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2041_3_lut_LC_13_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26312\,
            in2 => \N__27915\,
            in3 => \N__26339\,
            lcout => \eeprom.n3117\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2032_3_lut_LC_13_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26594\,
            in2 => \N__26561\,
            in3 => \N__27902\,
            lcout => \eeprom.n3108\,
            ltout => \eeprom.n3108_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2099_3_lut_LC_13_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21356\,
            in2 => \N__21347\,
            in3 => \N__21764\,
            lcout => \eeprom.n3207\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2029_3_lut_LC_13_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26468\,
            in2 => \N__26444\,
            in3 => \N__27903\,
            lcout => \eeprom.n3105\,
            ltout => \eeprom.n3105_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2096_3_lut_LC_13_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21326\,
            in2 => \N__21314\,
            in3 => \N__21763\,
            lcout => \eeprom.n3204\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2103_3_lut_LC_13_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23221\,
            in2 => \N__21278\,
            in3 => \N__21765\,
            lcout => \eeprom.n3211\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2039_3_lut_LC_13_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27874\,
            in2 => \N__26213\,
            in3 => \N__26245\,
            lcout => \eeprom.n3115\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2093_3_lut_LC_13_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__21593\,
            in1 => \N__21428\,
            in2 => \_gnd_net_\,
            in3 => \N__21776\,
            lcout => \eeprom.n3201\,
            ltout => \eeprom.n3201_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i9_4_lut_adj_93_LC_13_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__21876\,
            in1 => \N__21552\,
            in2 => \N__21536\,
            in3 => \N__21912\,
            lcout => \eeprom.n24_adj_481\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2038_3_lut_LC_13_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__26165\,
            in1 => \_gnd_net_\,
            in2 => \N__27908\,
            in3 => \N__26191\,
            lcout => \eeprom.n3114\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1960_3_lut_LC_13_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21494\,
            in2 => \N__21470\,
            in3 => \N__24763\,
            lcout => \eeprom.n3004\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2042_3_lut_LC_13_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26354\,
            in2 => \N__27907\,
            in3 => \N__26390\,
            lcout => \eeprom.n3118\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i8_4_lut_adj_42_LC_13_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__26418\,
            in1 => \N__26460\,
            in2 => \N__28030\,
            in3 => \N__28062\,
            lcout => \eeprom.n21_adj_422\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2026_3_lut_LC_13_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28026\,
            in2 => \N__27910\,
            in3 => \N__28010\,
            lcout => \eeprom.n3102\,
            ltout => \eeprom.n3102_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i8_4_lut_adj_67_LC_13_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__27805\,
            in1 => \N__23139\,
            in2 => \N__21416\,
            in3 => \N__22038\,
            lcout => \eeprom.n22_adj_465\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2028_3_lut_LC_13_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__26419\,
            in1 => \_gnd_net_\,
            in2 => \N__28091\,
            in3 => \N__27890\,
            lcout => \eeprom.n3104\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i7_3_lut_LC_13_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111010"
        )
    port map (
            in0 => \N__26703\,
            in1 => \_gnd_net_\,
            in2 => \N__27943\,
            in3 => \N__27987\,
            lcout => \eeprom.n20_adj_423\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2094_3_lut_LC_13_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21932\,
            in2 => \N__21794\,
            in3 => \N__23140\,
            lcout => \eeprom.n3202\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2092_3_lut_LC_13_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21896\,
            in2 => \N__22043\,
            in3 => \N__21784\,
            lcout => \eeprom.n3200\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1971_3_lut_LC_13_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21860\,
            in2 => \N__21848\,
            in3 => \N__24737\,
            lcout => \eeprom.n3015\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2030_3_lut_LC_13_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__27889\,
            in1 => \_gnd_net_\,
            in2 => \N__26483\,
            in3 => \N__26512\,
            lcout => \eeprom.n3106\,
            ltout => \eeprom.n3106_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2097_3_lut_LC_13_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21803\,
            in2 => \N__21797\,
            in3 => \N__21788\,
            lcout => \eeprom.n3205\,
            ltout => \eeprom.n3205_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i1_2_lut_adj_92_LC_13_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__21653\,
            in3 => \N__21643\,
            lcout => \eeprom.n16_adj_479\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1962_3_lut_LC_13_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22127\,
            in2 => \N__22100\,
            in3 => \N__24741\,
            lcout => \eeprom.n3006\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1969_3_lut_LC_13_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22085\,
            in2 => \N__24759\,
            in3 => \N__22055\,
            lcout => \eeprom.n3013\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2025_3_lut_LC_13_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27994\,
            in2 => \N__27965\,
            in3 => \N__27888\,
            lcout => \eeprom.n3101\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2290_2_lut_LC_14_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23425\,
            in2 => \_gnd_net_\,
            in3 => \N__22025\,
            lcout => \eeprom.n3486\,
            ltout => OPEN,
            carryin => \bfn_14_17_0_\,
            carryout => \eeprom.n3727\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2290_3_lut_LC_14_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27781\,
            in2 => \N__23078\,
            in3 => \N__22022\,
            lcout => \eeprom.n3485\,
            ltout => OPEN,
            carryin => \eeprom.n3727\,
            carryout => \eeprom.n3728\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2290_4_lut_LC_14_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__23113\,
            in3 => \N__22019\,
            lcout => \eeprom.n3484_adj_406\,
            ltout => OPEN,
            carryin => \eeprom.n3728\,
            carryout => \eeprom.n3729\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2290_5_lut_LC_14_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__23036\,
            in3 => \N__22016\,
            lcout => \eeprom.n3483_adj_404\,
            ltout => OPEN,
            carryin => \eeprom.n3729\,
            carryout => \eeprom.n3730\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2290_6_lut_LC_14_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__22013\,
            in3 => \N__21980\,
            lcout => \eeprom.n3482_adj_401\,
            ltout => OPEN,
            carryin => \eeprom.n3730\,
            carryout => \eeprom.n3731\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2290_7_lut_LC_14_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21977\,
            in2 => \_gnd_net_\,
            in3 => \N__21956\,
            lcout => \eeprom.n3481_adj_399\,
            ltout => OPEN,
            carryin => \eeprom.n3731\,
            carryout => \eeprom.n3732\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2290_8_lut_LC_14_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__22405\,
            in3 => \N__22379\,
            lcout => \eeprom.n3480_adj_398\,
            ltout => OPEN,
            carryin => \eeprom.n3732\,
            carryout => \eeprom.n3733\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2290_9_lut_LC_14_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27782\,
            in2 => \N__22376\,
            in3 => \N__22343\,
            lcout => \eeprom.n3479_adj_394\,
            ltout => OPEN,
            carryin => \eeprom.n3733\,
            carryout => \eeprom.n3734\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2290_10_lut_LC_14_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27708\,
            in2 => \N__22340\,
            in3 => \N__22307\,
            lcout => \eeprom.n3478_adj_393\,
            ltout => OPEN,
            carryin => \bfn_14_18_0_\,
            carryout => \eeprom.n3735\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2290_11_lut_LC_14_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27712\,
            in2 => \N__22304\,
            in3 => \N__22277\,
            lcout => \eeprom.n3477_adj_392\,
            ltout => OPEN,
            carryin => \eeprom.n3735\,
            carryout => \eeprom.n3736\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2290_12_lut_LC_14_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27709\,
            in2 => \N__22274\,
            in3 => \N__22244\,
            lcout => \eeprom.n3476_adj_391\,
            ltout => OPEN,
            carryin => \eeprom.n3736\,
            carryout => \eeprom.n3737\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2290_13_lut_LC_14_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27713\,
            in2 => \N__22241\,
            in3 => \N__22202\,
            lcout => \eeprom.n3475_adj_390\,
            ltout => OPEN,
            carryin => \eeprom.n3737\,
            carryout => \eeprom.n3738\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2290_14_lut_LC_14_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27710\,
            in2 => \N__22199\,
            in3 => \N__22169\,
            lcout => \eeprom.n3474_adj_389\,
            ltout => OPEN,
            carryin => \eeprom.n3738\,
            carryout => \eeprom.n3739\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2290_15_lut_LC_14_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27714\,
            in2 => \N__22166\,
            in3 => \N__22130\,
            lcout => \eeprom.n3473_adj_388\,
            ltout => OPEN,
            carryin => \eeprom.n3739\,
            carryout => \eeprom.n3740\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2290_16_lut_LC_14_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27711\,
            in2 => \N__22685\,
            in3 => \N__22652\,
            lcout => \eeprom.n3472_adj_387\,
            ltout => OPEN,
            carryin => \eeprom.n3740\,
            carryout => \eeprom.n3741\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2290_17_lut_LC_14_18_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27715\,
            in2 => \N__23255\,
            in3 => \N__22649\,
            lcout => \eeprom.n3471_adj_386\,
            ltout => OPEN,
            carryin => \eeprom.n3741\,
            carryout => \eeprom.n3742\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2290_18_lut_LC_14_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27509\,
            in2 => \N__22646\,
            in3 => \N__22613\,
            lcout => \eeprom.n3470_adj_385\,
            ltout => OPEN,
            carryin => \bfn_14_19_0_\,
            carryout => \eeprom.n3743\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2290_19_lut_LC_14_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22610\,
            in2 => \N__27706\,
            in3 => \N__22577\,
            lcout => \eeprom.n3469_adj_384\,
            ltout => OPEN,
            carryin => \eeprom.n3743\,
            carryout => \eeprom.n3744\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2290_20_lut_LC_14_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27513\,
            in2 => \N__22574\,
            in3 => \N__22532\,
            lcout => \eeprom.n3468_adj_383\,
            ltout => OPEN,
            carryin => \eeprom.n3744\,
            carryout => \eeprom.n3745\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2290_21_lut_LC_14_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27518\,
            in2 => \N__22529\,
            in3 => \N__22493\,
            lcout => \eeprom.n3467_adj_382\,
            ltout => OPEN,
            carryin => \eeprom.n3745\,
            carryout => \eeprom.n3746\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2290_22_lut_LC_14_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27514\,
            in2 => \N__22490\,
            in3 => \N__22448\,
            lcout => \eeprom.n3466_adj_381\,
            ltout => OPEN,
            carryin => \eeprom.n3746\,
            carryout => \eeprom.n3747\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2290_23_lut_LC_14_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22444\,
            in2 => \N__27707\,
            in3 => \N__22736\,
            lcout => \eeprom.n3465_adj_380\,
            ltout => OPEN,
            carryin => \eeprom.n3747\,
            carryout => \eeprom.n3748\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2290_24_lut_LC_14_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001000001100000"
        )
    port map (
            in0 => \N__27519\,
            in1 => \N__22733\,
            in2 => \N__23369\,
            in3 => \N__22712\,
            lcout => \eeprom.n3496\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i1_2_lut_adj_58_LC_14_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__26056\,
            in3 => \N__25525\,
            lcout => \eeprom.n4619\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i1_4_lut_adj_56_LC_14_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111100"
        )
    port map (
            in0 => \N__25445\,
            in1 => \N__25466\,
            in2 => \N__22709\,
            in3 => \N__25663\,
            lcout => OPEN,
            ltout => \eeprom.n31_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i1_4_lut_adj_62_LC_14_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__26014\,
            in1 => \N__22691\,
            in2 => \N__22700\,
            in3 => \N__22697\,
            lcout => \eeprom.n4567\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2445_3_lut_LC_14_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000000111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25478\,
            in2 => \N__25832\,
            in3 => \N__25502\,
            lcout => \eeprom.n3713_adj_443\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2362_3_lut_LC_14_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__25662\,
            in1 => \_gnd_net_\,
            in2 => \N__25217\,
            in3 => \N__25239\,
            lcout => \eeprom.n3598_adj_452\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2376_3_lut_LC_14_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25139\,
            in2 => \N__25175\,
            in3 => \N__25661\,
            lcout => \eeprom.n3612_adj_339\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2444_3_lut_LC_14_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26055\,
            in2 => \N__26033\,
            in3 => \N__25817\,
            lcout => \eeprom.n3712_adj_444\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2360_3_lut_LC_14_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__25664\,
            in1 => \_gnd_net_\,
            in2 => \N__25766\,
            in3 => \N__25739\,
            lcout => \eeprom.n3596_adj_454\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_mux_3_i3_3_lut_LC_14_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101010101"
        )
    port map (
            in0 => \N__23845\,
            in1 => \N__23003\,
            in2 => \_gnd_net_\,
            in3 => \N__22991\,
            lcout => \eeprom.n3723_adj_334\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i4077_1_lut_LC_14_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24091\,
            lcout => \eeprom.n4921\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i4080_1_lut_2_lut_LC_14_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25952\,
            in2 => \_gnd_net_\,
            in3 => \N__25833\,
            lcout => \eeprom.n4924\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i10_4_lut_adj_66_LC_14_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__24201\,
            in1 => \N__24231\,
            in2 => \N__24273\,
            in3 => \N__24171\,
            lcout => \eeprom.n24_adj_459\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i1_2_lut_adj_39_LC_14_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__26092\,
            in3 => \N__26184\,
            lcout => OPEN,
            ltout => \eeprom.n4559_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i1_4_lut_adj_40_LC_14_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__26244\,
            in1 => \N__26145\,
            in2 => \N__22760\,
            in3 => \N__26293\,
            lcout => OPEN,
            ltout => \eeprom.n4563_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i4_4_lut_adj_41_LC_14_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011101010"
        )
    port map (
            in0 => \N__26513\,
            in1 => \N__26385\,
            in2 => \N__22757\,
            in3 => \N__26331\,
            lcout => OPEN,
            ltout => \eeprom.n17_adj_421_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i11_4_lut_adj_43_LC_14_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__22754\,
            in1 => \N__26539\,
            in2 => \N__22748\,
            in3 => \N__26593\,
            lcout => OPEN,
            ltout => \eeprom.n24_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i12_4_lut_LC_14_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__26667\,
            in1 => \N__26635\,
            in2 => \N__22745\,
            in3 => \N__22742\,
            lcout => \eeprom.n3034\,
            ltout => \eeprom.n3034_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2036_3_lut_LC_14_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26088\,
            in2 => \N__23225\,
            in3 => \N__26069\,
            lcout => \eeprom.n3112\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1967_3_lut_LC_14_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23189\,
            in2 => \N__23159\,
            in3 => \N__24762\,
            lcout => \eeprom.n3011\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2027_3_lut_LC_14_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28072\,
            in2 => \N__28049\,
            in3 => \N__27887\,
            lcout => \eeprom.n3103\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i1_4_lut_adj_115_LC_15_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000000000000"
        )
    port map (
            in0 => \N__24600\,
            in1 => \N__24658\,
            in2 => \N__23435\,
            in3 => \N__23042\,
            lcout => \eeprom.n4137\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2312_3_lut_LC_15_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23114\,
            in2 => \N__23087\,
            in3 => \N__23372\,
            lcout => \eeprom.n3516_adj_372\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2380_3_lut_LC_15_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__24560\,
            in1 => \_gnd_net_\,
            in2 => \N__25705\,
            in3 => \N__24574\,
            lcout => \eeprom.n3616_adj_345\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2313_3_lut_LC_15_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23077\,
            in2 => \N__23054\,
            in3 => \N__23374\,
            lcout => \eeprom.n3517_adj_374\,
            ltout => \eeprom.n3517_adj_374_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i1_3_lut_adj_114_LC_15_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24483\,
            in2 => \N__23045\,
            in3 => \N__24543\,
            lcout => \eeprom.n4729\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2311_3_lut_LC_15_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23035\,
            in2 => \N__23012\,
            in3 => \N__23373\,
            lcout => \eeprom.n3515_adj_370\,
            ltout => \eeprom.n3515_adj_370_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i1_2_lut_adj_111_LC_15_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__23438\,
            in3 => \N__25161\,
            lcout => \eeprom.n4727\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2378_3_lut_LC_15_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24517\,
            in2 => \N__24503\,
            in3 => \N__25696\,
            lcout => \eeprom.n3614_adj_343\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2314_3_lut_LC_15_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__23426\,
            in1 => \N__23387\,
            in2 => \_gnd_net_\,
            in3 => \N__23365\,
            lcout => \eeprom.n3518_adj_376\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2299_3_lut_LC_15_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23381\,
            in2 => \N__23375\,
            in3 => \N__23254\,
            lcout => \eeprom.n3503\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2369_3_lut_LC_15_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24857\,
            in2 => \N__25704\,
            in3 => \N__24884\,
            lcout => \eeprom.n3605_adj_453\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2379_3_lut_LC_15_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24527\,
            in2 => \N__24551\,
            in3 => \N__25689\,
            lcout => \eeprom.n3615_adj_344\,
            ltout => \eeprom.n3615_adj_344_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2446_3_lut_LC_15_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25514\,
            in2 => \N__23231\,
            in3 => \N__25816\,
            lcout => \eeprom.n3714_adj_442\,
            ltout => \eeprom.n3714_adj_442_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i4071_1_lut_LC_15_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__23228\,
            in3 => \_gnd_net_\,
            lcout => \eeprom.n4915\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2381_3_lut_LC_15_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__24584\,
            in1 => \_gnd_net_\,
            in2 => \N__25703\,
            in3 => \N__24604\,
            lcout => \eeprom.n3617_adj_346\,
            ltout => \eeprom.n3617_adj_346_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i1_4_lut_adj_59_LC_15_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__25494\,
            in1 => \N__25980\,
            in2 => \N__23555\,
            in3 => \N__23552\,
            lcout => \eeprom.n4623\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i1_4_lut_adj_61_LC_15_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111100010"
        )
    port map (
            in0 => \N__25349\,
            in1 => \N__25684\,
            in2 => \N__25328\,
            in3 => \N__23507\,
            lcout => OPEN,
            ltout => \eeprom.n4427_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i1_4_lut_adj_63_LC_15_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110111111000"
        )
    port map (
            in0 => \N__25685\,
            in1 => \N__25775\,
            in2 => \N__23546\,
            in3 => \N__25199\,
            lcout => OPEN,
            ltout => \eeprom.n28_adj_455_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i1_4_lut_adj_64_LC_15_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__25571\,
            in1 => \N__23543\,
            in2 => \N__23537\,
            in3 => \N__23534\,
            lcout => \eeprom.n3628_adj_437\,
            ltout => \eeprom.n3628_adj_437_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2448_3_lut_LC_15_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000000111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25544\,
            in2 => \N__23528\,
            in3 => \N__25558\,
            lcout => \eeprom.n3716_adj_439\,
            ltout => \eeprom.n3716_adj_439_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i4065_1_lut_LC_15_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__23525\,
            in3 => \_gnd_net_\,
            lcout => \eeprom.n4909\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2382_3_lut_LC_15_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__24620\,
            in1 => \N__24654\,
            in2 => \_gnd_net_\,
            in3 => \N__25683\,
            lcout => \eeprom.n3618_adj_350\,
            ltout => \eeprom.n3618_adj_350_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i1_4_lut_adj_60_LC_15_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011001100"
        )
    port map (
            in0 => \N__25876\,
            in1 => \N__23522\,
            in2 => \N__23516\,
            in3 => \N__23513\,
            lcout => \eeprom.n4425\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2473_2_lut_LC_15_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101110111000"
        )
    port map (
            in0 => \N__23501\,
            in1 => \N__24062\,
            in2 => \N__23459\,
            in3 => \N__23441\,
            lcout => \eeprom.number_of_bytes_7_N_68_0\,
            ltout => OPEN,
            carryin => \bfn_15_20_0_\,
            carryout => \eeprom.n3772\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2473_3_lut_LC_15_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__23912\,
            in1 => \N__23867\,
            in2 => \N__24075\,
            in3 => \N__23855\,
            lcout => \eeprom.number_of_bytes_7_N_68_1\,
            ltout => OPEN,
            carryin => \eeprom.n3772\,
            carryout => \eeprom.n3773\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2473_4_lut_LC_15_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101110111000"
        )
    port map (
            in0 => \N__23852\,
            in1 => \N__24066\,
            in2 => \N__23804\,
            in3 => \N__23792\,
            lcout => \eeprom.number_of_bytes_7_N_68_2\,
            ltout => OPEN,
            carryin => \eeprom.n3773\,
            carryout => \eeprom.n3774\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2473_5_lut_LC_15_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__23789\,
            in1 => \N__23747\,
            in2 => \N__24076\,
            in3 => \N__23729\,
            lcout => \eeprom.number_of_bytes_7_N_68_3\,
            ltout => OPEN,
            carryin => \eeprom.n3774\,
            carryout => \eeprom.n3775\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2473_6_lut_LC_15_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101110111000"
        )
    port map (
            in0 => \N__23726\,
            in1 => \N__24070\,
            in2 => \N__23687\,
            in3 => \N__23675\,
            lcout => \eeprom.number_of_bytes_7_N_68_4\,
            ltout => OPEN,
            carryin => \eeprom.n3775\,
            carryout => \eeprom.n3776\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2473_7_lut_LC_15_20_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__23672\,
            in1 => \N__23630\,
            in2 => \N__24077\,
            in3 => \N__23621\,
            lcout => \eeprom.number_of_bytes_7_N_68_5\,
            ltout => OPEN,
            carryin => \eeprom.n3776\,
            carryout => \eeprom.n3777\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2473_8_lut_LC_15_20_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101110111000"
        )
    port map (
            in0 => \N__23618\,
            in1 => \N__24074\,
            in2 => \N__23579\,
            in3 => \N__23564\,
            lcout => \eeprom.number_of_bytes_7_N_68_6\,
            ltout => OPEN,
            carryin => \eeprom.n3777\,
            carryout => \eeprom.n3778\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2473_9_lut_LC_15_20_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101110111000"
        )
    port map (
            in0 => \N__26396\,
            in1 => \N__24059\,
            in2 => \N__25784\,
            in3 => \N__23561\,
            lcout => \eeprom.number_of_bytes_7_N_68_7\,
            ltout => OPEN,
            carryin => \eeprom.n3778\,
            carryout => \eeprom.n3779\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2473_10_lut_LC_15_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101110111000"
        )
    port map (
            in0 => \N__25889\,
            in1 => \N__24043\,
            in2 => \N__25901\,
            in3 => \N__23558\,
            lcout => \eeprom.number_of_bytes_7_N_68_8\,
            ltout => OPEN,
            carryin => \bfn_15_21_0_\,
            carryout => \eeprom.n3780\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2473_11_lut_LC_15_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101110111000"
        )
    port map (
            in0 => \N__24155\,
            in1 => \N__24033\,
            in2 => \N__24146\,
            in3 => \N__24134\,
            lcout => \eeprom.number_of_bytes_7_N_68_9\,
            ltout => OPEN,
            carryin => \eeprom.n3780\,
            carryout => \eeprom.n3781\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2473_12_lut_LC_15_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__25958\,
            in1 => \N__25967\,
            in2 => \N__24060\,
            in3 => \N__24131\,
            lcout => \eeprom.number_of_bytes_7_N_68_10\,
            ltout => OPEN,
            carryin => \eeprom.n3781\,
            carryout => \eeprom.n3782\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2473_13_lut_LC_15_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101110111000"
        )
    port map (
            in0 => \N__24128\,
            in1 => \N__24037\,
            in2 => \N__24119\,
            in3 => \N__24107\,
            lcout => \eeprom.number_of_bytes_7_N_68_11\,
            ltout => OPEN,
            carryin => \eeprom.n3782\,
            carryout => \eeprom.n3783\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2473_14_lut_LC_15_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__23948\,
            in1 => \N__23959\,
            in2 => \N__24061\,
            in3 => \N__24104\,
            lcout => \eeprom.number_of_bytes_7_N_68_12\,
            ltout => OPEN,
            carryin => \eeprom.n3783\,
            carryout => \eeprom.n3784\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2473_15_lut_LC_15_21_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101110111000"
        )
    port map (
            in0 => \N__24101\,
            in1 => \N__24041\,
            in2 => \N__24095\,
            in3 => \N__24080\,
            lcout => \eeprom.number_of_bytes_7_N_68_13\,
            ltout => OPEN,
            carryin => \eeprom.n3784\,
            carryout => \eeprom.n3785\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2473_16_lut_LC_15_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000110111011000"
        )
    port map (
            in0 => \N__24042\,
            in1 => \N__23969\,
            in2 => \N__25934\,
            in3 => \N__23963\,
            lcout => \eeprom.number_of_bytes_7_N_68_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i4074_1_lut_LC_15_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__23960\,
            in3 => \_gnd_net_\,
            lcout => \eeprom.n4918\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i1_4_lut_adj_113_LC_15_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__23942\,
            in1 => \N__23933\,
            in2 => \N__23924\,
            in3 => \N__24290\,
            lcout => OPEN,
            ltout => \eeprom.n4301_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i1_4_lut_adj_119_LC_15_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__24443\,
            in1 => \N__24434\,
            in2 => \N__24428\,
            in3 => \N__24425\,
            lcout => OPEN,
            ltout => \eeprom.n4307_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i1_4_lut_adj_120_LC_15_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__24416\,
            in1 => \N__24410\,
            in2 => \N__24404\,
            in3 => \N__24401\,
            lcout => OPEN,
            ltout => \eeprom.n4313_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.ena_12_LC_15_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__24395\,
            in1 => \N__24389\,
            in2 => \N__24383\,
            in3 => \N__24380\,
            lcout => sda_enable,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24349\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i1_3_lut_adj_112_LC_15_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__24317\,
            in1 => \N__24308\,
            in2 => \_gnd_net_\,
            in3 => \N__24299\,
            lcout => \eeprom.n4295\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2035_3_lut_LC_15_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26681\,
            in2 => \N__27909\,
            in3 => \N__26704\,
            lcout => \eeprom.n3111\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2033_3_lut_LC_15_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26639\,
            in2 => \N__26606\,
            in3 => \N__27882\,
            lcout => \eeprom.n3109\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2034_3_lut_LC_15_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26671\,
            in2 => \N__26651\,
            in3 => \N__27881\,
            lcout => \eeprom.n3110\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2031_3_lut_LC_15_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__26522\,
            in1 => \_gnd_net_\,
            in2 => \N__26543\,
            in3 => \N__27886\,
            lcout => \eeprom.n3107\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1974_3_lut_LC_15_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__24848\,
            in1 => \N__24836\,
            in2 => \_gnd_net_\,
            in3 => \N__24760\,
            lcout => \eeprom.n3018\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1964_3_lut_LC_15_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__24796\,
            in1 => \N__24776\,
            in2 => \_gnd_net_\,
            in3 => \N__24761\,
            lcout => \eeprom.n3008\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2357_2_lut_LC_16_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24659\,
            in2 => \_gnd_net_\,
            in3 => \N__24608\,
            lcout => \eeprom.n3586_adj_378\,
            ltout => OPEN,
            carryin => \bfn_16_17_0_\,
            carryout => \eeprom.n3749\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2357_3_lut_LC_16_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27024\,
            in2 => \N__24605\,
            in3 => \N__24578\,
            lcout => \eeprom.n3585_adj_375\,
            ltout => OPEN,
            carryin => \eeprom.n3749\,
            carryout => \eeprom.n3750\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2357_4_lut_LC_16_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__24575\,
            in3 => \N__24554\,
            lcout => \eeprom.n3584_adj_373\,
            ltout => OPEN,
            carryin => \eeprom.n3750\,
            carryout => \eeprom.n3751\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2357_5_lut_LC_16_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__24550\,
            in3 => \N__24521\,
            lcout => \eeprom.n3583_adj_371\,
            ltout => OPEN,
            carryin => \eeprom.n3751\,
            carryout => \eeprom.n3752\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2357_6_lut_LC_16_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__24518\,
            in3 => \N__24494\,
            lcout => \eeprom.n3582_adj_369\,
            ltout => OPEN,
            carryin => \eeprom.n3752\,
            carryout => \eeprom.n3753\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2357_7_lut_LC_16_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__24491\,
            in3 => \N__24446\,
            lcout => \eeprom.n3581_adj_367\,
            ltout => OPEN,
            carryin => \eeprom.n3753\,
            carryout => \eeprom.n3754\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2357_8_lut_LC_16_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__25174\,
            in3 => \N__25127\,
            lcout => \eeprom.n3580_adj_365\,
            ltout => OPEN,
            carryin => \eeprom.n3754\,
            carryout => \eeprom.n3755\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2357_9_lut_LC_16_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27025\,
            in2 => \N__25124\,
            in3 => \N__25082\,
            lcout => \eeprom.n3579_adj_363\,
            ltout => OPEN,
            carryin => \eeprom.n3755\,
            carryout => \eeprom.n3756\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2357_10_lut_LC_16_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27008\,
            in2 => \N__25079\,
            in3 => \N__25040\,
            lcout => \eeprom.n3578_adj_361\,
            ltout => OPEN,
            carryin => \bfn_16_18_0_\,
            carryout => \eeprom.n3757\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2357_11_lut_LC_16_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27016\,
            in2 => \N__25037\,
            in3 => \N__25001\,
            lcout => \eeprom.n3577_adj_359\,
            ltout => OPEN,
            carryin => \eeprom.n3757\,
            carryout => \eeprom.n3758\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2357_12_lut_LC_16_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27009\,
            in2 => \N__24998\,
            in3 => \N__24956\,
            lcout => \eeprom.n3576_adj_358\,
            ltout => OPEN,
            carryin => \eeprom.n3758\,
            carryout => \eeprom.n3759\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2357_13_lut_LC_16_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27017\,
            in2 => \N__24953\,
            in3 => \N__24926\,
            lcout => \eeprom.n3575_adj_357\,
            ltout => OPEN,
            carryin => \eeprom.n3759\,
            carryout => \eeprom.n3760\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2357_14_lut_LC_16_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24923\,
            in2 => \N__27194\,
            in3 => \N__24887\,
            lcout => \eeprom.n3574_adj_356\,
            ltout => OPEN,
            carryin => \eeprom.n3760\,
            carryout => \eeprom.n3761\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2357_15_lut_LC_16_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24883\,
            in2 => \N__27192\,
            in3 => \N__24851\,
            lcout => \eeprom.n3573_adj_355\,
            ltout => OPEN,
            carryin => \eeprom.n3761\,
            carryout => \eeprom.n3762\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2357_16_lut_LC_16_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25462\,
            in2 => \N__27195\,
            in3 => \N__25433\,
            lcout => \eeprom.n3572_adj_354\,
            ltout => OPEN,
            carryin => \eeprom.n3762\,
            carryout => \eeprom.n3763\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2357_17_lut_LC_16_18_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25430\,
            in2 => \N__27193\,
            in3 => \N__25397\,
            lcout => \eeprom.n3571_adj_353\,
            ltout => OPEN,
            carryin => \eeprom.n3763\,
            carryout => \eeprom.n3764\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2357_18_lut_LC_16_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26988\,
            in2 => \N__25389\,
            in3 => \N__25352\,
            lcout => \eeprom.n3570_adj_349\,
            ltout => OPEN,
            carryin => \bfn_16_19_0_\,
            carryout => \eeprom.n3765\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2357_19_lut_LC_16_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25348\,
            in2 => \N__27186\,
            in3 => \N__25319\,
            lcout => \eeprom.n3569_adj_348\,
            ltout => OPEN,
            carryin => \eeprom.n3765\,
            carryout => \eeprom.n3766\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2357_20_lut_LC_16_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25316\,
            in2 => \N__27189\,
            in3 => \N__25280\,
            lcout => \eeprom.n3568_adj_347\,
            ltout => OPEN,
            carryin => \eeprom.n3766\,
            carryout => \eeprom.n3767\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2357_21_lut_LC_16_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25277\,
            in2 => \N__27187\,
            in3 => \N__25244\,
            lcout => \eeprom.n3567_adj_341\,
            ltout => OPEN,
            carryin => \eeprom.n3767\,
            carryout => \eeprom.n3768\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2357_22_lut_LC_16_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25241\,
            in2 => \N__27190\,
            in3 => \N__25202\,
            lcout => \eeprom.n3566_adj_340\,
            ltout => OPEN,
            carryin => \eeprom.n3768\,
            carryout => \eeprom.n3769\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2357_23_lut_LC_16_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25198\,
            in2 => \N__27188\,
            in3 => \N__25769\,
            lcout => \eeprom.n3565_adj_338\,
            ltout => OPEN,
            carryin => \eeprom.n3769\,
            carryout => \eeprom.n3770\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2357_24_lut_LC_16_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25762\,
            in2 => \N__27191\,
            in3 => \N__25727\,
            lcout => \eeprom.n3564_adj_337\,
            ltout => OPEN,
            carryin => \eeprom.n3770\,
            carryout => \eeprom.n3771\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2357_25_lut_LC_16_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001000001100000"
        )
    port map (
            in0 => \N__26998\,
            in1 => \N__25724\,
            in2 => \N__25706\,
            in3 => \N__25574\,
            lcout => \eeprom.n4765\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.add_938_2_lut_LC_16_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25877\,
            in2 => \_gnd_net_\,
            in3 => \N__25565\,
            lcout => \eeprom.n1353\,
            ltout => OPEN,
            carryin => \bfn_16_20_0_\,
            carryout => \eeprom.n3510\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.add_938_3_lut_LC_16_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25912\,
            in2 => \N__27185\,
            in3 => \N__25562\,
            lcout => \eeprom.n1352\,
            ltout => OPEN,
            carryin => \eeprom.n3510\,
            carryout => \eeprom.n3511\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.add_938_4_lut_LC_16_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25559\,
            in2 => \_gnd_net_\,
            in3 => \N__25538\,
            lcout => \eeprom.n1351\,
            ltout => OPEN,
            carryin => \eeprom.n3511\,
            carryout => \eeprom.n3512\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.add_938_5_lut_LC_16_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__25993\,
            in3 => \N__25535\,
            lcout => \eeprom.n1350\,
            ltout => OPEN,
            carryin => \eeprom.n3512\,
            carryout => \eeprom.n3513\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.add_938_6_lut_LC_16_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__25532\,
            in3 => \N__25505\,
            lcout => \eeprom.n1349\,
            ltout => OPEN,
            carryin => \eeprom.n3513\,
            carryout => \eeprom.n3514\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.add_938_7_lut_LC_16_20_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25501\,
            in2 => \_gnd_net_\,
            in3 => \N__25469\,
            lcout => \eeprom.n1348\,
            ltout => OPEN,
            carryin => \eeprom.n3514\,
            carryout => \eeprom.n3515\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.add_938_8_lut_LC_16_20_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26057\,
            in2 => \_gnd_net_\,
            in3 => \N__26021\,
            lcout => \eeprom.n1347\,
            ltout => OPEN,
            carryin => \eeprom.n3515\,
            carryout => \eeprom.n3516\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.add_938_9_lut_LC_16_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__26987\,
            in1 => \N__26018\,
            in2 => \_gnd_net_\,
            in3 => \N__26003\,
            lcout => \eeprom.n1346\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2447_3_lut_LC_16_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000000111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26000\,
            in2 => \N__25834\,
            in3 => \N__25994\,
            lcout => \eeprom.n3715_adj_441\,
            ltout => \eeprom.n3715_adj_441_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i4068_1_lut_LC_16_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__25961\,
            in3 => \_gnd_net_\,
            lcout => \eeprom.n4912\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i4083_2_lut_LC_16_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__25835\,
            in3 => \N__25948\,
            lcout => \eeprom.n3711_adj_456\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2449_3_lut_LC_16_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25925\,
            in2 => \N__25919\,
            in3 => \N__25825\,
            lcout => \eeprom.n3717_adj_438\,
            ltout => \eeprom.n3717_adj_438_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i4062_1_lut_LC_16_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__25892\,
            in3 => \_gnd_net_\,
            lcout => \eeprom.n4906\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2450_rep_1_3_lut_LC_16_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100110011"
        )
    port map (
            in0 => \N__25883\,
            in1 => \N__25875\,
            in2 => \_gnd_net_\,
            in3 => \N__25824\,
            lcout => \eeprom.n4766\,
            ltout => \eeprom.n4766_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i4059_1_lut_LC_16_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__26399\,
            in3 => \_gnd_net_\,
            lcout => \eeprom.n4903\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2022_2_lut_LC_16_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26386\,
            in2 => \_gnd_net_\,
            in3 => \N__26342\,
            lcout => \eeprom.n3086\,
            ltout => OPEN,
            carryin => \bfn_16_23_0_\,
            carryout => \eeprom.n3649\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2022_3_lut_LC_16_23_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26936\,
            in2 => \N__26335\,
            in3 => \N__26300\,
            lcout => \eeprom.n3085\,
            ltout => OPEN,
            carryin => \eeprom.n3649\,
            carryout => \eeprom.n3650\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2022_4_lut_LC_16_23_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__26297\,
            in3 => \N__26252\,
            lcout => \eeprom.n3084\,
            ltout => OPEN,
            carryin => \eeprom.n3650\,
            carryout => \eeprom.n3651\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2022_5_lut_LC_16_23_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__26249\,
            in3 => \N__26198\,
            lcout => \eeprom.n3083\,
            ltout => OPEN,
            carryin => \eeprom.n3651\,
            carryout => \eeprom.n3652\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2022_6_lut_LC_16_23_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__26195\,
            in3 => \N__26153\,
            lcout => \eeprom.n3082\,
            ltout => OPEN,
            carryin => \eeprom.n3652\,
            carryout => \eeprom.n3653\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2022_7_lut_LC_16_23_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__26150\,
            in3 => \N__26099\,
            lcout => \eeprom.n3081\,
            ltout => OPEN,
            carryin => \eeprom.n3653\,
            carryout => \eeprom.n3654\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2022_8_lut_LC_16_23_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__26096\,
            in3 => \N__26060\,
            lcout => \eeprom.n3080\,
            ltout => OPEN,
            carryin => \eeprom.n3654\,
            carryout => \eeprom.n3655\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2022_9_lut_LC_16_23_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26937\,
            in2 => \N__26705\,
            in3 => \N__26675\,
            lcout => \eeprom.n3079\,
            ltout => OPEN,
            carryin => \eeprom.n3655\,
            carryout => \eeprom.n3656\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2022_10_lut_LC_16_24_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26672\,
            in2 => \N__27073\,
            in3 => \N__26642\,
            lcout => \eeprom.n3078\,
            ltout => OPEN,
            carryin => \bfn_16_24_0_\,
            carryout => \eeprom.n3657\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2022_11_lut_LC_16_24_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26885\,
            in2 => \N__26634\,
            in3 => \N__26597\,
            lcout => \eeprom.n3077\,
            ltout => OPEN,
            carryin => \eeprom.n3657\,
            carryout => \eeprom.n3658\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2022_12_lut_LC_16_24_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26586\,
            in2 => \N__27074\,
            in3 => \N__26546\,
            lcout => \eeprom.n3076\,
            ltout => OPEN,
            carryin => \eeprom.n3658\,
            carryout => \eeprom.n3659\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2022_13_lut_LC_16_24_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26538\,
            in2 => \N__27077\,
            in3 => \N__26516\,
            lcout => \eeprom.n3075\,
            ltout => OPEN,
            carryin => \eeprom.n3659\,
            carryout => \eeprom.n3660\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2022_14_lut_LC_16_24_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26511\,
            in2 => \N__27075\,
            in3 => \N__26471\,
            lcout => \eeprom.n3074\,
            ltout => OPEN,
            carryin => \eeprom.n3660\,
            carryout => \eeprom.n3661\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2022_15_lut_LC_16_24_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26467\,
            in2 => \N__27078\,
            in3 => \N__26429\,
            lcout => \eeprom.n3073\,
            ltout => OPEN,
            carryin => \eeprom.n3661\,
            carryout => \eeprom.n3662\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2022_16_lut_LC_16_24_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26426\,
            in2 => \N__27076\,
            in3 => \N__28076\,
            lcout => \eeprom.n3072\,
            ltout => OPEN,
            carryin => \eeprom.n3662\,
            carryout => \eeprom.n3663\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2022_17_lut_LC_16_24_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28073\,
            in2 => \N__27079\,
            in3 => \N__28037\,
            lcout => \eeprom.n3071\,
            ltout => OPEN,
            carryin => \eeprom.n3663\,
            carryout => \eeprom.n3664\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2022_18_lut_LC_16_25_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28034\,
            in2 => \N__26880\,
            in3 => \N__27998\,
            lcout => \eeprom.n3070\,
            ltout => OPEN,
            carryin => \bfn_16_25_0_\,
            carryout => \eeprom.n3665\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2022_19_lut_LC_16_25_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27995\,
            in2 => \N__26881\,
            in3 => \N__27950\,
            lcout => \eeprom.n3069\,
            ltout => OPEN,
            carryin => \eeprom.n3665\,
            carryout => \eeprom.n3666\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2022_20_lut_LC_16_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001000001100000"
        )
    port map (
            in0 => \N__26764\,
            in1 => \N__27947\,
            in2 => \N__27920\,
            in3 => \N__27809\,
            lcout => \eeprom.n3100\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_16_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;
